module basic_2500_25000_3000_125_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_463,In_95);
nor U1 (N_1,In_1342,In_1979);
or U2 (N_2,In_876,In_2279);
or U3 (N_3,In_592,In_416);
or U4 (N_4,In_2130,In_2220);
or U5 (N_5,In_1779,In_1075);
nor U6 (N_6,In_651,In_121);
nand U7 (N_7,In_787,In_1518);
nand U8 (N_8,In_679,In_1078);
or U9 (N_9,In_2188,In_1173);
and U10 (N_10,In_658,In_1437);
nor U11 (N_11,In_1562,In_469);
and U12 (N_12,In_803,In_271);
xor U13 (N_13,In_1899,In_1858);
xor U14 (N_14,In_2000,In_1586);
nand U15 (N_15,In_1423,In_1833);
xor U16 (N_16,In_2347,In_405);
or U17 (N_17,In_561,In_2266);
xnor U18 (N_18,In_1660,In_1553);
and U19 (N_19,In_602,In_638);
xor U20 (N_20,In_650,In_1972);
and U21 (N_21,In_1186,In_1396);
xnor U22 (N_22,In_1636,In_1961);
nor U23 (N_23,In_2428,In_599);
or U24 (N_24,In_2263,In_1687);
nand U25 (N_25,In_2245,In_2034);
xor U26 (N_26,In_2372,In_591);
or U27 (N_27,In_760,In_634);
and U28 (N_28,In_395,In_1294);
and U29 (N_29,In_1000,In_1135);
nor U30 (N_30,In_1603,In_1790);
and U31 (N_31,In_2168,In_472);
nand U32 (N_32,In_2275,In_1650);
and U33 (N_33,In_2499,In_2294);
nand U34 (N_34,In_1305,In_1669);
and U35 (N_35,In_117,In_988);
xnor U36 (N_36,In_179,In_1071);
or U37 (N_37,In_862,In_1450);
xnor U38 (N_38,In_105,In_1168);
nand U39 (N_39,In_805,In_826);
xor U40 (N_40,In_1814,In_114);
nand U41 (N_41,In_144,In_2274);
and U42 (N_42,In_1213,In_819);
or U43 (N_43,In_1343,In_1733);
nor U44 (N_44,In_1314,In_2158);
and U45 (N_45,In_727,In_1737);
or U46 (N_46,In_1479,In_1234);
nor U47 (N_47,In_1865,In_640);
and U48 (N_48,In_2196,In_1204);
xnor U49 (N_49,In_2169,In_484);
or U50 (N_50,In_198,In_1241);
nand U51 (N_51,In_1237,In_967);
or U52 (N_52,In_109,In_1292);
nand U53 (N_53,In_219,In_1582);
xor U54 (N_54,In_1291,In_2110);
nand U55 (N_55,In_1010,In_942);
xnor U56 (N_56,In_623,In_2173);
xor U57 (N_57,In_1409,In_2174);
or U58 (N_58,In_1716,In_2117);
or U59 (N_59,In_1220,In_995);
xor U60 (N_60,In_2067,In_2481);
and U61 (N_61,In_2309,In_549);
and U62 (N_62,In_2308,In_858);
and U63 (N_63,In_1963,In_196);
or U64 (N_64,In_2190,In_1251);
nand U65 (N_65,In_1609,In_936);
or U66 (N_66,In_1888,In_2445);
nor U67 (N_67,In_781,In_1602);
xnor U68 (N_68,In_2126,In_1550);
nand U69 (N_69,In_474,In_550);
nand U70 (N_70,In_2370,In_1465);
nor U71 (N_71,In_1785,In_1478);
nor U72 (N_72,In_361,In_2446);
nand U73 (N_73,In_2082,In_2291);
and U74 (N_74,In_353,In_2064);
nand U75 (N_75,In_1723,In_820);
nor U76 (N_76,In_1784,In_1049);
or U77 (N_77,In_1086,In_1445);
xor U78 (N_78,In_1548,In_149);
or U79 (N_79,In_1613,In_300);
and U80 (N_80,In_991,In_2120);
xor U81 (N_81,In_835,In_1632);
xor U82 (N_82,In_6,In_465);
and U83 (N_83,In_1530,In_2185);
and U84 (N_84,In_236,In_517);
nor U85 (N_85,In_1404,In_918);
or U86 (N_86,In_990,In_50);
xor U87 (N_87,In_148,In_122);
and U88 (N_88,In_1015,In_2334);
and U89 (N_89,In_2475,In_2189);
nand U90 (N_90,In_2198,In_1832);
nor U91 (N_91,In_1845,In_1317);
nor U92 (N_92,In_2460,In_1035);
and U93 (N_93,In_277,In_2332);
and U94 (N_94,In_884,In_2268);
xnor U95 (N_95,In_16,In_2039);
nand U96 (N_96,In_132,In_1993);
or U97 (N_97,In_230,In_718);
and U98 (N_98,In_2212,In_2097);
xnor U99 (N_99,In_719,In_2447);
nor U100 (N_100,In_130,In_863);
nor U101 (N_101,In_630,In_2317);
and U102 (N_102,In_245,In_1389);
nand U103 (N_103,In_272,In_1561);
nand U104 (N_104,In_226,In_362);
and U105 (N_105,In_1934,In_1635);
nand U106 (N_106,In_2214,In_2250);
and U107 (N_107,In_2001,In_204);
and U108 (N_108,In_1432,In_331);
and U109 (N_109,In_22,In_2116);
or U110 (N_110,In_808,In_2339);
or U111 (N_111,In_2006,In_1647);
nand U112 (N_112,In_1822,In_323);
or U113 (N_113,In_1643,In_986);
or U114 (N_114,In_1120,In_1202);
or U115 (N_115,In_2399,In_1672);
nor U116 (N_116,In_427,In_294);
xnor U117 (N_117,In_1750,In_984);
or U118 (N_118,In_1796,In_276);
or U119 (N_119,In_1986,In_770);
or U120 (N_120,In_346,In_1108);
nor U121 (N_121,In_2397,In_2432);
and U122 (N_122,In_2345,In_406);
and U123 (N_123,In_491,In_1286);
or U124 (N_124,In_1394,In_1703);
xnor U125 (N_125,In_481,In_1744);
or U126 (N_126,In_2218,In_1329);
or U127 (N_127,In_1434,In_921);
nand U128 (N_128,In_1803,In_1982);
and U129 (N_129,In_588,In_1715);
nor U130 (N_130,In_291,In_1365);
nand U131 (N_131,In_716,In_264);
xor U132 (N_132,In_2192,In_2316);
xnor U133 (N_133,In_227,In_2127);
xnor U134 (N_134,In_1501,In_1459);
and U135 (N_135,In_1496,In_573);
nor U136 (N_136,In_2155,In_486);
nand U137 (N_137,In_1084,In_115);
or U138 (N_138,In_2139,In_2448);
or U139 (N_139,In_1908,In_1812);
and U140 (N_140,In_2145,In_1416);
xor U141 (N_141,In_213,In_315);
or U142 (N_142,In_313,In_1136);
xor U143 (N_143,In_120,In_2299);
nor U144 (N_144,In_2438,In_170);
and U145 (N_145,In_2202,In_962);
nand U146 (N_146,In_440,In_2012);
nand U147 (N_147,In_2068,In_1412);
and U148 (N_148,In_2377,In_4);
nor U149 (N_149,In_1658,In_2051);
and U150 (N_150,In_1405,In_1217);
or U151 (N_151,In_1439,In_153);
nand U152 (N_152,In_721,In_206);
nor U153 (N_153,In_2261,In_37);
xnor U154 (N_154,In_1142,In_1903);
and U155 (N_155,In_1639,In_1770);
or U156 (N_156,In_521,In_1064);
and U157 (N_157,In_586,In_1990);
and U158 (N_158,In_2231,In_1746);
xnor U159 (N_159,In_2426,In_1567);
xor U160 (N_160,In_1355,In_1034);
or U161 (N_161,In_1498,In_375);
nor U162 (N_162,In_1623,In_838);
nor U163 (N_163,In_377,In_2376);
and U164 (N_164,In_365,In_169);
and U165 (N_165,In_2048,In_2373);
nand U166 (N_166,In_669,In_1181);
nand U167 (N_167,In_1483,In_1490);
or U168 (N_168,In_135,In_1066);
nor U169 (N_169,In_2137,In_1977);
and U170 (N_170,In_1360,In_1257);
xnor U171 (N_171,In_2490,In_767);
nor U172 (N_172,In_870,In_1742);
or U173 (N_173,In_828,In_608);
or U174 (N_174,In_1766,In_857);
and U175 (N_175,In_1968,In_1644);
nor U176 (N_176,In_2153,In_580);
or U177 (N_177,In_1587,In_703);
or U178 (N_178,In_1575,In_1617);
nand U179 (N_179,In_848,In_2161);
nand U180 (N_180,In_35,In_341);
nor U181 (N_181,In_1863,In_2437);
or U182 (N_182,In_1067,In_273);
and U183 (N_183,In_1208,In_1776);
xor U184 (N_184,In_2364,In_840);
nand U185 (N_185,In_418,In_419);
and U186 (N_186,In_2076,In_384);
xnor U187 (N_187,In_801,In_495);
nand U188 (N_188,In_2285,In_951);
or U189 (N_189,In_2369,In_1420);
and U190 (N_190,In_374,In_1390);
xor U191 (N_191,In_1093,In_185);
and U192 (N_192,In_2482,In_454);
or U193 (N_193,In_885,In_434);
and U194 (N_194,In_1585,In_947);
xor U195 (N_195,In_112,In_756);
and U196 (N_196,In_1267,In_1943);
nor U197 (N_197,In_17,In_940);
nand U198 (N_198,In_255,In_1134);
nor U199 (N_199,In_2394,In_1905);
and U200 (N_200,In_2464,In_846);
nor U201 (N_201,In_916,In_1451);
or U202 (N_202,In_1333,N_34);
nor U203 (N_203,In_500,In_261);
xnor U204 (N_204,In_758,In_184);
or U205 (N_205,In_2343,In_39);
nor U206 (N_206,In_1807,In_501);
or U207 (N_207,N_66,N_128);
nand U208 (N_208,In_2203,In_139);
nand U209 (N_209,In_1144,In_373);
nand U210 (N_210,In_973,N_78);
or U211 (N_211,In_1763,In_1732);
or U212 (N_212,In_642,In_794);
nor U213 (N_213,In_1211,In_1370);
xor U214 (N_214,In_1953,In_1873);
and U215 (N_215,In_359,In_391);
nor U216 (N_216,In_2409,In_665);
nand U217 (N_217,N_18,N_23);
nand U218 (N_218,In_1101,In_1275);
nand U219 (N_219,In_1346,In_730);
nand U220 (N_220,In_1053,In_1191);
or U221 (N_221,In_1788,In_1449);
and U222 (N_222,In_2259,In_2170);
and U223 (N_223,In_534,In_2270);
nor U224 (N_224,In_2267,In_287);
nand U225 (N_225,N_79,In_1826);
nor U226 (N_226,In_1328,In_620);
or U227 (N_227,In_2472,In_1726);
xnor U228 (N_228,In_919,In_161);
and U229 (N_229,In_337,In_1594);
xor U230 (N_230,In_1569,In_2183);
nor U231 (N_231,N_180,In_351);
or U232 (N_232,In_2111,In_285);
or U233 (N_233,N_61,In_1901);
or U234 (N_234,In_1523,In_2234);
nor U235 (N_235,In_1640,In_1062);
or U236 (N_236,In_2453,In_2119);
nor U237 (N_237,In_2427,In_2430);
nand U238 (N_238,N_71,In_1162);
nand U239 (N_239,In_1227,In_2027);
nor U240 (N_240,In_893,In_2099);
nor U241 (N_241,In_334,N_42);
or U242 (N_242,In_2381,In_1127);
or U243 (N_243,In_997,N_145);
xor U244 (N_244,In_507,In_177);
nand U245 (N_245,In_1487,In_1040);
or U246 (N_246,In_1852,In_660);
nand U247 (N_247,In_1590,In_448);
and U248 (N_248,In_663,In_2113);
and U249 (N_249,In_688,In_1753);
or U250 (N_250,In_1327,In_2239);
xor U251 (N_251,In_1301,In_2422);
nand U252 (N_252,In_254,In_1068);
and U253 (N_253,In_1502,In_1089);
xnor U254 (N_254,In_576,In_143);
and U255 (N_255,In_1731,In_720);
or U256 (N_256,In_666,In_1696);
nor U257 (N_257,In_766,In_1270);
xnor U258 (N_258,In_1942,In_456);
nor U259 (N_259,In_583,In_1676);
nand U260 (N_260,In_307,In_1201);
or U261 (N_261,In_60,In_248);
and U262 (N_262,N_171,In_2050);
nand U263 (N_263,In_1433,In_233);
xor U264 (N_264,In_2295,In_452);
nor U265 (N_265,In_386,N_104);
nand U266 (N_266,N_39,In_2433);
and U267 (N_267,In_1929,In_1051);
xnor U268 (N_268,In_1399,In_852);
nor U269 (N_269,In_1094,In_649);
or U270 (N_270,In_2181,In_2069);
xor U271 (N_271,In_1545,In_1386);
nand U272 (N_272,In_1453,In_606);
or U273 (N_273,In_853,In_1046);
xnor U274 (N_274,In_1568,In_306);
nand U275 (N_275,N_59,In_554);
xor U276 (N_276,In_2093,In_1005);
nand U277 (N_277,In_321,In_1098);
and U278 (N_278,In_626,In_1271);
nor U279 (N_279,In_447,In_2213);
nor U280 (N_280,In_843,In_625);
nor U281 (N_281,In_2491,In_30);
and U282 (N_282,N_101,In_529);
and U283 (N_283,In_311,In_281);
nand U284 (N_284,In_1383,In_1214);
or U285 (N_285,In_1302,In_2455);
xor U286 (N_286,N_65,In_1976);
nor U287 (N_287,In_43,In_1456);
and U288 (N_288,In_804,In_2469);
or U289 (N_289,N_27,In_818);
nand U290 (N_290,In_1016,In_1843);
or U291 (N_291,In_2028,In_1713);
nor U292 (N_292,In_2016,In_1427);
and U293 (N_293,In_251,In_1242);
or U294 (N_294,In_1042,In_222);
xnor U295 (N_295,In_1277,In_2289);
nor U296 (N_296,In_88,In_1447);
or U297 (N_297,In_1472,In_1653);
and U298 (N_298,In_1984,In_1893);
nand U299 (N_299,In_1930,In_968);
and U300 (N_300,In_2272,In_829);
or U301 (N_301,In_1918,In_119);
nand U302 (N_302,In_250,In_193);
xor U303 (N_303,In_1531,In_1368);
nor U304 (N_304,In_2303,In_1323);
nor U305 (N_305,In_1714,In_772);
and U306 (N_306,In_127,In_1679);
and U307 (N_307,In_157,In_303);
or U308 (N_308,In_1077,In_1555);
nor U309 (N_309,N_105,In_1824);
and U310 (N_310,In_1406,In_466);
and U311 (N_311,In_1090,In_1532);
and U312 (N_312,In_1648,In_1978);
and U313 (N_313,In_935,In_546);
nor U314 (N_314,In_1563,In_1526);
nand U315 (N_315,In_2252,In_570);
and U316 (N_316,In_1738,In_1190);
and U317 (N_317,In_24,In_417);
xnor U318 (N_318,In_1441,In_902);
nand U319 (N_319,In_302,In_851);
xnor U320 (N_320,In_1484,In_837);
xnor U321 (N_321,In_2121,N_26);
and U322 (N_322,In_154,In_113);
and U323 (N_323,In_1137,In_979);
xnor U324 (N_324,In_64,In_2312);
xor U325 (N_325,In_431,In_1158);
and U326 (N_326,In_2049,In_1400);
nor U327 (N_327,In_1810,In_423);
and U328 (N_328,In_1797,In_52);
nor U329 (N_329,In_559,In_1897);
or U330 (N_330,In_971,In_1678);
and U331 (N_331,In_2166,N_146);
nand U332 (N_332,In_2434,In_522);
xnor U333 (N_333,In_2487,In_2304);
nand U334 (N_334,In_1900,In_668);
nand U335 (N_335,In_933,In_2114);
and U336 (N_336,In_1611,In_998);
or U337 (N_337,In_1988,In_1265);
xnor U338 (N_338,In_1761,In_1534);
or U339 (N_339,In_698,N_87);
and U340 (N_340,In_1019,In_502);
and U341 (N_341,In_393,In_2260);
nand U342 (N_342,In_569,In_2389);
or U343 (N_343,In_49,N_60);
nor U344 (N_344,In_2492,In_1290);
xor U345 (N_345,In_430,In_761);
and U346 (N_346,N_142,In_404);
nand U347 (N_347,In_350,N_115);
nor U348 (N_348,In_1140,N_25);
nand U349 (N_349,In_2371,In_1172);
and U350 (N_350,In_367,In_795);
nand U351 (N_351,In_643,In_1350);
nor U352 (N_352,In_408,In_1730);
and U353 (N_353,N_117,In_86);
nor U354 (N_354,In_2219,In_260);
nor U355 (N_355,In_145,In_2305);
and U356 (N_356,In_344,In_1461);
or U357 (N_357,In_1004,In_2342);
xnor U358 (N_358,In_499,In_709);
or U359 (N_359,In_13,In_907);
nand U360 (N_360,In_1454,In_2094);
nand U361 (N_361,In_1503,In_478);
or U362 (N_362,In_1114,In_2329);
nand U363 (N_363,In_1741,In_1076);
nand U364 (N_364,In_519,In_2243);
and U365 (N_365,N_58,In_2035);
xor U366 (N_366,In_1970,In_221);
and U367 (N_367,In_2463,In_1092);
and U368 (N_368,In_778,In_1618);
and U369 (N_369,In_1673,In_924);
nor U370 (N_370,N_141,In_96);
or U371 (N_371,In_1957,In_195);
nor U372 (N_372,In_187,N_160);
xnor U373 (N_373,In_1707,In_518);
or U374 (N_374,N_24,In_1119);
nor U375 (N_375,In_619,In_687);
and U376 (N_376,In_232,In_1827);
nand U377 (N_377,In_1711,In_1748);
xor U378 (N_378,In_2497,In_2468);
xor U379 (N_379,In_305,In_326);
and U380 (N_380,In_125,In_26);
nand U381 (N_381,In_1388,In_832);
and U382 (N_382,In_777,N_32);
nor U383 (N_383,In_1682,In_791);
xnor U384 (N_384,N_197,In_163);
xnor U385 (N_385,In_107,In_711);
nand U386 (N_386,In_1699,In_201);
and U387 (N_387,In_963,In_2406);
or U388 (N_388,In_1991,In_1233);
or U389 (N_389,In_2178,In_2106);
and U390 (N_390,N_97,In_1219);
or U391 (N_391,In_1837,In_542);
and U392 (N_392,In_2040,In_1309);
xnor U393 (N_393,In_2199,In_1973);
nor U394 (N_394,In_81,In_1922);
or U395 (N_395,In_887,In_2375);
nand U396 (N_396,In_2327,In_1584);
xor U397 (N_397,In_2205,In_58);
xor U398 (N_398,In_2473,In_1250);
xor U399 (N_399,In_1727,In_1870);
xor U400 (N_400,In_2353,In_182);
xor U401 (N_401,In_1014,In_2314);
and U402 (N_402,In_2368,In_1285);
or U403 (N_403,In_68,N_127);
xor U404 (N_404,In_1011,In_1133);
nand U405 (N_405,In_2144,N_69);
nand U406 (N_406,N_229,In_732);
nor U407 (N_407,N_323,N_309);
xnor U408 (N_408,In_627,In_745);
and U409 (N_409,In_2379,In_1146);
xnor U410 (N_410,In_2336,In_156);
nand U411 (N_411,In_594,N_129);
nand U412 (N_412,N_5,In_2095);
nand U413 (N_413,N_98,In_845);
xor U414 (N_414,In_235,N_159);
nor U415 (N_415,In_1180,In_1818);
or U416 (N_416,In_1107,N_396);
or U417 (N_417,In_2156,In_771);
and U418 (N_418,In_1952,In_764);
and U419 (N_419,In_2367,In_1780);
xor U420 (N_420,In_864,N_370);
nand U421 (N_421,In_1598,In_1628);
xor U422 (N_422,In_2378,In_263);
nor U423 (N_423,In_681,N_14);
and U424 (N_424,In_253,In_1965);
or U425 (N_425,In_2032,In_783);
nand U426 (N_426,N_272,N_319);
nand U427 (N_427,N_174,In_661);
nand U428 (N_428,In_1507,N_364);
nand U429 (N_429,In_2200,In_8);
nand U430 (N_430,In_992,In_2385);
nand U431 (N_431,In_1698,N_243);
and U432 (N_432,In_2388,N_10);
and U433 (N_433,N_148,In_978);
xnor U434 (N_434,In_1911,N_17);
xnor U435 (N_435,In_1633,In_581);
and U436 (N_436,In_1994,In_409);
or U437 (N_437,In_1947,In_715);
nand U438 (N_438,N_390,In_538);
and U439 (N_439,In_2087,In_953);
or U440 (N_440,In_136,In_1709);
nand U441 (N_441,In_274,In_1356);
nand U442 (N_442,In_2123,In_1033);
and U443 (N_443,In_1684,In_487);
or U444 (N_444,In_1683,In_129);
nor U445 (N_445,In_2280,N_111);
nor U446 (N_446,In_1874,In_1504);
xnor U447 (N_447,In_584,In_1558);
or U448 (N_448,In_1996,In_1031);
or U449 (N_449,In_1573,In_1956);
xor U450 (N_450,In_1806,In_1815);
nor U451 (N_451,In_536,In_1228);
nor U452 (N_452,In_1247,In_1467);
xnor U453 (N_453,In_2459,In_2151);
or U454 (N_454,In_116,N_155);
and U455 (N_455,N_382,In_1123);
and U456 (N_456,In_1969,N_339);
nor U457 (N_457,In_2154,In_1366);
nor U458 (N_458,In_2056,In_684);
and U459 (N_459,In_2301,In_2357);
and U460 (N_460,In_901,In_1777);
nand U461 (N_461,In_2298,In_567);
and U462 (N_462,In_692,N_261);
or U463 (N_463,In_282,In_1869);
xnor U464 (N_464,In_1606,In_1909);
or U465 (N_465,In_1872,N_40);
or U466 (N_466,In_167,In_566);
nor U467 (N_467,In_1566,In_445);
xor U468 (N_468,N_336,In_457);
and U469 (N_469,In_2177,N_114);
and U470 (N_470,In_1725,In_289);
or U471 (N_471,In_1236,N_322);
and U472 (N_472,In_421,N_143);
nand U473 (N_473,In_937,In_724);
xnor U474 (N_474,In_241,In_2152);
nand U475 (N_475,In_2062,In_2398);
nand U476 (N_476,In_2251,In_1184);
nor U477 (N_477,In_357,In_1293);
and U478 (N_478,In_308,In_755);
and U479 (N_479,In_691,In_1087);
xnor U480 (N_480,In_2148,In_74);
xor U481 (N_481,In_2486,In_980);
nor U482 (N_482,In_1923,In_1167);
and U483 (N_483,N_247,In_2079);
or U484 (N_484,N_328,In_664);
or U485 (N_485,In_1549,In_2248);
xnor U486 (N_486,In_540,In_917);
xnor U487 (N_487,In_714,In_957);
xor U488 (N_488,In_1557,In_780);
nor U489 (N_489,In_891,In_338);
and U490 (N_490,In_200,In_1884);
or U491 (N_491,In_2090,N_321);
nor U492 (N_492,In_2017,N_140);
xnor U493 (N_493,N_90,N_244);
or U494 (N_494,In_733,In_865);
xnor U495 (N_495,In_19,In_1331);
or U496 (N_496,In_2282,In_2004);
xor U497 (N_497,In_390,In_2057);
nor U498 (N_498,In_1649,In_2041);
nand U499 (N_499,In_742,N_192);
xnor U500 (N_500,In_1050,In_762);
or U501 (N_501,In_356,In_2337);
and U502 (N_502,N_359,In_1896);
or U503 (N_503,In_2058,N_337);
nor U504 (N_504,In_180,In_1283);
nor U505 (N_505,In_2454,In_1686);
nand U506 (N_506,In_304,In_1332);
nor U507 (N_507,N_367,In_2403);
and U508 (N_508,In_1778,In_1511);
nand U509 (N_509,In_2391,In_1183);
xnor U510 (N_510,In_1515,In_1579);
nor U511 (N_511,In_2488,In_220);
xor U512 (N_512,In_2133,In_320);
or U513 (N_513,In_1048,In_1680);
or U514 (N_514,In_69,In_1565);
and U515 (N_515,N_214,In_2466);
xor U516 (N_516,In_1431,In_355);
xor U517 (N_517,In_1659,In_535);
and U518 (N_518,In_1297,N_80);
xnor U519 (N_519,In_1351,In_779);
nor U520 (N_520,In_218,In_1410);
and U521 (N_521,In_246,In_2390);
and U522 (N_522,N_208,In_1408);
nor U523 (N_523,In_782,In_674);
nor U524 (N_524,In_2351,In_1637);
nand U525 (N_525,In_1799,In_2201);
and U526 (N_526,In_1058,In_2);
or U527 (N_527,In_1912,In_1069);
nor U528 (N_528,In_676,In_1921);
nor U529 (N_529,N_9,In_577);
or U530 (N_530,In_2167,N_266);
and U531 (N_531,In_1085,In_1898);
xnor U532 (N_532,In_397,In_635);
nor U533 (N_533,In_2410,In_1185);
xor U534 (N_534,N_184,In_605);
and U535 (N_535,N_37,N_7);
nor U536 (N_536,In_1828,In_533);
nand U537 (N_537,In_1196,In_283);
nand U538 (N_538,In_1559,In_823);
nand U539 (N_539,In_1032,N_294);
xor U540 (N_540,In_1691,In_1831);
and U541 (N_541,In_799,In_568);
and U542 (N_542,In_2011,In_475);
nor U543 (N_543,In_747,N_63);
nor U544 (N_544,In_1794,In_1460);
and U545 (N_545,In_280,In_886);
nand U546 (N_546,N_151,N_385);
nand U547 (N_547,In_2414,N_162);
nand U548 (N_548,In_2227,In_671);
nand U549 (N_549,In_1268,N_394);
and U550 (N_550,In_1599,In_1139);
nor U551 (N_551,N_347,In_562);
nand U552 (N_552,In_1955,In_1189);
and U553 (N_553,In_1152,In_1306);
xor U554 (N_554,In_1195,In_257);
nor U555 (N_555,In_2240,In_631);
nor U556 (N_556,In_752,In_1436);
nor U557 (N_557,N_248,N_371);
xnor U558 (N_558,In_2101,In_1174);
or U559 (N_559,N_373,In_435);
nor U560 (N_560,In_1103,In_67);
nand U561 (N_561,N_303,In_1153);
xor U562 (N_562,In_25,N_259);
xor U563 (N_563,In_212,In_1206);
or U564 (N_564,In_76,N_195);
nand U565 (N_565,In_890,N_122);
nor U566 (N_566,In_1933,In_90);
nand U567 (N_567,In_55,N_222);
xnor U568 (N_568,In_1809,In_2271);
or U569 (N_569,In_523,In_217);
nor U570 (N_570,In_1348,N_113);
nand U571 (N_571,In_1052,In_722);
or U572 (N_572,N_284,In_1061);
xnor U573 (N_573,N_77,In_728);
nor U574 (N_574,In_493,N_103);
nand U575 (N_575,In_2187,In_892);
and U576 (N_576,In_1786,In_1890);
or U577 (N_577,In_1607,In_146);
nor U578 (N_578,In_616,In_92);
or U579 (N_579,In_525,In_2283);
and U580 (N_580,N_199,N_341);
xor U581 (N_581,In_482,In_1421);
nor U582 (N_582,In_1844,In_2075);
nor U583 (N_583,In_1194,In_1312);
nor U584 (N_584,In_806,In_2318);
nor U585 (N_585,In_172,In_270);
xor U586 (N_586,N_31,In_1857);
nand U587 (N_587,In_633,N_331);
nor U588 (N_588,In_464,In_2365);
nand U589 (N_589,In_1122,In_1508);
or U590 (N_590,In_75,In_1198);
xor U591 (N_591,In_2425,N_209);
nand U592 (N_592,In_726,N_262);
nor U593 (N_593,In_800,In_912);
xor U594 (N_594,In_909,In_821);
and U595 (N_595,In_2384,In_2191);
xor U596 (N_596,N_279,In_2055);
xor U597 (N_597,In_1111,In_1958);
or U598 (N_598,N_277,In_2023);
nor U599 (N_599,N_67,In_1871);
xor U600 (N_600,N_400,In_1308);
xnor U601 (N_601,In_1088,In_815);
nand U602 (N_602,N_177,In_2440);
nor U603 (N_603,In_2241,In_552);
or U604 (N_604,In_1316,In_1916);
nor U605 (N_605,In_216,N_325);
and U606 (N_606,In_332,N_70);
or U607 (N_607,N_297,N_235);
or U608 (N_608,N_278,In_1513);
or U609 (N_609,In_2419,N_399);
or U610 (N_610,In_1554,In_2043);
and U611 (N_611,In_2441,N_596);
nand U612 (N_612,In_1020,In_258);
or U613 (N_613,In_1597,In_1610);
xor U614 (N_614,In_2306,N_216);
and U615 (N_615,N_374,In_1097);
nand U616 (N_616,In_1413,N_476);
nand U617 (N_617,N_549,In_2045);
or U618 (N_618,In_1387,N_76);
nand U619 (N_619,In_428,In_1514);
xnor U620 (N_620,N_217,In_2341);
or U621 (N_621,In_2143,In_2211);
nand U622 (N_622,N_74,In_1941);
xnor U623 (N_623,In_85,In_1059);
nor U624 (N_624,In_1735,In_2207);
or U625 (N_625,In_994,N_354);
nor U626 (N_626,N_547,In_494);
and U627 (N_627,In_531,In_336);
nand U628 (N_628,N_91,In_1210);
xor U629 (N_629,N_249,In_2208);
or U630 (N_630,N_483,In_1262);
or U631 (N_631,N_273,In_1802);
nor U632 (N_632,N_6,In_784);
nor U633 (N_633,N_107,N_123);
and U634 (N_634,N_558,In_1330);
nand U635 (N_635,In_497,N_22);
nor U636 (N_636,N_241,In_656);
or U637 (N_637,In_966,In_952);
nand U638 (N_638,In_974,N_437);
nand U639 (N_639,N_546,In_1435);
or U640 (N_640,N_85,N_398);
and U641 (N_641,In_1712,N_454);
or U642 (N_642,In_166,N_254);
or U643 (N_643,N_417,In_1462);
nand U644 (N_644,In_1595,N_298);
xor U645 (N_645,In_571,In_1248);
or U646 (N_646,N_330,N_471);
nor U647 (N_647,In_1274,In_2401);
or U648 (N_648,In_1154,N_583);
nor U649 (N_649,In_792,N_94);
nand U650 (N_650,In_2476,In_1616);
xor U651 (N_651,In_1856,In_1516);
xnor U652 (N_652,In_2175,In_565);
and U653 (N_653,In_1021,In_483);
and U654 (N_654,In_444,In_2147);
nand U655 (N_655,In_983,In_436);
and U656 (N_656,In_961,In_1664);
xnor U657 (N_657,In_645,N_132);
nor U658 (N_658,N_2,N_86);
nor U659 (N_659,In_2254,In_1155);
xnor U660 (N_660,N_281,In_938);
nor U661 (N_661,N_242,In_451);
and U662 (N_662,In_1944,N_38);
nand U663 (N_663,In_48,In_1102);
and U664 (N_664,N_490,In_1263);
nand U665 (N_665,In_964,In_1480);
and U666 (N_666,In_1117,In_364);
xnor U667 (N_667,N_395,In_228);
nor U668 (N_668,N_551,In_1212);
and U669 (N_669,N_460,In_575);
xor U670 (N_670,In_789,N_486);
nand U671 (N_671,In_811,In_1129);
nand U672 (N_672,In_611,N_541);
nor U673 (N_673,In_2286,In_657);
and U674 (N_674,In_470,N_492);
or U675 (N_675,N_548,N_384);
nor U676 (N_676,In_2313,N_484);
or U677 (N_677,N_440,In_1626);
or U678 (N_678,In_2109,In_1876);
and U679 (N_679,In_1830,In_2338);
or U680 (N_680,N_335,In_1528);
and U681 (N_681,In_729,N_527);
or U682 (N_682,In_2408,In_705);
nand U683 (N_683,N_567,In_237);
xor U684 (N_684,In_2330,In_293);
and U685 (N_685,N_62,In_1564);
or U686 (N_686,In_2005,In_2416);
nor U687 (N_687,In_358,In_1338);
or U688 (N_688,In_1859,N_432);
nor U689 (N_689,In_1057,In_600);
nand U690 (N_690,N_168,In_813);
nand U691 (N_691,N_89,N_542);
xnor U692 (N_692,In_1288,In_1373);
and U693 (N_693,In_2074,In_520);
nor U694 (N_694,In_2081,In_1188);
and U695 (N_695,In_2080,In_1576);
or U696 (N_696,In_1006,N_334);
nor U697 (N_697,N_540,In_1159);
xor U698 (N_698,N_489,In_181);
nand U699 (N_699,In_1043,In_888);
xor U700 (N_700,In_1200,In_1700);
or U701 (N_701,In_1667,In_757);
nand U702 (N_702,In_1245,N_116);
or U703 (N_703,In_1842,In_441);
xnor U704 (N_704,In_131,In_1657);
nor U705 (N_705,In_1920,N_574);
nand U706 (N_706,In_1074,In_399);
and U707 (N_707,N_391,In_2065);
nand U708 (N_708,In_324,In_2323);
or U709 (N_709,In_242,In_29);
nand U710 (N_710,In_225,In_2479);
and U711 (N_711,In_1754,In_99);
xnor U712 (N_712,In_2417,N_196);
xnor U713 (N_713,N_207,In_1734);
nor U714 (N_714,N_267,N_16);
nand U715 (N_715,In_2423,In_7);
nor U716 (N_716,N_263,In_2439);
or U717 (N_717,In_1708,In_387);
nor U718 (N_718,In_2465,N_75);
or U719 (N_719,N_439,In_1891);
nand U720 (N_720,In_1936,N_53);
or U721 (N_721,In_2293,N_575);
nand U722 (N_722,In_1692,In_735);
and U723 (N_723,N_315,In_73);
xor U724 (N_724,In_1751,In_530);
or U725 (N_725,In_810,In_2396);
xor U726 (N_726,In_459,N_498);
and U727 (N_727,In_1358,N_478);
nor U728 (N_728,In_2072,In_1083);
and U729 (N_729,N_555,In_103);
nor U730 (N_730,In_388,In_950);
nand U731 (N_731,N_201,In_1710);
nor U732 (N_732,N_280,N_598);
nand U733 (N_733,In_1282,In_1887);
nor U734 (N_734,In_1345,In_941);
or U735 (N_735,N_48,N_172);
and U736 (N_736,In_1615,In_1975);
nand U737 (N_737,In_597,N_239);
xnor U738 (N_738,In_1645,In_1820);
xor U739 (N_739,N_213,In_713);
nor U740 (N_740,In_898,In_717);
xor U741 (N_741,In_1104,In_1150);
xor U742 (N_742,In_238,N_584);
or U743 (N_743,In_1885,N_255);
nor U744 (N_744,In_706,In_593);
and U745 (N_745,In_1166,In_763);
or U746 (N_746,N_438,N_528);
nand U747 (N_747,In_1688,N_220);
xor U748 (N_748,In_1224,In_1469);
nand U749 (N_749,N_83,N_212);
nor U750 (N_750,N_327,In_2392);
xor U751 (N_751,In_618,In_1971);
nor U752 (N_752,In_1047,In_1601);
or U753 (N_753,In_1017,In_712);
xnor U754 (N_754,In_2235,In_1470);
or U755 (N_755,In_1321,N_534);
or U756 (N_756,In_1864,In_1913);
xnor U757 (N_757,N_186,In_1854);
or U758 (N_758,In_595,N_1);
and U759 (N_759,In_1231,In_3);
and U760 (N_760,In_1027,In_1529);
or U761 (N_761,N_158,In_1962);
and U762 (N_762,In_2164,In_197);
nor U763 (N_763,In_309,In_2405);
nand U764 (N_764,In_557,N_218);
or U765 (N_765,In_844,In_505);
or U766 (N_766,N_379,In_348);
or U767 (N_767,N_451,N_543);
xor U768 (N_768,In_349,In_985);
and U769 (N_769,In_1605,In_1209);
xor U770 (N_770,In_686,In_678);
xor U771 (N_771,In_1266,In_1007);
or U772 (N_772,N_120,In_809);
or U773 (N_773,In_1974,In_895);
xor U774 (N_774,In_298,In_1574);
or U775 (N_775,In_598,In_2484);
xnor U776 (N_776,In_1774,N_501);
or U777 (N_777,In_1337,In_183);
xor U778 (N_778,In_1334,N_500);
nor U779 (N_779,In_1458,In_1823);
nand U780 (N_780,In_2457,In_14);
nand U781 (N_781,In_2326,In_1745);
xnor U782 (N_782,N_175,In_134);
nand U783 (N_783,In_299,N_588);
and U784 (N_784,In_1612,In_925);
xor U785 (N_785,In_1720,N_353);
and U786 (N_786,In_707,In_1197);
nor U787 (N_787,In_1536,In_2321);
or U788 (N_788,In_1319,In_693);
nor U789 (N_789,In_41,In_473);
and U790 (N_790,In_1235,In_877);
nor U791 (N_791,In_2435,N_571);
or U792 (N_792,In_1989,In_1940);
and U793 (N_793,In_316,N_593);
nor U794 (N_794,In_880,In_223);
nand U795 (N_795,In_609,In_585);
or U796 (N_796,In_151,N_301);
or U797 (N_797,In_582,In_190);
nand U798 (N_798,In_84,In_1654);
xor U799 (N_799,In_2400,In_2054);
nand U800 (N_800,In_1295,In_882);
and U801 (N_801,In_551,N_748);
or U802 (N_802,In_989,In_1499);
or U803 (N_803,In_490,In_2228);
or U804 (N_804,In_1258,N_788);
nor U805 (N_805,N_502,In_1199);
nor U806 (N_806,In_284,In_371);
and U807 (N_807,In_1425,N_314);
nand U808 (N_808,N_481,In_10);
nand U809 (N_809,N_453,In_401);
nand U810 (N_810,N_477,In_168);
and U811 (N_811,In_2162,In_443);
and U812 (N_812,N_651,In_2102);
nand U813 (N_813,In_1651,In_244);
nor U814 (N_814,In_1419,In_696);
nand U815 (N_815,In_18,In_1430);
nor U816 (N_816,In_2284,In_370);
nand U817 (N_817,In_2221,In_1882);
and U818 (N_818,In_1718,N_789);
or U819 (N_819,N_436,In_1877);
nand U820 (N_820,N_416,N_595);
nand U821 (N_821,In_310,In_72);
nor U822 (N_822,In_174,In_2044);
or U823 (N_823,N_529,In_1577);
nand U824 (N_824,In_2229,N_0);
nor U825 (N_825,N_45,In_1341);
nor U826 (N_826,In_867,In_330);
nand U827 (N_827,In_1771,N_721);
nor U828 (N_828,In_2141,In_753);
and U829 (N_829,In_834,In_40);
nor U830 (N_830,In_2358,N_348);
and U831 (N_831,N_317,In_1500);
and U832 (N_832,N_705,In_1226);
nand U833 (N_833,In_930,In_2470);
and U834 (N_834,In_1817,N_658);
nand U835 (N_835,N_776,N_568);
and U836 (N_836,In_2216,N_517);
nand U837 (N_837,In_2310,In_2022);
or U838 (N_838,In_2493,In_1642);
nor U839 (N_839,In_477,In_949);
or U840 (N_840,In_926,In_1685);
xnor U841 (N_841,In_2225,N_797);
nand U842 (N_842,In_2138,In_252);
nand U843 (N_843,In_1752,N_522);
nor U844 (N_844,In_1749,N_92);
xor U845 (N_845,N_412,In_328);
xnor U846 (N_846,In_1415,N_313);
or U847 (N_847,N_246,In_689);
or U848 (N_848,In_1438,In_825);
or U849 (N_849,In_931,In_1668);
nor U850 (N_850,In_2471,In_1284);
nand U851 (N_851,In_1866,In_2415);
nand U852 (N_852,In_171,In_1624);
xor U853 (N_853,In_704,In_1729);
nor U854 (N_854,In_637,N_250);
xor U855 (N_855,N_680,In_999);
nor U856 (N_856,N_796,In_1324);
or U857 (N_857,In_2063,N_232);
xnor U858 (N_858,N_223,N_691);
xnor U859 (N_859,In_725,In_2146);
nand U860 (N_860,In_1254,In_1375);
xor U861 (N_861,N_554,N_84);
and U862 (N_862,N_750,N_402);
nand U863 (N_863,In_203,N_702);
nor U864 (N_864,In_2354,In_972);
nand U865 (N_865,In_612,In_1801);
nand U866 (N_866,In_292,N_465);
nor U867 (N_867,N_689,In_2204);
nor U868 (N_868,N_43,N_761);
xor U869 (N_869,In_796,In_1805);
and U870 (N_870,In_1850,N_770);
nand U871 (N_871,N_50,In_1395);
nor U872 (N_872,N_553,In_1398);
nor U873 (N_873,N_134,In_2452);
and U874 (N_874,In_53,N_35);
or U875 (N_875,N_388,In_2150);
or U876 (N_876,In_2186,N_131);
and U877 (N_877,In_215,In_1792);
xor U878 (N_878,In_2325,In_133);
nand U879 (N_879,In_2236,In_2038);
xor U880 (N_880,N_530,In_948);
xor U881 (N_881,In_1464,N_444);
or U882 (N_882,In_841,In_2206);
and U883 (N_883,In_108,N_165);
and U884 (N_884,N_178,In_2073);
nand U885 (N_885,In_1661,In_1374);
xnor U886 (N_886,N_719,N_648);
xor U887 (N_887,N_4,N_739);
or U888 (N_888,In_32,In_413);
xor U889 (N_889,In_1821,In_1243);
or U890 (N_890,In_61,N_764);
nor U891 (N_891,N_552,In_424);
or U892 (N_892,N_283,In_1497);
and U893 (N_893,N_579,In_1652);
xnor U894 (N_894,N_652,N_520);
nor U895 (N_895,In_2349,N_227);
and U896 (N_896,N_638,In_1895);
nand U897 (N_897,In_1029,N_445);
nor U898 (N_898,N_711,In_1037);
or U899 (N_899,N_487,N_560);
nor U900 (N_900,N_147,In_1759);
nand U901 (N_901,N_318,N_350);
and U902 (N_902,In_955,In_2421);
nor U903 (N_903,In_1945,In_1663);
nor U904 (N_904,N_647,N_130);
nand U905 (N_905,In_1491,In_1697);
xnor U906 (N_906,N_755,In_2412);
or U907 (N_907,In_164,In_543);
and U908 (N_908,N_468,N_641);
nor U909 (N_909,In_2352,N_230);
xnor U910 (N_910,In_2010,N_302);
or U911 (N_911,In_563,In_208);
nand U912 (N_912,In_1148,In_553);
and U913 (N_913,In_2066,In_1393);
xnor U914 (N_914,N_642,In_814);
or U915 (N_915,N_99,N_170);
xnor U916 (N_916,N_545,N_669);
and U917 (N_917,N_310,N_611);
and U918 (N_918,In_439,In_1353);
and U919 (N_919,N_740,In_1681);
nor U920 (N_920,In_859,In_1442);
nand U921 (N_921,In_1272,In_1130);
xor U922 (N_922,In_1596,In_515);
nand U923 (N_923,In_460,In_1315);
and U924 (N_924,N_779,In_1036);
or U925 (N_925,In_194,In_1849);
or U926 (N_926,In_1177,N_271);
nor U927 (N_927,In_1105,In_1787);
nor U928 (N_928,In_1848,In_905);
nor U929 (N_929,In_1403,In_1473);
xnor U930 (N_930,In_1325,In_1666);
nand U931 (N_931,In_827,N_506);
nor U932 (N_932,In_2424,N_572);
and U933 (N_933,In_1429,In_2360);
and U934 (N_934,In_1717,In_1937);
or U935 (N_935,In_389,In_548);
nor U936 (N_936,In_1704,In_775);
nor U937 (N_937,N_735,N_224);
or U938 (N_938,N_590,N_707);
nand U939 (N_939,In_1391,In_2256);
nor U940 (N_940,In_871,In_38);
xnor U941 (N_941,N_621,In_1999);
nor U942 (N_942,In_2224,In_2197);
and U943 (N_943,N_509,In_296);
nor U944 (N_944,In_1326,N_765);
nor U945 (N_945,In_2031,In_2359);
xor U946 (N_946,In_1948,N_139);
nand U947 (N_947,N_634,N_717);
nand U948 (N_948,In_266,N_154);
or U949 (N_949,N_179,In_1378);
nand U950 (N_950,In_1182,In_1767);
nand U951 (N_951,N_592,N_767);
xor U952 (N_952,In_1363,In_2230);
or U953 (N_953,In_532,N_674);
or U954 (N_954,N_698,N_290);
and U955 (N_955,In_1512,N_210);
or U956 (N_956,In_954,In_265);
or U957 (N_957,In_489,In_1722);
nor U958 (N_958,In_503,N_383);
nand U959 (N_959,N_166,In_1287);
xnor U960 (N_960,In_476,In_743);
xnor U961 (N_961,In_2363,In_123);
xor U962 (N_962,In_2386,In_1187);
xor U963 (N_963,N_668,In_2135);
or U964 (N_964,In_1540,In_2046);
or U965 (N_965,In_1935,N_288);
and U966 (N_966,In_1060,In_2346);
xor U967 (N_967,In_2160,N_375);
xnor U968 (N_968,In_1482,N_410);
nand U969 (N_969,In_124,In_2193);
nand U970 (N_970,N_408,In_56);
nor U971 (N_971,In_1264,In_2418);
or U972 (N_972,In_1592,In_2356);
nor U973 (N_973,In_297,N_57);
nor U974 (N_974,N_724,In_1485);
nor U975 (N_975,In_1521,In_339);
or U976 (N_976,N_363,In_672);
nor U977 (N_977,In_1538,In_239);
or U978 (N_978,N_617,In_202);
nand U979 (N_979,N_311,In_2140);
nor U980 (N_980,N_741,In_402);
nand U981 (N_981,N_704,In_1377);
and U982 (N_982,In_1740,In_2276);
xor U983 (N_983,In_2292,In_644);
nand U984 (N_984,In_977,In_407);
nor U985 (N_985,In_1702,N_640);
or U986 (N_986,N_219,In_1892);
nand U987 (N_987,In_1303,In_2264);
nand U988 (N_988,N_633,In_2029);
nand U989 (N_989,In_2118,N_118);
nor U990 (N_990,In_150,In_790);
and U991 (N_991,N_609,N_673);
or U992 (N_992,In_1846,In_288);
nand U993 (N_993,N_386,In_1448);
xor U994 (N_994,N_358,In_1906);
and U995 (N_995,In_15,N_497);
and U996 (N_996,In_2210,N_36);
nand U997 (N_997,In_1392,N_329);
nor U998 (N_998,In_508,N_762);
xnor U999 (N_999,N_474,In_822);
nand U1000 (N_1000,In_2387,In_1881);
nor U1001 (N_1001,In_1560,In_1875);
nor U1002 (N_1002,In_207,In_824);
and U1003 (N_1003,In_2483,N_892);
nor U1004 (N_1004,In_400,N_389);
and U1005 (N_1005,In_802,In_1580);
and U1006 (N_1006,In_511,In_1340);
or U1007 (N_1007,N_108,N_926);
or U1008 (N_1008,In_438,In_1747);
xnor U1009 (N_1009,N_845,In_2171);
or U1010 (N_1010,In_1954,In_415);
xor U1011 (N_1011,N_756,In_906);
and U1012 (N_1012,N_996,In_1269);
xnor U1013 (N_1013,In_1589,In_2322);
nor U1014 (N_1014,N_992,In_2025);
or U1015 (N_1015,N_752,N_205);
nor U1016 (N_1016,N_100,In_1867);
nor U1017 (N_1017,N_630,N_690);
nand U1018 (N_1018,In_1525,In_697);
xnor U1019 (N_1019,In_1443,In_1834);
and U1020 (N_1020,N_275,In_1765);
and U1021 (N_1021,N_932,In_327);
xor U1022 (N_1022,N_714,In_1300);
xnor U1023 (N_1023,In_2003,In_1192);
xor U1024 (N_1024,In_2269,N_404);
and U1025 (N_1025,In_1125,In_394);
or U1026 (N_1026,N_185,N_708);
xnor U1027 (N_1027,N_692,In_2103);
nor U1028 (N_1028,N_226,In_1418);
xor U1029 (N_1029,N_780,N_204);
nor U1030 (N_1030,In_2007,In_2443);
or U1031 (N_1031,N_33,In_1024);
nor U1032 (N_1032,In_622,In_2474);
or U1033 (N_1033,In_682,In_1878);
nand U1034 (N_1034,In_1919,In_749);
or U1035 (N_1035,In_1115,N_886);
nand U1036 (N_1036,N_988,In_2036);
and U1037 (N_1037,In_2281,In_1925);
and U1038 (N_1038,N_744,In_1614);
or U1039 (N_1039,N_54,In_2495);
or U1040 (N_1040,N_215,N_345);
or U1041 (N_1041,N_121,N_734);
and U1042 (N_1042,In_2179,In_1656);
and U1043 (N_1043,In_1246,In_736);
xnor U1044 (N_1044,In_589,N_745);
nor U1045 (N_1045,In_2176,In_2024);
xnor U1046 (N_1046,In_433,In_1772);
xor U1047 (N_1047,In_2496,In_1889);
xnor U1048 (N_1048,In_1492,N_975);
xnor U1049 (N_1049,In_1018,In_209);
xnor U1050 (N_1050,N_955,In_1001);
and U1051 (N_1051,In_175,In_442);
and U1052 (N_1052,In_1466,In_2450);
xnor U1053 (N_1053,In_1694,N_809);
xor U1054 (N_1054,In_2431,In_71);
nor U1055 (N_1055,N_774,In_2296);
nand U1056 (N_1056,N_850,In_2478);
nand U1057 (N_1057,N_581,In_572);
nand U1058 (N_1058,N_282,In_1755);
nand U1059 (N_1059,In_2311,N_418);
xnor U1060 (N_1060,In_1,In_2420);
or U1061 (N_1061,In_788,N_591);
or U1062 (N_1062,N_922,N_434);
and U1063 (N_1063,N_644,In_2458);
nand U1064 (N_1064,In_2456,In_162);
or U1065 (N_1065,In_1987,In_914);
or U1066 (N_1066,N_995,N_51);
nor U1067 (N_1067,In_574,N_873);
nor U1068 (N_1068,In_1604,N_657);
and U1069 (N_1069,In_2249,In_63);
nor U1070 (N_1070,N_268,In_1463);
xor U1071 (N_1071,N_531,In_539);
and U1072 (N_1072,In_1904,In_1216);
nand U1073 (N_1073,In_89,In_410);
nand U1074 (N_1074,In_1543,N_614);
nand U1075 (N_1075,In_768,In_1862);
xnor U1076 (N_1076,N_916,In_652);
and U1077 (N_1077,N_790,N_608);
xnor U1078 (N_1078,In_969,In_51);
or U1079 (N_1079,N_167,In_396);
nor U1080 (N_1080,In_210,N_401);
nand U1081 (N_1081,In_0,In_667);
xnor U1082 (N_1082,In_587,In_249);
nor U1083 (N_1083,In_1571,N_963);
and U1084 (N_1084,N_931,N_562);
xor U1085 (N_1085,N_929,N_927);
xnor U1086 (N_1086,In_102,N_585);
and U1087 (N_1087,N_923,N_646);
and U1088 (N_1088,In_2100,N_666);
and U1089 (N_1089,N_360,N_95);
xnor U1090 (N_1090,In_915,In_1313);
and U1091 (N_1091,N_954,In_1578);
nor U1092 (N_1092,In_2242,In_2324);
xor U1093 (N_1093,In_1428,In_158);
and U1094 (N_1094,In_646,N_650);
and U1095 (N_1095,In_2157,N_786);
or U1096 (N_1096,N_989,In_2402);
xor U1097 (N_1097,In_1203,N_518);
xor U1098 (N_1098,In_329,N_978);
or U1099 (N_1099,In_928,In_458);
nand U1100 (N_1100,In_911,In_1939);
nor U1101 (N_1101,In_36,In_1915);
xnor U1102 (N_1102,N_28,N_183);
nand U1103 (N_1103,In_1665,In_831);
nand U1104 (N_1104,N_686,In_1768);
nand U1105 (N_1105,In_1621,N_912);
nand U1106 (N_1106,In_1157,N_512);
or U1107 (N_1107,N_966,In_98);
nor U1108 (N_1108,In_2307,In_1494);
xor U1109 (N_1109,In_488,N_820);
and U1110 (N_1110,N_754,N_663);
nand U1111 (N_1111,In_104,N_836);
nor U1112 (N_1112,In_278,In_2340);
nor U1113 (N_1113,In_2195,N_485);
xnor U1114 (N_1114,In_191,In_830);
or U1115 (N_1115,N_956,N_775);
nand U1116 (N_1116,N_415,N_157);
or U1117 (N_1117,In_1070,N_900);
nor U1118 (N_1118,N_269,In_186);
or U1119 (N_1119,N_378,N_948);
nor U1120 (N_1120,N_447,N_917);
nor U1121 (N_1121,N_971,N_253);
xnor U1122 (N_1122,N_897,In_1927);
nand U1123 (N_1123,In_2088,In_1143);
nor U1124 (N_1124,In_1230,In_1091);
nand U1125 (N_1125,N_326,In_1121);
nand U1126 (N_1126,In_462,In_773);
or U1127 (N_1127,In_1522,In_1072);
nor U1128 (N_1128,In_879,In_1960);
and U1129 (N_1129,In_1022,In_1128);
nor U1130 (N_1130,N_287,N_426);
nor U1131 (N_1131,In_54,In_934);
nand U1132 (N_1132,In_1855,In_1539);
and U1133 (N_1133,In_617,In_290);
nor U1134 (N_1134,N_868,In_1381);
and U1135 (N_1135,N_882,N_815);
nand U1136 (N_1136,In_1695,N_816);
and U1137 (N_1137,In_1252,N_312);
or U1138 (N_1138,In_468,In_2098);
nand U1139 (N_1139,N_307,In_1171);
and U1140 (N_1140,In_785,N_643);
or U1141 (N_1141,In_751,In_812);
nand U1142 (N_1142,N_576,N_612);
and U1143 (N_1143,In_100,In_793);
nand U1144 (N_1144,In_1588,N_499);
nand U1145 (N_1145,In_2180,In_883);
nor U1146 (N_1146,In_453,In_1489);
nor U1147 (N_1147,In_1112,In_138);
nand U1148 (N_1148,In_2047,In_77);
nand U1149 (N_1149,In_613,In_368);
xor U1150 (N_1150,In_379,In_1481);
nand U1151 (N_1151,N_627,N_928);
and U1152 (N_1152,N_305,In_2226);
nand U1153 (N_1153,In_1310,N_894);
nor U1154 (N_1154,N_939,N_938);
nand U1155 (N_1155,N_872,In_5);
xor U1156 (N_1156,In_1013,N_96);
xor U1157 (N_1157,N_746,In_1980);
nor U1158 (N_1158,N_962,In_286);
xnor U1159 (N_1159,In_1622,In_2018);
xor U1160 (N_1160,N_709,In_817);
xnor U1161 (N_1161,In_741,In_987);
xor U1162 (N_1162,N_781,In_1608);
and U1163 (N_1163,N_716,In_224);
xor U1164 (N_1164,N_366,In_231);
and U1165 (N_1165,N_722,N_812);
xor U1166 (N_1166,In_2013,N_356);
and U1167 (N_1167,In_1533,N_732);
nor U1168 (N_1168,N_523,In_2361);
nor U1169 (N_1169,In_1853,N_725);
or U1170 (N_1170,N_64,In_2132);
and U1171 (N_1171,In_240,In_1756);
nor U1172 (N_1172,In_1840,N_773);
or U1173 (N_1173,N_925,N_449);
and U1174 (N_1174,In_1964,N_747);
and U1175 (N_1175,N_427,In_128);
xor U1176 (N_1176,N_972,N_623);
or U1177 (N_1177,In_1426,In_873);
and U1178 (N_1178,In_754,N_135);
nand U1179 (N_1179,In_869,N_667);
or U1180 (N_1180,N_693,N_860);
nor U1181 (N_1181,In_33,In_739);
nor U1182 (N_1182,In_2159,N_480);
or U1183 (N_1183,N_306,N_924);
xor U1184 (N_1184,N_846,In_1907);
nand U1185 (N_1185,In_996,N_783);
and U1186 (N_1186,N_44,In_1424);
nor U1187 (N_1187,In_636,N_700);
xnor U1188 (N_1188,In_1452,N_604);
nor U1189 (N_1189,In_1992,In_1030);
or U1190 (N_1190,N_164,In_1364);
nor U1191 (N_1191,In_1556,In_1336);
nor U1192 (N_1192,In_744,In_2020);
nand U1193 (N_1193,In_683,In_1997);
or U1194 (N_1194,In_1379,N_981);
nor U1195 (N_1195,N_794,N_842);
nor U1196 (N_1196,N_908,N_959);
nand U1197 (N_1197,N_605,N_821);
or U1198 (N_1198,In_2125,In_1371);
nor U1199 (N_1199,In_740,N_169);
nor U1200 (N_1200,N_913,N_1034);
xnor U1201 (N_1201,N_544,N_519);
and U1202 (N_1202,In_1161,In_1347);
nand U1203 (N_1203,In_188,N_793);
xnor U1204 (N_1204,In_1367,In_1931);
xnor U1205 (N_1205,In_471,N_1042);
and U1206 (N_1206,N_569,N_1028);
xnor U1207 (N_1207,N_73,N_1133);
or U1208 (N_1208,In_1401,N_1087);
xnor U1209 (N_1209,In_1838,N_905);
nand U1210 (N_1210,N_653,N_977);
nor U1211 (N_1211,N_421,N_856);
nor U1212 (N_1212,N_1090,N_624);
and U1213 (N_1213,N_52,N_718);
nor U1214 (N_1214,In_45,In_1417);
nor U1215 (N_1215,N_274,In_2115);
and U1216 (N_1216,In_1414,N_881);
and U1217 (N_1217,In_2030,In_2037);
or U1218 (N_1218,In_1894,In_450);
or U1219 (N_1219,In_1836,In_2467);
nand U1220 (N_1220,N_655,N_1129);
and U1221 (N_1221,In_234,In_2257);
nand U1222 (N_1222,In_1382,In_1760);
xor U1223 (N_1223,In_1861,In_1783);
or U1224 (N_1224,In_1023,In_199);
xnor U1225 (N_1225,In_2061,In_614);
nand U1226 (N_1226,In_621,In_1141);
nand U1227 (N_1227,N_738,N_1019);
xor U1228 (N_1228,In_78,N_296);
nor U1229 (N_1229,In_1384,In_1674);
and U1230 (N_1230,In_2096,In_1041);
or U1231 (N_1231,N_332,In_2021);
or U1232 (N_1232,N_1075,N_430);
or U1233 (N_1233,N_696,N_1060);
and U1234 (N_1234,In_1151,In_509);
nor U1235 (N_1235,N_163,In_1537);
nand U1236 (N_1236,In_1476,In_1156);
nand U1237 (N_1237,N_837,N_730);
or U1238 (N_1238,In_723,In_1106);
and U1239 (N_1239,In_2042,N_1004);
nand U1240 (N_1240,In_449,N_1144);
or U1241 (N_1241,N_898,N_1114);
and U1242 (N_1242,In_527,N_441);
nor U1243 (N_1243,N_830,N_125);
xor U1244 (N_1244,N_715,In_2461);
xor U1245 (N_1245,In_2233,N_884);
nor U1246 (N_1246,N_503,N_1103);
nand U1247 (N_1247,N_1180,In_836);
nand U1248 (N_1248,N_276,In_913);
nand U1249 (N_1249,N_1195,N_636);
nand U1250 (N_1250,N_137,N_936);
nor U1251 (N_1251,N_893,In_1176);
and U1252 (N_1252,N_1011,N_839);
and U1253 (N_1253,N_456,In_83);
and U1254 (N_1254,N_411,N_1068);
and U1255 (N_1255,In_2350,In_380);
or U1256 (N_1256,In_1318,N_728);
xnor U1257 (N_1257,In_1256,N_619);
or U1258 (N_1258,In_2009,In_1721);
and U1259 (N_1259,N_757,N_1179);
xnor U1260 (N_1260,In_1813,N_1062);
nand U1261 (N_1261,In_685,N_629);
nor U1262 (N_1262,N_688,N_866);
nand U1263 (N_1263,In_1175,N_225);
nand U1264 (N_1264,N_1052,In_629);
xnor U1265 (N_1265,N_1001,In_2237);
or U1266 (N_1266,N_1056,In_479);
and U1267 (N_1267,In_2319,N_324);
nand U1268 (N_1268,In_2232,N_671);
or U1269 (N_1269,In_1223,In_155);
and U1270 (N_1270,N_742,In_2104);
or U1271 (N_1271,N_818,N_1085);
nand U1272 (N_1272,In_2122,In_774);
or U1273 (N_1273,In_579,N_994);
and U1274 (N_1274,In_1804,In_1003);
nand U1275 (N_1275,In_243,In_653);
nor U1276 (N_1276,In_1240,N_3);
xor U1277 (N_1277,In_866,In_960);
nor U1278 (N_1278,N_833,In_604);
or U1279 (N_1279,N_862,N_902);
nand U1280 (N_1280,N_865,In_2083);
or U1281 (N_1281,N_906,In_1782);
or U1282 (N_1282,In_1376,N_749);
nor U1283 (N_1283,In_1619,N_656);
nor U1284 (N_1284,In_849,In_354);
and U1285 (N_1285,In_57,In_2129);
nand U1286 (N_1286,In_2315,N_351);
and U1287 (N_1287,N_349,N_161);
nand U1288 (N_1288,N_606,In_363);
nor U1289 (N_1289,N_1099,N_1119);
and U1290 (N_1290,N_406,N_890);
nor U1291 (N_1291,N_763,N_814);
nor U1292 (N_1292,In_12,In_526);
nor U1293 (N_1293,N_413,In_21);
or U1294 (N_1294,N_510,In_1505);
or U1295 (N_1295,In_376,N_152);
and U1296 (N_1296,In_345,N_808);
nand U1297 (N_1297,In_1739,In_694);
nand U1298 (N_1298,N_431,N_414);
nor U1299 (N_1299,N_1140,In_1572);
and U1300 (N_1300,In_214,In_11);
nand U1301 (N_1301,N_587,In_455);
and U1302 (N_1302,In_1446,N_799);
nand U1303 (N_1303,N_878,In_654);
nand U1304 (N_1304,N_448,N_990);
nor U1305 (N_1305,In_27,In_1829);
nor U1306 (N_1306,In_1690,N_190);
nand U1307 (N_1307,N_1115,In_1207);
or U1308 (N_1308,In_23,In_662);
nand U1309 (N_1309,In_1719,N_804);
nand U1310 (N_1310,N_934,In_1546);
xnor U1311 (N_1311,In_411,N_1162);
nor U1312 (N_1312,In_1811,N_1137);
nor U1313 (N_1313,In_2383,In_1847);
nor U1314 (N_1314,N_802,N_577);
xnor U1315 (N_1315,In_1260,In_920);
nor U1316 (N_1316,In_847,N_852);
and U1317 (N_1317,N_425,In_516);
or U1318 (N_1318,In_641,In_110);
nand U1319 (N_1319,In_648,N_877);
and U1320 (N_1320,In_1253,In_2380);
xor U1321 (N_1321,In_446,In_1179);
or U1322 (N_1322,In_2320,N_909);
and U1323 (N_1323,N_144,N_1136);
nand U1324 (N_1324,N_1024,N_1177);
or U1325 (N_1325,N_1008,In_2086);
nor U1326 (N_1326,N_387,N_494);
nor U1327 (N_1327,In_956,N_236);
xnor U1328 (N_1328,N_475,N_819);
or U1329 (N_1329,In_2393,N_1108);
and U1330 (N_1330,N_683,N_823);
xor U1331 (N_1331,N_782,In_59);
nand U1332 (N_1332,N_206,In_2462);
and U1333 (N_1333,In_1998,In_70);
nor U1334 (N_1334,N_397,N_983);
or U1335 (N_1335,In_2084,N_1181);
nor U1336 (N_1336,N_600,In_850);
or U1337 (N_1337,In_42,N_1097);
nor U1338 (N_1338,In_335,In_1113);
or U1339 (N_1339,In_1039,N_760);
or U1340 (N_1340,In_414,In_537);
or U1341 (N_1341,In_1630,In_603);
nor U1342 (N_1342,In_318,In_965);
or U1343 (N_1343,In_2489,N_563);
nand U1344 (N_1344,In_1544,In_2085);
nor U1345 (N_1345,In_2278,In_2344);
xor U1346 (N_1346,In_2436,N_1196);
nor U1347 (N_1347,N_240,In_615);
xnor U1348 (N_1348,In_1026,N_153);
and U1349 (N_1349,N_703,N_1039);
xnor U1350 (N_1350,N_443,N_423);
nand U1351 (N_1351,N_1061,N_1054);
nand U1352 (N_1352,N_880,N_461);
nor U1353 (N_1353,In_1841,N_631);
nand U1354 (N_1354,N_496,In_1924);
or U1355 (N_1355,In_1474,N_903);
xor U1356 (N_1356,In_624,N_1116);
nor U1357 (N_1357,N_1030,In_342);
and U1358 (N_1358,In_748,In_734);
and U1359 (N_1359,N_943,N_967);
nor U1360 (N_1360,In_1009,N_1049);
and U1361 (N_1361,In_1255,In_2413);
xnor U1362 (N_1362,In_142,N_597);
nand U1363 (N_1363,In_944,N_1175);
nand U1364 (N_1364,N_333,N_594);
and U1365 (N_1365,N_863,In_982);
and U1366 (N_1366,N_234,N_701);
xor U1367 (N_1367,In_2265,N_920);
xnor U1368 (N_1368,N_889,N_1026);
nor U1369 (N_1369,N_811,In_392);
nor U1370 (N_1370,In_1096,In_94);
and U1371 (N_1371,N_1104,In_2300);
nand U1372 (N_1372,In_993,N_446);
or U1373 (N_1373,In_165,N_1045);
nor U1374 (N_1374,N_29,N_30);
and U1375 (N_1375,N_15,N_403);
and U1376 (N_1376,N_472,In_383);
nand U1377 (N_1377,N_295,In_319);
xor U1378 (N_1378,N_947,N_467);
and U1379 (N_1379,N_1048,In_2273);
nor U1380 (N_1380,In_701,N_1134);
xnor U1381 (N_1381,N_1092,In_673);
xor U1382 (N_1382,N_1084,N_376);
xor U1383 (N_1383,N_377,N_557);
nor U1384 (N_1384,N_733,N_1122);
xor U1385 (N_1385,N_1120,N_813);
and U1386 (N_1386,N_953,N_1183);
and U1387 (N_1387,In_590,In_1372);
and U1388 (N_1388,In_1535,In_1163);
xor U1389 (N_1389,N_13,In_1397);
xnor U1390 (N_1390,N_899,In_2015);
and U1391 (N_1391,N_109,In_301);
or U1392 (N_1392,In_2366,In_426);
nor U1393 (N_1393,In_1063,In_1527);
xnor U1394 (N_1394,N_1066,In_126);
xor U1395 (N_1395,In_1509,In_632);
or U1396 (N_1396,In_1160,In_875);
and U1397 (N_1397,In_2026,N_1172);
and U1398 (N_1398,In_422,In_2355);
nand U1399 (N_1399,N_1138,N_615);
and U1400 (N_1400,N_613,N_831);
xor U1401 (N_1401,N_429,In_1706);
nand U1402 (N_1402,In_899,N_1245);
nor U1403 (N_1403,N_56,In_1055);
xnor U1404 (N_1404,N_1069,In_1932);
xnor U1405 (N_1405,In_1359,In_737);
xnor U1406 (N_1406,N_875,N_1394);
nand U1407 (N_1407,In_152,N_570);
xor U1408 (N_1408,N_1031,N_987);
and U1409 (N_1409,N_320,In_2498);
and U1410 (N_1410,N_68,N_1249);
nor U1411 (N_1411,N_539,N_731);
nand U1412 (N_1412,In_1118,N_1235);
and U1413 (N_1413,N_1218,In_510);
nand U1414 (N_1414,N_1296,In_1299);
xor U1415 (N_1415,N_1078,In_1471);
nand U1416 (N_1416,In_1440,N_784);
xor U1417 (N_1417,N_365,N_968);
nor U1418 (N_1418,N_524,In_932);
xnor U1419 (N_1419,N_855,N_1258);
nand U1420 (N_1420,N_1343,N_664);
nand U1421 (N_1421,In_1320,N_685);
or U1422 (N_1422,N_589,In_1361);
or U1423 (N_1423,In_1296,In_564);
and U1424 (N_1424,In_1638,N_825);
or U1425 (N_1425,In_1880,N_1186);
nor U1426 (N_1426,N_1255,In_1457);
nand U1427 (N_1427,In_1165,N_1370);
xor U1428 (N_1428,N_993,N_1324);
xnor U1429 (N_1429,N_251,N_1389);
or U1430 (N_1430,N_1164,N_1037);
nor U1431 (N_1431,N_1157,In_1126);
nor U1432 (N_1432,N_1237,In_2253);
and U1433 (N_1433,N_507,N_133);
and U1434 (N_1434,N_1349,N_1150);
nor U1435 (N_1435,In_2223,N_1307);
or U1436 (N_1436,N_381,In_378);
or U1437 (N_1437,In_1625,N_1333);
nand U1438 (N_1438,In_65,N_424);
and U1439 (N_1439,In_759,N_649);
or U1440 (N_1440,In_1839,In_1791);
xnor U1441 (N_1441,N_941,N_1274);
and U1442 (N_1442,In_1056,In_1600);
nor U1443 (N_1443,N_136,In_607);
xnor U1444 (N_1444,In_1132,In_1225);
and U1445 (N_1445,In_670,N_1364);
nor U1446 (N_1446,In_1218,N_1041);
xor U1447 (N_1447,N_515,N_1348);
xnor U1448 (N_1448,In_1493,N_1141);
xor U1449 (N_1449,In_492,In_111);
and U1450 (N_1450,N_1050,N_442);
xor U1451 (N_1451,N_1340,In_506);
nor U1452 (N_1452,N_1003,In_1289);
xor U1453 (N_1453,In_118,N_1309);
nand U1454 (N_1454,N_1142,In_1517);
nor U1455 (N_1455,N_1101,In_1671);
nor U1456 (N_1456,N_455,N_338);
nor U1457 (N_1457,N_713,In_1116);
and U1458 (N_1458,N_661,In_2258);
nor U1459 (N_1459,N_1146,In_1444);
and U1460 (N_1460,In_1816,N_1329);
nand U1461 (N_1461,In_2184,N_407);
xnor U1462 (N_1462,N_409,N_1250);
and U1463 (N_1463,In_2108,In_1670);
and U1464 (N_1464,In_1914,N_47);
or U1465 (N_1465,In_2382,N_1178);
or U1466 (N_1466,N_1378,In_2328);
nor U1467 (N_1467,N_176,N_124);
nand U1468 (N_1468,In_504,N_1027);
or U1469 (N_1469,N_1165,N_957);
and U1470 (N_1470,In_2238,In_1232);
xor U1471 (N_1471,In_20,In_2078);
nand U1472 (N_1472,N_965,N_1055);
nor U1473 (N_1473,In_106,In_2008);
xnor U1474 (N_1474,N_660,N_602);
or U1475 (N_1475,In_1583,In_314);
nand U1476 (N_1476,In_1769,In_1627);
and U1477 (N_1477,In_959,N_874);
xor U1478 (N_1478,In_325,In_2217);
xnor U1479 (N_1479,In_1825,N_795);
and U1480 (N_1480,N_1190,N_1367);
nand U1481 (N_1481,N_1282,N_645);
or U1482 (N_1482,In_922,In_833);
nor U1483 (N_1483,N_1273,N_777);
xor U1484 (N_1484,N_1184,N_918);
nor U1485 (N_1485,N_829,In_1519);
or U1486 (N_1486,N_1362,N_822);
nand U1487 (N_1487,In_340,In_369);
nand U1488 (N_1488,N_1058,N_1156);
or U1489 (N_1489,N_1166,N_1013);
and U1490 (N_1490,N_1269,In_1025);
nand U1491 (N_1491,N_864,N_564);
nor U1492 (N_1492,N_1093,N_675);
xor U1493 (N_1493,N_1356,N_1336);
nand U1494 (N_1494,N_1070,In_1983);
nand U1495 (N_1495,N_1149,N_1118);
and U1496 (N_1496,In_699,N_488);
nand U1497 (N_1497,In_2131,N_466);
xor U1498 (N_1498,N_999,In_1138);
nor U1499 (N_1499,In_647,In_1249);
xor U1500 (N_1500,N_1395,In_929);
or U1501 (N_1501,N_1154,N_1295);
nand U1502 (N_1502,N_580,N_433);
or U1503 (N_1503,N_768,In_1757);
nand U1504 (N_1504,N_901,In_601);
or U1505 (N_1505,N_119,N_550);
or U1506 (N_1506,N_867,N_626);
xor U1507 (N_1507,In_2194,In_1349);
nand U1508 (N_1508,N_1167,N_1310);
or U1509 (N_1509,N_697,N_970);
and U1510 (N_1510,N_759,N_308);
nand U1511 (N_1511,N_1241,In_860);
and U1512 (N_1512,N_844,In_1045);
xnor U1513 (N_1513,N_620,N_1182);
xor U1514 (N_1514,N_858,In_1938);
and U1515 (N_1515,N_1322,N_792);
nand U1516 (N_1516,N_817,N_1006);
and U1517 (N_1517,In_1758,In_2060);
or U1518 (N_1518,In_1524,N_1229);
or U1519 (N_1519,In_1808,In_1008);
and U1520 (N_1520,N_1155,N_1063);
xnor U1521 (N_1521,N_1159,In_894);
nand U1522 (N_1522,N_72,N_933);
xor U1523 (N_1523,N_727,N_514);
xnor U1524 (N_1524,N_1073,In_544);
and U1525 (N_1525,N_1239,N_264);
nor U1526 (N_1526,N_1216,In_975);
nand U1527 (N_1527,In_2407,In_385);
nor U1528 (N_1528,N_1171,N_1192);
nor U1529 (N_1529,In_2112,N_1360);
nor U1530 (N_1530,In_173,N_202);
nor U1531 (N_1531,N_603,N_869);
nand U1532 (N_1532,N_1091,In_786);
nand U1533 (N_1533,In_101,In_1205);
xor U1534 (N_1534,N_1242,In_480);
nand U1535 (N_1535,N_1256,In_205);
nand U1536 (N_1536,In_970,N_607);
and U1537 (N_1537,N_930,In_769);
nor U1538 (N_1538,N_1176,In_1949);
xnor U1539 (N_1539,N_1106,N_1366);
nand U1540 (N_1540,N_459,N_997);
nand U1541 (N_1541,N_1015,N_188);
or U1542 (N_1542,In_874,N_19);
xnor U1543 (N_1543,N_1147,In_269);
nor U1544 (N_1544,In_1357,N_743);
and U1545 (N_1545,In_2077,N_1079);
xnor U1546 (N_1546,In_1239,N_961);
nor U1547 (N_1547,In_1170,N_1224);
or U1548 (N_1548,N_848,In_1280);
or U1549 (N_1549,In_312,In_578);
nand U1550 (N_1550,N_800,In_2411);
xnor U1551 (N_1551,In_1926,N_228);
nand U1552 (N_1552,In_1883,In_160);
nand U1553 (N_1553,In_1164,In_2277);
nor U1554 (N_1554,N_8,N_1368);
nor U1555 (N_1555,N_1189,In_904);
or U1556 (N_1556,In_2335,N_1346);
nand U1557 (N_1557,N_810,In_868);
nand U1558 (N_1558,N_1072,N_21);
or U1559 (N_1559,N_1327,N_1376);
xnor U1560 (N_1560,In_1147,N_1374);
xnor U1561 (N_1561,N_1117,N_368);
xnor U1562 (N_1562,N_986,N_504);
and U1563 (N_1563,In_1701,N_679);
and U1564 (N_1564,In_908,N_952);
nand U1565 (N_1565,N_1314,N_1332);
and U1566 (N_1566,N_1217,In_2255);
nor U1567 (N_1567,N_695,In_1728);
and U1568 (N_1568,N_1025,In_382);
or U1569 (N_1569,N_1319,N_1230);
nor U1570 (N_1570,In_1073,In_547);
xor U1571 (N_1571,N_1279,N_1014);
xnor U1572 (N_1572,In_856,N_945);
nand U1573 (N_1573,N_1173,N_1247);
xnor U1574 (N_1574,In_1110,N_1263);
xor U1575 (N_1575,N_1040,N_112);
and U1576 (N_1576,In_1724,In_360);
nand U1577 (N_1577,N_420,N_1163);
or U1578 (N_1578,In_1835,N_1188);
or U1579 (N_1579,N_601,N_1391);
or U1580 (N_1580,N_944,N_1193);
nor U1581 (N_1581,In_2348,In_596);
nor U1582 (N_1582,N_344,In_872);
nand U1583 (N_1583,In_512,N_915);
nand U1584 (N_1584,In_333,In_556);
nand U1585 (N_1585,In_1800,In_347);
nor U1586 (N_1586,N_1002,In_211);
nor U1587 (N_1587,N_1278,N_1194);
and U1588 (N_1588,In_2290,N_1215);
or U1589 (N_1589,N_578,In_1795);
or U1590 (N_1590,N_1209,N_616);
and U1591 (N_1591,N_1276,In_46);
and U1592 (N_1592,In_1570,In_2480);
or U1593 (N_1593,In_1468,N_801);
and U1594 (N_1594,N_1299,In_1109);
or U1595 (N_1595,N_632,N_960);
nor U1596 (N_1596,N_1021,N_238);
and U1597 (N_1597,In_854,N_1232);
and U1598 (N_1598,In_1065,In_1221);
xnor U1599 (N_1599,In_247,N_729);
nor U1600 (N_1600,In_1981,N_1145);
nand U1601 (N_1601,N_1516,N_149);
and U1602 (N_1602,N_513,N_1029);
or U1603 (N_1603,N_1345,In_1402);
nand U1604 (N_1604,N_1412,N_1538);
nor U1605 (N_1605,N_1480,N_1405);
nand U1606 (N_1606,N_1569,N_1561);
xor U1607 (N_1607,In_28,N_1521);
xnor U1608 (N_1608,In_1344,N_189);
nand U1609 (N_1609,In_910,N_1572);
nand U1610 (N_1610,N_1047,In_66);
xor U1611 (N_1611,N_1135,N_1306);
and U1612 (N_1612,In_381,N_1431);
nor U1613 (N_1613,In_700,In_1520);
or U1614 (N_1614,In_192,N_1483);
nor U1615 (N_1615,N_857,N_896);
xor U1616 (N_1616,N_1507,N_491);
nor U1617 (N_1617,N_1419,N_1531);
and U1618 (N_1618,In_2142,N_508);
nor U1619 (N_1619,N_1240,N_1017);
and U1620 (N_1620,In_1354,N_1086);
xor U1621 (N_1621,In_432,N_1568);
and U1622 (N_1622,N_1284,N_1131);
or U1623 (N_1623,N_49,In_437);
and U1624 (N_1624,In_1917,N_1459);
or U1625 (N_1625,N_1560,N_1410);
or U1626 (N_1626,N_1577,N_1403);
xor U1627 (N_1627,N_1158,N_710);
and U1628 (N_1628,N_1341,N_723);
nor U1629 (N_1629,N_1185,In_710);
and U1630 (N_1630,N_1100,In_731);
or U1631 (N_1631,N_859,N_1124);
nand U1632 (N_1632,N_187,N_1160);
nand U1633 (N_1633,N_1265,N_1536);
or U1634 (N_1634,In_558,N_1375);
or U1635 (N_1635,In_1380,In_1477);
or U1636 (N_1636,In_1488,N_1468);
nand U1637 (N_1637,N_622,N_463);
nor U1638 (N_1638,In_639,N_1563);
and U1639 (N_1639,N_1291,N_292);
and U1640 (N_1640,N_726,N_1077);
or U1641 (N_1641,N_1585,In_1966);
nand U1642 (N_1642,N_1498,In_2172);
nor U1643 (N_1643,In_923,N_1201);
nor U1644 (N_1644,N_1202,In_1631);
xor U1645 (N_1645,N_1334,N_372);
nand U1646 (N_1646,In_738,N_921);
xor U1647 (N_1647,In_903,N_55);
nor U1648 (N_1648,In_1879,N_285);
nor U1649 (N_1649,In_47,In_1510);
nor U1650 (N_1650,N_1225,N_851);
or U1651 (N_1651,N_1557,N_1511);
nand U1652 (N_1652,N_1462,N_1268);
or U1653 (N_1653,In_1781,N_300);
or U1654 (N_1654,N_1490,In_2053);
nor U1655 (N_1655,In_1541,In_2182);
nand U1656 (N_1656,N_526,N_1233);
or U1657 (N_1657,In_279,N_1484);
xor U1658 (N_1658,N_556,In_176);
nand U1659 (N_1659,N_1386,N_1552);
nand U1660 (N_1660,N_1413,N_1472);
or U1661 (N_1661,In_498,In_958);
and U1662 (N_1662,N_1443,N_1323);
or U1663 (N_1663,N_1244,In_1475);
nand U1664 (N_1664,N_1452,N_1238);
and U1665 (N_1665,N_1302,N_221);
and U1666 (N_1666,N_1358,N_1456);
nor U1667 (N_1667,N_1574,N_200);
nand U1668 (N_1668,N_355,N_1294);
xor U1669 (N_1669,N_1281,N_1046);
nand U1670 (N_1670,N_1280,N_265);
or U1671 (N_1671,N_380,N_876);
or U1672 (N_1672,N_511,In_765);
nand U1673 (N_1673,N_1153,N_1525);
or U1674 (N_1674,In_229,N_93);
xnor U1675 (N_1675,In_1298,N_885);
nand U1676 (N_1676,In_2395,In_1950);
or U1677 (N_1677,N_1081,N_982);
or U1678 (N_1678,In_1736,N_911);
or U1679 (N_1679,N_1204,In_680);
nand U1680 (N_1680,N_1303,N_1305);
nor U1681 (N_1681,N_1488,In_1547);
nand U1682 (N_1682,N_1286,In_900);
and U1683 (N_1683,In_861,N_958);
nand U1684 (N_1684,N_1365,In_1145);
and U1685 (N_1685,N_1369,In_275);
nor U1686 (N_1686,In_1629,N_935);
and U1687 (N_1687,N_469,N_1257);
nand U1688 (N_1688,N_1074,In_44);
nand U1689 (N_1689,N_694,N_1082);
or U1690 (N_1690,N_1283,N_1473);
and U1691 (N_1691,N_505,N_678);
or U1692 (N_1692,In_946,N_1466);
nand U1693 (N_1693,N_1036,N_393);
xnor U1694 (N_1694,N_1328,N_1293);
nand U1695 (N_1695,N_835,In_1215);
nor U1696 (N_1696,N_1290,N_535);
or U1697 (N_1697,N_495,In_750);
or U1698 (N_1698,In_2105,N_1300);
nor U1699 (N_1699,N_1493,N_361);
and U1700 (N_1700,N_1565,N_521);
or U1701 (N_1701,N_1562,N_1515);
or U1702 (N_1702,N_1475,In_2297);
nor U1703 (N_1703,N_1355,N_677);
and U1704 (N_1704,N_1555,N_879);
and U1705 (N_1705,N_1009,N_1226);
nand U1706 (N_1706,N_1344,In_1407);
or U1707 (N_1707,N_1471,N_1353);
or U1708 (N_1708,In_2374,N_1148);
xor U1709 (N_1709,N_346,N_1556);
nor U1710 (N_1710,N_1254,In_1764);
xnor U1711 (N_1711,N_1298,N_1380);
xor U1712 (N_1712,N_1430,In_1910);
and U1713 (N_1713,N_1000,N_1297);
nor U1714 (N_1714,N_1486,In_1928);
nand U1715 (N_1715,In_1124,N_1465);
and U1716 (N_1716,N_1083,N_198);
and U1717 (N_1717,In_1081,In_2442);
nand U1718 (N_1718,N_1575,N_1464);
xnor U1719 (N_1719,N_1513,N_1308);
or U1720 (N_1720,N_1379,N_1205);
xor U1721 (N_1721,N_1357,N_803);
or U1722 (N_1722,In_1773,N_1098);
or U1723 (N_1723,N_493,In_702);
or U1724 (N_1724,N_1285,In_1038);
and U1725 (N_1725,N_1421,N_1112);
nor U1726 (N_1726,In_897,N_834);
and U1727 (N_1727,N_766,In_1641);
or U1728 (N_1728,N_1438,N_1442);
nor U1729 (N_1729,N_904,In_1193);
and U1730 (N_1730,In_1542,N_1126);
nand U1731 (N_1731,N_1385,N_1330);
or U1732 (N_1732,N_1203,N_1044);
nand U1733 (N_1733,N_1542,N_1482);
and U1734 (N_1734,In_1675,In_1860);
nor U1735 (N_1735,In_147,In_1276);
or U1736 (N_1736,N_843,In_372);
or U1737 (N_1737,N_470,In_798);
or U1738 (N_1738,In_1551,In_87);
and U1739 (N_1739,In_91,N_1110);
and U1740 (N_1740,N_1064,In_2244);
and U1741 (N_1741,N_561,In_141);
xnor U1742 (N_1742,In_513,N_891);
xor U1743 (N_1743,N_482,N_173);
xor U1744 (N_1744,N_798,In_1705);
xor U1745 (N_1745,In_2477,N_237);
nand U1746 (N_1746,N_1502,N_1304);
and U1747 (N_1747,N_1080,N_565);
nand U1748 (N_1748,N_1351,In_1995);
and U1749 (N_1749,N_1287,N_369);
and U1750 (N_1750,In_1793,N_1467);
nand U1751 (N_1751,N_1549,N_1530);
and U1752 (N_1752,In_1278,N_1059);
and U1753 (N_1753,In_34,N_1331);
and U1754 (N_1754,N_193,N_1517);
nand U1755 (N_1755,N_1010,N_1477);
xor U1756 (N_1756,N_699,In_1079);
nand U1757 (N_1757,N_1023,N_778);
nor U1758 (N_1758,N_1559,In_2494);
nor U1759 (N_1759,N_1262,N_973);
and U1760 (N_1760,N_736,N_1169);
and U1761 (N_1761,N_1527,N_252);
and U1762 (N_1762,N_1018,N_1236);
nor U1763 (N_1763,N_964,N_1455);
nand U1764 (N_1764,In_1012,N_1445);
and U1765 (N_1765,N_1253,In_352);
and U1766 (N_1766,N_1453,N_1325);
xor U1767 (N_1767,N_1210,N_405);
or U1768 (N_1768,In_1495,In_295);
nor U1769 (N_1769,N_1383,In_1028);
nor U1770 (N_1770,In_945,N_1554);
or U1771 (N_1771,N_1359,N_1251);
nand U1772 (N_1772,N_1474,N_1596);
nand U1773 (N_1773,In_1281,N_1424);
and U1774 (N_1774,N_1399,N_1267);
xnor U1775 (N_1775,N_979,N_1252);
nor U1776 (N_1776,N_1537,In_2002);
and U1777 (N_1777,N_1415,N_769);
nor U1778 (N_1778,N_1546,In_1620);
nand U1779 (N_1779,N_1460,N_1387);
or U1780 (N_1780,N_985,N_1506);
or U1781 (N_1781,N_1503,In_2091);
nor U1782 (N_1782,In_366,N_1487);
xnor U1783 (N_1783,In_981,N_1500);
nor U1784 (N_1784,In_2485,N_150);
nand U1785 (N_1785,In_1662,N_1558);
and U1786 (N_1786,In_878,N_1350);
and U1787 (N_1787,N_464,N_1441);
xnor U1788 (N_1788,N_662,N_1220);
nand U1789 (N_1789,N_639,N_1544);
or U1790 (N_1790,In_268,N_1398);
or U1791 (N_1791,N_1005,N_1067);
or U1792 (N_1792,N_1588,N_940);
and U1793 (N_1793,N_1512,N_1371);
and U1794 (N_1794,N_1520,N_807);
xnor U1795 (N_1795,N_1213,N_887);
and U1796 (N_1796,In_398,In_1798);
nand U1797 (N_1797,N_610,N_942);
or U1798 (N_1798,N_824,In_1149);
and U1799 (N_1799,N_81,N_1377);
or U1800 (N_1800,N_785,N_687);
xor U1801 (N_1801,N_772,N_1645);
xnor U1802 (N_1802,N_1121,N_628);
nand U1803 (N_1803,N_256,N_1695);
or U1804 (N_1804,N_1598,In_2222);
or U1805 (N_1805,N_110,N_1635);
or U1806 (N_1806,N_1339,N_258);
xor U1807 (N_1807,N_1783,In_545);
nor U1808 (N_1808,N_566,In_976);
and U1809 (N_1809,In_267,N_1616);
nor U1810 (N_1810,N_462,N_1611);
or U1811 (N_1811,N_304,N_245);
and U1812 (N_1812,N_1676,N_1672);
nand U1813 (N_1813,In_159,In_2262);
nor U1814 (N_1814,N_1102,N_1681);
or U1815 (N_1815,N_1151,N_1657);
and U1816 (N_1816,N_1043,N_1685);
or U1817 (N_1817,In_1222,N_1505);
and U1818 (N_1818,N_1794,N_654);
and U1819 (N_1819,N_419,N_976);
or U1820 (N_1820,N_1168,N_1763);
nand U1821 (N_1821,In_1677,N_342);
xor U1822 (N_1822,In_1339,In_1259);
nor U1823 (N_1823,N_1449,N_233);
and U1824 (N_1824,In_816,N_479);
or U1825 (N_1825,N_1687,N_536);
nand U1826 (N_1826,N_672,In_2128);
nand U1827 (N_1827,In_496,N_1495);
nand U1828 (N_1828,N_826,N_1016);
nor U1829 (N_1829,N_1663,In_610);
xor U1830 (N_1830,N_1715,N_194);
and U1831 (N_1831,N_1388,N_1289);
or U1832 (N_1832,N_1790,N_1277);
xnor U1833 (N_1833,In_776,N_937);
and U1834 (N_1834,N_1650,N_1605);
nand U1835 (N_1835,N_1646,N_1765);
or U1836 (N_1836,N_1658,N_1423);
or U1837 (N_1837,N_191,In_1959);
nor U1838 (N_1838,N_1458,N_1701);
or U1839 (N_1839,N_1602,N_1592);
xnor U1840 (N_1840,N_1476,N_1797);
and U1841 (N_1841,N_1750,N_1677);
or U1842 (N_1842,N_1723,In_2429);
nor U1843 (N_1843,In_2071,N_1407);
or U1844 (N_1844,N_910,N_1670);
nor U1845 (N_1845,N_853,In_2451);
xor U1846 (N_1846,N_1187,N_1533);
and U1847 (N_1847,N_991,N_1347);
nor U1848 (N_1848,N_1579,N_1744);
nand U1849 (N_1849,N_1626,In_1352);
and U1850 (N_1850,In_1095,N_1751);
nor U1851 (N_1851,N_1393,N_1796);
and U1852 (N_1852,N_1524,N_1128);
xnor U1853 (N_1853,N_1724,N_1649);
or U1854 (N_1854,N_1710,N_1633);
nor U1855 (N_1855,N_599,In_1689);
nand U1856 (N_1856,N_625,N_805);
nor U1857 (N_1857,N_1582,N_1694);
xnor U1858 (N_1858,N_1778,N_1746);
or U1859 (N_1859,N_1665,N_1668);
nor U1860 (N_1860,N_1313,N_1450);
xor U1861 (N_1861,In_93,N_635);
nor U1862 (N_1862,N_1640,N_1402);
xor U1863 (N_1863,N_1214,In_412);
or U1864 (N_1864,In_1082,N_182);
nand U1865 (N_1865,In_1002,N_1338);
nor U1866 (N_1866,In_429,N_1491);
nand U1867 (N_1867,In_514,N_1311);
or U1868 (N_1868,N_1704,In_2302);
nand U1869 (N_1869,N_1461,N_1779);
nor U1870 (N_1870,N_457,N_706);
nand U1871 (N_1871,N_1752,N_1447);
or U1872 (N_1872,In_1775,In_82);
xor U1873 (N_1873,N_1729,N_758);
or U1874 (N_1874,In_746,N_586);
xor U1875 (N_1875,N_1113,In_659);
and U1876 (N_1876,N_1606,N_1095);
xor U1877 (N_1877,N_1381,N_1094);
xor U1878 (N_1878,N_1489,N_1444);
or U1879 (N_1879,N_1767,In_2404);
and U1880 (N_1880,N_1734,N_1326);
xor U1881 (N_1881,N_1706,In_2247);
nor U1882 (N_1882,In_889,N_1799);
or U1883 (N_1883,In_80,N_1161);
xor U1884 (N_1884,N_1020,N_1578);
nand U1885 (N_1885,N_1659,N_1035);
nand U1886 (N_1886,N_1433,N_299);
nor U1887 (N_1887,In_2333,In_1851);
and U1888 (N_1888,In_31,N_1361);
nor U1889 (N_1889,N_1526,N_532);
nor U1890 (N_1890,N_1548,In_1743);
nand U1891 (N_1891,N_980,N_1599);
xnor U1892 (N_1892,N_1739,N_1508);
nor U1893 (N_1893,In_1099,N_270);
nand U1894 (N_1894,In_1552,N_1228);
xor U1895 (N_1895,In_485,N_1691);
nand U1896 (N_1896,N_1197,N_1221);
and U1897 (N_1897,In_1967,N_1152);
nor U1898 (N_1898,N_138,N_435);
or U1899 (N_1899,N_573,In_2059);
nor U1900 (N_1900,N_1781,In_79);
nor U1901 (N_1901,In_1385,N_1553);
and U1902 (N_1902,N_1780,N_1261);
or U1903 (N_1903,N_1680,N_1697);
xor U1904 (N_1904,N_1636,N_1411);
xnor U1905 (N_1905,In_1868,N_984);
xor U1906 (N_1906,In_1307,In_62);
nor U1907 (N_1907,N_231,N_1545);
nand U1908 (N_1908,In_178,N_1586);
xnor U1909 (N_1909,N_1688,N_1373);
nand U1910 (N_1910,N_1089,N_1396);
nand U1911 (N_1911,N_1567,N_1429);
nor U1912 (N_1912,In_1655,N_1768);
nor U1913 (N_1913,N_854,N_1535);
or U1914 (N_1914,N_1497,N_1745);
nand U1915 (N_1915,In_1261,N_1470);
or U1916 (N_1916,In_1591,In_797);
xnor U1917 (N_1917,N_974,N_1634);
xnor U1918 (N_1918,N_1726,N_1454);
nand U1919 (N_1919,N_1107,N_11);
or U1920 (N_1920,N_1532,N_1076);
nand U1921 (N_1921,N_1427,In_1044);
and U1922 (N_1922,N_525,N_1620);
xnor U1923 (N_1923,N_1719,N_1566);
xnor U1924 (N_1924,N_753,In_1100);
nand U1925 (N_1925,N_1481,N_1469);
and U1926 (N_1926,N_260,N_1621);
nand U1927 (N_1927,N_1492,In_1335);
nor U1928 (N_1928,N_473,N_1275);
or U1929 (N_1929,In_2331,N_1730);
nor U1930 (N_1930,N_1440,In_675);
xor U1931 (N_1931,N_791,N_1321);
nand U1932 (N_1932,N_1266,N_787);
and U1933 (N_1933,N_1600,In_1486);
xor U1934 (N_1934,N_428,N_1212);
or U1935 (N_1935,N_946,In_1054);
xnor U1936 (N_1936,N_1312,In_420);
or U1937 (N_1937,N_712,N_362);
nand U1938 (N_1938,N_1501,N_1451);
nor U1939 (N_1939,N_1777,In_1369);
nand U1940 (N_1940,In_896,N_1661);
nand U1941 (N_1941,In_343,N_1753);
nor U1942 (N_1942,N_1591,N_1594);
and U1943 (N_1943,N_1742,N_1038);
or U1944 (N_1944,N_969,N_156);
nand U1945 (N_1945,N_357,N_1696);
xnor U1946 (N_1946,N_1479,In_1506);
and U1947 (N_1947,In_322,In_2070);
or U1948 (N_1948,In_708,N_1581);
or U1949 (N_1949,N_1784,N_1335);
nor U1950 (N_1950,N_1624,In_1322);
and U1951 (N_1951,In_1362,N_1234);
nor U1952 (N_1952,N_1669,N_343);
and U1953 (N_1953,N_1264,N_1732);
nand U1954 (N_1954,N_1774,N_1651);
nand U1955 (N_1955,N_1539,In_2014);
xnor U1956 (N_1956,N_1426,In_690);
xor U1957 (N_1957,N_1711,N_1718);
xnor U1958 (N_1958,N_1609,N_1416);
nor U1959 (N_1959,N_1573,In_1762);
and U1960 (N_1960,N_1514,N_1666);
nand U1961 (N_1961,N_392,N_1655);
nand U1962 (N_1962,N_1485,N_1728);
xnor U1963 (N_1963,N_1769,In_2165);
xnor U1964 (N_1964,In_1169,In_2052);
and U1965 (N_1965,N_1637,N_676);
nand U1966 (N_1966,N_352,N_1793);
and U1967 (N_1967,In_881,N_1625);
nor U1968 (N_1968,N_1703,In_1946);
or U1969 (N_1969,In_2209,N_1408);
xnor U1970 (N_1970,In_461,In_2246);
xnor U1971 (N_1971,N_1654,N_1628);
nor U1972 (N_1972,N_1200,N_1684);
and U1973 (N_1973,N_1764,N_582);
nand U1974 (N_1974,N_1519,In_628);
nand U1975 (N_1975,In_1131,N_1644);
and U1976 (N_1976,N_895,N_537);
nand U1977 (N_1977,N_1648,N_1643);
or U1978 (N_1978,N_1589,N_1617);
nand U1979 (N_1979,N_102,N_1317);
nor U1980 (N_1980,In_317,N_1522);
xnor U1981 (N_1981,N_1708,N_1656);
or U1982 (N_1982,N_1420,N_840);
or U1983 (N_1983,N_1692,N_1771);
nor U1984 (N_1984,N_211,In_2362);
xor U1985 (N_1985,N_1105,In_2163);
xnor U1986 (N_1986,In_259,N_1721);
nand U1987 (N_1987,N_1641,N_1406);
or U1988 (N_1988,N_1478,N_1630);
and U1989 (N_1989,N_422,In_1238);
nand U1990 (N_1990,N_1288,N_1259);
or U1991 (N_1991,In_943,N_289);
nand U1992 (N_1992,In_1273,N_1798);
xor U1993 (N_1993,N_257,N_1595);
nand U1994 (N_1994,N_1143,N_46);
nor U1995 (N_1995,N_1571,N_1773);
and U1996 (N_1996,N_1698,N_1610);
nand U1997 (N_1997,N_1570,N_847);
and U1998 (N_1998,N_1523,N_1702);
nand U1999 (N_1999,N_1418,N_1401);
nand U2000 (N_2000,N_1985,N_1132);
and U2001 (N_2001,N_1738,N_1812);
nand U2002 (N_2002,N_1065,N_88);
nor U2003 (N_2003,N_951,In_2107);
nand U2004 (N_2004,N_1935,N_458);
or U2005 (N_2005,N_1856,N_1088);
nand U2006 (N_2006,N_1766,In_2136);
xnor U2007 (N_2007,N_1873,In_555);
xor U2008 (N_2008,N_1564,N_1936);
and U2009 (N_2009,N_659,In_2092);
or U2010 (N_2010,N_1918,N_1968);
nand U2011 (N_2011,N_1912,N_1975);
or U2012 (N_2012,N_1436,N_450);
nor U2013 (N_2013,N_637,N_1587);
nand U2014 (N_2014,N_1979,N_771);
nor U2015 (N_2015,N_1758,N_1788);
nand U2016 (N_2016,N_1896,In_1229);
nand U2017 (N_2017,N_1550,N_1925);
nor U2018 (N_2018,N_1820,N_1866);
or U2019 (N_2019,N_1978,N_1805);
nand U2020 (N_2020,N_1987,N_1853);
xnor U2021 (N_2021,N_1930,N_1953);
or U2022 (N_2022,N_1583,N_1826);
or U2023 (N_2023,N_1053,N_1825);
xnor U2024 (N_2024,N_1816,N_1690);
nand U2025 (N_2025,N_1888,N_1660);
nor U2026 (N_2026,N_1754,N_1755);
nand U2027 (N_2027,N_1786,N_1824);
and U2028 (N_2028,N_1908,N_1905);
or U2029 (N_2029,In_403,N_1707);
xor U2030 (N_2030,N_1971,N_670);
nand U2031 (N_2031,N_1422,N_1384);
nand U2032 (N_2032,In_1634,N_516);
xnor U2033 (N_2033,N_998,N_1007);
xor U2034 (N_2034,N_1638,N_1910);
nand U2035 (N_2035,N_1727,N_1872);
xnor U2036 (N_2036,N_1913,N_1980);
or U2037 (N_2037,N_1604,N_1540);
and U2038 (N_2038,N_1770,N_1960);
nand U2039 (N_2039,N_1404,N_1869);
or U2040 (N_2040,N_1863,In_1886);
or U2041 (N_2041,N_1852,N_1997);
xor U2042 (N_2042,N_1400,N_1881);
nand U2043 (N_2043,N_1607,N_1884);
xnor U2044 (N_2044,N_1915,N_1921);
xor U2045 (N_2045,N_1808,N_1722);
or U2046 (N_2046,N_1109,N_1923);
nand U2047 (N_2047,N_1518,N_1885);
or U2048 (N_2048,N_1622,N_1875);
and U2049 (N_2049,N_1759,N_1686);
xor U2050 (N_2050,In_1951,N_538);
and U2051 (N_2051,N_1463,N_1528);
xnor U2052 (N_2052,N_1917,In_1422);
and U2053 (N_2053,N_1874,N_203);
or U2054 (N_2054,N_1998,In_528);
and U2055 (N_2055,N_883,N_1022);
xnor U2056 (N_2056,N_1850,N_1822);
or U2057 (N_2057,N_1689,N_1270);
nand U2058 (N_2058,N_1301,In_2449);
nor U2059 (N_2059,N_1206,N_1725);
and U2060 (N_2060,In_1304,In_855);
nand U2061 (N_2061,N_888,N_1352);
nor U2062 (N_2062,N_1409,N_1776);
and U2063 (N_2063,N_1819,N_1748);
xnor U2064 (N_2064,N_1841,N_316);
xor U2065 (N_2065,N_1977,N_1815);
nor U2066 (N_2066,N_1509,N_1846);
nor U2067 (N_2067,N_1804,N_1961);
and U2068 (N_2068,N_1337,In_560);
xnor U2069 (N_2069,In_1178,N_1584);
nand U2070 (N_2070,N_1551,N_1828);
nor U2071 (N_2071,N_1760,N_1966);
xnor U2072 (N_2072,N_950,N_1929);
or U2073 (N_2073,N_20,N_1123);
nand U2074 (N_2074,N_1807,N_1832);
or U2075 (N_2075,N_1614,N_1747);
nand U2076 (N_2076,N_1191,N_1623);
or U2077 (N_2077,N_1207,N_1861);
nand U2078 (N_2078,N_1897,N_1843);
nand U2079 (N_2079,N_1911,N_1830);
nor U2080 (N_2080,N_1889,N_1955);
or U2081 (N_2081,N_737,N_1900);
and U2082 (N_2082,N_1700,In_1693);
xnor U2083 (N_2083,N_1683,In_655);
nor U2084 (N_2084,N_1821,N_1833);
nand U2085 (N_2085,N_1877,N_1868);
xnor U2086 (N_2086,N_1982,N_1954);
nand U2087 (N_2087,N_1962,N_1792);
xnor U2088 (N_2088,N_1292,N_1615);
or U2089 (N_2089,N_1227,N_1757);
nor U2090 (N_2090,N_1899,N_681);
or U2091 (N_2091,N_1392,In_425);
and U2092 (N_2092,N_1397,N_907);
xor U2093 (N_2093,N_1716,N_452);
and U2094 (N_2094,N_1504,In_2124);
nand U2095 (N_2095,N_870,N_1943);
or U2096 (N_2096,N_1879,N_1272);
nand U2097 (N_2097,N_1248,N_1741);
xor U2098 (N_2098,N_1880,N_1597);
nand U2099 (N_2099,N_1772,N_1906);
nand U2100 (N_2100,N_1231,In_695);
xor U2101 (N_2101,N_1051,N_1639);
nor U2102 (N_2102,N_1886,N_1496);
nor U2103 (N_2103,N_1803,In_1902);
xor U2104 (N_2104,N_1994,N_1895);
nor U2105 (N_2105,N_1999,N_1740);
nor U2106 (N_2106,N_1414,N_293);
and U2107 (N_2107,N_665,N_1878);
or U2108 (N_2108,In_842,N_1827);
or U2109 (N_2109,In_839,N_1848);
nand U2110 (N_2110,N_1731,N_1125);
or U2111 (N_2111,N_1909,N_1838);
or U2112 (N_2112,In_1455,N_1933);
and U2113 (N_2113,N_1801,N_1847);
xor U2114 (N_2114,N_1939,N_41);
nor U2115 (N_2115,N_1806,N_1845);
and U2116 (N_2116,In_1411,N_1984);
xor U2117 (N_2117,In_137,In_2287);
nand U2118 (N_2118,N_1632,N_1762);
nor U2119 (N_2119,N_919,N_1810);
nand U2120 (N_2120,N_1432,N_1919);
and U2121 (N_2121,N_1457,N_1316);
and U2122 (N_2122,N_126,In_2288);
or U2123 (N_2123,N_1800,In_927);
nand U2124 (N_2124,N_1749,N_832);
nand U2125 (N_2125,N_1876,N_1831);
and U2126 (N_2126,N_1219,N_1678);
and U2127 (N_2127,In_2149,N_751);
or U2128 (N_2128,N_1603,N_1989);
or U2129 (N_2129,N_1667,N_1958);
and U2130 (N_2130,N_1986,N_1499);
nor U2131 (N_2131,N_1926,N_1934);
nand U2132 (N_2132,N_1970,N_1817);
nand U2133 (N_2133,N_1260,N_1947);
and U2134 (N_2134,N_1743,In_1279);
nor U2135 (N_2135,N_1855,N_1756);
and U2136 (N_2136,N_1271,N_1942);
nor U2137 (N_2137,N_1995,N_1618);
nand U2138 (N_2138,In_807,N_871);
nor U2139 (N_2139,N_618,N_1950);
and U2140 (N_2140,N_1834,N_1653);
xor U2141 (N_2141,N_1674,N_1883);
xor U2142 (N_2142,N_1836,N_1705);
nand U2143 (N_2143,N_1775,N_1096);
or U2144 (N_2144,N_1829,N_1647);
nand U2145 (N_2145,N_1627,N_1945);
nor U2146 (N_2146,N_1964,N_181);
xnor U2147 (N_2147,N_1898,N_1837);
nand U2148 (N_2148,N_1679,In_524);
nand U2149 (N_2149,In_1593,N_1996);
or U2150 (N_2150,N_1320,N_1033);
or U2151 (N_2151,N_1782,In_262);
xor U2152 (N_2152,N_1682,N_1787);
nand U2153 (N_2153,N_1543,N_291);
or U2154 (N_2154,N_1435,N_1437);
nor U2155 (N_2155,N_1417,N_1693);
and U2156 (N_2156,N_1318,In_541);
nor U2157 (N_2157,N_1991,N_1811);
or U2158 (N_2158,N_1901,N_1547);
or U2159 (N_2159,N_1071,N_914);
or U2160 (N_2160,N_720,N_1671);
nand U2161 (N_2161,N_1946,N_1860);
or U2162 (N_2162,N_949,N_1174);
nand U2163 (N_2163,In_189,N_827);
or U2164 (N_2164,N_1887,N_1211);
xor U2165 (N_2165,N_1903,N_1892);
and U2166 (N_2166,In_1789,In_1581);
nand U2167 (N_2167,N_1529,N_1941);
and U2168 (N_2168,N_1642,N_1354);
nand U2169 (N_2169,N_1840,N_1949);
xor U2170 (N_2170,N_1717,N_106);
nor U2171 (N_2171,N_1951,In_939);
and U2172 (N_2172,N_1448,N_1814);
and U2173 (N_2173,N_1714,N_1720);
or U2174 (N_2174,N_1363,N_1931);
nand U2175 (N_2175,N_1809,N_1871);
or U2176 (N_2176,N_12,N_1372);
xor U2177 (N_2177,N_806,N_1315);
nor U2178 (N_2178,In_1819,N_1904);
and U2179 (N_2179,N_1791,N_1541);
xnor U2180 (N_2180,In_2089,N_1601);
or U2181 (N_2181,N_1130,N_1613);
nand U2182 (N_2182,N_1246,N_1425);
xnor U2183 (N_2183,N_1382,N_1170);
xor U2184 (N_2184,N_1673,In_2019);
nor U2185 (N_2185,N_1631,N_838);
and U2186 (N_2186,N_1733,N_1057);
nand U2187 (N_2187,N_1510,N_1854);
and U2188 (N_2188,N_1844,N_1963);
nand U2189 (N_2189,N_1835,In_2134);
nor U2190 (N_2190,In_677,N_1222);
nor U2191 (N_2191,N_1608,N_1859);
xnor U2192 (N_2192,N_1920,N_1223);
nand U2193 (N_2193,N_1851,N_1818);
or U2194 (N_2194,N_1969,N_1914);
or U2195 (N_2195,N_1736,N_1590);
nand U2196 (N_2196,N_1619,N_1785);
xnor U2197 (N_2197,N_1882,N_1823);
and U2198 (N_2198,N_1864,N_1894);
and U2199 (N_2199,N_1737,N_1972);
or U2200 (N_2200,N_2090,N_2037);
or U2201 (N_2201,N_2070,N_2033);
and U2202 (N_2202,N_2125,N_1938);
nor U2203 (N_2203,N_2049,N_2130);
xnor U2204 (N_2204,N_2139,N_2088);
or U2205 (N_2205,N_1937,N_2013);
nand U2206 (N_2206,N_1857,N_2054);
or U2207 (N_2207,N_2092,N_2136);
nor U2208 (N_2208,N_2069,N_1849);
nor U2209 (N_2209,N_2132,In_1985);
nor U2210 (N_2210,N_2095,N_1983);
xor U2211 (N_2211,N_1870,N_2005);
nor U2212 (N_2212,N_2034,N_2190);
xnor U2213 (N_2213,N_2015,N_2039);
nand U2214 (N_2214,N_2177,N_2166);
or U2215 (N_2215,In_467,N_1922);
nor U2216 (N_2216,N_1927,N_2111);
nor U2217 (N_2217,N_2179,N_1993);
nor U2218 (N_2218,N_2170,N_2060);
xor U2219 (N_2219,N_1111,N_2145);
or U2220 (N_2220,N_2147,N_1208);
and U2221 (N_2221,N_2083,N_1944);
and U2222 (N_2222,N_1924,N_2189);
or U2223 (N_2223,N_2064,N_684);
nor U2224 (N_2224,N_2178,N_1956);
and U2225 (N_2225,N_2063,N_2097);
nor U2226 (N_2226,N_1865,N_2146);
nor U2227 (N_2227,N_1990,N_1957);
xor U2228 (N_2228,N_2086,N_1974);
nor U2229 (N_2229,N_2161,N_2058);
or U2230 (N_2230,N_2142,N_2062);
and U2231 (N_2231,N_2038,N_2183);
nand U2232 (N_2232,N_1867,N_2100);
or U2233 (N_2233,N_1858,N_2074);
or U2234 (N_2234,N_2109,N_1699);
and U2235 (N_2235,N_1959,N_2162);
nor U2236 (N_2236,N_2067,N_1434);
or U2237 (N_2237,N_1439,In_2444);
xor U2238 (N_2238,N_1712,N_1675);
or U2239 (N_2239,N_2157,N_2078);
xnor U2240 (N_2240,N_1662,N_2126);
or U2241 (N_2241,N_2027,N_2112);
nand U2242 (N_2242,N_1713,N_2003);
xnor U2243 (N_2243,N_1390,N_2061);
nor U2244 (N_2244,N_2007,N_2047);
nor U2245 (N_2245,N_533,N_340);
or U2246 (N_2246,N_2175,N_2023);
nor U2247 (N_2247,N_2030,N_2093);
xnor U2248 (N_2248,N_2152,N_1928);
nor U2249 (N_2249,N_1789,N_1139);
or U2250 (N_2250,N_2169,N_2068);
nand U2251 (N_2251,N_2050,N_2123);
nand U2252 (N_2252,N_559,N_2022);
xor U2253 (N_2253,N_2160,N_2087);
and U2254 (N_2254,N_2052,N_2041);
nor U2255 (N_2255,N_2148,N_1967);
xor U2256 (N_2256,N_1916,N_2188);
nand U2257 (N_2257,N_2104,N_2153);
nand U2258 (N_2258,N_2131,N_1342);
and U2259 (N_2259,N_2105,N_2017);
or U2260 (N_2260,N_2110,N_2138);
nor U2261 (N_2261,N_2091,N_2133);
nor U2262 (N_2262,N_2084,N_1243);
xnor U2263 (N_2263,N_2102,N_1902);
nand U2264 (N_2264,N_2118,N_1629);
nor U2265 (N_2265,N_2071,N_2024);
and U2266 (N_2266,N_2196,N_1981);
nor U2267 (N_2267,N_2099,N_2122);
xor U2268 (N_2268,N_2186,N_2141);
nor U2269 (N_2269,N_2085,N_828);
nor U2270 (N_2270,N_2168,N_2075);
nand U2271 (N_2271,N_1952,N_2098);
nand U2272 (N_2272,N_1795,N_2001);
or U2273 (N_2273,N_2018,In_97);
xnor U2274 (N_2274,N_2040,N_2191);
xor U2275 (N_2275,N_2020,N_2029);
or U2276 (N_2276,N_2011,N_2171);
and U2277 (N_2277,N_1976,N_1127);
or U2278 (N_2278,N_841,In_1080);
xnor U2279 (N_2279,N_2077,N_2006);
xor U2280 (N_2280,N_2094,N_2198);
and U2281 (N_2281,N_1198,N_2158);
or U2282 (N_2282,N_2080,N_2000);
nand U2283 (N_2283,N_2009,N_2172);
xnor U2284 (N_2284,N_2036,N_1664);
nand U2285 (N_2285,N_2032,N_2079);
xor U2286 (N_2286,N_2159,N_2059);
or U2287 (N_2287,N_1032,N_2180);
nand U2288 (N_2288,N_1652,N_2140);
nor U2289 (N_2289,N_2010,N_2115);
nand U2290 (N_2290,N_2025,N_2002);
xnor U2291 (N_2291,N_2154,N_2117);
nand U2292 (N_2292,N_2127,N_2045);
nor U2293 (N_2293,N_2046,In_1244);
nor U2294 (N_2294,N_1012,N_286);
nor U2295 (N_2295,N_2103,N_2164);
nand U2296 (N_2296,In_1646,N_2173);
nor U2297 (N_2297,N_2129,N_2012);
xor U2298 (N_2298,N_1992,In_140);
xor U2299 (N_2299,N_861,N_2134);
nand U2300 (N_2300,N_2081,N_1940);
nor U2301 (N_2301,N_2185,N_2195);
or U2302 (N_2302,N_2113,N_682);
and U2303 (N_2303,N_2187,N_1890);
or U2304 (N_2304,N_2128,N_2014);
xnor U2305 (N_2305,N_2051,N_2016);
nor U2306 (N_2306,N_82,N_2026);
or U2307 (N_2307,N_1965,In_256);
and U2308 (N_2308,N_1893,N_1761);
and U2309 (N_2309,N_2124,N_2082);
nand U2310 (N_2310,N_2116,N_2199);
xnor U2311 (N_2311,N_2072,N_2055);
nor U2312 (N_2312,N_2031,N_2021);
nor U2313 (N_2313,N_2076,N_2089);
xnor U2314 (N_2314,N_2065,N_1948);
nand U2315 (N_2315,N_1709,N_2008);
nand U2316 (N_2316,N_2119,N_2053);
nor U2317 (N_2317,N_2106,N_2004);
nor U2318 (N_2318,N_2197,N_2121);
xor U2319 (N_2319,N_2042,N_2056);
or U2320 (N_2320,N_2035,N_2107);
xor U2321 (N_2321,N_2167,N_1576);
or U2322 (N_2322,N_1534,N_2028);
or U2323 (N_2323,In_2215,N_2156);
nor U2324 (N_2324,N_2163,N_2019);
and U2325 (N_2325,N_2108,N_1593);
xnor U2326 (N_2326,N_1428,N_2066);
nor U2327 (N_2327,N_1862,N_2150);
nand U2328 (N_2328,N_1494,N_2144);
xnor U2329 (N_2329,N_2048,N_1802);
nand U2330 (N_2330,N_2184,N_1932);
nor U2331 (N_2331,N_1988,N_1735);
xnor U2332 (N_2332,N_2114,In_1311);
or U2333 (N_2333,N_1891,N_2192);
and U2334 (N_2334,N_2143,N_1580);
nand U2335 (N_2335,N_2101,N_1612);
xor U2336 (N_2336,N_2135,N_2043);
nand U2337 (N_2337,N_2044,N_1842);
and U2338 (N_2338,N_2182,N_2193);
and U2339 (N_2339,N_2176,N_2096);
xnor U2340 (N_2340,N_1907,N_2174);
nor U2341 (N_2341,N_2165,N_2137);
or U2342 (N_2342,N_1813,N_2120);
nor U2343 (N_2343,N_1199,N_2194);
or U2344 (N_2344,N_2073,N_2149);
xor U2345 (N_2345,In_2033,In_9);
nor U2346 (N_2346,N_849,N_2151);
xnor U2347 (N_2347,N_1839,N_2057);
nor U2348 (N_2348,N_2181,N_1973);
xor U2349 (N_2349,N_1446,N_2155);
nand U2350 (N_2350,N_2123,N_1712);
nor U2351 (N_2351,N_2165,N_1940);
xnor U2352 (N_2352,N_2148,N_2039);
nand U2353 (N_2353,N_2045,N_2194);
xor U2354 (N_2354,N_1593,N_2198);
nand U2355 (N_2355,N_2166,N_2043);
xor U2356 (N_2356,N_1111,N_1446);
nand U2357 (N_2357,N_2097,N_2001);
and U2358 (N_2358,N_2187,N_2035);
xor U2359 (N_2359,N_2086,N_1576);
or U2360 (N_2360,N_1937,N_2017);
or U2361 (N_2361,N_286,N_2079);
or U2362 (N_2362,N_2189,N_2140);
and U2363 (N_2363,N_2097,N_2127);
or U2364 (N_2364,N_1675,N_2130);
xor U2365 (N_2365,N_2132,N_1902);
xnor U2366 (N_2366,N_2130,N_2188);
nand U2367 (N_2367,N_2198,N_2092);
nand U2368 (N_2368,N_2188,N_2015);
nor U2369 (N_2369,N_1802,N_1612);
nand U2370 (N_2370,N_2115,N_2085);
and U2371 (N_2371,N_2167,N_1428);
xor U2372 (N_2372,N_2058,N_1795);
xnor U2373 (N_2373,N_2085,N_2093);
nor U2374 (N_2374,N_2091,N_2191);
nor U2375 (N_2375,N_2103,N_2173);
and U2376 (N_2376,N_1870,N_1439);
xor U2377 (N_2377,N_2170,N_2134);
and U2378 (N_2378,N_828,N_2126);
nor U2379 (N_2379,N_2079,N_1652);
nand U2380 (N_2380,N_2127,In_1985);
nand U2381 (N_2381,N_2123,N_2186);
and U2382 (N_2382,N_2198,N_2187);
xnor U2383 (N_2383,N_2071,N_2155);
nor U2384 (N_2384,N_2052,In_2215);
nor U2385 (N_2385,N_2038,N_2142);
nor U2386 (N_2386,N_1439,N_2183);
and U2387 (N_2387,In_1985,N_2023);
nand U2388 (N_2388,N_1208,N_2158);
nand U2389 (N_2389,N_2031,N_2099);
xnor U2390 (N_2390,N_2135,N_2138);
or U2391 (N_2391,N_2077,N_2141);
or U2392 (N_2392,N_2067,N_2175);
or U2393 (N_2393,N_2087,N_1629);
nand U2394 (N_2394,N_2102,N_2084);
xnor U2395 (N_2395,N_1494,N_2188);
and U2396 (N_2396,N_2049,N_2124);
xnor U2397 (N_2397,N_2199,N_1890);
nor U2398 (N_2398,N_2068,N_1993);
xnor U2399 (N_2399,N_1967,N_2016);
nor U2400 (N_2400,N_2276,N_2340);
or U2401 (N_2401,N_2300,N_2361);
or U2402 (N_2402,N_2239,N_2255);
and U2403 (N_2403,N_2253,N_2345);
nand U2404 (N_2404,N_2307,N_2346);
and U2405 (N_2405,N_2310,N_2221);
and U2406 (N_2406,N_2257,N_2210);
and U2407 (N_2407,N_2241,N_2291);
or U2408 (N_2408,N_2285,N_2201);
nor U2409 (N_2409,N_2322,N_2295);
nor U2410 (N_2410,N_2288,N_2242);
nand U2411 (N_2411,N_2219,N_2353);
nor U2412 (N_2412,N_2309,N_2213);
or U2413 (N_2413,N_2258,N_2304);
and U2414 (N_2414,N_2364,N_2232);
and U2415 (N_2415,N_2325,N_2256);
xor U2416 (N_2416,N_2370,N_2344);
or U2417 (N_2417,N_2275,N_2329);
or U2418 (N_2418,N_2296,N_2246);
and U2419 (N_2419,N_2342,N_2243);
xnor U2420 (N_2420,N_2223,N_2200);
xor U2421 (N_2421,N_2204,N_2284);
or U2422 (N_2422,N_2394,N_2281);
xor U2423 (N_2423,N_2220,N_2274);
and U2424 (N_2424,N_2366,N_2376);
nand U2425 (N_2425,N_2287,N_2374);
nand U2426 (N_2426,N_2356,N_2280);
or U2427 (N_2427,N_2397,N_2308);
nor U2428 (N_2428,N_2264,N_2278);
xnor U2429 (N_2429,N_2339,N_2266);
nor U2430 (N_2430,N_2244,N_2386);
or U2431 (N_2431,N_2251,N_2379);
xor U2432 (N_2432,N_2218,N_2225);
xor U2433 (N_2433,N_2289,N_2303);
nand U2434 (N_2434,N_2240,N_2282);
nand U2435 (N_2435,N_2294,N_2262);
and U2436 (N_2436,N_2252,N_2381);
xor U2437 (N_2437,N_2229,N_2235);
nand U2438 (N_2438,N_2270,N_2231);
nand U2439 (N_2439,N_2206,N_2211);
xnor U2440 (N_2440,N_2298,N_2377);
nand U2441 (N_2441,N_2385,N_2343);
nand U2442 (N_2442,N_2305,N_2348);
xor U2443 (N_2443,N_2317,N_2208);
or U2444 (N_2444,N_2334,N_2315);
nand U2445 (N_2445,N_2389,N_2222);
nor U2446 (N_2446,N_2362,N_2233);
or U2447 (N_2447,N_2354,N_2227);
or U2448 (N_2448,N_2267,N_2388);
nor U2449 (N_2449,N_2350,N_2369);
nand U2450 (N_2450,N_2358,N_2312);
or U2451 (N_2451,N_2203,N_2216);
and U2452 (N_2452,N_2328,N_2332);
or U2453 (N_2453,N_2224,N_2372);
nor U2454 (N_2454,N_2355,N_2230);
xnor U2455 (N_2455,N_2327,N_2269);
or U2456 (N_2456,N_2214,N_2337);
and U2457 (N_2457,N_2260,N_2399);
nor U2458 (N_2458,N_2202,N_2321);
or U2459 (N_2459,N_2387,N_2265);
nor U2460 (N_2460,N_2352,N_2368);
nor U2461 (N_2461,N_2272,N_2249);
xnor U2462 (N_2462,N_2301,N_2395);
nor U2463 (N_2463,N_2254,N_2283);
nor U2464 (N_2464,N_2378,N_2236);
nor U2465 (N_2465,N_2393,N_2293);
nand U2466 (N_2466,N_2326,N_2248);
nor U2467 (N_2467,N_2311,N_2299);
nor U2468 (N_2468,N_2363,N_2391);
or U2469 (N_2469,N_2347,N_2205);
and U2470 (N_2470,N_2318,N_2316);
nor U2471 (N_2471,N_2286,N_2259);
and U2472 (N_2472,N_2390,N_2207);
nand U2473 (N_2473,N_2212,N_2292);
nor U2474 (N_2474,N_2261,N_2373);
xor U2475 (N_2475,N_2263,N_2320);
nor U2476 (N_2476,N_2228,N_2277);
nor U2477 (N_2477,N_2306,N_2383);
xnor U2478 (N_2478,N_2382,N_2336);
nor U2479 (N_2479,N_2371,N_2359);
and U2480 (N_2480,N_2302,N_2331);
nand U2481 (N_2481,N_2338,N_2341);
and U2482 (N_2482,N_2250,N_2247);
or U2483 (N_2483,N_2319,N_2215);
nor U2484 (N_2484,N_2324,N_2380);
or U2485 (N_2485,N_2323,N_2268);
or U2486 (N_2486,N_2314,N_2271);
nand U2487 (N_2487,N_2384,N_2217);
or U2488 (N_2488,N_2333,N_2357);
and U2489 (N_2489,N_2273,N_2360);
or U2490 (N_2490,N_2234,N_2365);
nor U2491 (N_2491,N_2209,N_2335);
nor U2492 (N_2492,N_2245,N_2290);
and U2493 (N_2493,N_2226,N_2351);
nand U2494 (N_2494,N_2349,N_2375);
xor U2495 (N_2495,N_2297,N_2330);
or U2496 (N_2496,N_2313,N_2396);
or U2497 (N_2497,N_2367,N_2279);
nor U2498 (N_2498,N_2392,N_2237);
xor U2499 (N_2499,N_2398,N_2238);
or U2500 (N_2500,N_2235,N_2250);
or U2501 (N_2501,N_2213,N_2242);
nor U2502 (N_2502,N_2326,N_2383);
or U2503 (N_2503,N_2309,N_2273);
or U2504 (N_2504,N_2242,N_2201);
xnor U2505 (N_2505,N_2257,N_2262);
nor U2506 (N_2506,N_2311,N_2284);
xnor U2507 (N_2507,N_2270,N_2278);
nor U2508 (N_2508,N_2392,N_2210);
nor U2509 (N_2509,N_2305,N_2328);
nor U2510 (N_2510,N_2251,N_2216);
or U2511 (N_2511,N_2350,N_2363);
xnor U2512 (N_2512,N_2231,N_2338);
nand U2513 (N_2513,N_2395,N_2220);
or U2514 (N_2514,N_2348,N_2219);
or U2515 (N_2515,N_2362,N_2306);
nand U2516 (N_2516,N_2295,N_2238);
xor U2517 (N_2517,N_2334,N_2311);
xor U2518 (N_2518,N_2288,N_2204);
nor U2519 (N_2519,N_2262,N_2219);
xnor U2520 (N_2520,N_2210,N_2319);
and U2521 (N_2521,N_2394,N_2233);
xnor U2522 (N_2522,N_2259,N_2308);
or U2523 (N_2523,N_2281,N_2294);
and U2524 (N_2524,N_2322,N_2313);
nor U2525 (N_2525,N_2343,N_2316);
and U2526 (N_2526,N_2329,N_2285);
nor U2527 (N_2527,N_2268,N_2383);
nand U2528 (N_2528,N_2360,N_2376);
nor U2529 (N_2529,N_2340,N_2358);
and U2530 (N_2530,N_2217,N_2395);
nand U2531 (N_2531,N_2299,N_2208);
and U2532 (N_2532,N_2345,N_2378);
xnor U2533 (N_2533,N_2211,N_2245);
and U2534 (N_2534,N_2328,N_2397);
and U2535 (N_2535,N_2275,N_2216);
xor U2536 (N_2536,N_2290,N_2376);
and U2537 (N_2537,N_2287,N_2335);
nor U2538 (N_2538,N_2255,N_2241);
and U2539 (N_2539,N_2284,N_2218);
or U2540 (N_2540,N_2246,N_2284);
xor U2541 (N_2541,N_2268,N_2200);
xnor U2542 (N_2542,N_2269,N_2389);
nand U2543 (N_2543,N_2360,N_2257);
and U2544 (N_2544,N_2299,N_2291);
xnor U2545 (N_2545,N_2302,N_2334);
or U2546 (N_2546,N_2391,N_2305);
xor U2547 (N_2547,N_2298,N_2276);
xor U2548 (N_2548,N_2240,N_2231);
nor U2549 (N_2549,N_2331,N_2260);
nand U2550 (N_2550,N_2255,N_2291);
xnor U2551 (N_2551,N_2398,N_2229);
or U2552 (N_2552,N_2255,N_2344);
nand U2553 (N_2553,N_2202,N_2216);
nand U2554 (N_2554,N_2280,N_2320);
xor U2555 (N_2555,N_2266,N_2265);
nor U2556 (N_2556,N_2337,N_2261);
or U2557 (N_2557,N_2217,N_2394);
and U2558 (N_2558,N_2353,N_2321);
and U2559 (N_2559,N_2380,N_2314);
or U2560 (N_2560,N_2329,N_2240);
or U2561 (N_2561,N_2295,N_2324);
xnor U2562 (N_2562,N_2239,N_2302);
xnor U2563 (N_2563,N_2215,N_2245);
nor U2564 (N_2564,N_2207,N_2258);
xnor U2565 (N_2565,N_2347,N_2203);
nand U2566 (N_2566,N_2282,N_2316);
or U2567 (N_2567,N_2248,N_2348);
xor U2568 (N_2568,N_2289,N_2371);
nand U2569 (N_2569,N_2334,N_2333);
and U2570 (N_2570,N_2215,N_2202);
xnor U2571 (N_2571,N_2263,N_2227);
nand U2572 (N_2572,N_2253,N_2213);
or U2573 (N_2573,N_2246,N_2359);
or U2574 (N_2574,N_2267,N_2375);
or U2575 (N_2575,N_2329,N_2226);
nor U2576 (N_2576,N_2281,N_2346);
nand U2577 (N_2577,N_2351,N_2289);
xnor U2578 (N_2578,N_2221,N_2279);
and U2579 (N_2579,N_2260,N_2207);
or U2580 (N_2580,N_2283,N_2378);
nand U2581 (N_2581,N_2301,N_2265);
xor U2582 (N_2582,N_2384,N_2344);
nor U2583 (N_2583,N_2328,N_2247);
nor U2584 (N_2584,N_2374,N_2312);
xnor U2585 (N_2585,N_2306,N_2231);
or U2586 (N_2586,N_2208,N_2372);
nor U2587 (N_2587,N_2377,N_2385);
and U2588 (N_2588,N_2222,N_2234);
and U2589 (N_2589,N_2229,N_2237);
and U2590 (N_2590,N_2228,N_2342);
and U2591 (N_2591,N_2284,N_2389);
nor U2592 (N_2592,N_2378,N_2273);
nand U2593 (N_2593,N_2235,N_2219);
nand U2594 (N_2594,N_2360,N_2220);
or U2595 (N_2595,N_2394,N_2241);
xor U2596 (N_2596,N_2338,N_2297);
nand U2597 (N_2597,N_2272,N_2242);
or U2598 (N_2598,N_2350,N_2323);
or U2599 (N_2599,N_2330,N_2371);
or U2600 (N_2600,N_2555,N_2486);
and U2601 (N_2601,N_2409,N_2509);
or U2602 (N_2602,N_2417,N_2469);
and U2603 (N_2603,N_2551,N_2490);
xnor U2604 (N_2604,N_2597,N_2405);
nand U2605 (N_2605,N_2543,N_2418);
xnor U2606 (N_2606,N_2514,N_2493);
xor U2607 (N_2607,N_2477,N_2431);
xnor U2608 (N_2608,N_2588,N_2488);
or U2609 (N_2609,N_2408,N_2422);
nor U2610 (N_2610,N_2519,N_2424);
xor U2611 (N_2611,N_2532,N_2578);
nor U2612 (N_2612,N_2451,N_2448);
or U2613 (N_2613,N_2446,N_2492);
nand U2614 (N_2614,N_2536,N_2548);
xnor U2615 (N_2615,N_2564,N_2458);
nor U2616 (N_2616,N_2423,N_2464);
nand U2617 (N_2617,N_2554,N_2472);
and U2618 (N_2618,N_2414,N_2452);
and U2619 (N_2619,N_2552,N_2589);
xnor U2620 (N_2620,N_2593,N_2474);
or U2621 (N_2621,N_2419,N_2599);
nand U2622 (N_2622,N_2429,N_2416);
xnor U2623 (N_2623,N_2504,N_2468);
nor U2624 (N_2624,N_2583,N_2459);
nand U2625 (N_2625,N_2497,N_2539);
and U2626 (N_2626,N_2595,N_2523);
or U2627 (N_2627,N_2455,N_2527);
nand U2628 (N_2628,N_2515,N_2473);
and U2629 (N_2629,N_2550,N_2565);
nand U2630 (N_2630,N_2412,N_2450);
or U2631 (N_2631,N_2436,N_2503);
and U2632 (N_2632,N_2498,N_2547);
nor U2633 (N_2633,N_2462,N_2502);
or U2634 (N_2634,N_2542,N_2584);
nor U2635 (N_2635,N_2563,N_2401);
nor U2636 (N_2636,N_2546,N_2513);
nand U2637 (N_2637,N_2591,N_2495);
or U2638 (N_2638,N_2454,N_2561);
xnor U2639 (N_2639,N_2425,N_2580);
or U2640 (N_2640,N_2471,N_2537);
xor U2641 (N_2641,N_2512,N_2475);
nand U2642 (N_2642,N_2438,N_2559);
and U2643 (N_2643,N_2541,N_2587);
xor U2644 (N_2644,N_2510,N_2480);
nor U2645 (N_2645,N_2406,N_2421);
xor U2646 (N_2646,N_2441,N_2444);
and U2647 (N_2647,N_2501,N_2427);
nor U2648 (N_2648,N_2411,N_2534);
or U2649 (N_2649,N_2579,N_2439);
nor U2650 (N_2650,N_2598,N_2483);
and U2651 (N_2651,N_2413,N_2590);
or U2652 (N_2652,N_2531,N_2538);
and U2653 (N_2653,N_2573,N_2567);
or U2654 (N_2654,N_2432,N_2505);
nor U2655 (N_2655,N_2434,N_2463);
and U2656 (N_2656,N_2467,N_2585);
xor U2657 (N_2657,N_2568,N_2443);
and U2658 (N_2658,N_2465,N_2592);
nand U2659 (N_2659,N_2478,N_2571);
nand U2660 (N_2660,N_2521,N_2400);
nand U2661 (N_2661,N_2572,N_2506);
xor U2662 (N_2662,N_2576,N_2440);
nor U2663 (N_2663,N_2586,N_2524);
xnor U2664 (N_2664,N_2508,N_2403);
or U2665 (N_2665,N_2499,N_2470);
nand U2666 (N_2666,N_2535,N_2447);
or U2667 (N_2667,N_2544,N_2420);
nand U2668 (N_2668,N_2496,N_2453);
or U2669 (N_2669,N_2553,N_2560);
and U2670 (N_2670,N_2569,N_2460);
and U2671 (N_2671,N_2556,N_2402);
or U2672 (N_2672,N_2575,N_2482);
nand U2673 (N_2673,N_2549,N_2407);
or U2674 (N_2674,N_2442,N_2461);
xor U2675 (N_2675,N_2433,N_2529);
nor U2676 (N_2676,N_2530,N_2511);
and U2677 (N_2677,N_2570,N_2518);
nor U2678 (N_2678,N_2540,N_2494);
or U2679 (N_2679,N_2526,N_2557);
or U2680 (N_2680,N_2581,N_2404);
nor U2681 (N_2681,N_2479,N_2566);
and U2682 (N_2682,N_2430,N_2415);
or U2683 (N_2683,N_2476,N_2426);
or U2684 (N_2684,N_2574,N_2485);
nand U2685 (N_2685,N_2487,N_2445);
or U2686 (N_2686,N_2517,N_2466);
and U2687 (N_2687,N_2507,N_2562);
nor U2688 (N_2688,N_2533,N_2500);
xnor U2689 (N_2689,N_2449,N_2484);
and U2690 (N_2690,N_2577,N_2528);
or U2691 (N_2691,N_2516,N_2558);
nand U2692 (N_2692,N_2437,N_2435);
nor U2693 (N_2693,N_2545,N_2520);
and U2694 (N_2694,N_2428,N_2582);
nor U2695 (N_2695,N_2489,N_2481);
xnor U2696 (N_2696,N_2491,N_2522);
or U2697 (N_2697,N_2410,N_2525);
nor U2698 (N_2698,N_2457,N_2456);
and U2699 (N_2699,N_2596,N_2594);
and U2700 (N_2700,N_2598,N_2506);
and U2701 (N_2701,N_2553,N_2528);
or U2702 (N_2702,N_2507,N_2584);
and U2703 (N_2703,N_2542,N_2578);
nor U2704 (N_2704,N_2501,N_2471);
nor U2705 (N_2705,N_2568,N_2427);
nor U2706 (N_2706,N_2563,N_2556);
and U2707 (N_2707,N_2544,N_2403);
nand U2708 (N_2708,N_2425,N_2443);
xnor U2709 (N_2709,N_2590,N_2472);
nand U2710 (N_2710,N_2439,N_2440);
nand U2711 (N_2711,N_2533,N_2597);
and U2712 (N_2712,N_2532,N_2486);
nand U2713 (N_2713,N_2416,N_2468);
xnor U2714 (N_2714,N_2581,N_2577);
or U2715 (N_2715,N_2599,N_2441);
or U2716 (N_2716,N_2449,N_2468);
and U2717 (N_2717,N_2463,N_2487);
or U2718 (N_2718,N_2499,N_2502);
xnor U2719 (N_2719,N_2437,N_2555);
xnor U2720 (N_2720,N_2418,N_2439);
nor U2721 (N_2721,N_2441,N_2478);
xor U2722 (N_2722,N_2572,N_2461);
nand U2723 (N_2723,N_2516,N_2585);
and U2724 (N_2724,N_2485,N_2430);
nand U2725 (N_2725,N_2470,N_2548);
nand U2726 (N_2726,N_2574,N_2591);
nor U2727 (N_2727,N_2497,N_2413);
nand U2728 (N_2728,N_2466,N_2545);
nor U2729 (N_2729,N_2562,N_2506);
xor U2730 (N_2730,N_2449,N_2530);
or U2731 (N_2731,N_2592,N_2439);
nand U2732 (N_2732,N_2413,N_2430);
and U2733 (N_2733,N_2537,N_2556);
or U2734 (N_2734,N_2464,N_2453);
or U2735 (N_2735,N_2432,N_2497);
or U2736 (N_2736,N_2420,N_2497);
xor U2737 (N_2737,N_2544,N_2570);
or U2738 (N_2738,N_2442,N_2559);
nand U2739 (N_2739,N_2401,N_2482);
xnor U2740 (N_2740,N_2451,N_2574);
or U2741 (N_2741,N_2417,N_2459);
xor U2742 (N_2742,N_2591,N_2496);
or U2743 (N_2743,N_2426,N_2436);
nand U2744 (N_2744,N_2546,N_2405);
nor U2745 (N_2745,N_2434,N_2408);
or U2746 (N_2746,N_2417,N_2539);
nor U2747 (N_2747,N_2434,N_2538);
and U2748 (N_2748,N_2537,N_2451);
or U2749 (N_2749,N_2478,N_2554);
or U2750 (N_2750,N_2506,N_2411);
or U2751 (N_2751,N_2578,N_2479);
nand U2752 (N_2752,N_2414,N_2544);
nor U2753 (N_2753,N_2585,N_2430);
xor U2754 (N_2754,N_2428,N_2536);
nand U2755 (N_2755,N_2460,N_2410);
nand U2756 (N_2756,N_2532,N_2422);
xnor U2757 (N_2757,N_2473,N_2552);
nand U2758 (N_2758,N_2518,N_2559);
and U2759 (N_2759,N_2586,N_2435);
xor U2760 (N_2760,N_2567,N_2475);
xnor U2761 (N_2761,N_2575,N_2473);
or U2762 (N_2762,N_2531,N_2499);
nand U2763 (N_2763,N_2443,N_2456);
nand U2764 (N_2764,N_2411,N_2404);
and U2765 (N_2765,N_2506,N_2494);
xnor U2766 (N_2766,N_2514,N_2499);
nor U2767 (N_2767,N_2490,N_2419);
xor U2768 (N_2768,N_2471,N_2587);
nor U2769 (N_2769,N_2521,N_2407);
nor U2770 (N_2770,N_2535,N_2574);
xnor U2771 (N_2771,N_2408,N_2449);
nor U2772 (N_2772,N_2432,N_2592);
nor U2773 (N_2773,N_2468,N_2458);
and U2774 (N_2774,N_2441,N_2481);
nor U2775 (N_2775,N_2514,N_2418);
or U2776 (N_2776,N_2499,N_2591);
nor U2777 (N_2777,N_2479,N_2431);
nand U2778 (N_2778,N_2584,N_2402);
or U2779 (N_2779,N_2513,N_2578);
nor U2780 (N_2780,N_2506,N_2553);
xor U2781 (N_2781,N_2582,N_2491);
xor U2782 (N_2782,N_2448,N_2575);
nand U2783 (N_2783,N_2555,N_2592);
or U2784 (N_2784,N_2473,N_2457);
nand U2785 (N_2785,N_2429,N_2575);
xnor U2786 (N_2786,N_2462,N_2450);
nor U2787 (N_2787,N_2491,N_2450);
or U2788 (N_2788,N_2587,N_2523);
xnor U2789 (N_2789,N_2448,N_2438);
or U2790 (N_2790,N_2562,N_2587);
nand U2791 (N_2791,N_2539,N_2529);
or U2792 (N_2792,N_2499,N_2586);
and U2793 (N_2793,N_2460,N_2404);
and U2794 (N_2794,N_2534,N_2457);
nor U2795 (N_2795,N_2453,N_2471);
nand U2796 (N_2796,N_2402,N_2410);
xor U2797 (N_2797,N_2559,N_2496);
xnor U2798 (N_2798,N_2510,N_2458);
xnor U2799 (N_2799,N_2470,N_2430);
and U2800 (N_2800,N_2602,N_2798);
and U2801 (N_2801,N_2634,N_2614);
xnor U2802 (N_2802,N_2727,N_2760);
nand U2803 (N_2803,N_2646,N_2768);
or U2804 (N_2804,N_2712,N_2678);
nand U2805 (N_2805,N_2746,N_2615);
or U2806 (N_2806,N_2639,N_2669);
nand U2807 (N_2807,N_2717,N_2604);
nand U2808 (N_2808,N_2790,N_2704);
or U2809 (N_2809,N_2780,N_2605);
nand U2810 (N_2810,N_2799,N_2774);
or U2811 (N_2811,N_2680,N_2733);
nor U2812 (N_2812,N_2784,N_2688);
or U2813 (N_2813,N_2761,N_2679);
and U2814 (N_2814,N_2729,N_2611);
xor U2815 (N_2815,N_2792,N_2745);
or U2816 (N_2816,N_2601,N_2707);
nor U2817 (N_2817,N_2762,N_2734);
xor U2818 (N_2818,N_2748,N_2642);
nand U2819 (N_2819,N_2624,N_2721);
and U2820 (N_2820,N_2657,N_2663);
nand U2821 (N_2821,N_2718,N_2786);
nor U2822 (N_2822,N_2626,N_2695);
xor U2823 (N_2823,N_2608,N_2728);
nand U2824 (N_2824,N_2747,N_2777);
and U2825 (N_2825,N_2703,N_2710);
nand U2826 (N_2826,N_2654,N_2765);
or U2827 (N_2827,N_2606,N_2672);
nand U2828 (N_2828,N_2737,N_2755);
nand U2829 (N_2829,N_2648,N_2693);
nor U2830 (N_2830,N_2714,N_2656);
nor U2831 (N_2831,N_2686,N_2667);
xor U2832 (N_2832,N_2711,N_2740);
xor U2833 (N_2833,N_2771,N_2676);
nor U2834 (N_2834,N_2732,N_2702);
nor U2835 (N_2835,N_2754,N_2730);
nor U2836 (N_2836,N_2757,N_2769);
xor U2837 (N_2837,N_2795,N_2778);
or U2838 (N_2838,N_2675,N_2785);
xnor U2839 (N_2839,N_2649,N_2724);
or U2840 (N_2840,N_2751,N_2715);
and U2841 (N_2841,N_2622,N_2677);
xor U2842 (N_2842,N_2632,N_2643);
and U2843 (N_2843,N_2600,N_2690);
nand U2844 (N_2844,N_2696,N_2618);
and U2845 (N_2845,N_2650,N_2770);
nand U2846 (N_2846,N_2674,N_2658);
or U2847 (N_2847,N_2779,N_2759);
nor U2848 (N_2848,N_2743,N_2753);
xnor U2849 (N_2849,N_2756,N_2640);
and U2850 (N_2850,N_2735,N_2694);
nand U2851 (N_2851,N_2668,N_2700);
and U2852 (N_2852,N_2791,N_2662);
nand U2853 (N_2853,N_2665,N_2691);
or U2854 (N_2854,N_2797,N_2713);
xor U2855 (N_2855,N_2758,N_2738);
nand U2856 (N_2856,N_2722,N_2775);
or U2857 (N_2857,N_2630,N_2720);
xor U2858 (N_2858,N_2772,N_2788);
and U2859 (N_2859,N_2623,N_2763);
xnor U2860 (N_2860,N_2682,N_2766);
and U2861 (N_2861,N_2628,N_2612);
and U2862 (N_2862,N_2636,N_2645);
and U2863 (N_2863,N_2699,N_2776);
nand U2864 (N_2864,N_2641,N_2767);
nor U2865 (N_2865,N_2644,N_2789);
xnor U2866 (N_2866,N_2603,N_2671);
and U2867 (N_2867,N_2698,N_2683);
nor U2868 (N_2868,N_2681,N_2664);
or U2869 (N_2869,N_2726,N_2651);
nand U2870 (N_2870,N_2706,N_2773);
nand U2871 (N_2871,N_2782,N_2744);
nand U2872 (N_2872,N_2647,N_2692);
or U2873 (N_2873,N_2617,N_2652);
nor U2874 (N_2874,N_2749,N_2625);
and U2875 (N_2875,N_2627,N_2689);
nand U2876 (N_2876,N_2701,N_2633);
nand U2877 (N_2877,N_2736,N_2609);
nand U2878 (N_2878,N_2666,N_2607);
and U2879 (N_2879,N_2739,N_2719);
xnor U2880 (N_2880,N_2629,N_2741);
xnor U2881 (N_2881,N_2742,N_2635);
nor U2882 (N_2882,N_2638,N_2670);
nor U2883 (N_2883,N_2610,N_2794);
and U2884 (N_2884,N_2659,N_2716);
or U2885 (N_2885,N_2685,N_2616);
nand U2886 (N_2886,N_2783,N_2731);
nor U2887 (N_2887,N_2621,N_2684);
or U2888 (N_2888,N_2655,N_2673);
or U2889 (N_2889,N_2637,N_2752);
xor U2890 (N_2890,N_2781,N_2687);
nor U2891 (N_2891,N_2697,N_2660);
xor U2892 (N_2892,N_2631,N_2750);
or U2893 (N_2893,N_2661,N_2764);
and U2894 (N_2894,N_2793,N_2723);
or U2895 (N_2895,N_2709,N_2620);
or U2896 (N_2896,N_2653,N_2787);
nand U2897 (N_2897,N_2796,N_2725);
xor U2898 (N_2898,N_2613,N_2619);
or U2899 (N_2899,N_2708,N_2705);
xor U2900 (N_2900,N_2622,N_2726);
xnor U2901 (N_2901,N_2653,N_2632);
xnor U2902 (N_2902,N_2744,N_2749);
and U2903 (N_2903,N_2741,N_2699);
nand U2904 (N_2904,N_2790,N_2736);
and U2905 (N_2905,N_2604,N_2738);
xor U2906 (N_2906,N_2694,N_2766);
nor U2907 (N_2907,N_2766,N_2634);
or U2908 (N_2908,N_2672,N_2602);
or U2909 (N_2909,N_2603,N_2771);
nand U2910 (N_2910,N_2639,N_2687);
xor U2911 (N_2911,N_2709,N_2671);
or U2912 (N_2912,N_2679,N_2734);
nor U2913 (N_2913,N_2606,N_2671);
and U2914 (N_2914,N_2755,N_2730);
or U2915 (N_2915,N_2611,N_2683);
nor U2916 (N_2916,N_2632,N_2639);
or U2917 (N_2917,N_2664,N_2608);
or U2918 (N_2918,N_2714,N_2796);
xnor U2919 (N_2919,N_2630,N_2665);
nor U2920 (N_2920,N_2646,N_2627);
nor U2921 (N_2921,N_2730,N_2684);
and U2922 (N_2922,N_2753,N_2655);
nand U2923 (N_2923,N_2649,N_2607);
or U2924 (N_2924,N_2646,N_2645);
or U2925 (N_2925,N_2608,N_2717);
xnor U2926 (N_2926,N_2665,N_2716);
xnor U2927 (N_2927,N_2679,N_2793);
or U2928 (N_2928,N_2617,N_2784);
or U2929 (N_2929,N_2631,N_2653);
xor U2930 (N_2930,N_2652,N_2724);
and U2931 (N_2931,N_2623,N_2688);
xor U2932 (N_2932,N_2796,N_2606);
or U2933 (N_2933,N_2724,N_2610);
and U2934 (N_2934,N_2782,N_2724);
xnor U2935 (N_2935,N_2786,N_2614);
nor U2936 (N_2936,N_2731,N_2661);
nor U2937 (N_2937,N_2789,N_2648);
nor U2938 (N_2938,N_2625,N_2796);
nand U2939 (N_2939,N_2769,N_2645);
and U2940 (N_2940,N_2606,N_2649);
or U2941 (N_2941,N_2751,N_2740);
nand U2942 (N_2942,N_2738,N_2782);
or U2943 (N_2943,N_2627,N_2622);
nor U2944 (N_2944,N_2735,N_2737);
and U2945 (N_2945,N_2799,N_2601);
xor U2946 (N_2946,N_2729,N_2646);
xnor U2947 (N_2947,N_2626,N_2670);
nand U2948 (N_2948,N_2764,N_2753);
nand U2949 (N_2949,N_2643,N_2748);
nand U2950 (N_2950,N_2797,N_2755);
xnor U2951 (N_2951,N_2783,N_2637);
xnor U2952 (N_2952,N_2628,N_2746);
nand U2953 (N_2953,N_2604,N_2628);
and U2954 (N_2954,N_2665,N_2768);
nor U2955 (N_2955,N_2673,N_2725);
nand U2956 (N_2956,N_2752,N_2681);
and U2957 (N_2957,N_2604,N_2781);
or U2958 (N_2958,N_2708,N_2619);
and U2959 (N_2959,N_2773,N_2638);
nand U2960 (N_2960,N_2694,N_2740);
xnor U2961 (N_2961,N_2694,N_2789);
nand U2962 (N_2962,N_2788,N_2695);
and U2963 (N_2963,N_2731,N_2626);
nand U2964 (N_2964,N_2686,N_2796);
or U2965 (N_2965,N_2734,N_2745);
or U2966 (N_2966,N_2632,N_2774);
nand U2967 (N_2967,N_2740,N_2656);
nand U2968 (N_2968,N_2677,N_2631);
xnor U2969 (N_2969,N_2749,N_2781);
nand U2970 (N_2970,N_2738,N_2611);
nand U2971 (N_2971,N_2770,N_2689);
xnor U2972 (N_2972,N_2767,N_2680);
nor U2973 (N_2973,N_2773,N_2612);
nand U2974 (N_2974,N_2793,N_2786);
xor U2975 (N_2975,N_2745,N_2654);
or U2976 (N_2976,N_2603,N_2752);
nor U2977 (N_2977,N_2622,N_2637);
and U2978 (N_2978,N_2749,N_2754);
and U2979 (N_2979,N_2724,N_2798);
xor U2980 (N_2980,N_2756,N_2773);
or U2981 (N_2981,N_2641,N_2754);
or U2982 (N_2982,N_2703,N_2708);
or U2983 (N_2983,N_2644,N_2735);
and U2984 (N_2984,N_2629,N_2758);
nand U2985 (N_2985,N_2790,N_2664);
nor U2986 (N_2986,N_2757,N_2616);
nand U2987 (N_2987,N_2689,N_2662);
xnor U2988 (N_2988,N_2624,N_2687);
xnor U2989 (N_2989,N_2689,N_2730);
nand U2990 (N_2990,N_2688,N_2618);
nor U2991 (N_2991,N_2733,N_2650);
or U2992 (N_2992,N_2609,N_2697);
and U2993 (N_2993,N_2607,N_2672);
and U2994 (N_2994,N_2711,N_2607);
nor U2995 (N_2995,N_2677,N_2789);
nor U2996 (N_2996,N_2717,N_2633);
nor U2997 (N_2997,N_2699,N_2665);
and U2998 (N_2998,N_2753,N_2653);
xnor U2999 (N_2999,N_2689,N_2761);
xor U3000 (N_3000,N_2870,N_2990);
nor U3001 (N_3001,N_2921,N_2895);
xor U3002 (N_3002,N_2855,N_2953);
or U3003 (N_3003,N_2962,N_2801);
and U3004 (N_3004,N_2919,N_2971);
or U3005 (N_3005,N_2903,N_2922);
xnor U3006 (N_3006,N_2970,N_2917);
or U3007 (N_3007,N_2829,N_2897);
or U3008 (N_3008,N_2983,N_2908);
xor U3009 (N_3009,N_2934,N_2861);
nor U3010 (N_3010,N_2816,N_2853);
nor U3011 (N_3011,N_2849,N_2914);
xnor U3012 (N_3012,N_2927,N_2891);
or U3013 (N_3013,N_2833,N_2982);
xor U3014 (N_3014,N_2856,N_2898);
xor U3015 (N_3015,N_2862,N_2832);
and U3016 (N_3016,N_2810,N_2872);
and U3017 (N_3017,N_2991,N_2915);
xnor U3018 (N_3018,N_2886,N_2893);
or U3019 (N_3019,N_2865,N_2941);
nand U3020 (N_3020,N_2975,N_2819);
or U3021 (N_3021,N_2884,N_2815);
xnor U3022 (N_3022,N_2844,N_2987);
and U3023 (N_3023,N_2916,N_2882);
nand U3024 (N_3024,N_2986,N_2948);
and U3025 (N_3025,N_2998,N_2878);
nor U3026 (N_3026,N_2912,N_2969);
xnor U3027 (N_3027,N_2952,N_2894);
or U3028 (N_3028,N_2814,N_2946);
xnor U3029 (N_3029,N_2824,N_2845);
xor U3030 (N_3030,N_2977,N_2993);
or U3031 (N_3031,N_2812,N_2978);
or U3032 (N_3032,N_2883,N_2847);
or U3033 (N_3033,N_2939,N_2877);
xor U3034 (N_3034,N_2825,N_2803);
nand U3035 (N_3035,N_2944,N_2858);
or U3036 (N_3036,N_2863,N_2857);
nor U3037 (N_3037,N_2918,N_2822);
xnor U3038 (N_3038,N_2959,N_2956);
xnor U3039 (N_3039,N_2938,N_2836);
xnor U3040 (N_3040,N_2820,N_2831);
xnor U3041 (N_3041,N_2997,N_2867);
and U3042 (N_3042,N_2967,N_2830);
xor U3043 (N_3043,N_2900,N_2910);
or U3044 (N_3044,N_2935,N_2926);
nand U3045 (N_3045,N_2839,N_2920);
nor U3046 (N_3046,N_2907,N_2923);
nor U3047 (N_3047,N_2851,N_2880);
and U3048 (N_3048,N_2841,N_2995);
nor U3049 (N_3049,N_2838,N_2901);
and U3050 (N_3050,N_2864,N_2823);
xor U3051 (N_3051,N_2818,N_2848);
nor U3052 (N_3052,N_2888,N_2874);
or U3053 (N_3053,N_2988,N_2945);
xor U3054 (N_3054,N_2964,N_2984);
xnor U3055 (N_3055,N_2968,N_2890);
or U3056 (N_3056,N_2972,N_2854);
and U3057 (N_3057,N_2868,N_2911);
nor U3058 (N_3058,N_2965,N_2846);
and U3059 (N_3059,N_2979,N_2899);
and U3060 (N_3060,N_2954,N_2802);
and U3061 (N_3061,N_2813,N_2834);
nand U3062 (N_3062,N_2892,N_2992);
or U3063 (N_3063,N_2980,N_2936);
and U3064 (N_3064,N_2973,N_2902);
nand U3065 (N_3065,N_2860,N_2835);
nand U3066 (N_3066,N_2960,N_2976);
xor U3067 (N_3067,N_2828,N_2974);
xor U3068 (N_3068,N_2885,N_2871);
or U3069 (N_3069,N_2994,N_2817);
nand U3070 (N_3070,N_2806,N_2940);
and U3071 (N_3071,N_2924,N_2951);
xor U3072 (N_3072,N_2807,N_2932);
xor U3073 (N_3073,N_2805,N_2942);
or U3074 (N_3074,N_2840,N_2881);
nor U3075 (N_3075,N_2947,N_2985);
or U3076 (N_3076,N_2852,N_2906);
or U3077 (N_3077,N_2955,N_2875);
nand U3078 (N_3078,N_2957,N_2937);
xnor U3079 (N_3079,N_2804,N_2961);
xor U3080 (N_3080,N_2981,N_2925);
and U3081 (N_3081,N_2966,N_2905);
nor U3082 (N_3082,N_2887,N_2896);
or U3083 (N_3083,N_2930,N_2928);
and U3084 (N_3084,N_2879,N_2933);
nand U3085 (N_3085,N_2821,N_2811);
xor U3086 (N_3086,N_2949,N_2873);
nand U3087 (N_3087,N_2842,N_2889);
nor U3088 (N_3088,N_2989,N_2904);
nor U3089 (N_3089,N_2943,N_2963);
nand U3090 (N_3090,N_2843,N_2950);
nor U3091 (N_3091,N_2808,N_2929);
nand U3092 (N_3092,N_2859,N_2931);
nand U3093 (N_3093,N_2850,N_2826);
nand U3094 (N_3094,N_2996,N_2999);
xnor U3095 (N_3095,N_2866,N_2909);
and U3096 (N_3096,N_2869,N_2827);
xor U3097 (N_3097,N_2809,N_2913);
nor U3098 (N_3098,N_2800,N_2837);
xor U3099 (N_3099,N_2958,N_2876);
nand U3100 (N_3100,N_2944,N_2989);
nor U3101 (N_3101,N_2823,N_2989);
and U3102 (N_3102,N_2838,N_2849);
xnor U3103 (N_3103,N_2973,N_2908);
xor U3104 (N_3104,N_2836,N_2829);
and U3105 (N_3105,N_2833,N_2929);
or U3106 (N_3106,N_2819,N_2933);
nand U3107 (N_3107,N_2917,N_2805);
nand U3108 (N_3108,N_2872,N_2859);
nand U3109 (N_3109,N_2943,N_2877);
nand U3110 (N_3110,N_2906,N_2935);
or U3111 (N_3111,N_2880,N_2945);
nand U3112 (N_3112,N_2934,N_2989);
nand U3113 (N_3113,N_2980,N_2834);
and U3114 (N_3114,N_2806,N_2801);
or U3115 (N_3115,N_2899,N_2818);
nand U3116 (N_3116,N_2922,N_2944);
or U3117 (N_3117,N_2862,N_2947);
xor U3118 (N_3118,N_2817,N_2822);
nor U3119 (N_3119,N_2812,N_2892);
or U3120 (N_3120,N_2950,N_2982);
and U3121 (N_3121,N_2867,N_2827);
or U3122 (N_3122,N_2805,N_2955);
nor U3123 (N_3123,N_2995,N_2851);
or U3124 (N_3124,N_2922,N_2998);
nor U3125 (N_3125,N_2876,N_2922);
nor U3126 (N_3126,N_2825,N_2912);
and U3127 (N_3127,N_2834,N_2977);
or U3128 (N_3128,N_2953,N_2988);
and U3129 (N_3129,N_2967,N_2981);
nand U3130 (N_3130,N_2940,N_2864);
and U3131 (N_3131,N_2853,N_2946);
nand U3132 (N_3132,N_2809,N_2937);
and U3133 (N_3133,N_2897,N_2833);
and U3134 (N_3134,N_2912,N_2967);
nand U3135 (N_3135,N_2979,N_2934);
xor U3136 (N_3136,N_2952,N_2958);
nand U3137 (N_3137,N_2901,N_2977);
or U3138 (N_3138,N_2870,N_2841);
nand U3139 (N_3139,N_2828,N_2843);
nor U3140 (N_3140,N_2834,N_2916);
and U3141 (N_3141,N_2849,N_2841);
or U3142 (N_3142,N_2819,N_2806);
or U3143 (N_3143,N_2993,N_2923);
xor U3144 (N_3144,N_2856,N_2996);
or U3145 (N_3145,N_2875,N_2897);
and U3146 (N_3146,N_2971,N_2922);
and U3147 (N_3147,N_2931,N_2996);
and U3148 (N_3148,N_2979,N_2996);
or U3149 (N_3149,N_2925,N_2874);
nor U3150 (N_3150,N_2837,N_2840);
and U3151 (N_3151,N_2966,N_2848);
or U3152 (N_3152,N_2869,N_2858);
xor U3153 (N_3153,N_2940,N_2881);
xnor U3154 (N_3154,N_2913,N_2807);
nor U3155 (N_3155,N_2931,N_2900);
or U3156 (N_3156,N_2823,N_2896);
nor U3157 (N_3157,N_2904,N_2826);
nand U3158 (N_3158,N_2992,N_2935);
and U3159 (N_3159,N_2921,N_2858);
xor U3160 (N_3160,N_2903,N_2888);
nand U3161 (N_3161,N_2980,N_2960);
nor U3162 (N_3162,N_2942,N_2990);
nor U3163 (N_3163,N_2832,N_2927);
xnor U3164 (N_3164,N_2832,N_2984);
nor U3165 (N_3165,N_2992,N_2870);
and U3166 (N_3166,N_2971,N_2867);
and U3167 (N_3167,N_2947,N_2946);
xor U3168 (N_3168,N_2869,N_2964);
nand U3169 (N_3169,N_2857,N_2934);
xnor U3170 (N_3170,N_2920,N_2960);
and U3171 (N_3171,N_2852,N_2970);
nor U3172 (N_3172,N_2846,N_2823);
or U3173 (N_3173,N_2984,N_2971);
nor U3174 (N_3174,N_2868,N_2881);
and U3175 (N_3175,N_2917,N_2929);
or U3176 (N_3176,N_2903,N_2822);
and U3177 (N_3177,N_2841,N_2969);
and U3178 (N_3178,N_2873,N_2909);
nand U3179 (N_3179,N_2837,N_2935);
nor U3180 (N_3180,N_2919,N_2800);
or U3181 (N_3181,N_2965,N_2934);
or U3182 (N_3182,N_2969,N_2809);
and U3183 (N_3183,N_2912,N_2896);
xnor U3184 (N_3184,N_2957,N_2939);
nand U3185 (N_3185,N_2996,N_2907);
xnor U3186 (N_3186,N_2909,N_2958);
xnor U3187 (N_3187,N_2818,N_2958);
nand U3188 (N_3188,N_2987,N_2913);
or U3189 (N_3189,N_2998,N_2891);
and U3190 (N_3190,N_2984,N_2858);
xnor U3191 (N_3191,N_2973,N_2959);
nor U3192 (N_3192,N_2800,N_2830);
and U3193 (N_3193,N_2987,N_2890);
or U3194 (N_3194,N_2974,N_2928);
nor U3195 (N_3195,N_2932,N_2995);
nand U3196 (N_3196,N_2970,N_2842);
or U3197 (N_3197,N_2887,N_2853);
nor U3198 (N_3198,N_2886,N_2963);
and U3199 (N_3199,N_2855,N_2984);
nand U3200 (N_3200,N_3100,N_3180);
or U3201 (N_3201,N_3175,N_3093);
and U3202 (N_3202,N_3131,N_3030);
xnor U3203 (N_3203,N_3060,N_3087);
or U3204 (N_3204,N_3125,N_3144);
nand U3205 (N_3205,N_3021,N_3011);
nand U3206 (N_3206,N_3171,N_3101);
nor U3207 (N_3207,N_3023,N_3188);
xor U3208 (N_3208,N_3183,N_3046);
and U3209 (N_3209,N_3031,N_3035);
xnor U3210 (N_3210,N_3070,N_3017);
xor U3211 (N_3211,N_3128,N_3120);
nor U3212 (N_3212,N_3064,N_3028);
xnor U3213 (N_3213,N_3066,N_3004);
nor U3214 (N_3214,N_3166,N_3049);
and U3215 (N_3215,N_3081,N_3122);
or U3216 (N_3216,N_3062,N_3147);
or U3217 (N_3217,N_3140,N_3037);
or U3218 (N_3218,N_3136,N_3138);
or U3219 (N_3219,N_3165,N_3098);
and U3220 (N_3220,N_3112,N_3095);
or U3221 (N_3221,N_3013,N_3045);
nand U3222 (N_3222,N_3126,N_3182);
nor U3223 (N_3223,N_3152,N_3111);
xor U3224 (N_3224,N_3186,N_3119);
nand U3225 (N_3225,N_3072,N_3056);
xnor U3226 (N_3226,N_3092,N_3083);
xor U3227 (N_3227,N_3099,N_3003);
and U3228 (N_3228,N_3157,N_3002);
and U3229 (N_3229,N_3041,N_3109);
or U3230 (N_3230,N_3074,N_3055);
and U3231 (N_3231,N_3127,N_3159);
or U3232 (N_3232,N_3061,N_3179);
nor U3233 (N_3233,N_3088,N_3016);
nor U3234 (N_3234,N_3156,N_3103);
nor U3235 (N_3235,N_3089,N_3130);
or U3236 (N_3236,N_3199,N_3008);
xor U3237 (N_3237,N_3192,N_3090);
and U3238 (N_3238,N_3150,N_3190);
nor U3239 (N_3239,N_3075,N_3038);
nor U3240 (N_3240,N_3094,N_3177);
nand U3241 (N_3241,N_3198,N_3184);
xnor U3242 (N_3242,N_3104,N_3151);
and U3243 (N_3243,N_3012,N_3033);
and U3244 (N_3244,N_3197,N_3052);
nor U3245 (N_3245,N_3153,N_3086);
nor U3246 (N_3246,N_3148,N_3113);
or U3247 (N_3247,N_3071,N_3169);
or U3248 (N_3248,N_3118,N_3080);
or U3249 (N_3249,N_3133,N_3024);
or U3250 (N_3250,N_3026,N_3007);
nor U3251 (N_3251,N_3196,N_3123);
xor U3252 (N_3252,N_3173,N_3077);
and U3253 (N_3253,N_3051,N_3027);
xnor U3254 (N_3254,N_3163,N_3142);
nor U3255 (N_3255,N_3124,N_3115);
and U3256 (N_3256,N_3000,N_3063);
nand U3257 (N_3257,N_3161,N_3143);
xnor U3258 (N_3258,N_3058,N_3069);
nor U3259 (N_3259,N_3191,N_3110);
or U3260 (N_3260,N_3195,N_3034);
and U3261 (N_3261,N_3187,N_3057);
or U3262 (N_3262,N_3139,N_3121);
nor U3263 (N_3263,N_3054,N_3048);
or U3264 (N_3264,N_3149,N_3076);
or U3265 (N_3265,N_3167,N_3014);
and U3266 (N_3266,N_3042,N_3006);
and U3267 (N_3267,N_3059,N_3025);
xor U3268 (N_3268,N_3162,N_3039);
or U3269 (N_3269,N_3194,N_3085);
nand U3270 (N_3270,N_3178,N_3044);
and U3271 (N_3271,N_3102,N_3068);
nand U3272 (N_3272,N_3107,N_3155);
xnor U3273 (N_3273,N_3091,N_3082);
and U3274 (N_3274,N_3174,N_3032);
nand U3275 (N_3275,N_3116,N_3015);
and U3276 (N_3276,N_3073,N_3129);
xnor U3277 (N_3277,N_3065,N_3160);
or U3278 (N_3278,N_3067,N_3135);
xor U3279 (N_3279,N_3043,N_3108);
nand U3280 (N_3280,N_3009,N_3010);
nand U3281 (N_3281,N_3097,N_3117);
or U3282 (N_3282,N_3145,N_3020);
nand U3283 (N_3283,N_3170,N_3079);
and U3284 (N_3284,N_3132,N_3105);
nor U3285 (N_3285,N_3001,N_3029);
nor U3286 (N_3286,N_3078,N_3158);
xor U3287 (N_3287,N_3168,N_3154);
nand U3288 (N_3288,N_3084,N_3053);
nor U3289 (N_3289,N_3096,N_3172);
xor U3290 (N_3290,N_3047,N_3185);
xnor U3291 (N_3291,N_3106,N_3040);
or U3292 (N_3292,N_3005,N_3134);
nand U3293 (N_3293,N_3164,N_3193);
or U3294 (N_3294,N_3022,N_3146);
or U3295 (N_3295,N_3189,N_3036);
nor U3296 (N_3296,N_3181,N_3141);
nor U3297 (N_3297,N_3019,N_3050);
nor U3298 (N_3298,N_3114,N_3018);
or U3299 (N_3299,N_3137,N_3176);
nor U3300 (N_3300,N_3151,N_3081);
and U3301 (N_3301,N_3106,N_3188);
nand U3302 (N_3302,N_3131,N_3005);
nand U3303 (N_3303,N_3009,N_3039);
nor U3304 (N_3304,N_3037,N_3093);
nand U3305 (N_3305,N_3070,N_3199);
or U3306 (N_3306,N_3084,N_3192);
nand U3307 (N_3307,N_3141,N_3043);
or U3308 (N_3308,N_3018,N_3130);
nand U3309 (N_3309,N_3031,N_3064);
xor U3310 (N_3310,N_3116,N_3016);
nor U3311 (N_3311,N_3197,N_3107);
and U3312 (N_3312,N_3130,N_3198);
and U3313 (N_3313,N_3100,N_3150);
nand U3314 (N_3314,N_3146,N_3007);
nand U3315 (N_3315,N_3002,N_3188);
and U3316 (N_3316,N_3022,N_3145);
and U3317 (N_3317,N_3011,N_3130);
nand U3318 (N_3318,N_3143,N_3042);
xnor U3319 (N_3319,N_3007,N_3122);
and U3320 (N_3320,N_3104,N_3035);
or U3321 (N_3321,N_3099,N_3199);
nand U3322 (N_3322,N_3095,N_3002);
nand U3323 (N_3323,N_3139,N_3074);
nand U3324 (N_3324,N_3169,N_3027);
xnor U3325 (N_3325,N_3037,N_3105);
nor U3326 (N_3326,N_3199,N_3040);
xor U3327 (N_3327,N_3033,N_3047);
nor U3328 (N_3328,N_3039,N_3062);
xor U3329 (N_3329,N_3081,N_3168);
or U3330 (N_3330,N_3146,N_3074);
or U3331 (N_3331,N_3076,N_3137);
and U3332 (N_3332,N_3160,N_3078);
nand U3333 (N_3333,N_3092,N_3198);
or U3334 (N_3334,N_3172,N_3063);
xor U3335 (N_3335,N_3186,N_3016);
and U3336 (N_3336,N_3005,N_3062);
nor U3337 (N_3337,N_3046,N_3180);
nand U3338 (N_3338,N_3003,N_3189);
nand U3339 (N_3339,N_3115,N_3149);
nor U3340 (N_3340,N_3123,N_3091);
nor U3341 (N_3341,N_3188,N_3060);
xnor U3342 (N_3342,N_3030,N_3143);
and U3343 (N_3343,N_3112,N_3029);
nand U3344 (N_3344,N_3061,N_3160);
nand U3345 (N_3345,N_3182,N_3107);
and U3346 (N_3346,N_3133,N_3092);
nand U3347 (N_3347,N_3044,N_3092);
nand U3348 (N_3348,N_3196,N_3047);
nor U3349 (N_3349,N_3073,N_3087);
or U3350 (N_3350,N_3119,N_3023);
nand U3351 (N_3351,N_3001,N_3057);
nand U3352 (N_3352,N_3053,N_3066);
nor U3353 (N_3353,N_3030,N_3092);
xnor U3354 (N_3354,N_3152,N_3191);
nor U3355 (N_3355,N_3106,N_3111);
nor U3356 (N_3356,N_3031,N_3134);
nand U3357 (N_3357,N_3054,N_3181);
or U3358 (N_3358,N_3114,N_3101);
and U3359 (N_3359,N_3144,N_3091);
and U3360 (N_3360,N_3070,N_3186);
or U3361 (N_3361,N_3183,N_3108);
or U3362 (N_3362,N_3180,N_3061);
xnor U3363 (N_3363,N_3153,N_3010);
xnor U3364 (N_3364,N_3159,N_3091);
xor U3365 (N_3365,N_3187,N_3163);
nor U3366 (N_3366,N_3080,N_3112);
or U3367 (N_3367,N_3047,N_3170);
xor U3368 (N_3368,N_3176,N_3167);
nor U3369 (N_3369,N_3076,N_3068);
xnor U3370 (N_3370,N_3147,N_3007);
and U3371 (N_3371,N_3011,N_3017);
or U3372 (N_3372,N_3096,N_3099);
nor U3373 (N_3373,N_3064,N_3048);
xnor U3374 (N_3374,N_3103,N_3118);
or U3375 (N_3375,N_3145,N_3043);
nand U3376 (N_3376,N_3063,N_3019);
nand U3377 (N_3377,N_3136,N_3015);
xor U3378 (N_3378,N_3042,N_3088);
nor U3379 (N_3379,N_3173,N_3112);
or U3380 (N_3380,N_3079,N_3193);
nand U3381 (N_3381,N_3060,N_3172);
nand U3382 (N_3382,N_3163,N_3091);
or U3383 (N_3383,N_3027,N_3162);
or U3384 (N_3384,N_3045,N_3103);
nor U3385 (N_3385,N_3063,N_3025);
nor U3386 (N_3386,N_3054,N_3167);
and U3387 (N_3387,N_3132,N_3117);
xor U3388 (N_3388,N_3034,N_3186);
xor U3389 (N_3389,N_3001,N_3048);
xnor U3390 (N_3390,N_3138,N_3058);
nor U3391 (N_3391,N_3199,N_3193);
and U3392 (N_3392,N_3186,N_3073);
nor U3393 (N_3393,N_3071,N_3012);
xor U3394 (N_3394,N_3115,N_3188);
or U3395 (N_3395,N_3168,N_3065);
xnor U3396 (N_3396,N_3143,N_3063);
and U3397 (N_3397,N_3073,N_3077);
nand U3398 (N_3398,N_3024,N_3181);
nand U3399 (N_3399,N_3176,N_3050);
and U3400 (N_3400,N_3223,N_3234);
or U3401 (N_3401,N_3387,N_3396);
nand U3402 (N_3402,N_3240,N_3232);
xor U3403 (N_3403,N_3349,N_3276);
nor U3404 (N_3404,N_3311,N_3369);
xnor U3405 (N_3405,N_3318,N_3213);
nand U3406 (N_3406,N_3281,N_3365);
nand U3407 (N_3407,N_3221,N_3344);
nor U3408 (N_3408,N_3378,N_3388);
xnor U3409 (N_3409,N_3353,N_3341);
nor U3410 (N_3410,N_3391,N_3266);
xnor U3411 (N_3411,N_3201,N_3210);
xnor U3412 (N_3412,N_3254,N_3329);
xor U3413 (N_3413,N_3324,N_3309);
xor U3414 (N_3414,N_3268,N_3306);
xor U3415 (N_3415,N_3299,N_3323);
nand U3416 (N_3416,N_3204,N_3383);
nand U3417 (N_3417,N_3345,N_3308);
nand U3418 (N_3418,N_3314,N_3262);
nor U3419 (N_3419,N_3357,N_3363);
and U3420 (N_3420,N_3284,N_3360);
xnor U3421 (N_3421,N_3233,N_3313);
and U3422 (N_3422,N_3216,N_3297);
and U3423 (N_3423,N_3257,N_3265);
or U3424 (N_3424,N_3261,N_3352);
and U3425 (N_3425,N_3279,N_3200);
and U3426 (N_3426,N_3244,N_3250);
or U3427 (N_3427,N_3251,N_3248);
or U3428 (N_3428,N_3272,N_3399);
nor U3429 (N_3429,N_3390,N_3290);
nor U3430 (N_3430,N_3245,N_3212);
and U3431 (N_3431,N_3348,N_3338);
and U3432 (N_3432,N_3382,N_3325);
or U3433 (N_3433,N_3370,N_3303);
nand U3434 (N_3434,N_3226,N_3280);
nor U3435 (N_3435,N_3243,N_3298);
nor U3436 (N_3436,N_3332,N_3236);
nor U3437 (N_3437,N_3368,N_3249);
nor U3438 (N_3438,N_3277,N_3220);
nand U3439 (N_3439,N_3205,N_3230);
and U3440 (N_3440,N_3337,N_3334);
nand U3441 (N_3441,N_3289,N_3207);
and U3442 (N_3442,N_3376,N_3287);
xnor U3443 (N_3443,N_3218,N_3231);
or U3444 (N_3444,N_3260,N_3291);
xor U3445 (N_3445,N_3300,N_3385);
xnor U3446 (N_3446,N_3274,N_3393);
or U3447 (N_3447,N_3347,N_3229);
and U3448 (N_3448,N_3307,N_3356);
or U3449 (N_3449,N_3346,N_3215);
nand U3450 (N_3450,N_3367,N_3246);
xor U3451 (N_3451,N_3288,N_3374);
nand U3452 (N_3452,N_3342,N_3361);
or U3453 (N_3453,N_3371,N_3331);
xnor U3454 (N_3454,N_3312,N_3253);
or U3455 (N_3455,N_3259,N_3269);
xnor U3456 (N_3456,N_3235,N_3214);
xor U3457 (N_3457,N_3294,N_3238);
and U3458 (N_3458,N_3362,N_3217);
and U3459 (N_3459,N_3270,N_3228);
nand U3460 (N_3460,N_3310,N_3319);
xor U3461 (N_3461,N_3282,N_3258);
nor U3462 (N_3462,N_3327,N_3242);
nor U3463 (N_3463,N_3392,N_3364);
nor U3464 (N_3464,N_3389,N_3315);
xor U3465 (N_3465,N_3225,N_3267);
xnor U3466 (N_3466,N_3285,N_3203);
nor U3467 (N_3467,N_3380,N_3386);
and U3468 (N_3468,N_3255,N_3321);
or U3469 (N_3469,N_3275,N_3320);
nand U3470 (N_3470,N_3209,N_3273);
nor U3471 (N_3471,N_3379,N_3358);
nand U3472 (N_3472,N_3224,N_3283);
xnor U3473 (N_3473,N_3295,N_3278);
or U3474 (N_3474,N_3286,N_3301);
and U3475 (N_3475,N_3256,N_3293);
and U3476 (N_3476,N_3373,N_3271);
or U3477 (N_3477,N_3219,N_3394);
xor U3478 (N_3478,N_3375,N_3206);
nor U3479 (N_3479,N_3398,N_3354);
or U3480 (N_3480,N_3372,N_3366);
xor U3481 (N_3481,N_3330,N_3322);
nand U3482 (N_3482,N_3237,N_3395);
or U3483 (N_3483,N_3340,N_3326);
xor U3484 (N_3484,N_3208,N_3222);
nand U3485 (N_3485,N_3316,N_3302);
or U3486 (N_3486,N_3305,N_3202);
nand U3487 (N_3487,N_3351,N_3336);
nand U3488 (N_3488,N_3239,N_3350);
nand U3489 (N_3489,N_3343,N_3335);
or U3490 (N_3490,N_3263,N_3339);
xnor U3491 (N_3491,N_3211,N_3252);
xnor U3492 (N_3492,N_3241,N_3384);
and U3493 (N_3493,N_3333,N_3355);
or U3494 (N_3494,N_3292,N_3264);
xnor U3495 (N_3495,N_3227,N_3247);
or U3496 (N_3496,N_3397,N_3317);
nand U3497 (N_3497,N_3359,N_3296);
nor U3498 (N_3498,N_3328,N_3377);
and U3499 (N_3499,N_3304,N_3381);
or U3500 (N_3500,N_3318,N_3355);
nand U3501 (N_3501,N_3208,N_3359);
and U3502 (N_3502,N_3342,N_3301);
and U3503 (N_3503,N_3249,N_3318);
nand U3504 (N_3504,N_3339,N_3209);
nor U3505 (N_3505,N_3214,N_3252);
xnor U3506 (N_3506,N_3370,N_3296);
and U3507 (N_3507,N_3255,N_3266);
nor U3508 (N_3508,N_3347,N_3394);
nand U3509 (N_3509,N_3293,N_3384);
and U3510 (N_3510,N_3200,N_3216);
xor U3511 (N_3511,N_3397,N_3352);
and U3512 (N_3512,N_3304,N_3219);
and U3513 (N_3513,N_3205,N_3268);
nor U3514 (N_3514,N_3341,N_3363);
nand U3515 (N_3515,N_3292,N_3250);
nand U3516 (N_3516,N_3220,N_3386);
xnor U3517 (N_3517,N_3297,N_3258);
or U3518 (N_3518,N_3244,N_3213);
xnor U3519 (N_3519,N_3373,N_3235);
nand U3520 (N_3520,N_3283,N_3379);
xnor U3521 (N_3521,N_3316,N_3348);
or U3522 (N_3522,N_3374,N_3336);
nand U3523 (N_3523,N_3241,N_3217);
or U3524 (N_3524,N_3203,N_3246);
or U3525 (N_3525,N_3240,N_3375);
xnor U3526 (N_3526,N_3372,N_3333);
nor U3527 (N_3527,N_3316,N_3360);
nand U3528 (N_3528,N_3370,N_3255);
and U3529 (N_3529,N_3359,N_3383);
nand U3530 (N_3530,N_3362,N_3209);
nor U3531 (N_3531,N_3235,N_3286);
nor U3532 (N_3532,N_3292,N_3237);
xnor U3533 (N_3533,N_3278,N_3242);
and U3534 (N_3534,N_3235,N_3314);
and U3535 (N_3535,N_3216,N_3324);
nand U3536 (N_3536,N_3317,N_3205);
or U3537 (N_3537,N_3251,N_3380);
nand U3538 (N_3538,N_3384,N_3335);
xor U3539 (N_3539,N_3289,N_3322);
xnor U3540 (N_3540,N_3354,N_3213);
nor U3541 (N_3541,N_3246,N_3250);
or U3542 (N_3542,N_3305,N_3352);
and U3543 (N_3543,N_3304,N_3352);
nor U3544 (N_3544,N_3202,N_3343);
and U3545 (N_3545,N_3285,N_3332);
xnor U3546 (N_3546,N_3249,N_3289);
or U3547 (N_3547,N_3354,N_3360);
xnor U3548 (N_3548,N_3228,N_3267);
nand U3549 (N_3549,N_3332,N_3364);
xnor U3550 (N_3550,N_3394,N_3291);
xnor U3551 (N_3551,N_3377,N_3249);
and U3552 (N_3552,N_3272,N_3214);
nor U3553 (N_3553,N_3301,N_3386);
nand U3554 (N_3554,N_3213,N_3267);
xor U3555 (N_3555,N_3333,N_3217);
or U3556 (N_3556,N_3217,N_3393);
xor U3557 (N_3557,N_3324,N_3377);
xor U3558 (N_3558,N_3329,N_3360);
nand U3559 (N_3559,N_3388,N_3267);
nor U3560 (N_3560,N_3352,N_3282);
and U3561 (N_3561,N_3397,N_3311);
and U3562 (N_3562,N_3243,N_3373);
or U3563 (N_3563,N_3279,N_3271);
xnor U3564 (N_3564,N_3235,N_3329);
nor U3565 (N_3565,N_3385,N_3264);
xnor U3566 (N_3566,N_3363,N_3295);
or U3567 (N_3567,N_3399,N_3306);
nor U3568 (N_3568,N_3252,N_3301);
nand U3569 (N_3569,N_3306,N_3215);
or U3570 (N_3570,N_3364,N_3346);
and U3571 (N_3571,N_3201,N_3315);
nor U3572 (N_3572,N_3350,N_3311);
nor U3573 (N_3573,N_3223,N_3250);
and U3574 (N_3574,N_3387,N_3287);
and U3575 (N_3575,N_3264,N_3361);
and U3576 (N_3576,N_3287,N_3392);
xnor U3577 (N_3577,N_3381,N_3350);
or U3578 (N_3578,N_3291,N_3358);
xnor U3579 (N_3579,N_3356,N_3358);
nand U3580 (N_3580,N_3286,N_3323);
xor U3581 (N_3581,N_3342,N_3380);
or U3582 (N_3582,N_3321,N_3384);
nor U3583 (N_3583,N_3255,N_3385);
nand U3584 (N_3584,N_3344,N_3380);
and U3585 (N_3585,N_3217,N_3215);
and U3586 (N_3586,N_3248,N_3304);
xnor U3587 (N_3587,N_3380,N_3335);
or U3588 (N_3588,N_3271,N_3358);
xor U3589 (N_3589,N_3342,N_3224);
nor U3590 (N_3590,N_3387,N_3243);
nor U3591 (N_3591,N_3267,N_3354);
or U3592 (N_3592,N_3362,N_3221);
xor U3593 (N_3593,N_3361,N_3203);
or U3594 (N_3594,N_3237,N_3270);
nand U3595 (N_3595,N_3325,N_3320);
nand U3596 (N_3596,N_3284,N_3273);
or U3597 (N_3597,N_3346,N_3312);
or U3598 (N_3598,N_3283,N_3355);
xnor U3599 (N_3599,N_3387,N_3286);
or U3600 (N_3600,N_3499,N_3534);
and U3601 (N_3601,N_3578,N_3476);
or U3602 (N_3602,N_3408,N_3516);
and U3603 (N_3603,N_3531,N_3466);
nand U3604 (N_3604,N_3450,N_3519);
xnor U3605 (N_3605,N_3539,N_3412);
nor U3606 (N_3606,N_3564,N_3555);
xor U3607 (N_3607,N_3436,N_3455);
or U3608 (N_3608,N_3494,N_3416);
xnor U3609 (N_3609,N_3544,N_3524);
nor U3610 (N_3610,N_3532,N_3421);
nor U3611 (N_3611,N_3487,N_3521);
nor U3612 (N_3612,N_3439,N_3549);
nand U3613 (N_3613,N_3481,N_3420);
and U3614 (N_3614,N_3590,N_3495);
xnor U3615 (N_3615,N_3468,N_3536);
nor U3616 (N_3616,N_3509,N_3489);
or U3617 (N_3617,N_3520,N_3484);
nor U3618 (N_3618,N_3570,N_3542);
and U3619 (N_3619,N_3458,N_3589);
and U3620 (N_3620,N_3454,N_3418);
or U3621 (N_3621,N_3559,N_3488);
or U3622 (N_3622,N_3596,N_3514);
nor U3623 (N_3623,N_3429,N_3551);
nor U3624 (N_3624,N_3535,N_3417);
nor U3625 (N_3625,N_3594,N_3441);
and U3626 (N_3626,N_3595,N_3410);
nor U3627 (N_3627,N_3548,N_3471);
and U3628 (N_3628,N_3401,N_3546);
nand U3629 (N_3629,N_3486,N_3438);
nand U3630 (N_3630,N_3558,N_3496);
or U3631 (N_3631,N_3586,N_3437);
nor U3632 (N_3632,N_3423,N_3428);
or U3633 (N_3633,N_3477,N_3587);
xor U3634 (N_3634,N_3561,N_3527);
or U3635 (N_3635,N_3550,N_3599);
nand U3636 (N_3636,N_3427,N_3498);
nand U3637 (N_3637,N_3407,N_3442);
nand U3638 (N_3638,N_3537,N_3465);
or U3639 (N_3639,N_3447,N_3591);
nand U3640 (N_3640,N_3434,N_3457);
nor U3641 (N_3641,N_3577,N_3492);
nor U3642 (N_3642,N_3545,N_3448);
xnor U3643 (N_3643,N_3409,N_3568);
or U3644 (N_3644,N_3581,N_3517);
nor U3645 (N_3645,N_3403,N_3415);
and U3646 (N_3646,N_3430,N_3422);
nor U3647 (N_3647,N_3400,N_3593);
nand U3648 (N_3648,N_3583,N_3552);
nor U3649 (N_3649,N_3510,N_3449);
nand U3650 (N_3650,N_3435,N_3526);
xnor U3651 (N_3651,N_3523,N_3515);
or U3652 (N_3652,N_3553,N_3574);
or U3653 (N_3653,N_3431,N_3480);
or U3654 (N_3654,N_3563,N_3529);
or U3655 (N_3655,N_3566,N_3585);
xor U3656 (N_3656,N_3597,N_3541);
and U3657 (N_3657,N_3575,N_3459);
nor U3658 (N_3658,N_3470,N_3413);
or U3659 (N_3659,N_3445,N_3525);
or U3660 (N_3660,N_3567,N_3414);
nor U3661 (N_3661,N_3402,N_3560);
or U3662 (N_3662,N_3497,N_3503);
xnor U3663 (N_3663,N_3440,N_3513);
and U3664 (N_3664,N_3461,N_3571);
nor U3665 (N_3665,N_3547,N_3543);
nand U3666 (N_3666,N_3556,N_3576);
xor U3667 (N_3667,N_3491,N_3404);
xor U3668 (N_3668,N_3530,N_3528);
and U3669 (N_3669,N_3507,N_3554);
nor U3670 (N_3670,N_3467,N_3478);
nor U3671 (N_3671,N_3452,N_3518);
nor U3672 (N_3672,N_3501,N_3573);
or U3673 (N_3673,N_3598,N_3474);
nor U3674 (N_3674,N_3584,N_3579);
xor U3675 (N_3675,N_3490,N_3562);
or U3676 (N_3676,N_3504,N_3592);
xor U3677 (N_3677,N_3572,N_3565);
nor U3678 (N_3678,N_3426,N_3469);
nor U3679 (N_3679,N_3453,N_3512);
nand U3680 (N_3680,N_3482,N_3500);
nor U3681 (N_3681,N_3580,N_3462);
or U3682 (N_3682,N_3432,N_3569);
xnor U3683 (N_3683,N_3444,N_3485);
nor U3684 (N_3684,N_3464,N_3463);
or U3685 (N_3685,N_3582,N_3472);
or U3686 (N_3686,N_3424,N_3540);
nor U3687 (N_3687,N_3511,N_3446);
and U3688 (N_3688,N_3405,N_3479);
xor U3689 (N_3689,N_3493,N_3443);
and U3690 (N_3690,N_3451,N_3406);
nand U3691 (N_3691,N_3508,N_3411);
or U3692 (N_3692,N_3538,N_3475);
nand U3693 (N_3693,N_3473,N_3483);
xnor U3694 (N_3694,N_3425,N_3419);
nor U3695 (N_3695,N_3433,N_3456);
and U3696 (N_3696,N_3505,N_3557);
nor U3697 (N_3697,N_3460,N_3502);
or U3698 (N_3698,N_3588,N_3506);
and U3699 (N_3699,N_3522,N_3533);
nor U3700 (N_3700,N_3404,N_3406);
xnor U3701 (N_3701,N_3468,N_3489);
nand U3702 (N_3702,N_3557,N_3403);
xnor U3703 (N_3703,N_3483,N_3580);
and U3704 (N_3704,N_3459,N_3452);
or U3705 (N_3705,N_3494,N_3569);
nor U3706 (N_3706,N_3479,N_3520);
xor U3707 (N_3707,N_3524,N_3558);
nand U3708 (N_3708,N_3465,N_3495);
xnor U3709 (N_3709,N_3539,N_3478);
or U3710 (N_3710,N_3413,N_3556);
nand U3711 (N_3711,N_3577,N_3559);
and U3712 (N_3712,N_3578,N_3445);
and U3713 (N_3713,N_3527,N_3436);
or U3714 (N_3714,N_3592,N_3561);
nand U3715 (N_3715,N_3510,N_3430);
or U3716 (N_3716,N_3505,N_3543);
and U3717 (N_3717,N_3428,N_3582);
or U3718 (N_3718,N_3453,N_3592);
and U3719 (N_3719,N_3513,N_3481);
or U3720 (N_3720,N_3513,N_3473);
nand U3721 (N_3721,N_3563,N_3571);
or U3722 (N_3722,N_3439,N_3567);
nand U3723 (N_3723,N_3547,N_3402);
or U3724 (N_3724,N_3495,N_3573);
nand U3725 (N_3725,N_3452,N_3553);
and U3726 (N_3726,N_3527,N_3449);
xnor U3727 (N_3727,N_3445,N_3533);
xnor U3728 (N_3728,N_3456,N_3587);
xor U3729 (N_3729,N_3469,N_3546);
and U3730 (N_3730,N_3462,N_3571);
or U3731 (N_3731,N_3501,N_3551);
and U3732 (N_3732,N_3479,N_3565);
or U3733 (N_3733,N_3544,N_3538);
or U3734 (N_3734,N_3587,N_3594);
or U3735 (N_3735,N_3500,N_3564);
and U3736 (N_3736,N_3596,N_3413);
nand U3737 (N_3737,N_3574,N_3409);
nor U3738 (N_3738,N_3482,N_3462);
xor U3739 (N_3739,N_3549,N_3416);
xnor U3740 (N_3740,N_3481,N_3594);
or U3741 (N_3741,N_3511,N_3582);
and U3742 (N_3742,N_3448,N_3425);
or U3743 (N_3743,N_3513,N_3514);
nor U3744 (N_3744,N_3541,N_3496);
nand U3745 (N_3745,N_3583,N_3465);
nand U3746 (N_3746,N_3488,N_3496);
nand U3747 (N_3747,N_3490,N_3487);
nor U3748 (N_3748,N_3543,N_3427);
nand U3749 (N_3749,N_3429,N_3489);
nand U3750 (N_3750,N_3514,N_3456);
and U3751 (N_3751,N_3550,N_3577);
xor U3752 (N_3752,N_3400,N_3526);
or U3753 (N_3753,N_3594,N_3540);
nand U3754 (N_3754,N_3491,N_3538);
and U3755 (N_3755,N_3409,N_3425);
and U3756 (N_3756,N_3416,N_3595);
xnor U3757 (N_3757,N_3461,N_3430);
nand U3758 (N_3758,N_3536,N_3428);
or U3759 (N_3759,N_3570,N_3505);
nor U3760 (N_3760,N_3538,N_3552);
and U3761 (N_3761,N_3574,N_3560);
or U3762 (N_3762,N_3583,N_3566);
nand U3763 (N_3763,N_3515,N_3451);
nor U3764 (N_3764,N_3518,N_3561);
nand U3765 (N_3765,N_3560,N_3428);
and U3766 (N_3766,N_3468,N_3404);
nor U3767 (N_3767,N_3529,N_3459);
and U3768 (N_3768,N_3441,N_3468);
nor U3769 (N_3769,N_3477,N_3553);
nand U3770 (N_3770,N_3467,N_3428);
and U3771 (N_3771,N_3450,N_3426);
nor U3772 (N_3772,N_3445,N_3597);
or U3773 (N_3773,N_3482,N_3505);
or U3774 (N_3774,N_3570,N_3559);
or U3775 (N_3775,N_3407,N_3439);
xor U3776 (N_3776,N_3454,N_3577);
or U3777 (N_3777,N_3510,N_3514);
and U3778 (N_3778,N_3431,N_3522);
and U3779 (N_3779,N_3450,N_3588);
nand U3780 (N_3780,N_3525,N_3544);
xor U3781 (N_3781,N_3529,N_3571);
and U3782 (N_3782,N_3503,N_3562);
nand U3783 (N_3783,N_3545,N_3498);
or U3784 (N_3784,N_3439,N_3531);
nand U3785 (N_3785,N_3543,N_3572);
or U3786 (N_3786,N_3476,N_3450);
xnor U3787 (N_3787,N_3400,N_3434);
nor U3788 (N_3788,N_3451,N_3575);
nor U3789 (N_3789,N_3550,N_3487);
nor U3790 (N_3790,N_3571,N_3436);
xnor U3791 (N_3791,N_3522,N_3457);
or U3792 (N_3792,N_3541,N_3425);
and U3793 (N_3793,N_3571,N_3448);
nor U3794 (N_3794,N_3428,N_3415);
or U3795 (N_3795,N_3403,N_3574);
or U3796 (N_3796,N_3410,N_3573);
or U3797 (N_3797,N_3417,N_3517);
and U3798 (N_3798,N_3421,N_3471);
nor U3799 (N_3799,N_3452,N_3437);
xor U3800 (N_3800,N_3683,N_3647);
or U3801 (N_3801,N_3741,N_3621);
xnor U3802 (N_3802,N_3617,N_3654);
nor U3803 (N_3803,N_3673,N_3783);
and U3804 (N_3804,N_3678,N_3752);
nor U3805 (N_3805,N_3750,N_3653);
nand U3806 (N_3806,N_3727,N_3793);
nand U3807 (N_3807,N_3724,N_3706);
and U3808 (N_3808,N_3627,N_3603);
or U3809 (N_3809,N_3639,N_3662);
nor U3810 (N_3810,N_3782,N_3762);
xor U3811 (N_3811,N_3642,N_3784);
xnor U3812 (N_3812,N_3710,N_3643);
and U3813 (N_3813,N_3666,N_3791);
xor U3814 (N_3814,N_3624,N_3789);
xnor U3815 (N_3815,N_3798,N_3708);
and U3816 (N_3816,N_3799,N_3797);
nor U3817 (N_3817,N_3615,N_3610);
and U3818 (N_3818,N_3619,N_3732);
nor U3819 (N_3819,N_3601,N_3764);
xor U3820 (N_3820,N_3620,N_3770);
or U3821 (N_3821,N_3622,N_3777);
nor U3822 (N_3822,N_3700,N_3664);
nand U3823 (N_3823,N_3690,N_3759);
or U3824 (N_3824,N_3614,N_3788);
nor U3825 (N_3825,N_3736,N_3696);
or U3826 (N_3826,N_3697,N_3607);
nor U3827 (N_3827,N_3787,N_3689);
xnor U3828 (N_3828,N_3719,N_3748);
xor U3829 (N_3829,N_3657,N_3716);
and U3830 (N_3830,N_3705,N_3723);
nor U3831 (N_3831,N_3794,N_3667);
xnor U3832 (N_3832,N_3650,N_3681);
nand U3833 (N_3833,N_3611,N_3633);
nor U3834 (N_3834,N_3602,N_3780);
nand U3835 (N_3835,N_3648,N_3746);
and U3836 (N_3836,N_3720,N_3671);
xor U3837 (N_3837,N_3790,N_3768);
nor U3838 (N_3838,N_3684,N_3652);
xor U3839 (N_3839,N_3767,N_3707);
and U3840 (N_3840,N_3781,N_3682);
or U3841 (N_3841,N_3663,N_3651);
xnor U3842 (N_3842,N_3747,N_3628);
nand U3843 (N_3843,N_3718,N_3763);
or U3844 (N_3844,N_3743,N_3735);
nor U3845 (N_3845,N_3731,N_3668);
nand U3846 (N_3846,N_3795,N_3641);
xnor U3847 (N_3847,N_3618,N_3659);
nand U3848 (N_3848,N_3665,N_3769);
and U3849 (N_3849,N_3677,N_3728);
xor U3850 (N_3850,N_3629,N_3771);
nor U3851 (N_3851,N_3632,N_3729);
and U3852 (N_3852,N_3714,N_3608);
and U3853 (N_3853,N_3649,N_3715);
and U3854 (N_3854,N_3712,N_3721);
nand U3855 (N_3855,N_3775,N_3703);
xor U3856 (N_3856,N_3717,N_3645);
and U3857 (N_3857,N_3630,N_3740);
nand U3858 (N_3858,N_3695,N_3637);
and U3859 (N_3859,N_3766,N_3745);
nand U3860 (N_3860,N_3757,N_3711);
and U3861 (N_3861,N_3686,N_3744);
and U3862 (N_3862,N_3606,N_3680);
nor U3863 (N_3863,N_3774,N_3704);
or U3864 (N_3864,N_3730,N_3760);
xor U3865 (N_3865,N_3609,N_3698);
nor U3866 (N_3866,N_3604,N_3679);
xnor U3867 (N_3867,N_3638,N_3772);
and U3868 (N_3868,N_3623,N_3733);
xnor U3869 (N_3869,N_3792,N_3640);
nand U3870 (N_3870,N_3613,N_3674);
xor U3871 (N_3871,N_3687,N_3634);
nand U3872 (N_3872,N_3636,N_3786);
nor U3873 (N_3873,N_3656,N_3778);
and U3874 (N_3874,N_3693,N_3773);
and U3875 (N_3875,N_3753,N_3694);
nor U3876 (N_3876,N_3699,N_3761);
or U3877 (N_3877,N_3702,N_3749);
and U3878 (N_3878,N_3672,N_3765);
or U3879 (N_3879,N_3644,N_3658);
nand U3880 (N_3880,N_3692,N_3726);
nand U3881 (N_3881,N_3779,N_3612);
or U3882 (N_3882,N_3756,N_3655);
nand U3883 (N_3883,N_3616,N_3709);
and U3884 (N_3884,N_3701,N_3605);
or U3885 (N_3885,N_3661,N_3758);
or U3886 (N_3886,N_3737,N_3625);
nor U3887 (N_3887,N_3742,N_3751);
nand U3888 (N_3888,N_3685,N_3676);
and U3889 (N_3889,N_3600,N_3785);
or U3890 (N_3890,N_3635,N_3754);
xnor U3891 (N_3891,N_3725,N_3660);
xor U3892 (N_3892,N_3755,N_3631);
nor U3893 (N_3893,N_3713,N_3669);
and U3894 (N_3894,N_3675,N_3739);
and U3895 (N_3895,N_3688,N_3776);
nor U3896 (N_3896,N_3734,N_3646);
nand U3897 (N_3897,N_3722,N_3670);
nand U3898 (N_3898,N_3691,N_3796);
nor U3899 (N_3899,N_3738,N_3626);
and U3900 (N_3900,N_3668,N_3707);
nor U3901 (N_3901,N_3640,N_3715);
nand U3902 (N_3902,N_3751,N_3658);
and U3903 (N_3903,N_3633,N_3784);
nand U3904 (N_3904,N_3639,N_3605);
or U3905 (N_3905,N_3710,N_3783);
nand U3906 (N_3906,N_3642,N_3763);
or U3907 (N_3907,N_3650,N_3799);
nand U3908 (N_3908,N_3633,N_3674);
or U3909 (N_3909,N_3604,N_3697);
nor U3910 (N_3910,N_3731,N_3602);
and U3911 (N_3911,N_3716,N_3691);
xor U3912 (N_3912,N_3728,N_3701);
and U3913 (N_3913,N_3701,N_3786);
xor U3914 (N_3914,N_3670,N_3736);
xor U3915 (N_3915,N_3717,N_3691);
nor U3916 (N_3916,N_3730,N_3609);
nand U3917 (N_3917,N_3696,N_3729);
or U3918 (N_3918,N_3692,N_3732);
or U3919 (N_3919,N_3738,N_3791);
and U3920 (N_3920,N_3758,N_3637);
or U3921 (N_3921,N_3741,N_3677);
nand U3922 (N_3922,N_3648,N_3736);
or U3923 (N_3923,N_3782,N_3675);
nor U3924 (N_3924,N_3618,N_3704);
nand U3925 (N_3925,N_3716,N_3698);
or U3926 (N_3926,N_3676,N_3615);
nor U3927 (N_3927,N_3753,N_3631);
xnor U3928 (N_3928,N_3674,N_3799);
or U3929 (N_3929,N_3610,N_3628);
nand U3930 (N_3930,N_3678,N_3708);
xor U3931 (N_3931,N_3637,N_3748);
xnor U3932 (N_3932,N_3699,N_3648);
nand U3933 (N_3933,N_3664,N_3697);
and U3934 (N_3934,N_3755,N_3776);
and U3935 (N_3935,N_3740,N_3632);
nor U3936 (N_3936,N_3645,N_3635);
and U3937 (N_3937,N_3616,N_3750);
nand U3938 (N_3938,N_3743,N_3733);
or U3939 (N_3939,N_3760,N_3601);
and U3940 (N_3940,N_3746,N_3697);
nand U3941 (N_3941,N_3793,N_3627);
and U3942 (N_3942,N_3764,N_3777);
nor U3943 (N_3943,N_3696,N_3746);
nand U3944 (N_3944,N_3735,N_3722);
xnor U3945 (N_3945,N_3681,N_3729);
or U3946 (N_3946,N_3768,N_3758);
xor U3947 (N_3947,N_3641,N_3758);
and U3948 (N_3948,N_3716,N_3708);
nor U3949 (N_3949,N_3695,N_3639);
and U3950 (N_3950,N_3609,N_3629);
nand U3951 (N_3951,N_3614,N_3709);
or U3952 (N_3952,N_3736,N_3701);
or U3953 (N_3953,N_3627,N_3761);
xnor U3954 (N_3954,N_3653,N_3607);
xor U3955 (N_3955,N_3630,N_3774);
nand U3956 (N_3956,N_3703,N_3750);
or U3957 (N_3957,N_3652,N_3648);
nand U3958 (N_3958,N_3625,N_3671);
or U3959 (N_3959,N_3633,N_3645);
xor U3960 (N_3960,N_3746,N_3625);
and U3961 (N_3961,N_3772,N_3609);
xnor U3962 (N_3962,N_3626,N_3624);
and U3963 (N_3963,N_3679,N_3729);
nor U3964 (N_3964,N_3677,N_3614);
nor U3965 (N_3965,N_3689,N_3696);
nor U3966 (N_3966,N_3707,N_3608);
nor U3967 (N_3967,N_3700,N_3616);
xnor U3968 (N_3968,N_3721,N_3672);
and U3969 (N_3969,N_3715,N_3656);
and U3970 (N_3970,N_3724,N_3699);
and U3971 (N_3971,N_3639,N_3674);
and U3972 (N_3972,N_3794,N_3605);
or U3973 (N_3973,N_3658,N_3633);
nand U3974 (N_3974,N_3769,N_3648);
nor U3975 (N_3975,N_3793,N_3707);
or U3976 (N_3976,N_3664,N_3630);
nand U3977 (N_3977,N_3688,N_3637);
nor U3978 (N_3978,N_3770,N_3778);
or U3979 (N_3979,N_3690,N_3641);
nand U3980 (N_3980,N_3609,N_3720);
and U3981 (N_3981,N_3614,N_3799);
nand U3982 (N_3982,N_3757,N_3759);
or U3983 (N_3983,N_3769,N_3788);
or U3984 (N_3984,N_3732,N_3601);
xnor U3985 (N_3985,N_3764,N_3723);
and U3986 (N_3986,N_3714,N_3616);
and U3987 (N_3987,N_3663,N_3618);
nand U3988 (N_3988,N_3786,N_3729);
nand U3989 (N_3989,N_3642,N_3778);
nand U3990 (N_3990,N_3642,N_3618);
and U3991 (N_3991,N_3736,N_3659);
xor U3992 (N_3992,N_3749,N_3689);
nand U3993 (N_3993,N_3717,N_3657);
nand U3994 (N_3994,N_3632,N_3685);
and U3995 (N_3995,N_3618,N_3649);
nor U3996 (N_3996,N_3648,N_3645);
or U3997 (N_3997,N_3779,N_3650);
xor U3998 (N_3998,N_3745,N_3710);
nand U3999 (N_3999,N_3790,N_3724);
or U4000 (N_4000,N_3891,N_3812);
nor U4001 (N_4001,N_3938,N_3928);
xor U4002 (N_4002,N_3948,N_3914);
nor U4003 (N_4003,N_3964,N_3994);
nand U4004 (N_4004,N_3830,N_3820);
and U4005 (N_4005,N_3906,N_3963);
and U4006 (N_4006,N_3806,N_3946);
nand U4007 (N_4007,N_3924,N_3886);
nor U4008 (N_4008,N_3917,N_3930);
or U4009 (N_4009,N_3856,N_3945);
nor U4010 (N_4010,N_3915,N_3801);
and U4011 (N_4011,N_3933,N_3846);
nor U4012 (N_4012,N_3921,N_3864);
nor U4013 (N_4013,N_3923,N_3976);
or U4014 (N_4014,N_3985,N_3872);
nand U4015 (N_4015,N_3977,N_3890);
and U4016 (N_4016,N_3983,N_3868);
nand U4017 (N_4017,N_3804,N_3925);
nor U4018 (N_4018,N_3822,N_3813);
xor U4019 (N_4019,N_3950,N_3800);
nor U4020 (N_4020,N_3805,N_3995);
or U4021 (N_4021,N_3972,N_3823);
or U4022 (N_4022,N_3902,N_3997);
and U4023 (N_4023,N_3895,N_3929);
or U4024 (N_4024,N_3952,N_3847);
nor U4025 (N_4025,N_3918,N_3942);
nand U4026 (N_4026,N_3838,N_3852);
and U4027 (N_4027,N_3877,N_3888);
and U4028 (N_4028,N_3878,N_3916);
nor U4029 (N_4029,N_3885,N_3957);
nand U4030 (N_4030,N_3880,N_3871);
or U4031 (N_4031,N_3892,N_3810);
or U4032 (N_4032,N_3870,N_3966);
or U4033 (N_4033,N_3807,N_3862);
nor U4034 (N_4034,N_3958,N_3860);
nand U4035 (N_4035,N_3980,N_3910);
or U4036 (N_4036,N_3881,N_3836);
or U4037 (N_4037,N_3959,N_3855);
nand U4038 (N_4038,N_3819,N_3841);
nor U4039 (N_4039,N_3986,N_3940);
nor U4040 (N_4040,N_3951,N_3889);
or U4041 (N_4041,N_3832,N_3999);
nor U4042 (N_4042,N_3908,N_3996);
nand U4043 (N_4043,N_3935,N_3874);
or U4044 (N_4044,N_3834,N_3947);
xor U4045 (N_4045,N_3939,N_3802);
or U4046 (N_4046,N_3825,N_3894);
and U4047 (N_4047,N_3936,N_3816);
nand U4048 (N_4048,N_3967,N_3949);
and U4049 (N_4049,N_3861,N_3919);
xor U4050 (N_4050,N_3865,N_3858);
nor U4051 (N_4051,N_3960,N_3969);
or U4052 (N_4052,N_3845,N_3992);
xnor U4053 (N_4053,N_3884,N_3851);
nor U4054 (N_4054,N_3844,N_3943);
nor U4055 (N_4055,N_3989,N_3835);
and U4056 (N_4056,N_3912,N_3991);
nor U4057 (N_4057,N_3934,N_3809);
xor U4058 (N_4058,N_3965,N_3887);
xor U4059 (N_4059,N_3837,N_3876);
nor U4060 (N_4060,N_3828,N_3955);
nand U4061 (N_4061,N_3897,N_3900);
and U4062 (N_4062,N_3869,N_3998);
or U4063 (N_4063,N_3824,N_3867);
nand U4064 (N_4064,N_3941,N_3873);
and U4065 (N_4065,N_3931,N_3843);
nor U4066 (N_4066,N_3982,N_3909);
or U4067 (N_4067,N_3815,N_3905);
nand U4068 (N_4068,N_3883,N_3866);
or U4069 (N_4069,N_3975,N_3882);
and U4070 (N_4070,N_3808,N_3829);
and U4071 (N_4071,N_3961,N_3944);
xor U4072 (N_4072,N_3970,N_3833);
nor U4073 (N_4073,N_3899,N_3978);
nor U4074 (N_4074,N_3971,N_3839);
xor U4075 (N_4075,N_3849,N_3973);
nor U4076 (N_4076,N_3831,N_3875);
or U4077 (N_4077,N_3811,N_3842);
nand U4078 (N_4078,N_3953,N_3974);
xor U4079 (N_4079,N_3893,N_3968);
and U4080 (N_4080,N_3913,N_3927);
xnor U4081 (N_4081,N_3954,N_3898);
nor U4082 (N_4082,N_3907,N_3854);
nand U4083 (N_4083,N_3937,N_3904);
xnor U4084 (N_4084,N_3990,N_3981);
xnor U4085 (N_4085,N_3818,N_3850);
or U4086 (N_4086,N_3817,N_3920);
and U4087 (N_4087,N_3863,N_3879);
xor U4088 (N_4088,N_3853,N_3821);
nand U4089 (N_4089,N_3903,N_3896);
xor U4090 (N_4090,N_3993,N_3848);
or U4091 (N_4091,N_3988,N_3962);
nand U4092 (N_4092,N_3911,N_3901);
nor U4093 (N_4093,N_3803,N_3857);
xor U4094 (N_4094,N_3926,N_3932);
and U4095 (N_4095,N_3956,N_3814);
xnor U4096 (N_4096,N_3826,N_3859);
nor U4097 (N_4097,N_3979,N_3827);
nand U4098 (N_4098,N_3987,N_3840);
nand U4099 (N_4099,N_3984,N_3922);
or U4100 (N_4100,N_3814,N_3839);
nand U4101 (N_4101,N_3918,N_3876);
xor U4102 (N_4102,N_3803,N_3921);
xor U4103 (N_4103,N_3905,N_3858);
nor U4104 (N_4104,N_3996,N_3808);
xnor U4105 (N_4105,N_3996,N_3899);
or U4106 (N_4106,N_3815,N_3940);
nand U4107 (N_4107,N_3974,N_3841);
or U4108 (N_4108,N_3992,N_3843);
nor U4109 (N_4109,N_3981,N_3845);
nor U4110 (N_4110,N_3867,N_3835);
or U4111 (N_4111,N_3867,N_3964);
nand U4112 (N_4112,N_3934,N_3860);
nand U4113 (N_4113,N_3915,N_3967);
or U4114 (N_4114,N_3975,N_3857);
xnor U4115 (N_4115,N_3820,N_3956);
nand U4116 (N_4116,N_3935,N_3961);
nor U4117 (N_4117,N_3923,N_3953);
nor U4118 (N_4118,N_3998,N_3948);
and U4119 (N_4119,N_3971,N_3832);
nand U4120 (N_4120,N_3958,N_3819);
or U4121 (N_4121,N_3949,N_3853);
or U4122 (N_4122,N_3804,N_3989);
xor U4123 (N_4123,N_3858,N_3837);
nor U4124 (N_4124,N_3935,N_3881);
xnor U4125 (N_4125,N_3985,N_3802);
nand U4126 (N_4126,N_3813,N_3986);
or U4127 (N_4127,N_3903,N_3942);
and U4128 (N_4128,N_3944,N_3833);
xnor U4129 (N_4129,N_3909,N_3905);
xor U4130 (N_4130,N_3848,N_3802);
or U4131 (N_4131,N_3923,N_3972);
nand U4132 (N_4132,N_3891,N_3849);
nor U4133 (N_4133,N_3808,N_3928);
xor U4134 (N_4134,N_3952,N_3816);
and U4135 (N_4135,N_3883,N_3906);
xnor U4136 (N_4136,N_3880,N_3995);
nand U4137 (N_4137,N_3865,N_3862);
nor U4138 (N_4138,N_3841,N_3910);
nand U4139 (N_4139,N_3937,N_3883);
and U4140 (N_4140,N_3894,N_3916);
or U4141 (N_4141,N_3904,N_3802);
nand U4142 (N_4142,N_3894,N_3818);
xor U4143 (N_4143,N_3806,N_3826);
or U4144 (N_4144,N_3859,N_3981);
nand U4145 (N_4145,N_3946,N_3881);
nand U4146 (N_4146,N_3863,N_3817);
and U4147 (N_4147,N_3998,N_3908);
nand U4148 (N_4148,N_3912,N_3988);
nor U4149 (N_4149,N_3967,N_3856);
xor U4150 (N_4150,N_3894,N_3900);
and U4151 (N_4151,N_3805,N_3913);
nor U4152 (N_4152,N_3838,N_3991);
xnor U4153 (N_4153,N_3939,N_3837);
nor U4154 (N_4154,N_3818,N_3900);
xnor U4155 (N_4155,N_3946,N_3955);
nand U4156 (N_4156,N_3861,N_3936);
nor U4157 (N_4157,N_3801,N_3825);
nor U4158 (N_4158,N_3995,N_3900);
nor U4159 (N_4159,N_3914,N_3904);
nor U4160 (N_4160,N_3906,N_3960);
xnor U4161 (N_4161,N_3932,N_3836);
or U4162 (N_4162,N_3990,N_3892);
nand U4163 (N_4163,N_3979,N_3987);
or U4164 (N_4164,N_3818,N_3914);
xor U4165 (N_4165,N_3969,N_3881);
xor U4166 (N_4166,N_3928,N_3856);
nand U4167 (N_4167,N_3914,N_3889);
nand U4168 (N_4168,N_3924,N_3800);
and U4169 (N_4169,N_3871,N_3912);
or U4170 (N_4170,N_3947,N_3890);
nor U4171 (N_4171,N_3990,N_3875);
or U4172 (N_4172,N_3847,N_3908);
or U4173 (N_4173,N_3848,N_3913);
xor U4174 (N_4174,N_3930,N_3934);
and U4175 (N_4175,N_3845,N_3966);
xor U4176 (N_4176,N_3902,N_3804);
xor U4177 (N_4177,N_3997,N_3942);
and U4178 (N_4178,N_3922,N_3830);
xnor U4179 (N_4179,N_3886,N_3859);
and U4180 (N_4180,N_3889,N_3854);
nor U4181 (N_4181,N_3945,N_3848);
xor U4182 (N_4182,N_3962,N_3956);
xnor U4183 (N_4183,N_3964,N_3954);
nor U4184 (N_4184,N_3862,N_3957);
or U4185 (N_4185,N_3979,N_3801);
or U4186 (N_4186,N_3877,N_3937);
nand U4187 (N_4187,N_3885,N_3936);
nand U4188 (N_4188,N_3826,N_3903);
nor U4189 (N_4189,N_3905,N_3982);
nand U4190 (N_4190,N_3987,N_3894);
xor U4191 (N_4191,N_3819,N_3943);
xnor U4192 (N_4192,N_3914,N_3840);
xor U4193 (N_4193,N_3805,N_3825);
nor U4194 (N_4194,N_3930,N_3874);
nor U4195 (N_4195,N_3919,N_3831);
nand U4196 (N_4196,N_3930,N_3994);
nor U4197 (N_4197,N_3882,N_3814);
nor U4198 (N_4198,N_3910,N_3804);
xor U4199 (N_4199,N_3896,N_3928);
or U4200 (N_4200,N_4084,N_4058);
nor U4201 (N_4201,N_4191,N_4071);
xnor U4202 (N_4202,N_4102,N_4108);
nand U4203 (N_4203,N_4014,N_4109);
nand U4204 (N_4204,N_4164,N_4182);
xor U4205 (N_4205,N_4138,N_4124);
or U4206 (N_4206,N_4147,N_4028);
xnor U4207 (N_4207,N_4153,N_4050);
xor U4208 (N_4208,N_4094,N_4010);
nor U4209 (N_4209,N_4118,N_4085);
nand U4210 (N_4210,N_4125,N_4117);
nand U4211 (N_4211,N_4065,N_4072);
xnor U4212 (N_4212,N_4196,N_4089);
nand U4213 (N_4213,N_4185,N_4130);
nor U4214 (N_4214,N_4142,N_4063);
or U4215 (N_4215,N_4047,N_4045);
nor U4216 (N_4216,N_4007,N_4022);
nand U4217 (N_4217,N_4111,N_4016);
or U4218 (N_4218,N_4105,N_4175);
nand U4219 (N_4219,N_4123,N_4012);
xor U4220 (N_4220,N_4104,N_4120);
xor U4221 (N_4221,N_4139,N_4181);
xnor U4222 (N_4222,N_4027,N_4056);
and U4223 (N_4223,N_4031,N_4132);
nand U4224 (N_4224,N_4193,N_4140);
xnor U4225 (N_4225,N_4001,N_4005);
and U4226 (N_4226,N_4099,N_4115);
nand U4227 (N_4227,N_4129,N_4034);
xor U4228 (N_4228,N_4026,N_4006);
xnor U4229 (N_4229,N_4011,N_4039);
nand U4230 (N_4230,N_4070,N_4018);
xnor U4231 (N_4231,N_4192,N_4054);
xor U4232 (N_4232,N_4076,N_4144);
nor U4233 (N_4233,N_4101,N_4122);
or U4234 (N_4234,N_4145,N_4075);
xnor U4235 (N_4235,N_4074,N_4051);
and U4236 (N_4236,N_4003,N_4121);
or U4237 (N_4237,N_4095,N_4159);
and U4238 (N_4238,N_4148,N_4092);
nand U4239 (N_4239,N_4106,N_4177);
and U4240 (N_4240,N_4043,N_4146);
and U4241 (N_4241,N_4041,N_4136);
or U4242 (N_4242,N_4154,N_4096);
or U4243 (N_4243,N_4059,N_4152);
and U4244 (N_4244,N_4069,N_4021);
and U4245 (N_4245,N_4008,N_4165);
nand U4246 (N_4246,N_4168,N_4029);
and U4247 (N_4247,N_4093,N_4035);
nand U4248 (N_4248,N_4055,N_4067);
xnor U4249 (N_4249,N_4052,N_4066);
and U4250 (N_4250,N_4135,N_4013);
nor U4251 (N_4251,N_4020,N_4037);
and U4252 (N_4252,N_4033,N_4040);
nor U4253 (N_4253,N_4189,N_4017);
and U4254 (N_4254,N_4114,N_4080);
xor U4255 (N_4255,N_4170,N_4131);
and U4256 (N_4256,N_4048,N_4187);
or U4257 (N_4257,N_4155,N_4156);
nand U4258 (N_4258,N_4169,N_4097);
nor U4259 (N_4259,N_4090,N_4133);
or U4260 (N_4260,N_4128,N_4081);
nor U4261 (N_4261,N_4062,N_4126);
nor U4262 (N_4262,N_4044,N_4143);
and U4263 (N_4263,N_4110,N_4180);
or U4264 (N_4264,N_4015,N_4113);
xnor U4265 (N_4265,N_4174,N_4023);
nand U4266 (N_4266,N_4166,N_4195);
nand U4267 (N_4267,N_4100,N_4197);
xnor U4268 (N_4268,N_4088,N_4030);
or U4269 (N_4269,N_4002,N_4053);
xor U4270 (N_4270,N_4036,N_4078);
nand U4271 (N_4271,N_4186,N_4158);
nor U4272 (N_4272,N_4049,N_4183);
and U4273 (N_4273,N_4019,N_4091);
and U4274 (N_4274,N_4098,N_4061);
xnor U4275 (N_4275,N_4190,N_4046);
nor U4276 (N_4276,N_4087,N_4194);
and U4277 (N_4277,N_4079,N_4112);
and U4278 (N_4278,N_4173,N_4000);
nor U4279 (N_4279,N_4116,N_4057);
nor U4280 (N_4280,N_4162,N_4150);
and U4281 (N_4281,N_4137,N_4198);
or U4282 (N_4282,N_4032,N_4107);
nor U4283 (N_4283,N_4038,N_4163);
or U4284 (N_4284,N_4199,N_4119);
nor U4285 (N_4285,N_4073,N_4176);
and U4286 (N_4286,N_4024,N_4171);
xnor U4287 (N_4287,N_4157,N_4009);
nor U4288 (N_4288,N_4178,N_4141);
nor U4289 (N_4289,N_4161,N_4077);
nor U4290 (N_4290,N_4060,N_4179);
or U4291 (N_4291,N_4068,N_4149);
or U4292 (N_4292,N_4134,N_4188);
nand U4293 (N_4293,N_4167,N_4042);
and U4294 (N_4294,N_4184,N_4004);
nand U4295 (N_4295,N_4086,N_4127);
or U4296 (N_4296,N_4064,N_4103);
nand U4297 (N_4297,N_4172,N_4151);
nor U4298 (N_4298,N_4083,N_4082);
nand U4299 (N_4299,N_4160,N_4025);
xnor U4300 (N_4300,N_4077,N_4078);
nand U4301 (N_4301,N_4194,N_4109);
xor U4302 (N_4302,N_4071,N_4022);
xnor U4303 (N_4303,N_4172,N_4141);
nand U4304 (N_4304,N_4190,N_4142);
nor U4305 (N_4305,N_4111,N_4138);
nand U4306 (N_4306,N_4114,N_4011);
nor U4307 (N_4307,N_4007,N_4023);
nand U4308 (N_4308,N_4136,N_4000);
nand U4309 (N_4309,N_4195,N_4140);
nand U4310 (N_4310,N_4180,N_4182);
nand U4311 (N_4311,N_4186,N_4039);
nor U4312 (N_4312,N_4032,N_4184);
nand U4313 (N_4313,N_4169,N_4047);
or U4314 (N_4314,N_4017,N_4080);
nand U4315 (N_4315,N_4140,N_4076);
nor U4316 (N_4316,N_4095,N_4057);
or U4317 (N_4317,N_4158,N_4135);
nand U4318 (N_4318,N_4063,N_4010);
nor U4319 (N_4319,N_4129,N_4151);
and U4320 (N_4320,N_4164,N_4037);
nand U4321 (N_4321,N_4010,N_4039);
nand U4322 (N_4322,N_4149,N_4033);
nor U4323 (N_4323,N_4176,N_4005);
xnor U4324 (N_4324,N_4047,N_4062);
and U4325 (N_4325,N_4172,N_4161);
nand U4326 (N_4326,N_4012,N_4019);
xor U4327 (N_4327,N_4090,N_4119);
nand U4328 (N_4328,N_4072,N_4052);
xor U4329 (N_4329,N_4035,N_4194);
nor U4330 (N_4330,N_4180,N_4125);
nor U4331 (N_4331,N_4137,N_4013);
xnor U4332 (N_4332,N_4065,N_4056);
nand U4333 (N_4333,N_4198,N_4128);
nor U4334 (N_4334,N_4175,N_4015);
or U4335 (N_4335,N_4045,N_4059);
nor U4336 (N_4336,N_4004,N_4088);
xnor U4337 (N_4337,N_4150,N_4076);
and U4338 (N_4338,N_4047,N_4103);
xnor U4339 (N_4339,N_4109,N_4140);
nor U4340 (N_4340,N_4033,N_4021);
xnor U4341 (N_4341,N_4165,N_4063);
nand U4342 (N_4342,N_4072,N_4185);
nand U4343 (N_4343,N_4090,N_4069);
and U4344 (N_4344,N_4019,N_4055);
and U4345 (N_4345,N_4173,N_4128);
nand U4346 (N_4346,N_4173,N_4103);
or U4347 (N_4347,N_4063,N_4099);
or U4348 (N_4348,N_4048,N_4070);
xnor U4349 (N_4349,N_4092,N_4168);
nand U4350 (N_4350,N_4073,N_4133);
and U4351 (N_4351,N_4039,N_4130);
or U4352 (N_4352,N_4170,N_4125);
nand U4353 (N_4353,N_4058,N_4091);
or U4354 (N_4354,N_4118,N_4004);
and U4355 (N_4355,N_4050,N_4140);
nand U4356 (N_4356,N_4032,N_4123);
nand U4357 (N_4357,N_4070,N_4014);
nor U4358 (N_4358,N_4144,N_4188);
and U4359 (N_4359,N_4087,N_4014);
xor U4360 (N_4360,N_4144,N_4110);
xnor U4361 (N_4361,N_4123,N_4069);
and U4362 (N_4362,N_4027,N_4061);
or U4363 (N_4363,N_4000,N_4164);
and U4364 (N_4364,N_4042,N_4176);
nor U4365 (N_4365,N_4047,N_4063);
nand U4366 (N_4366,N_4194,N_4096);
nand U4367 (N_4367,N_4074,N_4129);
xnor U4368 (N_4368,N_4158,N_4141);
nor U4369 (N_4369,N_4191,N_4128);
nor U4370 (N_4370,N_4198,N_4179);
xnor U4371 (N_4371,N_4064,N_4062);
and U4372 (N_4372,N_4177,N_4199);
or U4373 (N_4373,N_4165,N_4116);
nor U4374 (N_4374,N_4021,N_4006);
nor U4375 (N_4375,N_4184,N_4081);
or U4376 (N_4376,N_4188,N_4129);
nand U4377 (N_4377,N_4047,N_4036);
or U4378 (N_4378,N_4061,N_4053);
nor U4379 (N_4379,N_4140,N_4031);
or U4380 (N_4380,N_4061,N_4015);
or U4381 (N_4381,N_4181,N_4195);
nand U4382 (N_4382,N_4167,N_4020);
xnor U4383 (N_4383,N_4052,N_4192);
or U4384 (N_4384,N_4167,N_4172);
xor U4385 (N_4385,N_4091,N_4142);
nor U4386 (N_4386,N_4049,N_4033);
xnor U4387 (N_4387,N_4105,N_4014);
or U4388 (N_4388,N_4135,N_4054);
xnor U4389 (N_4389,N_4112,N_4100);
nor U4390 (N_4390,N_4054,N_4118);
and U4391 (N_4391,N_4129,N_4021);
and U4392 (N_4392,N_4020,N_4140);
or U4393 (N_4393,N_4088,N_4115);
nor U4394 (N_4394,N_4111,N_4042);
nand U4395 (N_4395,N_4123,N_4077);
and U4396 (N_4396,N_4091,N_4175);
and U4397 (N_4397,N_4178,N_4143);
nand U4398 (N_4398,N_4087,N_4180);
and U4399 (N_4399,N_4097,N_4188);
nand U4400 (N_4400,N_4390,N_4294);
and U4401 (N_4401,N_4279,N_4348);
and U4402 (N_4402,N_4376,N_4258);
nand U4403 (N_4403,N_4296,N_4350);
nand U4404 (N_4404,N_4340,N_4388);
nor U4405 (N_4405,N_4347,N_4267);
and U4406 (N_4406,N_4394,N_4361);
nand U4407 (N_4407,N_4230,N_4215);
xor U4408 (N_4408,N_4327,N_4220);
and U4409 (N_4409,N_4362,N_4249);
nand U4410 (N_4410,N_4236,N_4341);
nor U4411 (N_4411,N_4202,N_4253);
or U4412 (N_4412,N_4268,N_4342);
or U4413 (N_4413,N_4306,N_4235);
nor U4414 (N_4414,N_4336,N_4315);
nor U4415 (N_4415,N_4317,N_4261);
nand U4416 (N_4416,N_4318,N_4262);
nand U4417 (N_4417,N_4324,N_4387);
or U4418 (N_4418,N_4397,N_4239);
xor U4419 (N_4419,N_4223,N_4365);
or U4420 (N_4420,N_4329,N_4281);
and U4421 (N_4421,N_4382,N_4240);
nand U4422 (N_4422,N_4391,N_4287);
and U4423 (N_4423,N_4205,N_4290);
nor U4424 (N_4424,N_4373,N_4251);
xor U4425 (N_4425,N_4218,N_4266);
nor U4426 (N_4426,N_4201,N_4278);
nor U4427 (N_4427,N_4320,N_4344);
xor U4428 (N_4428,N_4370,N_4386);
and U4429 (N_4429,N_4245,N_4284);
or U4430 (N_4430,N_4305,N_4309);
and U4431 (N_4431,N_4354,N_4204);
nor U4432 (N_4432,N_4207,N_4288);
xnor U4433 (N_4433,N_4285,N_4222);
nor U4434 (N_4434,N_4292,N_4375);
and U4435 (N_4435,N_4300,N_4369);
nand U4436 (N_4436,N_4217,N_4255);
nand U4437 (N_4437,N_4393,N_4367);
and U4438 (N_4438,N_4269,N_4241);
and U4439 (N_4439,N_4203,N_4242);
xnor U4440 (N_4440,N_4323,N_4257);
nand U4441 (N_4441,N_4297,N_4328);
nor U4442 (N_4442,N_4208,N_4228);
nand U4443 (N_4443,N_4247,N_4256);
nor U4444 (N_4444,N_4346,N_4263);
xnor U4445 (N_4445,N_4364,N_4310);
or U4446 (N_4446,N_4276,N_4304);
xor U4447 (N_4447,N_4248,N_4380);
and U4448 (N_4448,N_4334,N_4371);
or U4449 (N_4449,N_4272,N_4211);
xnor U4450 (N_4450,N_4254,N_4232);
xor U4451 (N_4451,N_4312,N_4377);
and U4452 (N_4452,N_4359,N_4384);
and U4453 (N_4453,N_4273,N_4293);
xnor U4454 (N_4454,N_4343,N_4338);
nor U4455 (N_4455,N_4383,N_4396);
nor U4456 (N_4456,N_4252,N_4289);
and U4457 (N_4457,N_4243,N_4358);
xor U4458 (N_4458,N_4385,N_4295);
xnor U4459 (N_4459,N_4234,N_4277);
nor U4460 (N_4460,N_4363,N_4280);
or U4461 (N_4461,N_4283,N_4399);
nor U4462 (N_4462,N_4302,N_4352);
or U4463 (N_4463,N_4206,N_4233);
nor U4464 (N_4464,N_4259,N_4351);
nand U4465 (N_4465,N_4260,N_4291);
or U4466 (N_4466,N_4337,N_4356);
nor U4467 (N_4467,N_4392,N_4286);
or U4468 (N_4468,N_4314,N_4270);
xor U4469 (N_4469,N_4216,N_4246);
or U4470 (N_4470,N_4331,N_4330);
or U4471 (N_4471,N_4298,N_4332);
and U4472 (N_4472,N_4357,N_4282);
or U4473 (N_4473,N_4265,N_4231);
nand U4474 (N_4474,N_4333,N_4303);
nor U4475 (N_4475,N_4299,N_4381);
or U4476 (N_4476,N_4313,N_4374);
nor U4477 (N_4477,N_4250,N_4368);
and U4478 (N_4478,N_4224,N_4210);
and U4479 (N_4479,N_4221,N_4322);
and U4480 (N_4480,N_4238,N_4321);
xnor U4481 (N_4481,N_4372,N_4244);
nand U4482 (N_4482,N_4335,N_4379);
nand U4483 (N_4483,N_4227,N_4355);
xor U4484 (N_4484,N_4237,N_4274);
or U4485 (N_4485,N_4225,N_4319);
xnor U4486 (N_4486,N_4325,N_4271);
or U4487 (N_4487,N_4214,N_4389);
nor U4488 (N_4488,N_4378,N_4345);
xnor U4489 (N_4489,N_4360,N_4311);
xnor U4490 (N_4490,N_4213,N_4308);
nand U4491 (N_4491,N_4366,N_4219);
nand U4492 (N_4492,N_4395,N_4212);
or U4493 (N_4493,N_4353,N_4349);
nand U4494 (N_4494,N_4301,N_4339);
or U4495 (N_4495,N_4200,N_4226);
nor U4496 (N_4496,N_4229,N_4264);
nand U4497 (N_4497,N_4209,N_4326);
or U4498 (N_4498,N_4307,N_4316);
and U4499 (N_4499,N_4398,N_4275);
and U4500 (N_4500,N_4273,N_4261);
nand U4501 (N_4501,N_4379,N_4275);
nand U4502 (N_4502,N_4284,N_4339);
or U4503 (N_4503,N_4375,N_4204);
nand U4504 (N_4504,N_4282,N_4216);
nor U4505 (N_4505,N_4248,N_4265);
nand U4506 (N_4506,N_4215,N_4286);
nand U4507 (N_4507,N_4329,N_4245);
nor U4508 (N_4508,N_4393,N_4275);
xor U4509 (N_4509,N_4360,N_4210);
nand U4510 (N_4510,N_4246,N_4375);
nor U4511 (N_4511,N_4291,N_4369);
nor U4512 (N_4512,N_4255,N_4206);
nand U4513 (N_4513,N_4329,N_4312);
or U4514 (N_4514,N_4212,N_4210);
or U4515 (N_4515,N_4364,N_4241);
or U4516 (N_4516,N_4359,N_4293);
or U4517 (N_4517,N_4277,N_4304);
nor U4518 (N_4518,N_4256,N_4229);
xnor U4519 (N_4519,N_4345,N_4206);
or U4520 (N_4520,N_4268,N_4258);
nor U4521 (N_4521,N_4202,N_4308);
or U4522 (N_4522,N_4307,N_4313);
nor U4523 (N_4523,N_4289,N_4352);
xor U4524 (N_4524,N_4397,N_4369);
or U4525 (N_4525,N_4291,N_4259);
and U4526 (N_4526,N_4296,N_4239);
and U4527 (N_4527,N_4398,N_4345);
or U4528 (N_4528,N_4310,N_4346);
or U4529 (N_4529,N_4269,N_4329);
and U4530 (N_4530,N_4386,N_4354);
nor U4531 (N_4531,N_4250,N_4204);
nor U4532 (N_4532,N_4347,N_4232);
and U4533 (N_4533,N_4313,N_4266);
and U4534 (N_4534,N_4274,N_4214);
xnor U4535 (N_4535,N_4200,N_4344);
xor U4536 (N_4536,N_4308,N_4265);
or U4537 (N_4537,N_4331,N_4358);
nand U4538 (N_4538,N_4377,N_4306);
or U4539 (N_4539,N_4364,N_4213);
xor U4540 (N_4540,N_4338,N_4254);
nor U4541 (N_4541,N_4353,N_4399);
nor U4542 (N_4542,N_4215,N_4279);
nand U4543 (N_4543,N_4258,N_4227);
nor U4544 (N_4544,N_4316,N_4292);
and U4545 (N_4545,N_4372,N_4213);
nor U4546 (N_4546,N_4377,N_4286);
xor U4547 (N_4547,N_4365,N_4276);
and U4548 (N_4548,N_4273,N_4240);
or U4549 (N_4549,N_4395,N_4210);
nand U4550 (N_4550,N_4392,N_4287);
nand U4551 (N_4551,N_4334,N_4201);
or U4552 (N_4552,N_4391,N_4355);
or U4553 (N_4553,N_4363,N_4226);
nor U4554 (N_4554,N_4269,N_4260);
nand U4555 (N_4555,N_4327,N_4362);
or U4556 (N_4556,N_4251,N_4302);
and U4557 (N_4557,N_4308,N_4336);
and U4558 (N_4558,N_4231,N_4358);
and U4559 (N_4559,N_4392,N_4376);
and U4560 (N_4560,N_4207,N_4392);
and U4561 (N_4561,N_4285,N_4317);
nand U4562 (N_4562,N_4221,N_4273);
xor U4563 (N_4563,N_4339,N_4233);
or U4564 (N_4564,N_4200,N_4319);
nand U4565 (N_4565,N_4353,N_4344);
nand U4566 (N_4566,N_4374,N_4261);
or U4567 (N_4567,N_4282,N_4267);
and U4568 (N_4568,N_4309,N_4347);
xnor U4569 (N_4569,N_4331,N_4340);
xnor U4570 (N_4570,N_4310,N_4321);
nand U4571 (N_4571,N_4213,N_4315);
nand U4572 (N_4572,N_4306,N_4352);
or U4573 (N_4573,N_4296,N_4313);
nand U4574 (N_4574,N_4218,N_4347);
xor U4575 (N_4575,N_4248,N_4324);
and U4576 (N_4576,N_4385,N_4310);
and U4577 (N_4577,N_4253,N_4213);
nand U4578 (N_4578,N_4236,N_4390);
nand U4579 (N_4579,N_4293,N_4254);
nand U4580 (N_4580,N_4373,N_4304);
and U4581 (N_4581,N_4379,N_4348);
and U4582 (N_4582,N_4344,N_4363);
or U4583 (N_4583,N_4305,N_4382);
nand U4584 (N_4584,N_4383,N_4262);
nor U4585 (N_4585,N_4286,N_4383);
and U4586 (N_4586,N_4348,N_4267);
or U4587 (N_4587,N_4301,N_4356);
or U4588 (N_4588,N_4343,N_4239);
nand U4589 (N_4589,N_4224,N_4217);
xor U4590 (N_4590,N_4240,N_4296);
and U4591 (N_4591,N_4396,N_4310);
nor U4592 (N_4592,N_4318,N_4336);
xor U4593 (N_4593,N_4358,N_4289);
or U4594 (N_4594,N_4278,N_4248);
xnor U4595 (N_4595,N_4200,N_4270);
and U4596 (N_4596,N_4277,N_4389);
xor U4597 (N_4597,N_4272,N_4348);
xor U4598 (N_4598,N_4202,N_4213);
nor U4599 (N_4599,N_4254,N_4344);
nor U4600 (N_4600,N_4571,N_4400);
and U4601 (N_4601,N_4492,N_4528);
and U4602 (N_4602,N_4413,N_4460);
and U4603 (N_4603,N_4402,N_4496);
nor U4604 (N_4604,N_4423,N_4527);
xor U4605 (N_4605,N_4552,N_4586);
nand U4606 (N_4606,N_4458,N_4559);
nor U4607 (N_4607,N_4462,N_4522);
and U4608 (N_4608,N_4551,N_4549);
nand U4609 (N_4609,N_4599,N_4510);
or U4610 (N_4610,N_4555,N_4450);
xor U4611 (N_4611,N_4419,N_4457);
nand U4612 (N_4612,N_4428,N_4445);
and U4613 (N_4613,N_4524,N_4414);
nand U4614 (N_4614,N_4403,N_4570);
xnor U4615 (N_4615,N_4447,N_4541);
xor U4616 (N_4616,N_4479,N_4515);
or U4617 (N_4617,N_4483,N_4585);
xor U4618 (N_4618,N_4500,N_4540);
xor U4619 (N_4619,N_4480,N_4475);
nor U4620 (N_4620,N_4566,N_4452);
xnor U4621 (N_4621,N_4521,N_4503);
nand U4622 (N_4622,N_4598,N_4514);
nand U4623 (N_4623,N_4487,N_4433);
nor U4624 (N_4624,N_4544,N_4567);
nor U4625 (N_4625,N_4516,N_4553);
or U4626 (N_4626,N_4424,N_4589);
xor U4627 (N_4627,N_4557,N_4554);
nand U4628 (N_4628,N_4578,N_4407);
or U4629 (N_4629,N_4563,N_4550);
and U4630 (N_4630,N_4469,N_4441);
or U4631 (N_4631,N_4468,N_4547);
or U4632 (N_4632,N_4591,N_4584);
or U4633 (N_4633,N_4427,N_4594);
nand U4634 (N_4634,N_4426,N_4512);
xor U4635 (N_4635,N_4471,N_4504);
xnor U4636 (N_4636,N_4558,N_4493);
nand U4637 (N_4637,N_4533,N_4435);
xnor U4638 (N_4638,N_4484,N_4560);
nand U4639 (N_4639,N_4411,N_4459);
nand U4640 (N_4640,N_4587,N_4443);
nor U4641 (N_4641,N_4532,N_4463);
nor U4642 (N_4642,N_4506,N_4530);
nor U4643 (N_4643,N_4431,N_4481);
or U4644 (N_4644,N_4417,N_4434);
xnor U4645 (N_4645,N_4509,N_4491);
and U4646 (N_4646,N_4579,N_4473);
nor U4647 (N_4647,N_4440,N_4499);
or U4648 (N_4648,N_4543,N_4505);
and U4649 (N_4649,N_4454,N_4437);
and U4650 (N_4650,N_4485,N_4456);
or U4651 (N_4651,N_4482,N_4581);
and U4652 (N_4652,N_4507,N_4561);
nand U4653 (N_4653,N_4576,N_4489);
or U4654 (N_4654,N_4474,N_4477);
nor U4655 (N_4655,N_4494,N_4430);
nand U4656 (N_4656,N_4596,N_4476);
nand U4657 (N_4657,N_4467,N_4531);
nand U4658 (N_4658,N_4465,N_4548);
or U4659 (N_4659,N_4588,N_4511);
nand U4660 (N_4660,N_4546,N_4573);
and U4661 (N_4661,N_4446,N_4595);
and U4662 (N_4662,N_4518,N_4451);
nand U4663 (N_4663,N_4535,N_4520);
and U4664 (N_4664,N_4406,N_4490);
and U4665 (N_4665,N_4517,N_4448);
nand U4666 (N_4666,N_4534,N_4575);
and U4667 (N_4667,N_4464,N_4453);
xor U4668 (N_4668,N_4568,N_4409);
and U4669 (N_4669,N_4569,N_4429);
xnor U4670 (N_4670,N_4502,N_4421);
or U4671 (N_4671,N_4495,N_4582);
and U4672 (N_4672,N_4536,N_4537);
nand U4673 (N_4673,N_4410,N_4416);
or U4674 (N_4674,N_4404,N_4442);
nor U4675 (N_4675,N_4538,N_4556);
nand U4676 (N_4676,N_4497,N_4564);
or U4677 (N_4677,N_4519,N_4478);
or U4678 (N_4678,N_4580,N_4401);
and U4679 (N_4679,N_4436,N_4574);
nand U4680 (N_4680,N_4472,N_4444);
or U4681 (N_4681,N_4592,N_4408);
nand U4682 (N_4682,N_4455,N_4418);
nor U4683 (N_4683,N_4523,N_4529);
and U4684 (N_4684,N_4405,N_4542);
xor U4685 (N_4685,N_4412,N_4466);
nor U4686 (N_4686,N_4488,N_4525);
and U4687 (N_4687,N_4425,N_4498);
or U4688 (N_4688,N_4501,N_4432);
xnor U4689 (N_4689,N_4583,N_4565);
xnor U4690 (N_4690,N_4539,N_4562);
nor U4691 (N_4691,N_4438,N_4593);
or U4692 (N_4692,N_4526,N_4513);
nand U4693 (N_4693,N_4486,N_4420);
nor U4694 (N_4694,N_4461,N_4415);
and U4695 (N_4695,N_4597,N_4470);
nor U4696 (N_4696,N_4545,N_4572);
nor U4697 (N_4697,N_4439,N_4449);
nor U4698 (N_4698,N_4422,N_4508);
or U4699 (N_4699,N_4577,N_4590);
nand U4700 (N_4700,N_4552,N_4544);
xor U4701 (N_4701,N_4583,N_4545);
nand U4702 (N_4702,N_4501,N_4495);
and U4703 (N_4703,N_4430,N_4443);
nand U4704 (N_4704,N_4474,N_4597);
and U4705 (N_4705,N_4525,N_4536);
xor U4706 (N_4706,N_4480,N_4525);
or U4707 (N_4707,N_4561,N_4477);
and U4708 (N_4708,N_4400,N_4590);
nand U4709 (N_4709,N_4554,N_4565);
nand U4710 (N_4710,N_4519,N_4531);
and U4711 (N_4711,N_4599,N_4506);
nand U4712 (N_4712,N_4549,N_4493);
xnor U4713 (N_4713,N_4442,N_4503);
nand U4714 (N_4714,N_4420,N_4483);
xnor U4715 (N_4715,N_4476,N_4570);
or U4716 (N_4716,N_4418,N_4545);
nand U4717 (N_4717,N_4405,N_4466);
xnor U4718 (N_4718,N_4402,N_4549);
nor U4719 (N_4719,N_4597,N_4564);
nand U4720 (N_4720,N_4551,N_4436);
and U4721 (N_4721,N_4485,N_4414);
nand U4722 (N_4722,N_4505,N_4510);
nand U4723 (N_4723,N_4526,N_4470);
xnor U4724 (N_4724,N_4497,N_4548);
and U4725 (N_4725,N_4438,N_4540);
and U4726 (N_4726,N_4553,N_4403);
xnor U4727 (N_4727,N_4555,N_4579);
or U4728 (N_4728,N_4473,N_4499);
nor U4729 (N_4729,N_4514,N_4482);
or U4730 (N_4730,N_4490,N_4550);
nor U4731 (N_4731,N_4571,N_4500);
xor U4732 (N_4732,N_4566,N_4572);
or U4733 (N_4733,N_4413,N_4421);
xnor U4734 (N_4734,N_4593,N_4583);
and U4735 (N_4735,N_4518,N_4584);
and U4736 (N_4736,N_4528,N_4584);
and U4737 (N_4737,N_4401,N_4591);
or U4738 (N_4738,N_4489,N_4587);
or U4739 (N_4739,N_4558,N_4588);
nor U4740 (N_4740,N_4498,N_4532);
nor U4741 (N_4741,N_4417,N_4429);
nor U4742 (N_4742,N_4521,N_4524);
or U4743 (N_4743,N_4468,N_4549);
and U4744 (N_4744,N_4500,N_4590);
nand U4745 (N_4745,N_4502,N_4568);
and U4746 (N_4746,N_4432,N_4557);
and U4747 (N_4747,N_4417,N_4509);
and U4748 (N_4748,N_4469,N_4443);
xor U4749 (N_4749,N_4413,N_4527);
xnor U4750 (N_4750,N_4468,N_4502);
nor U4751 (N_4751,N_4505,N_4493);
xor U4752 (N_4752,N_4416,N_4458);
or U4753 (N_4753,N_4581,N_4467);
or U4754 (N_4754,N_4536,N_4508);
or U4755 (N_4755,N_4502,N_4419);
nand U4756 (N_4756,N_4507,N_4556);
nor U4757 (N_4757,N_4457,N_4453);
nor U4758 (N_4758,N_4500,N_4560);
nor U4759 (N_4759,N_4585,N_4490);
xor U4760 (N_4760,N_4436,N_4506);
xnor U4761 (N_4761,N_4439,N_4437);
nand U4762 (N_4762,N_4545,N_4556);
or U4763 (N_4763,N_4510,N_4474);
or U4764 (N_4764,N_4493,N_4572);
or U4765 (N_4765,N_4421,N_4581);
nor U4766 (N_4766,N_4410,N_4589);
and U4767 (N_4767,N_4580,N_4575);
nand U4768 (N_4768,N_4408,N_4591);
xnor U4769 (N_4769,N_4564,N_4478);
and U4770 (N_4770,N_4502,N_4444);
xnor U4771 (N_4771,N_4518,N_4484);
nor U4772 (N_4772,N_4525,N_4404);
and U4773 (N_4773,N_4439,N_4434);
nand U4774 (N_4774,N_4507,N_4479);
and U4775 (N_4775,N_4403,N_4527);
xor U4776 (N_4776,N_4592,N_4500);
nand U4777 (N_4777,N_4418,N_4518);
and U4778 (N_4778,N_4438,N_4494);
or U4779 (N_4779,N_4430,N_4584);
nor U4780 (N_4780,N_4433,N_4551);
and U4781 (N_4781,N_4554,N_4476);
nand U4782 (N_4782,N_4449,N_4408);
nor U4783 (N_4783,N_4446,N_4551);
nand U4784 (N_4784,N_4567,N_4586);
and U4785 (N_4785,N_4528,N_4588);
or U4786 (N_4786,N_4559,N_4423);
xnor U4787 (N_4787,N_4561,N_4453);
nor U4788 (N_4788,N_4596,N_4561);
nor U4789 (N_4789,N_4529,N_4415);
and U4790 (N_4790,N_4471,N_4580);
nand U4791 (N_4791,N_4435,N_4477);
or U4792 (N_4792,N_4523,N_4581);
xor U4793 (N_4793,N_4542,N_4562);
or U4794 (N_4794,N_4512,N_4565);
and U4795 (N_4795,N_4439,N_4539);
or U4796 (N_4796,N_4470,N_4549);
and U4797 (N_4797,N_4406,N_4408);
nand U4798 (N_4798,N_4566,N_4407);
xor U4799 (N_4799,N_4598,N_4489);
and U4800 (N_4800,N_4728,N_4724);
nor U4801 (N_4801,N_4613,N_4797);
xor U4802 (N_4802,N_4693,N_4717);
xnor U4803 (N_4803,N_4622,N_4783);
or U4804 (N_4804,N_4705,N_4652);
nor U4805 (N_4805,N_4644,N_4642);
nor U4806 (N_4806,N_4645,N_4711);
xnor U4807 (N_4807,N_4625,N_4630);
xor U4808 (N_4808,N_4757,N_4621);
nor U4809 (N_4809,N_4703,N_4730);
nand U4810 (N_4810,N_4754,N_4742);
nand U4811 (N_4811,N_4773,N_4765);
or U4812 (N_4812,N_4637,N_4792);
and U4813 (N_4813,N_4736,N_4780);
xnor U4814 (N_4814,N_4658,N_4688);
xor U4815 (N_4815,N_4603,N_4734);
and U4816 (N_4816,N_4704,N_4627);
or U4817 (N_4817,N_4682,N_4798);
or U4818 (N_4818,N_4666,N_4737);
or U4819 (N_4819,N_4660,N_4782);
or U4820 (N_4820,N_4692,N_4675);
or U4821 (N_4821,N_4731,N_4710);
and U4822 (N_4822,N_4752,N_4691);
nor U4823 (N_4823,N_4775,N_4657);
nor U4824 (N_4824,N_4733,N_4680);
or U4825 (N_4825,N_4795,N_4655);
and U4826 (N_4826,N_4701,N_4651);
nand U4827 (N_4827,N_4776,N_4612);
and U4828 (N_4828,N_4722,N_4764);
nand U4829 (N_4829,N_4611,N_4650);
nand U4830 (N_4830,N_4709,N_4661);
nor U4831 (N_4831,N_4667,N_4602);
nand U4832 (N_4832,N_4656,N_4636);
or U4833 (N_4833,N_4609,N_4696);
nand U4834 (N_4834,N_4756,N_4659);
nor U4835 (N_4835,N_4649,N_4623);
nand U4836 (N_4836,N_4605,N_4790);
and U4837 (N_4837,N_4760,N_4647);
xnor U4838 (N_4838,N_4787,N_4715);
and U4839 (N_4839,N_4740,N_4750);
nand U4840 (N_4840,N_4683,N_4723);
nand U4841 (N_4841,N_4713,N_4654);
and U4842 (N_4842,N_4600,N_4706);
nor U4843 (N_4843,N_4772,N_4665);
nor U4844 (N_4844,N_4629,N_4751);
nand U4845 (N_4845,N_4759,N_4727);
and U4846 (N_4846,N_4628,N_4671);
nor U4847 (N_4847,N_4699,N_4771);
and U4848 (N_4848,N_4672,N_4674);
nor U4849 (N_4849,N_4668,N_4746);
nor U4850 (N_4850,N_4662,N_4770);
nor U4851 (N_4851,N_4690,N_4639);
or U4852 (N_4852,N_4604,N_4633);
nand U4853 (N_4853,N_4689,N_4778);
or U4854 (N_4854,N_4763,N_4606);
or U4855 (N_4855,N_4615,N_4747);
xnor U4856 (N_4856,N_4748,N_4753);
nand U4857 (N_4857,N_4617,N_4624);
xor U4858 (N_4858,N_4762,N_4694);
or U4859 (N_4859,N_4631,N_4726);
or U4860 (N_4860,N_4608,N_4745);
xnor U4861 (N_4861,N_4786,N_4610);
nor U4862 (N_4862,N_4784,N_4673);
nor U4863 (N_4863,N_4702,N_4601);
xor U4864 (N_4864,N_4677,N_4768);
xor U4865 (N_4865,N_4788,N_4669);
and U4866 (N_4866,N_4641,N_4719);
xor U4867 (N_4867,N_4695,N_4697);
or U4868 (N_4868,N_4758,N_4676);
nor U4869 (N_4869,N_4619,N_4769);
or U4870 (N_4870,N_4626,N_4721);
nand U4871 (N_4871,N_4681,N_4791);
nor U4872 (N_4872,N_4761,N_4712);
xor U4873 (N_4873,N_4714,N_4766);
and U4874 (N_4874,N_4678,N_4685);
nor U4875 (N_4875,N_4684,N_4781);
nor U4876 (N_4876,N_4799,N_4720);
and U4877 (N_4877,N_4744,N_4632);
nand U4878 (N_4878,N_4638,N_4725);
nor U4879 (N_4879,N_4732,N_4738);
and U4880 (N_4880,N_4687,N_4718);
and U4881 (N_4881,N_4749,N_4698);
xnor U4882 (N_4882,N_4634,N_4793);
or U4883 (N_4883,N_4741,N_4796);
nor U4884 (N_4884,N_4653,N_4716);
nand U4885 (N_4885,N_4664,N_4614);
or U4886 (N_4886,N_4785,N_4743);
or U4887 (N_4887,N_4794,N_4607);
or U4888 (N_4888,N_4640,N_4739);
xor U4889 (N_4889,N_4729,N_4618);
nor U4890 (N_4890,N_4774,N_4663);
xor U4891 (N_4891,N_4735,N_4670);
or U4892 (N_4892,N_4686,N_4646);
nand U4893 (N_4893,N_4767,N_4643);
nand U4894 (N_4894,N_4777,N_4700);
nand U4895 (N_4895,N_4648,N_4789);
and U4896 (N_4896,N_4679,N_4616);
and U4897 (N_4897,N_4708,N_4755);
nand U4898 (N_4898,N_4707,N_4635);
nand U4899 (N_4899,N_4620,N_4779);
and U4900 (N_4900,N_4726,N_4611);
or U4901 (N_4901,N_4755,N_4775);
or U4902 (N_4902,N_4612,N_4779);
nand U4903 (N_4903,N_4623,N_4738);
or U4904 (N_4904,N_4678,N_4666);
nor U4905 (N_4905,N_4742,N_4705);
and U4906 (N_4906,N_4715,N_4690);
and U4907 (N_4907,N_4772,N_4747);
xor U4908 (N_4908,N_4748,N_4671);
and U4909 (N_4909,N_4728,N_4731);
or U4910 (N_4910,N_4688,N_4771);
xor U4911 (N_4911,N_4784,N_4628);
or U4912 (N_4912,N_4624,N_4735);
nand U4913 (N_4913,N_4608,N_4722);
xnor U4914 (N_4914,N_4683,N_4648);
nor U4915 (N_4915,N_4769,N_4639);
or U4916 (N_4916,N_4775,N_4732);
or U4917 (N_4917,N_4613,N_4760);
and U4918 (N_4918,N_4612,N_4699);
and U4919 (N_4919,N_4749,N_4600);
xor U4920 (N_4920,N_4621,N_4772);
and U4921 (N_4921,N_4777,N_4790);
nand U4922 (N_4922,N_4757,N_4707);
and U4923 (N_4923,N_4665,N_4668);
and U4924 (N_4924,N_4609,N_4630);
nor U4925 (N_4925,N_4684,N_4637);
xnor U4926 (N_4926,N_4649,N_4689);
and U4927 (N_4927,N_4701,N_4675);
nand U4928 (N_4928,N_4776,N_4739);
or U4929 (N_4929,N_4706,N_4719);
or U4930 (N_4930,N_4768,N_4601);
xnor U4931 (N_4931,N_4669,N_4659);
nor U4932 (N_4932,N_4793,N_4765);
xor U4933 (N_4933,N_4742,N_4793);
nor U4934 (N_4934,N_4658,N_4682);
or U4935 (N_4935,N_4666,N_4768);
and U4936 (N_4936,N_4768,N_4631);
nand U4937 (N_4937,N_4786,N_4607);
and U4938 (N_4938,N_4711,N_4747);
nand U4939 (N_4939,N_4724,N_4691);
nor U4940 (N_4940,N_4687,N_4659);
nand U4941 (N_4941,N_4780,N_4798);
nand U4942 (N_4942,N_4779,N_4627);
nor U4943 (N_4943,N_4644,N_4669);
nand U4944 (N_4944,N_4602,N_4650);
xnor U4945 (N_4945,N_4708,N_4727);
or U4946 (N_4946,N_4605,N_4702);
nor U4947 (N_4947,N_4658,N_4624);
and U4948 (N_4948,N_4634,N_4711);
xor U4949 (N_4949,N_4724,N_4664);
xnor U4950 (N_4950,N_4771,N_4700);
xor U4951 (N_4951,N_4630,N_4602);
nand U4952 (N_4952,N_4728,N_4746);
and U4953 (N_4953,N_4623,N_4710);
and U4954 (N_4954,N_4620,N_4648);
nand U4955 (N_4955,N_4719,N_4783);
or U4956 (N_4956,N_4792,N_4626);
or U4957 (N_4957,N_4767,N_4600);
nand U4958 (N_4958,N_4694,N_4630);
nand U4959 (N_4959,N_4673,N_4735);
xnor U4960 (N_4960,N_4744,N_4662);
nand U4961 (N_4961,N_4673,N_4743);
and U4962 (N_4962,N_4620,N_4661);
xor U4963 (N_4963,N_4637,N_4765);
and U4964 (N_4964,N_4736,N_4663);
nand U4965 (N_4965,N_4633,N_4753);
xnor U4966 (N_4966,N_4647,N_4764);
or U4967 (N_4967,N_4770,N_4696);
nor U4968 (N_4968,N_4693,N_4753);
xnor U4969 (N_4969,N_4710,N_4620);
nand U4970 (N_4970,N_4665,N_4780);
xor U4971 (N_4971,N_4729,N_4725);
nand U4972 (N_4972,N_4612,N_4757);
nand U4973 (N_4973,N_4743,N_4675);
nand U4974 (N_4974,N_4632,N_4678);
and U4975 (N_4975,N_4615,N_4760);
or U4976 (N_4976,N_4633,N_4708);
nor U4977 (N_4977,N_4645,N_4670);
nor U4978 (N_4978,N_4670,N_4740);
and U4979 (N_4979,N_4640,N_4649);
nand U4980 (N_4980,N_4726,N_4765);
nand U4981 (N_4981,N_4709,N_4710);
nand U4982 (N_4982,N_4663,N_4646);
xor U4983 (N_4983,N_4614,N_4702);
and U4984 (N_4984,N_4706,N_4733);
or U4985 (N_4985,N_4696,N_4760);
nor U4986 (N_4986,N_4656,N_4644);
nor U4987 (N_4987,N_4655,N_4668);
nor U4988 (N_4988,N_4728,N_4604);
or U4989 (N_4989,N_4794,N_4723);
or U4990 (N_4990,N_4637,N_4621);
nand U4991 (N_4991,N_4710,N_4674);
xnor U4992 (N_4992,N_4615,N_4668);
nor U4993 (N_4993,N_4638,N_4699);
and U4994 (N_4994,N_4775,N_4787);
and U4995 (N_4995,N_4778,N_4688);
and U4996 (N_4996,N_4718,N_4647);
xor U4997 (N_4997,N_4796,N_4601);
and U4998 (N_4998,N_4659,N_4635);
nor U4999 (N_4999,N_4778,N_4649);
nand U5000 (N_5000,N_4839,N_4977);
nor U5001 (N_5001,N_4956,N_4818);
nor U5002 (N_5002,N_4937,N_4985);
xnor U5003 (N_5003,N_4935,N_4810);
or U5004 (N_5004,N_4885,N_4915);
xor U5005 (N_5005,N_4948,N_4876);
xnor U5006 (N_5006,N_4934,N_4833);
xor U5007 (N_5007,N_4815,N_4894);
and U5008 (N_5008,N_4846,N_4866);
nand U5009 (N_5009,N_4832,N_4962);
xor U5010 (N_5010,N_4931,N_4857);
nor U5011 (N_5011,N_4851,N_4946);
nor U5012 (N_5012,N_4979,N_4825);
and U5013 (N_5013,N_4940,N_4871);
and U5014 (N_5014,N_4995,N_4837);
xor U5015 (N_5015,N_4865,N_4801);
nand U5016 (N_5016,N_4811,N_4838);
or U5017 (N_5017,N_4941,N_4921);
nor U5018 (N_5018,N_4884,N_4972);
xor U5019 (N_5019,N_4895,N_4889);
xor U5020 (N_5020,N_4997,N_4848);
nand U5021 (N_5021,N_4953,N_4812);
and U5022 (N_5022,N_4869,N_4945);
and U5023 (N_5023,N_4904,N_4873);
xor U5024 (N_5024,N_4844,N_4809);
or U5025 (N_5025,N_4878,N_4847);
xor U5026 (N_5026,N_4969,N_4887);
nand U5027 (N_5027,N_4827,N_4918);
or U5028 (N_5028,N_4888,N_4830);
xnor U5029 (N_5029,N_4944,N_4881);
nor U5030 (N_5030,N_4978,N_4989);
and U5031 (N_5031,N_4882,N_4808);
or U5032 (N_5032,N_4816,N_4968);
or U5033 (N_5033,N_4843,N_4919);
or U5034 (N_5034,N_4817,N_4870);
nor U5035 (N_5035,N_4982,N_4981);
nor U5036 (N_5036,N_4975,N_4903);
or U5037 (N_5037,N_4858,N_4988);
and U5038 (N_5038,N_4917,N_4883);
xor U5039 (N_5039,N_4928,N_4983);
or U5040 (N_5040,N_4823,N_4892);
or U5041 (N_5041,N_4987,N_4834);
xor U5042 (N_5042,N_4856,N_4958);
nor U5043 (N_5043,N_4829,N_4850);
nor U5044 (N_5044,N_4853,N_4831);
nand U5045 (N_5045,N_4893,N_4936);
or U5046 (N_5046,N_4899,N_4820);
and U5047 (N_5047,N_4971,N_4932);
and U5048 (N_5048,N_4994,N_4993);
nor U5049 (N_5049,N_4841,N_4957);
xnor U5050 (N_5050,N_4901,N_4891);
nor U5051 (N_5051,N_4942,N_4947);
or U5052 (N_5052,N_4867,N_4986);
and U5053 (N_5053,N_4933,N_4807);
or U5054 (N_5054,N_4926,N_4907);
nand U5055 (N_5055,N_4970,N_4999);
nor U5056 (N_5056,N_4802,N_4880);
and U5057 (N_5057,N_4805,N_4821);
nand U5058 (N_5058,N_4992,N_4973);
xor U5059 (N_5059,N_4960,N_4991);
nand U5060 (N_5060,N_4949,N_4961);
nor U5061 (N_5061,N_4842,N_4912);
nor U5062 (N_5062,N_4840,N_4852);
or U5063 (N_5063,N_4913,N_4900);
xor U5064 (N_5064,N_4860,N_4898);
and U5065 (N_5065,N_4864,N_4855);
nand U5066 (N_5066,N_4954,N_4939);
nor U5067 (N_5067,N_4862,N_4925);
and U5068 (N_5068,N_4911,N_4861);
or U5069 (N_5069,N_4819,N_4826);
nand U5070 (N_5070,N_4890,N_4951);
nor U5071 (N_5071,N_4872,N_4950);
nor U5072 (N_5072,N_4943,N_4875);
nor U5073 (N_5073,N_4976,N_4905);
xnor U5074 (N_5074,N_4952,N_4984);
and U5075 (N_5075,N_4980,N_4849);
nand U5076 (N_5076,N_4906,N_4938);
and U5077 (N_5077,N_4965,N_4908);
nor U5078 (N_5078,N_4886,N_4877);
xor U5079 (N_5079,N_4824,N_4963);
or U5080 (N_5080,N_4806,N_4924);
nor U5081 (N_5081,N_4896,N_4916);
nand U5082 (N_5082,N_4974,N_4835);
or U5083 (N_5083,N_4996,N_4927);
xnor U5084 (N_5084,N_4813,N_4955);
nor U5085 (N_5085,N_4922,N_4800);
nor U5086 (N_5086,N_4828,N_4910);
nor U5087 (N_5087,N_4920,N_4914);
nor U5088 (N_5088,N_4967,N_4814);
nand U5089 (N_5089,N_4879,N_4990);
nand U5090 (N_5090,N_4923,N_4868);
nor U5091 (N_5091,N_4803,N_4909);
nor U5092 (N_5092,N_4845,N_4822);
nand U5093 (N_5093,N_4859,N_4902);
nand U5094 (N_5094,N_4998,N_4966);
nand U5095 (N_5095,N_4930,N_4897);
nand U5096 (N_5096,N_4874,N_4854);
nand U5097 (N_5097,N_4964,N_4863);
nor U5098 (N_5098,N_4959,N_4804);
xor U5099 (N_5099,N_4836,N_4929);
and U5100 (N_5100,N_4927,N_4864);
nand U5101 (N_5101,N_4823,N_4862);
and U5102 (N_5102,N_4829,N_4923);
nand U5103 (N_5103,N_4842,N_4942);
and U5104 (N_5104,N_4913,N_4942);
xor U5105 (N_5105,N_4924,N_4929);
nor U5106 (N_5106,N_4814,N_4986);
nand U5107 (N_5107,N_4875,N_4960);
xnor U5108 (N_5108,N_4960,N_4901);
nand U5109 (N_5109,N_4884,N_4896);
xor U5110 (N_5110,N_4978,N_4876);
and U5111 (N_5111,N_4974,N_4826);
nor U5112 (N_5112,N_4942,N_4870);
nand U5113 (N_5113,N_4958,N_4880);
and U5114 (N_5114,N_4937,N_4840);
xor U5115 (N_5115,N_4976,N_4921);
xnor U5116 (N_5116,N_4825,N_4874);
and U5117 (N_5117,N_4991,N_4938);
nor U5118 (N_5118,N_4895,N_4892);
xor U5119 (N_5119,N_4937,N_4969);
nand U5120 (N_5120,N_4850,N_4972);
nand U5121 (N_5121,N_4986,N_4895);
nor U5122 (N_5122,N_4969,N_4822);
and U5123 (N_5123,N_4991,N_4945);
nor U5124 (N_5124,N_4844,N_4853);
and U5125 (N_5125,N_4974,N_4864);
nor U5126 (N_5126,N_4846,N_4815);
and U5127 (N_5127,N_4926,N_4929);
or U5128 (N_5128,N_4896,N_4811);
or U5129 (N_5129,N_4980,N_4976);
xnor U5130 (N_5130,N_4938,N_4852);
and U5131 (N_5131,N_4841,N_4868);
or U5132 (N_5132,N_4926,N_4811);
xor U5133 (N_5133,N_4912,N_4818);
nand U5134 (N_5134,N_4829,N_4972);
xnor U5135 (N_5135,N_4910,N_4874);
nor U5136 (N_5136,N_4990,N_4891);
nand U5137 (N_5137,N_4856,N_4985);
xor U5138 (N_5138,N_4886,N_4922);
and U5139 (N_5139,N_4912,N_4976);
or U5140 (N_5140,N_4908,N_4861);
nand U5141 (N_5141,N_4876,N_4940);
nand U5142 (N_5142,N_4857,N_4947);
xnor U5143 (N_5143,N_4897,N_4828);
and U5144 (N_5144,N_4964,N_4928);
nor U5145 (N_5145,N_4899,N_4994);
or U5146 (N_5146,N_4995,N_4905);
xor U5147 (N_5147,N_4991,N_4912);
or U5148 (N_5148,N_4971,N_4924);
or U5149 (N_5149,N_4868,N_4803);
nor U5150 (N_5150,N_4879,N_4938);
or U5151 (N_5151,N_4900,N_4800);
xor U5152 (N_5152,N_4967,N_4969);
nor U5153 (N_5153,N_4954,N_4891);
nor U5154 (N_5154,N_4959,N_4943);
nand U5155 (N_5155,N_4856,N_4905);
and U5156 (N_5156,N_4933,N_4971);
or U5157 (N_5157,N_4803,N_4892);
xnor U5158 (N_5158,N_4839,N_4801);
nor U5159 (N_5159,N_4834,N_4862);
or U5160 (N_5160,N_4885,N_4973);
xor U5161 (N_5161,N_4837,N_4890);
and U5162 (N_5162,N_4866,N_4893);
xor U5163 (N_5163,N_4804,N_4812);
and U5164 (N_5164,N_4819,N_4890);
and U5165 (N_5165,N_4820,N_4892);
nand U5166 (N_5166,N_4823,N_4983);
xor U5167 (N_5167,N_4893,N_4943);
nand U5168 (N_5168,N_4854,N_4836);
and U5169 (N_5169,N_4808,N_4917);
nor U5170 (N_5170,N_4943,N_4812);
and U5171 (N_5171,N_4804,N_4856);
and U5172 (N_5172,N_4923,N_4897);
or U5173 (N_5173,N_4828,N_4909);
or U5174 (N_5174,N_4879,N_4839);
xor U5175 (N_5175,N_4982,N_4885);
xor U5176 (N_5176,N_4937,N_4813);
or U5177 (N_5177,N_4863,N_4859);
nand U5178 (N_5178,N_4808,N_4908);
nand U5179 (N_5179,N_4951,N_4922);
nand U5180 (N_5180,N_4967,N_4980);
or U5181 (N_5181,N_4986,N_4982);
or U5182 (N_5182,N_4939,N_4856);
and U5183 (N_5183,N_4865,N_4876);
xnor U5184 (N_5184,N_4819,N_4945);
or U5185 (N_5185,N_4831,N_4973);
xnor U5186 (N_5186,N_4862,N_4983);
and U5187 (N_5187,N_4884,N_4823);
and U5188 (N_5188,N_4976,N_4838);
nor U5189 (N_5189,N_4858,N_4901);
nand U5190 (N_5190,N_4832,N_4819);
xnor U5191 (N_5191,N_4860,N_4851);
xnor U5192 (N_5192,N_4961,N_4980);
nand U5193 (N_5193,N_4994,N_4997);
nor U5194 (N_5194,N_4992,N_4804);
or U5195 (N_5195,N_4930,N_4873);
nand U5196 (N_5196,N_4846,N_4997);
nor U5197 (N_5197,N_4805,N_4845);
nand U5198 (N_5198,N_4812,N_4832);
nand U5199 (N_5199,N_4841,N_4924);
nand U5200 (N_5200,N_5084,N_5066);
nor U5201 (N_5201,N_5141,N_5068);
nor U5202 (N_5202,N_5067,N_5086);
nand U5203 (N_5203,N_5000,N_5128);
nor U5204 (N_5204,N_5162,N_5168);
and U5205 (N_5205,N_5112,N_5182);
or U5206 (N_5206,N_5126,N_5058);
or U5207 (N_5207,N_5070,N_5136);
nor U5208 (N_5208,N_5073,N_5119);
nand U5209 (N_5209,N_5163,N_5090);
nor U5210 (N_5210,N_5094,N_5181);
and U5211 (N_5211,N_5172,N_5150);
or U5212 (N_5212,N_5178,N_5046);
or U5213 (N_5213,N_5075,N_5038);
xor U5214 (N_5214,N_5191,N_5185);
or U5215 (N_5215,N_5034,N_5044);
or U5216 (N_5216,N_5171,N_5199);
xor U5217 (N_5217,N_5057,N_5098);
or U5218 (N_5218,N_5133,N_5151);
nand U5219 (N_5219,N_5147,N_5180);
nand U5220 (N_5220,N_5155,N_5145);
or U5221 (N_5221,N_5148,N_5134);
nor U5222 (N_5222,N_5174,N_5161);
and U5223 (N_5223,N_5124,N_5158);
nand U5224 (N_5224,N_5184,N_5129);
and U5225 (N_5225,N_5096,N_5011);
or U5226 (N_5226,N_5052,N_5135);
nor U5227 (N_5227,N_5117,N_5104);
and U5228 (N_5228,N_5153,N_5010);
nand U5229 (N_5229,N_5054,N_5077);
xnor U5230 (N_5230,N_5197,N_5087);
xor U5231 (N_5231,N_5079,N_5101);
or U5232 (N_5232,N_5027,N_5091);
xor U5233 (N_5233,N_5173,N_5015);
and U5234 (N_5234,N_5029,N_5007);
nor U5235 (N_5235,N_5144,N_5021);
xnor U5236 (N_5236,N_5118,N_5022);
nor U5237 (N_5237,N_5009,N_5127);
nand U5238 (N_5238,N_5059,N_5140);
nor U5239 (N_5239,N_5092,N_5024);
nand U5240 (N_5240,N_5005,N_5045);
xnor U5241 (N_5241,N_5016,N_5142);
nand U5242 (N_5242,N_5165,N_5072);
or U5243 (N_5243,N_5008,N_5063);
and U5244 (N_5244,N_5049,N_5138);
or U5245 (N_5245,N_5196,N_5189);
or U5246 (N_5246,N_5107,N_5019);
nor U5247 (N_5247,N_5120,N_5111);
nor U5248 (N_5248,N_5047,N_5193);
xnor U5249 (N_5249,N_5042,N_5179);
nor U5250 (N_5250,N_5139,N_5035);
nor U5251 (N_5251,N_5017,N_5152);
or U5252 (N_5252,N_5025,N_5160);
nand U5253 (N_5253,N_5083,N_5146);
nor U5254 (N_5254,N_5082,N_5095);
xnor U5255 (N_5255,N_5100,N_5061);
nand U5256 (N_5256,N_5004,N_5078);
and U5257 (N_5257,N_5065,N_5037);
nor U5258 (N_5258,N_5137,N_5166);
xor U5259 (N_5259,N_5169,N_5114);
nor U5260 (N_5260,N_5113,N_5041);
nor U5261 (N_5261,N_5093,N_5051);
nor U5262 (N_5262,N_5060,N_5192);
nand U5263 (N_5263,N_5187,N_5050);
and U5264 (N_5264,N_5177,N_5186);
nand U5265 (N_5265,N_5014,N_5033);
and U5266 (N_5266,N_5183,N_5088);
and U5267 (N_5267,N_5110,N_5143);
or U5268 (N_5268,N_5125,N_5164);
nor U5269 (N_5269,N_5020,N_5188);
xnor U5270 (N_5270,N_5028,N_5089);
nor U5271 (N_5271,N_5003,N_5039);
nand U5272 (N_5272,N_5099,N_5159);
and U5273 (N_5273,N_5115,N_5056);
and U5274 (N_5274,N_5175,N_5102);
or U5275 (N_5275,N_5176,N_5030);
xor U5276 (N_5276,N_5130,N_5018);
xor U5277 (N_5277,N_5167,N_5062);
nor U5278 (N_5278,N_5123,N_5076);
nand U5279 (N_5279,N_5043,N_5001);
and U5280 (N_5280,N_5108,N_5132);
or U5281 (N_5281,N_5031,N_5080);
and U5282 (N_5282,N_5156,N_5040);
and U5283 (N_5283,N_5032,N_5122);
or U5284 (N_5284,N_5109,N_5170);
xnor U5285 (N_5285,N_5023,N_5053);
xor U5286 (N_5286,N_5116,N_5002);
xnor U5287 (N_5287,N_5012,N_5036);
and U5288 (N_5288,N_5154,N_5105);
or U5289 (N_5289,N_5106,N_5055);
or U5290 (N_5290,N_5026,N_5006);
nor U5291 (N_5291,N_5157,N_5121);
nor U5292 (N_5292,N_5198,N_5103);
xor U5293 (N_5293,N_5081,N_5097);
or U5294 (N_5294,N_5071,N_5190);
and U5295 (N_5295,N_5074,N_5013);
nor U5296 (N_5296,N_5131,N_5195);
xnor U5297 (N_5297,N_5069,N_5149);
xnor U5298 (N_5298,N_5048,N_5064);
and U5299 (N_5299,N_5194,N_5085);
or U5300 (N_5300,N_5184,N_5006);
and U5301 (N_5301,N_5058,N_5165);
nand U5302 (N_5302,N_5027,N_5110);
xnor U5303 (N_5303,N_5053,N_5190);
nor U5304 (N_5304,N_5125,N_5149);
xor U5305 (N_5305,N_5047,N_5151);
nor U5306 (N_5306,N_5180,N_5198);
nor U5307 (N_5307,N_5033,N_5176);
xnor U5308 (N_5308,N_5034,N_5126);
xor U5309 (N_5309,N_5106,N_5135);
xor U5310 (N_5310,N_5147,N_5046);
xnor U5311 (N_5311,N_5178,N_5039);
nand U5312 (N_5312,N_5145,N_5050);
nor U5313 (N_5313,N_5033,N_5072);
xor U5314 (N_5314,N_5076,N_5101);
or U5315 (N_5315,N_5059,N_5196);
xor U5316 (N_5316,N_5084,N_5057);
xnor U5317 (N_5317,N_5197,N_5041);
or U5318 (N_5318,N_5090,N_5108);
nor U5319 (N_5319,N_5026,N_5082);
or U5320 (N_5320,N_5011,N_5010);
and U5321 (N_5321,N_5059,N_5013);
and U5322 (N_5322,N_5008,N_5188);
or U5323 (N_5323,N_5193,N_5126);
xor U5324 (N_5324,N_5030,N_5135);
and U5325 (N_5325,N_5125,N_5097);
nand U5326 (N_5326,N_5063,N_5004);
and U5327 (N_5327,N_5166,N_5159);
or U5328 (N_5328,N_5152,N_5052);
and U5329 (N_5329,N_5105,N_5044);
xor U5330 (N_5330,N_5158,N_5030);
nor U5331 (N_5331,N_5039,N_5030);
or U5332 (N_5332,N_5122,N_5049);
or U5333 (N_5333,N_5152,N_5078);
nand U5334 (N_5334,N_5130,N_5116);
xor U5335 (N_5335,N_5023,N_5178);
nor U5336 (N_5336,N_5080,N_5131);
or U5337 (N_5337,N_5037,N_5060);
xnor U5338 (N_5338,N_5086,N_5049);
xor U5339 (N_5339,N_5173,N_5056);
nor U5340 (N_5340,N_5198,N_5176);
and U5341 (N_5341,N_5089,N_5151);
or U5342 (N_5342,N_5169,N_5194);
nand U5343 (N_5343,N_5112,N_5017);
and U5344 (N_5344,N_5088,N_5049);
nand U5345 (N_5345,N_5105,N_5109);
nand U5346 (N_5346,N_5155,N_5088);
and U5347 (N_5347,N_5040,N_5185);
nor U5348 (N_5348,N_5123,N_5073);
nor U5349 (N_5349,N_5053,N_5042);
xnor U5350 (N_5350,N_5092,N_5134);
xor U5351 (N_5351,N_5192,N_5111);
nor U5352 (N_5352,N_5104,N_5012);
or U5353 (N_5353,N_5037,N_5141);
nor U5354 (N_5354,N_5193,N_5042);
xor U5355 (N_5355,N_5101,N_5004);
nand U5356 (N_5356,N_5012,N_5122);
or U5357 (N_5357,N_5104,N_5195);
or U5358 (N_5358,N_5055,N_5026);
nor U5359 (N_5359,N_5120,N_5009);
or U5360 (N_5360,N_5054,N_5045);
nand U5361 (N_5361,N_5130,N_5026);
or U5362 (N_5362,N_5171,N_5022);
and U5363 (N_5363,N_5137,N_5169);
and U5364 (N_5364,N_5080,N_5183);
xnor U5365 (N_5365,N_5030,N_5008);
and U5366 (N_5366,N_5155,N_5157);
and U5367 (N_5367,N_5074,N_5010);
nor U5368 (N_5368,N_5042,N_5110);
xor U5369 (N_5369,N_5121,N_5021);
and U5370 (N_5370,N_5156,N_5049);
xnor U5371 (N_5371,N_5061,N_5010);
xor U5372 (N_5372,N_5009,N_5027);
or U5373 (N_5373,N_5089,N_5059);
nand U5374 (N_5374,N_5167,N_5057);
xor U5375 (N_5375,N_5002,N_5182);
nand U5376 (N_5376,N_5161,N_5076);
or U5377 (N_5377,N_5026,N_5117);
nand U5378 (N_5378,N_5162,N_5060);
xor U5379 (N_5379,N_5131,N_5190);
or U5380 (N_5380,N_5142,N_5035);
or U5381 (N_5381,N_5069,N_5062);
nor U5382 (N_5382,N_5055,N_5198);
xnor U5383 (N_5383,N_5150,N_5157);
nand U5384 (N_5384,N_5197,N_5075);
nor U5385 (N_5385,N_5048,N_5159);
xor U5386 (N_5386,N_5145,N_5172);
nand U5387 (N_5387,N_5160,N_5060);
xor U5388 (N_5388,N_5012,N_5171);
nor U5389 (N_5389,N_5164,N_5099);
xor U5390 (N_5390,N_5132,N_5023);
or U5391 (N_5391,N_5091,N_5196);
or U5392 (N_5392,N_5014,N_5008);
nor U5393 (N_5393,N_5033,N_5093);
or U5394 (N_5394,N_5172,N_5128);
or U5395 (N_5395,N_5044,N_5061);
or U5396 (N_5396,N_5056,N_5185);
or U5397 (N_5397,N_5116,N_5021);
xor U5398 (N_5398,N_5056,N_5086);
nor U5399 (N_5399,N_5005,N_5003);
or U5400 (N_5400,N_5377,N_5218);
and U5401 (N_5401,N_5301,N_5293);
and U5402 (N_5402,N_5336,N_5298);
nand U5403 (N_5403,N_5369,N_5323);
xor U5404 (N_5404,N_5292,N_5287);
xnor U5405 (N_5405,N_5355,N_5272);
nand U5406 (N_5406,N_5263,N_5212);
or U5407 (N_5407,N_5357,N_5279);
and U5408 (N_5408,N_5219,N_5305);
nor U5409 (N_5409,N_5278,N_5393);
or U5410 (N_5410,N_5353,N_5349);
xor U5411 (N_5411,N_5335,N_5379);
nor U5412 (N_5412,N_5259,N_5216);
nand U5413 (N_5413,N_5362,N_5304);
or U5414 (N_5414,N_5237,N_5289);
and U5415 (N_5415,N_5230,N_5367);
and U5416 (N_5416,N_5344,N_5217);
nand U5417 (N_5417,N_5275,N_5329);
nand U5418 (N_5418,N_5324,N_5284);
and U5419 (N_5419,N_5375,N_5372);
nand U5420 (N_5420,N_5249,N_5392);
or U5421 (N_5421,N_5331,N_5211);
xnor U5422 (N_5422,N_5226,N_5229);
xor U5423 (N_5423,N_5232,N_5273);
xnor U5424 (N_5424,N_5389,N_5370);
xor U5425 (N_5425,N_5363,N_5397);
xnor U5426 (N_5426,N_5347,N_5281);
and U5427 (N_5427,N_5398,N_5383);
and U5428 (N_5428,N_5277,N_5319);
and U5429 (N_5429,N_5310,N_5339);
and U5430 (N_5430,N_5228,N_5322);
nor U5431 (N_5431,N_5356,N_5387);
and U5432 (N_5432,N_5235,N_5303);
and U5433 (N_5433,N_5245,N_5286);
nand U5434 (N_5434,N_5334,N_5280);
or U5435 (N_5435,N_5296,N_5343);
nand U5436 (N_5436,N_5358,N_5200);
and U5437 (N_5437,N_5208,N_5290);
nor U5438 (N_5438,N_5233,N_5246);
and U5439 (N_5439,N_5396,N_5224);
xnor U5440 (N_5440,N_5271,N_5382);
or U5441 (N_5441,N_5395,N_5257);
and U5442 (N_5442,N_5210,N_5316);
nand U5443 (N_5443,N_5205,N_5307);
nand U5444 (N_5444,N_5352,N_5297);
or U5445 (N_5445,N_5328,N_5381);
xnor U5446 (N_5446,N_5221,N_5294);
xor U5447 (N_5447,N_5373,N_5223);
nor U5448 (N_5448,N_5380,N_5274);
and U5449 (N_5449,N_5253,N_5258);
nand U5450 (N_5450,N_5342,N_5309);
and U5451 (N_5451,N_5360,N_5209);
nand U5452 (N_5452,N_5231,N_5384);
nand U5453 (N_5453,N_5256,N_5222);
nand U5454 (N_5454,N_5325,N_5346);
and U5455 (N_5455,N_5260,N_5213);
nand U5456 (N_5456,N_5311,N_5268);
and U5457 (N_5457,N_5388,N_5348);
xnor U5458 (N_5458,N_5262,N_5390);
nor U5459 (N_5459,N_5320,N_5207);
nor U5460 (N_5460,N_5285,N_5201);
nand U5461 (N_5461,N_5354,N_5288);
or U5462 (N_5462,N_5265,N_5368);
or U5463 (N_5463,N_5299,N_5295);
and U5464 (N_5464,N_5255,N_5252);
nand U5465 (N_5465,N_5341,N_5337);
and U5466 (N_5466,N_5269,N_5374);
or U5467 (N_5467,N_5214,N_5266);
or U5468 (N_5468,N_5242,N_5248);
nor U5469 (N_5469,N_5361,N_5317);
or U5470 (N_5470,N_5378,N_5243);
or U5471 (N_5471,N_5312,N_5276);
nor U5472 (N_5472,N_5306,N_5315);
and U5473 (N_5473,N_5206,N_5282);
and U5474 (N_5474,N_5203,N_5399);
nor U5475 (N_5475,N_5239,N_5326);
nor U5476 (N_5476,N_5314,N_5215);
or U5477 (N_5477,N_5313,N_5338);
or U5478 (N_5478,N_5366,N_5236);
nand U5479 (N_5479,N_5283,N_5267);
nor U5480 (N_5480,N_5327,N_5364);
nand U5481 (N_5481,N_5264,N_5376);
nor U5482 (N_5482,N_5250,N_5220);
nand U5483 (N_5483,N_5302,N_5351);
and U5484 (N_5484,N_5254,N_5234);
xor U5485 (N_5485,N_5350,N_5318);
or U5486 (N_5486,N_5333,N_5340);
nor U5487 (N_5487,N_5241,N_5394);
nor U5488 (N_5488,N_5308,N_5371);
nand U5489 (N_5489,N_5251,N_5227);
xnor U5490 (N_5490,N_5202,N_5261);
nand U5491 (N_5491,N_5240,N_5270);
or U5492 (N_5492,N_5244,N_5345);
nor U5493 (N_5493,N_5385,N_5321);
xor U5494 (N_5494,N_5391,N_5386);
or U5495 (N_5495,N_5300,N_5330);
nor U5496 (N_5496,N_5247,N_5365);
nor U5497 (N_5497,N_5238,N_5332);
nand U5498 (N_5498,N_5359,N_5291);
xnor U5499 (N_5499,N_5225,N_5204);
or U5500 (N_5500,N_5278,N_5304);
xnor U5501 (N_5501,N_5335,N_5341);
and U5502 (N_5502,N_5298,N_5320);
nor U5503 (N_5503,N_5363,N_5223);
nand U5504 (N_5504,N_5259,N_5303);
nor U5505 (N_5505,N_5231,N_5387);
and U5506 (N_5506,N_5201,N_5222);
nor U5507 (N_5507,N_5289,N_5207);
and U5508 (N_5508,N_5378,N_5367);
nor U5509 (N_5509,N_5347,N_5391);
or U5510 (N_5510,N_5308,N_5312);
xnor U5511 (N_5511,N_5387,N_5390);
xnor U5512 (N_5512,N_5358,N_5224);
xnor U5513 (N_5513,N_5218,N_5310);
nor U5514 (N_5514,N_5264,N_5354);
or U5515 (N_5515,N_5306,N_5251);
xnor U5516 (N_5516,N_5394,N_5254);
nand U5517 (N_5517,N_5351,N_5214);
nor U5518 (N_5518,N_5343,N_5214);
nand U5519 (N_5519,N_5365,N_5334);
nand U5520 (N_5520,N_5362,N_5342);
and U5521 (N_5521,N_5263,N_5380);
xor U5522 (N_5522,N_5256,N_5338);
nand U5523 (N_5523,N_5368,N_5211);
xnor U5524 (N_5524,N_5240,N_5262);
nand U5525 (N_5525,N_5327,N_5289);
nand U5526 (N_5526,N_5362,N_5248);
xnor U5527 (N_5527,N_5367,N_5279);
xnor U5528 (N_5528,N_5215,N_5223);
nand U5529 (N_5529,N_5279,N_5237);
or U5530 (N_5530,N_5203,N_5367);
or U5531 (N_5531,N_5248,N_5238);
nor U5532 (N_5532,N_5238,N_5300);
and U5533 (N_5533,N_5352,N_5200);
and U5534 (N_5534,N_5291,N_5350);
or U5535 (N_5535,N_5385,N_5367);
nor U5536 (N_5536,N_5329,N_5203);
and U5537 (N_5537,N_5342,N_5385);
nand U5538 (N_5538,N_5254,N_5279);
and U5539 (N_5539,N_5344,N_5212);
nor U5540 (N_5540,N_5277,N_5314);
xnor U5541 (N_5541,N_5360,N_5222);
nor U5542 (N_5542,N_5364,N_5366);
or U5543 (N_5543,N_5369,N_5205);
nor U5544 (N_5544,N_5307,N_5242);
and U5545 (N_5545,N_5200,N_5285);
xor U5546 (N_5546,N_5276,N_5212);
xnor U5547 (N_5547,N_5264,N_5277);
or U5548 (N_5548,N_5361,N_5248);
nand U5549 (N_5549,N_5307,N_5292);
nor U5550 (N_5550,N_5362,N_5360);
or U5551 (N_5551,N_5340,N_5319);
xnor U5552 (N_5552,N_5370,N_5284);
or U5553 (N_5553,N_5389,N_5206);
nor U5554 (N_5554,N_5371,N_5342);
xnor U5555 (N_5555,N_5301,N_5315);
nand U5556 (N_5556,N_5384,N_5394);
and U5557 (N_5557,N_5246,N_5305);
and U5558 (N_5558,N_5264,N_5384);
nand U5559 (N_5559,N_5313,N_5331);
or U5560 (N_5560,N_5341,N_5283);
or U5561 (N_5561,N_5306,N_5350);
nor U5562 (N_5562,N_5231,N_5340);
nand U5563 (N_5563,N_5399,N_5364);
nand U5564 (N_5564,N_5312,N_5251);
xor U5565 (N_5565,N_5242,N_5239);
nor U5566 (N_5566,N_5358,N_5282);
xnor U5567 (N_5567,N_5322,N_5317);
nand U5568 (N_5568,N_5388,N_5289);
and U5569 (N_5569,N_5226,N_5386);
or U5570 (N_5570,N_5310,N_5263);
or U5571 (N_5571,N_5339,N_5248);
xor U5572 (N_5572,N_5387,N_5389);
or U5573 (N_5573,N_5394,N_5222);
and U5574 (N_5574,N_5214,N_5213);
xor U5575 (N_5575,N_5233,N_5245);
or U5576 (N_5576,N_5385,N_5234);
or U5577 (N_5577,N_5364,N_5202);
xor U5578 (N_5578,N_5265,N_5208);
or U5579 (N_5579,N_5245,N_5335);
and U5580 (N_5580,N_5280,N_5320);
nand U5581 (N_5581,N_5362,N_5235);
nand U5582 (N_5582,N_5265,N_5264);
xnor U5583 (N_5583,N_5373,N_5292);
or U5584 (N_5584,N_5309,N_5238);
and U5585 (N_5585,N_5201,N_5281);
nand U5586 (N_5586,N_5211,N_5388);
nor U5587 (N_5587,N_5357,N_5275);
xor U5588 (N_5588,N_5399,N_5243);
and U5589 (N_5589,N_5338,N_5387);
nor U5590 (N_5590,N_5286,N_5270);
nand U5591 (N_5591,N_5220,N_5266);
nand U5592 (N_5592,N_5373,N_5291);
and U5593 (N_5593,N_5220,N_5376);
or U5594 (N_5594,N_5227,N_5230);
xor U5595 (N_5595,N_5358,N_5269);
nor U5596 (N_5596,N_5285,N_5273);
xor U5597 (N_5597,N_5389,N_5375);
xnor U5598 (N_5598,N_5326,N_5317);
and U5599 (N_5599,N_5260,N_5241);
nand U5600 (N_5600,N_5486,N_5473);
and U5601 (N_5601,N_5514,N_5494);
nand U5602 (N_5602,N_5508,N_5447);
xor U5603 (N_5603,N_5597,N_5542);
or U5604 (N_5604,N_5594,N_5459);
nor U5605 (N_5605,N_5571,N_5506);
or U5606 (N_5606,N_5536,N_5461);
nor U5607 (N_5607,N_5468,N_5590);
xor U5608 (N_5608,N_5533,N_5527);
nand U5609 (N_5609,N_5568,N_5488);
and U5610 (N_5610,N_5462,N_5591);
nand U5611 (N_5611,N_5464,N_5589);
xnor U5612 (N_5612,N_5535,N_5439);
nand U5613 (N_5613,N_5565,N_5544);
nor U5614 (N_5614,N_5441,N_5557);
or U5615 (N_5615,N_5437,N_5550);
and U5616 (N_5616,N_5415,N_5418);
and U5617 (N_5617,N_5408,N_5496);
and U5618 (N_5618,N_5472,N_5541);
xnor U5619 (N_5619,N_5458,N_5519);
xor U5620 (N_5620,N_5445,N_5562);
or U5621 (N_5621,N_5561,N_5577);
or U5622 (N_5622,N_5526,N_5443);
or U5623 (N_5623,N_5442,N_5463);
and U5624 (N_5624,N_5517,N_5455);
and U5625 (N_5625,N_5466,N_5446);
xor U5626 (N_5626,N_5449,N_5503);
and U5627 (N_5627,N_5498,N_5593);
and U5628 (N_5628,N_5476,N_5406);
nor U5629 (N_5629,N_5483,N_5484);
xor U5630 (N_5630,N_5502,N_5559);
and U5631 (N_5631,N_5578,N_5429);
and U5632 (N_5632,N_5579,N_5487);
nor U5633 (N_5633,N_5420,N_5400);
nand U5634 (N_5634,N_5547,N_5428);
or U5635 (N_5635,N_5582,N_5529);
nand U5636 (N_5636,N_5478,N_5407);
xor U5637 (N_5637,N_5588,N_5583);
or U5638 (N_5638,N_5581,N_5467);
xnor U5639 (N_5639,N_5505,N_5523);
nor U5640 (N_5640,N_5491,N_5524);
nand U5641 (N_5641,N_5560,N_5518);
xor U5642 (N_5642,N_5564,N_5402);
or U5643 (N_5643,N_5580,N_5454);
nor U5644 (N_5644,N_5431,N_5510);
and U5645 (N_5645,N_5411,N_5501);
nand U5646 (N_5646,N_5599,N_5436);
nand U5647 (N_5647,N_5576,N_5471);
or U5648 (N_5648,N_5440,N_5525);
and U5649 (N_5649,N_5474,N_5497);
nand U5650 (N_5650,N_5465,N_5417);
xor U5651 (N_5651,N_5444,N_5433);
and U5652 (N_5652,N_5493,N_5574);
or U5653 (N_5653,N_5516,N_5425);
and U5654 (N_5654,N_5485,N_5522);
nand U5655 (N_5655,N_5534,N_5531);
and U5656 (N_5656,N_5570,N_5489);
or U5657 (N_5657,N_5512,N_5548);
xor U5658 (N_5658,N_5592,N_5586);
or U5659 (N_5659,N_5424,N_5584);
xor U5660 (N_5660,N_5587,N_5539);
nor U5661 (N_5661,N_5567,N_5413);
xor U5662 (N_5662,N_5515,N_5448);
and U5663 (N_5663,N_5521,N_5481);
or U5664 (N_5664,N_5509,N_5416);
nor U5665 (N_5665,N_5470,N_5530);
xor U5666 (N_5666,N_5403,N_5452);
xnor U5667 (N_5667,N_5457,N_5543);
nand U5668 (N_5668,N_5475,N_5549);
xnor U5669 (N_5669,N_5451,N_5546);
nand U5670 (N_5670,N_5573,N_5414);
nand U5671 (N_5671,N_5520,N_5499);
nand U5672 (N_5672,N_5495,N_5507);
nand U5673 (N_5673,N_5421,N_5595);
nand U5674 (N_5674,N_5585,N_5511);
xnor U5675 (N_5675,N_5469,N_5435);
nand U5676 (N_5676,N_5553,N_5412);
nor U5677 (N_5677,N_5540,N_5572);
and U5678 (N_5678,N_5423,N_5422);
xor U5679 (N_5679,N_5430,N_5427);
or U5680 (N_5680,N_5551,N_5545);
nor U5681 (N_5681,N_5405,N_5563);
xor U5682 (N_5682,N_5432,N_5456);
nor U5683 (N_5683,N_5532,N_5538);
and U5684 (N_5684,N_5426,N_5450);
nor U5685 (N_5685,N_5555,N_5537);
nor U5686 (N_5686,N_5410,N_5492);
or U5687 (N_5687,N_5552,N_5596);
xor U5688 (N_5688,N_5460,N_5419);
xor U5689 (N_5689,N_5598,N_5528);
nor U5690 (N_5690,N_5404,N_5401);
nand U5691 (N_5691,N_5453,N_5504);
nor U5692 (N_5692,N_5438,N_5500);
or U5693 (N_5693,N_5558,N_5434);
and U5694 (N_5694,N_5554,N_5409);
xnor U5695 (N_5695,N_5575,N_5482);
xnor U5696 (N_5696,N_5556,N_5490);
or U5697 (N_5697,N_5479,N_5566);
xnor U5698 (N_5698,N_5569,N_5513);
xor U5699 (N_5699,N_5477,N_5480);
nand U5700 (N_5700,N_5596,N_5558);
or U5701 (N_5701,N_5584,N_5450);
nor U5702 (N_5702,N_5510,N_5422);
and U5703 (N_5703,N_5492,N_5479);
xnor U5704 (N_5704,N_5593,N_5434);
and U5705 (N_5705,N_5508,N_5470);
nor U5706 (N_5706,N_5405,N_5460);
nand U5707 (N_5707,N_5537,N_5592);
and U5708 (N_5708,N_5499,N_5544);
nand U5709 (N_5709,N_5485,N_5460);
or U5710 (N_5710,N_5488,N_5407);
and U5711 (N_5711,N_5407,N_5479);
or U5712 (N_5712,N_5596,N_5430);
or U5713 (N_5713,N_5495,N_5422);
xor U5714 (N_5714,N_5507,N_5593);
nor U5715 (N_5715,N_5556,N_5528);
nor U5716 (N_5716,N_5439,N_5448);
and U5717 (N_5717,N_5474,N_5423);
and U5718 (N_5718,N_5586,N_5573);
or U5719 (N_5719,N_5401,N_5523);
or U5720 (N_5720,N_5499,N_5403);
xor U5721 (N_5721,N_5486,N_5510);
nor U5722 (N_5722,N_5404,N_5547);
or U5723 (N_5723,N_5416,N_5543);
or U5724 (N_5724,N_5494,N_5470);
nor U5725 (N_5725,N_5441,N_5496);
and U5726 (N_5726,N_5443,N_5453);
nand U5727 (N_5727,N_5502,N_5596);
xnor U5728 (N_5728,N_5467,N_5525);
nand U5729 (N_5729,N_5407,N_5551);
xnor U5730 (N_5730,N_5532,N_5448);
nor U5731 (N_5731,N_5506,N_5562);
nand U5732 (N_5732,N_5528,N_5459);
and U5733 (N_5733,N_5542,N_5499);
and U5734 (N_5734,N_5536,N_5415);
xnor U5735 (N_5735,N_5518,N_5573);
xor U5736 (N_5736,N_5462,N_5526);
and U5737 (N_5737,N_5542,N_5440);
nor U5738 (N_5738,N_5590,N_5482);
and U5739 (N_5739,N_5489,N_5567);
nor U5740 (N_5740,N_5553,N_5545);
nor U5741 (N_5741,N_5493,N_5484);
and U5742 (N_5742,N_5470,N_5411);
and U5743 (N_5743,N_5480,N_5430);
nor U5744 (N_5744,N_5453,N_5487);
and U5745 (N_5745,N_5444,N_5475);
nand U5746 (N_5746,N_5567,N_5438);
and U5747 (N_5747,N_5453,N_5580);
xnor U5748 (N_5748,N_5585,N_5523);
and U5749 (N_5749,N_5466,N_5598);
nand U5750 (N_5750,N_5589,N_5405);
and U5751 (N_5751,N_5521,N_5526);
nand U5752 (N_5752,N_5531,N_5479);
nor U5753 (N_5753,N_5499,N_5561);
xnor U5754 (N_5754,N_5525,N_5560);
nand U5755 (N_5755,N_5441,N_5490);
xnor U5756 (N_5756,N_5504,N_5596);
nor U5757 (N_5757,N_5447,N_5429);
or U5758 (N_5758,N_5503,N_5533);
nand U5759 (N_5759,N_5474,N_5452);
xnor U5760 (N_5760,N_5416,N_5539);
and U5761 (N_5761,N_5527,N_5553);
xor U5762 (N_5762,N_5486,N_5582);
nor U5763 (N_5763,N_5405,N_5510);
xnor U5764 (N_5764,N_5572,N_5493);
or U5765 (N_5765,N_5407,N_5598);
or U5766 (N_5766,N_5413,N_5424);
xnor U5767 (N_5767,N_5501,N_5575);
nor U5768 (N_5768,N_5417,N_5406);
and U5769 (N_5769,N_5549,N_5453);
and U5770 (N_5770,N_5461,N_5577);
nand U5771 (N_5771,N_5595,N_5470);
and U5772 (N_5772,N_5594,N_5423);
or U5773 (N_5773,N_5461,N_5473);
or U5774 (N_5774,N_5598,N_5509);
xor U5775 (N_5775,N_5482,N_5517);
nor U5776 (N_5776,N_5535,N_5543);
or U5777 (N_5777,N_5591,N_5510);
or U5778 (N_5778,N_5433,N_5521);
and U5779 (N_5779,N_5436,N_5587);
or U5780 (N_5780,N_5500,N_5596);
or U5781 (N_5781,N_5423,N_5413);
or U5782 (N_5782,N_5475,N_5463);
nor U5783 (N_5783,N_5542,N_5457);
and U5784 (N_5784,N_5476,N_5576);
or U5785 (N_5785,N_5519,N_5430);
xnor U5786 (N_5786,N_5582,N_5595);
nor U5787 (N_5787,N_5514,N_5558);
or U5788 (N_5788,N_5474,N_5467);
nor U5789 (N_5789,N_5432,N_5587);
nand U5790 (N_5790,N_5566,N_5469);
xnor U5791 (N_5791,N_5587,N_5598);
nor U5792 (N_5792,N_5484,N_5491);
nand U5793 (N_5793,N_5486,N_5597);
or U5794 (N_5794,N_5458,N_5597);
or U5795 (N_5795,N_5590,N_5489);
xnor U5796 (N_5796,N_5591,N_5458);
and U5797 (N_5797,N_5530,N_5554);
and U5798 (N_5798,N_5415,N_5599);
nand U5799 (N_5799,N_5459,N_5409);
and U5800 (N_5800,N_5634,N_5642);
nand U5801 (N_5801,N_5647,N_5601);
xor U5802 (N_5802,N_5717,N_5675);
and U5803 (N_5803,N_5697,N_5643);
xor U5804 (N_5804,N_5703,N_5769);
or U5805 (N_5805,N_5686,N_5748);
nand U5806 (N_5806,N_5670,N_5649);
nand U5807 (N_5807,N_5753,N_5684);
or U5808 (N_5808,N_5630,N_5696);
xor U5809 (N_5809,N_5676,N_5652);
nand U5810 (N_5810,N_5747,N_5673);
xor U5811 (N_5811,N_5688,N_5789);
nand U5812 (N_5812,N_5668,N_5700);
xnor U5813 (N_5813,N_5650,N_5632);
xnor U5814 (N_5814,N_5659,N_5743);
and U5815 (N_5815,N_5763,N_5623);
nand U5816 (N_5816,N_5691,N_5674);
nor U5817 (N_5817,N_5786,N_5774);
or U5818 (N_5818,N_5705,N_5683);
nor U5819 (N_5819,N_5790,N_5681);
xor U5820 (N_5820,N_5784,N_5605);
and U5821 (N_5821,N_5621,N_5692);
and U5822 (N_5822,N_5775,N_5766);
or U5823 (N_5823,N_5732,N_5754);
nand U5824 (N_5824,N_5730,N_5704);
xor U5825 (N_5825,N_5798,N_5685);
xor U5826 (N_5826,N_5612,N_5664);
and U5827 (N_5827,N_5609,N_5708);
and U5828 (N_5828,N_5667,N_5755);
and U5829 (N_5829,N_5633,N_5662);
or U5830 (N_5830,N_5735,N_5779);
nor U5831 (N_5831,N_5767,N_5600);
nand U5832 (N_5832,N_5738,N_5610);
nand U5833 (N_5833,N_5770,N_5602);
nor U5834 (N_5834,N_5603,N_5669);
or U5835 (N_5835,N_5648,N_5646);
and U5836 (N_5836,N_5733,N_5636);
or U5837 (N_5837,N_5617,N_5702);
nand U5838 (N_5838,N_5739,N_5611);
and U5839 (N_5839,N_5724,N_5785);
xnor U5840 (N_5840,N_5761,N_5654);
or U5841 (N_5841,N_5772,N_5663);
xor U5842 (N_5842,N_5768,N_5710);
or U5843 (N_5843,N_5628,N_5604);
nand U5844 (N_5844,N_5719,N_5764);
or U5845 (N_5845,N_5799,N_5728);
or U5846 (N_5846,N_5760,N_5797);
nor U5847 (N_5847,N_5695,N_5619);
nor U5848 (N_5848,N_5606,N_5655);
or U5849 (N_5849,N_5701,N_5639);
nand U5850 (N_5850,N_5627,N_5699);
nand U5851 (N_5851,N_5645,N_5677);
nor U5852 (N_5852,N_5720,N_5746);
nor U5853 (N_5853,N_5796,N_5776);
or U5854 (N_5854,N_5687,N_5638);
nor U5855 (N_5855,N_5783,N_5741);
and U5856 (N_5856,N_5788,N_5706);
and U5857 (N_5857,N_5765,N_5737);
xnor U5858 (N_5858,N_5742,N_5780);
xnor U5859 (N_5859,N_5672,N_5637);
nor U5860 (N_5860,N_5641,N_5608);
or U5861 (N_5861,N_5629,N_5757);
nor U5862 (N_5862,N_5625,N_5644);
nand U5863 (N_5863,N_5731,N_5758);
nor U5864 (N_5864,N_5750,N_5773);
nor U5865 (N_5865,N_5723,N_5736);
nor U5866 (N_5866,N_5626,N_5713);
nand U5867 (N_5867,N_5791,N_5661);
nor U5868 (N_5868,N_5759,N_5781);
nand U5869 (N_5869,N_5751,N_5726);
xor U5870 (N_5870,N_5745,N_5620);
xnor U5871 (N_5871,N_5665,N_5653);
and U5872 (N_5872,N_5718,N_5794);
nand U5873 (N_5873,N_5744,N_5716);
or U5874 (N_5874,N_5614,N_5678);
or U5875 (N_5875,N_5711,N_5782);
xnor U5876 (N_5876,N_5792,N_5658);
or U5877 (N_5877,N_5651,N_5712);
nor U5878 (N_5878,N_5752,N_5689);
nand U5879 (N_5879,N_5682,N_5734);
and U5880 (N_5880,N_5777,N_5715);
or U5881 (N_5881,N_5698,N_5607);
xor U5882 (N_5882,N_5635,N_5693);
or U5883 (N_5883,N_5727,N_5740);
nor U5884 (N_5884,N_5615,N_5725);
nor U5885 (N_5885,N_5624,N_5640);
xor U5886 (N_5886,N_5660,N_5690);
and U5887 (N_5887,N_5749,N_5694);
xor U5888 (N_5888,N_5756,N_5657);
nand U5889 (N_5889,N_5795,N_5618);
or U5890 (N_5890,N_5680,N_5721);
nand U5891 (N_5891,N_5631,N_5778);
xnor U5892 (N_5892,N_5709,N_5679);
or U5893 (N_5893,N_5793,N_5787);
nand U5894 (N_5894,N_5622,N_5671);
nor U5895 (N_5895,N_5707,N_5714);
xor U5896 (N_5896,N_5613,N_5666);
nand U5897 (N_5897,N_5616,N_5656);
and U5898 (N_5898,N_5762,N_5729);
xnor U5899 (N_5899,N_5771,N_5722);
nand U5900 (N_5900,N_5692,N_5707);
or U5901 (N_5901,N_5633,N_5748);
or U5902 (N_5902,N_5610,N_5775);
or U5903 (N_5903,N_5764,N_5739);
xor U5904 (N_5904,N_5765,N_5780);
xnor U5905 (N_5905,N_5752,N_5669);
nor U5906 (N_5906,N_5626,N_5708);
and U5907 (N_5907,N_5674,N_5631);
or U5908 (N_5908,N_5654,N_5642);
nor U5909 (N_5909,N_5742,N_5631);
or U5910 (N_5910,N_5768,N_5641);
or U5911 (N_5911,N_5771,N_5763);
nand U5912 (N_5912,N_5656,N_5762);
and U5913 (N_5913,N_5730,N_5681);
and U5914 (N_5914,N_5742,N_5641);
or U5915 (N_5915,N_5765,N_5778);
nand U5916 (N_5916,N_5689,N_5647);
xnor U5917 (N_5917,N_5756,N_5673);
nand U5918 (N_5918,N_5609,N_5653);
or U5919 (N_5919,N_5702,N_5689);
or U5920 (N_5920,N_5639,N_5630);
nor U5921 (N_5921,N_5620,N_5713);
and U5922 (N_5922,N_5780,N_5701);
and U5923 (N_5923,N_5603,N_5754);
xor U5924 (N_5924,N_5779,N_5673);
xnor U5925 (N_5925,N_5688,N_5622);
and U5926 (N_5926,N_5777,N_5761);
and U5927 (N_5927,N_5707,N_5676);
nor U5928 (N_5928,N_5771,N_5690);
or U5929 (N_5929,N_5796,N_5711);
and U5930 (N_5930,N_5774,N_5654);
nand U5931 (N_5931,N_5664,N_5721);
nand U5932 (N_5932,N_5701,N_5646);
nand U5933 (N_5933,N_5760,N_5790);
and U5934 (N_5934,N_5633,N_5720);
and U5935 (N_5935,N_5782,N_5748);
and U5936 (N_5936,N_5745,N_5769);
xnor U5937 (N_5937,N_5795,N_5793);
or U5938 (N_5938,N_5763,N_5758);
or U5939 (N_5939,N_5761,N_5795);
nand U5940 (N_5940,N_5708,N_5747);
or U5941 (N_5941,N_5771,N_5784);
and U5942 (N_5942,N_5776,N_5783);
nand U5943 (N_5943,N_5713,N_5785);
nand U5944 (N_5944,N_5714,N_5770);
xor U5945 (N_5945,N_5603,N_5666);
and U5946 (N_5946,N_5783,N_5699);
or U5947 (N_5947,N_5748,N_5621);
nand U5948 (N_5948,N_5679,N_5646);
xor U5949 (N_5949,N_5792,N_5688);
nor U5950 (N_5950,N_5668,N_5702);
or U5951 (N_5951,N_5629,N_5714);
xor U5952 (N_5952,N_5643,N_5678);
and U5953 (N_5953,N_5793,N_5669);
or U5954 (N_5954,N_5780,N_5665);
and U5955 (N_5955,N_5694,N_5771);
xor U5956 (N_5956,N_5695,N_5620);
xnor U5957 (N_5957,N_5720,N_5680);
xnor U5958 (N_5958,N_5700,N_5790);
or U5959 (N_5959,N_5692,N_5618);
nand U5960 (N_5960,N_5730,N_5670);
or U5961 (N_5961,N_5701,N_5666);
nor U5962 (N_5962,N_5737,N_5790);
and U5963 (N_5963,N_5792,N_5776);
nor U5964 (N_5964,N_5734,N_5747);
nand U5965 (N_5965,N_5632,N_5776);
or U5966 (N_5966,N_5691,N_5765);
xnor U5967 (N_5967,N_5632,N_5660);
xnor U5968 (N_5968,N_5611,N_5723);
nor U5969 (N_5969,N_5689,N_5600);
and U5970 (N_5970,N_5631,N_5741);
and U5971 (N_5971,N_5601,N_5688);
or U5972 (N_5972,N_5756,N_5784);
and U5973 (N_5973,N_5655,N_5761);
nor U5974 (N_5974,N_5707,N_5608);
nand U5975 (N_5975,N_5721,N_5798);
or U5976 (N_5976,N_5761,N_5644);
or U5977 (N_5977,N_5792,N_5606);
and U5978 (N_5978,N_5722,N_5616);
xor U5979 (N_5979,N_5600,N_5622);
xnor U5980 (N_5980,N_5613,N_5672);
and U5981 (N_5981,N_5712,N_5693);
nor U5982 (N_5982,N_5760,N_5761);
xnor U5983 (N_5983,N_5669,N_5601);
nor U5984 (N_5984,N_5781,N_5630);
xor U5985 (N_5985,N_5733,N_5743);
nor U5986 (N_5986,N_5627,N_5686);
nand U5987 (N_5987,N_5601,N_5663);
xnor U5988 (N_5988,N_5745,N_5783);
nand U5989 (N_5989,N_5795,N_5799);
xnor U5990 (N_5990,N_5669,N_5606);
xor U5991 (N_5991,N_5786,N_5684);
nor U5992 (N_5992,N_5699,N_5752);
nor U5993 (N_5993,N_5750,N_5698);
nor U5994 (N_5994,N_5783,N_5718);
xor U5995 (N_5995,N_5602,N_5617);
nor U5996 (N_5996,N_5733,N_5692);
nor U5997 (N_5997,N_5637,N_5686);
and U5998 (N_5998,N_5691,N_5777);
nand U5999 (N_5999,N_5699,N_5721);
nor U6000 (N_6000,N_5932,N_5840);
nand U6001 (N_6001,N_5970,N_5803);
nand U6002 (N_6002,N_5871,N_5869);
nor U6003 (N_6003,N_5819,N_5831);
or U6004 (N_6004,N_5815,N_5888);
nand U6005 (N_6005,N_5852,N_5913);
and U6006 (N_6006,N_5813,N_5996);
xnor U6007 (N_6007,N_5902,N_5889);
xor U6008 (N_6008,N_5984,N_5824);
and U6009 (N_6009,N_5873,N_5825);
nor U6010 (N_6010,N_5878,N_5905);
nand U6011 (N_6011,N_5926,N_5844);
nor U6012 (N_6012,N_5909,N_5924);
or U6013 (N_6013,N_5914,N_5884);
nand U6014 (N_6014,N_5904,N_5881);
nor U6015 (N_6015,N_5809,N_5939);
xor U6016 (N_6016,N_5928,N_5942);
and U6017 (N_6017,N_5858,N_5842);
nand U6018 (N_6018,N_5960,N_5965);
nor U6019 (N_6019,N_5916,N_5950);
or U6020 (N_6020,N_5816,N_5872);
or U6021 (N_6021,N_5846,N_5829);
nand U6022 (N_6022,N_5957,N_5836);
or U6023 (N_6023,N_5892,N_5862);
nand U6024 (N_6024,N_5901,N_5969);
nand U6025 (N_6025,N_5850,N_5808);
and U6026 (N_6026,N_5908,N_5987);
xor U6027 (N_6027,N_5810,N_5955);
or U6028 (N_6028,N_5857,N_5956);
nand U6029 (N_6029,N_5856,N_5976);
or U6030 (N_6030,N_5887,N_5870);
xnor U6031 (N_6031,N_5893,N_5922);
nand U6032 (N_6032,N_5993,N_5986);
nor U6033 (N_6033,N_5899,N_5860);
xnor U6034 (N_6034,N_5935,N_5938);
or U6035 (N_6035,N_5999,N_5863);
and U6036 (N_6036,N_5835,N_5900);
nor U6037 (N_6037,N_5898,N_5855);
nand U6038 (N_6038,N_5845,N_5992);
or U6039 (N_6039,N_5981,N_5934);
or U6040 (N_6040,N_5895,N_5927);
and U6041 (N_6041,N_5997,N_5826);
xnor U6042 (N_6042,N_5964,N_5915);
nand U6043 (N_6043,N_5804,N_5827);
and U6044 (N_6044,N_5838,N_5866);
nand U6045 (N_6045,N_5933,N_5874);
or U6046 (N_6046,N_5941,N_5975);
or U6047 (N_6047,N_5979,N_5807);
nor U6048 (N_6048,N_5943,N_5925);
nor U6049 (N_6049,N_5954,N_5973);
nor U6050 (N_6050,N_5920,N_5977);
nor U6051 (N_6051,N_5880,N_5944);
xnor U6052 (N_6052,N_5865,N_5822);
or U6053 (N_6053,N_5885,N_5991);
nand U6054 (N_6054,N_5919,N_5823);
xnor U6055 (N_6055,N_5994,N_5883);
nand U6056 (N_6056,N_5980,N_5995);
nor U6057 (N_6057,N_5875,N_5894);
nor U6058 (N_6058,N_5968,N_5886);
xnor U6059 (N_6059,N_5876,N_5990);
nor U6060 (N_6060,N_5832,N_5982);
nand U6061 (N_6061,N_5849,N_5974);
xor U6062 (N_6062,N_5949,N_5843);
xnor U6063 (N_6063,N_5814,N_5940);
or U6064 (N_6064,N_5821,N_5930);
and U6065 (N_6065,N_5983,N_5958);
or U6066 (N_6066,N_5962,N_5811);
xor U6067 (N_6067,N_5985,N_5910);
xnor U6068 (N_6068,N_5848,N_5967);
or U6069 (N_6069,N_5896,N_5882);
xor U6070 (N_6070,N_5989,N_5948);
nor U6071 (N_6071,N_5971,N_5929);
xor U6072 (N_6072,N_5918,N_5937);
nand U6073 (N_6073,N_5868,N_5951);
and U6074 (N_6074,N_5897,N_5828);
xnor U6075 (N_6075,N_5859,N_5998);
nor U6076 (N_6076,N_5817,N_5961);
nor U6077 (N_6077,N_5953,N_5959);
xor U6078 (N_6078,N_5923,N_5805);
and U6079 (N_6079,N_5945,N_5978);
nand U6080 (N_6080,N_5952,N_5877);
nand U6081 (N_6081,N_5800,N_5911);
xnor U6082 (N_6082,N_5820,N_5907);
nor U6083 (N_6083,N_5834,N_5921);
and U6084 (N_6084,N_5851,N_5864);
or U6085 (N_6085,N_5853,N_5801);
and U6086 (N_6086,N_5917,N_5837);
nand U6087 (N_6087,N_5839,N_5946);
or U6088 (N_6088,N_5988,N_5966);
xnor U6089 (N_6089,N_5867,N_5903);
xor U6090 (N_6090,N_5890,N_5912);
nand U6091 (N_6091,N_5963,N_5841);
xor U6092 (N_6092,N_5833,N_5947);
or U6093 (N_6093,N_5972,N_5854);
nor U6094 (N_6094,N_5906,N_5818);
xnor U6095 (N_6095,N_5936,N_5830);
and U6096 (N_6096,N_5812,N_5879);
and U6097 (N_6097,N_5861,N_5802);
or U6098 (N_6098,N_5931,N_5891);
and U6099 (N_6099,N_5847,N_5806);
nor U6100 (N_6100,N_5923,N_5803);
nand U6101 (N_6101,N_5870,N_5801);
nand U6102 (N_6102,N_5934,N_5863);
nand U6103 (N_6103,N_5839,N_5921);
and U6104 (N_6104,N_5956,N_5947);
nor U6105 (N_6105,N_5971,N_5852);
nor U6106 (N_6106,N_5858,N_5863);
and U6107 (N_6107,N_5834,N_5974);
nor U6108 (N_6108,N_5907,N_5942);
nand U6109 (N_6109,N_5904,N_5839);
nand U6110 (N_6110,N_5975,N_5857);
and U6111 (N_6111,N_5851,N_5894);
xnor U6112 (N_6112,N_5966,N_5927);
and U6113 (N_6113,N_5833,N_5918);
nor U6114 (N_6114,N_5895,N_5858);
xor U6115 (N_6115,N_5839,N_5906);
nor U6116 (N_6116,N_5882,N_5934);
or U6117 (N_6117,N_5999,N_5947);
and U6118 (N_6118,N_5969,N_5951);
nor U6119 (N_6119,N_5899,N_5961);
nor U6120 (N_6120,N_5836,N_5821);
nor U6121 (N_6121,N_5963,N_5990);
xnor U6122 (N_6122,N_5910,N_5865);
nand U6123 (N_6123,N_5809,N_5916);
nand U6124 (N_6124,N_5809,N_5959);
and U6125 (N_6125,N_5908,N_5959);
or U6126 (N_6126,N_5926,N_5807);
and U6127 (N_6127,N_5911,N_5849);
and U6128 (N_6128,N_5941,N_5921);
xor U6129 (N_6129,N_5846,N_5929);
nand U6130 (N_6130,N_5918,N_5960);
and U6131 (N_6131,N_5960,N_5955);
xor U6132 (N_6132,N_5809,N_5839);
or U6133 (N_6133,N_5873,N_5830);
and U6134 (N_6134,N_5863,N_5975);
and U6135 (N_6135,N_5921,N_5915);
nand U6136 (N_6136,N_5929,N_5956);
or U6137 (N_6137,N_5906,N_5834);
and U6138 (N_6138,N_5807,N_5927);
xor U6139 (N_6139,N_5844,N_5967);
xor U6140 (N_6140,N_5847,N_5843);
nand U6141 (N_6141,N_5965,N_5922);
nand U6142 (N_6142,N_5906,N_5902);
or U6143 (N_6143,N_5828,N_5822);
or U6144 (N_6144,N_5988,N_5940);
and U6145 (N_6145,N_5980,N_5969);
xnor U6146 (N_6146,N_5879,N_5891);
xor U6147 (N_6147,N_5968,N_5909);
and U6148 (N_6148,N_5838,N_5990);
xor U6149 (N_6149,N_5958,N_5982);
or U6150 (N_6150,N_5936,N_5911);
nor U6151 (N_6151,N_5898,N_5800);
nand U6152 (N_6152,N_5858,N_5882);
nor U6153 (N_6153,N_5838,N_5924);
or U6154 (N_6154,N_5839,N_5908);
nand U6155 (N_6155,N_5879,N_5996);
xor U6156 (N_6156,N_5959,N_5932);
xor U6157 (N_6157,N_5816,N_5851);
nor U6158 (N_6158,N_5874,N_5824);
nand U6159 (N_6159,N_5983,N_5909);
nor U6160 (N_6160,N_5854,N_5984);
and U6161 (N_6161,N_5913,N_5908);
and U6162 (N_6162,N_5977,N_5992);
xor U6163 (N_6163,N_5986,N_5808);
xnor U6164 (N_6164,N_5954,N_5804);
and U6165 (N_6165,N_5837,N_5825);
or U6166 (N_6166,N_5997,N_5937);
and U6167 (N_6167,N_5971,N_5903);
or U6168 (N_6168,N_5807,N_5822);
or U6169 (N_6169,N_5959,N_5905);
xor U6170 (N_6170,N_5964,N_5933);
nor U6171 (N_6171,N_5931,N_5973);
nand U6172 (N_6172,N_5911,N_5828);
nand U6173 (N_6173,N_5873,N_5940);
or U6174 (N_6174,N_5993,N_5846);
nor U6175 (N_6175,N_5919,N_5816);
and U6176 (N_6176,N_5907,N_5969);
or U6177 (N_6177,N_5843,N_5832);
and U6178 (N_6178,N_5811,N_5950);
xor U6179 (N_6179,N_5955,N_5989);
nand U6180 (N_6180,N_5919,N_5812);
nand U6181 (N_6181,N_5938,N_5907);
nor U6182 (N_6182,N_5939,N_5945);
or U6183 (N_6183,N_5807,N_5924);
xnor U6184 (N_6184,N_5960,N_5878);
nor U6185 (N_6185,N_5814,N_5998);
and U6186 (N_6186,N_5893,N_5801);
nor U6187 (N_6187,N_5884,N_5949);
xor U6188 (N_6188,N_5802,N_5805);
or U6189 (N_6189,N_5991,N_5874);
nor U6190 (N_6190,N_5937,N_5856);
or U6191 (N_6191,N_5957,N_5992);
xnor U6192 (N_6192,N_5835,N_5912);
nand U6193 (N_6193,N_5956,N_5888);
or U6194 (N_6194,N_5914,N_5996);
nand U6195 (N_6195,N_5919,N_5911);
or U6196 (N_6196,N_5917,N_5979);
or U6197 (N_6197,N_5924,N_5995);
xor U6198 (N_6198,N_5803,N_5956);
and U6199 (N_6199,N_5915,N_5893);
or U6200 (N_6200,N_6082,N_6179);
nand U6201 (N_6201,N_6198,N_6064);
nand U6202 (N_6202,N_6123,N_6006);
or U6203 (N_6203,N_6152,N_6197);
or U6204 (N_6204,N_6007,N_6132);
nor U6205 (N_6205,N_6157,N_6090);
nor U6206 (N_6206,N_6009,N_6033);
nand U6207 (N_6207,N_6170,N_6185);
xor U6208 (N_6208,N_6094,N_6074);
xnor U6209 (N_6209,N_6072,N_6057);
xor U6210 (N_6210,N_6115,N_6168);
xnor U6211 (N_6211,N_6018,N_6138);
nand U6212 (N_6212,N_6174,N_6036);
nand U6213 (N_6213,N_6026,N_6095);
nand U6214 (N_6214,N_6004,N_6188);
nor U6215 (N_6215,N_6088,N_6141);
and U6216 (N_6216,N_6024,N_6003);
nand U6217 (N_6217,N_6013,N_6031);
nand U6218 (N_6218,N_6124,N_6130);
and U6219 (N_6219,N_6010,N_6142);
and U6220 (N_6220,N_6032,N_6187);
xnor U6221 (N_6221,N_6114,N_6101);
or U6222 (N_6222,N_6085,N_6107);
and U6223 (N_6223,N_6149,N_6139);
nand U6224 (N_6224,N_6190,N_6028);
and U6225 (N_6225,N_6155,N_6102);
or U6226 (N_6226,N_6086,N_6106);
nand U6227 (N_6227,N_6080,N_6076);
or U6228 (N_6228,N_6005,N_6183);
xor U6229 (N_6229,N_6098,N_6159);
or U6230 (N_6230,N_6062,N_6103);
nor U6231 (N_6231,N_6025,N_6070);
nand U6232 (N_6232,N_6023,N_6069);
nor U6233 (N_6233,N_6056,N_6035);
nor U6234 (N_6234,N_6058,N_6049);
nor U6235 (N_6235,N_6131,N_6161);
xnor U6236 (N_6236,N_6136,N_6078);
and U6237 (N_6237,N_6117,N_6121);
nor U6238 (N_6238,N_6084,N_6104);
nand U6239 (N_6239,N_6175,N_6111);
or U6240 (N_6240,N_6027,N_6011);
nand U6241 (N_6241,N_6193,N_6030);
nor U6242 (N_6242,N_6119,N_6001);
xor U6243 (N_6243,N_6040,N_6148);
nor U6244 (N_6244,N_6195,N_6039);
or U6245 (N_6245,N_6063,N_6044);
nor U6246 (N_6246,N_6118,N_6050);
xnor U6247 (N_6247,N_6037,N_6177);
nand U6248 (N_6248,N_6060,N_6077);
nand U6249 (N_6249,N_6191,N_6120);
xnor U6250 (N_6250,N_6017,N_6163);
xor U6251 (N_6251,N_6066,N_6065);
or U6252 (N_6252,N_6158,N_6015);
xor U6253 (N_6253,N_6012,N_6048);
or U6254 (N_6254,N_6046,N_6097);
nand U6255 (N_6255,N_6092,N_6068);
and U6256 (N_6256,N_6112,N_6165);
xnor U6257 (N_6257,N_6184,N_6162);
xnor U6258 (N_6258,N_6172,N_6180);
xnor U6259 (N_6259,N_6091,N_6109);
or U6260 (N_6260,N_6153,N_6176);
and U6261 (N_6261,N_6075,N_6129);
nor U6262 (N_6262,N_6083,N_6002);
nand U6263 (N_6263,N_6038,N_6099);
xnor U6264 (N_6264,N_6016,N_6116);
nand U6265 (N_6265,N_6008,N_6182);
and U6266 (N_6266,N_6087,N_6053);
nor U6267 (N_6267,N_6043,N_6105);
nor U6268 (N_6268,N_6071,N_6178);
and U6269 (N_6269,N_6100,N_6199);
nand U6270 (N_6270,N_6156,N_6171);
xnor U6271 (N_6271,N_6145,N_6192);
nand U6272 (N_6272,N_6093,N_6143);
nor U6273 (N_6273,N_6079,N_6167);
nand U6274 (N_6274,N_6181,N_6144);
xnor U6275 (N_6275,N_6122,N_6021);
and U6276 (N_6276,N_6173,N_6096);
and U6277 (N_6277,N_6042,N_6089);
and U6278 (N_6278,N_6169,N_6000);
or U6279 (N_6279,N_6051,N_6127);
and U6280 (N_6280,N_6019,N_6081);
nand U6281 (N_6281,N_6113,N_6164);
nand U6282 (N_6282,N_6128,N_6135);
or U6283 (N_6283,N_6014,N_6146);
xor U6284 (N_6284,N_6022,N_6047);
and U6285 (N_6285,N_6140,N_6134);
xnor U6286 (N_6286,N_6125,N_6186);
xor U6287 (N_6287,N_6189,N_6067);
and U6288 (N_6288,N_6110,N_6052);
or U6289 (N_6289,N_6126,N_6147);
and U6290 (N_6290,N_6055,N_6133);
nor U6291 (N_6291,N_6160,N_6073);
and U6292 (N_6292,N_6041,N_6020);
or U6293 (N_6293,N_6137,N_6054);
nand U6294 (N_6294,N_6154,N_6045);
nor U6295 (N_6295,N_6150,N_6059);
and U6296 (N_6296,N_6151,N_6166);
or U6297 (N_6297,N_6034,N_6108);
nor U6298 (N_6298,N_6029,N_6194);
xor U6299 (N_6299,N_6061,N_6196);
xnor U6300 (N_6300,N_6006,N_6041);
nand U6301 (N_6301,N_6093,N_6073);
or U6302 (N_6302,N_6124,N_6043);
nand U6303 (N_6303,N_6049,N_6107);
nand U6304 (N_6304,N_6144,N_6108);
nand U6305 (N_6305,N_6118,N_6003);
or U6306 (N_6306,N_6027,N_6160);
nor U6307 (N_6307,N_6018,N_6066);
or U6308 (N_6308,N_6026,N_6060);
nand U6309 (N_6309,N_6187,N_6101);
and U6310 (N_6310,N_6021,N_6034);
xnor U6311 (N_6311,N_6163,N_6148);
and U6312 (N_6312,N_6142,N_6067);
or U6313 (N_6313,N_6074,N_6137);
or U6314 (N_6314,N_6057,N_6007);
nor U6315 (N_6315,N_6135,N_6186);
and U6316 (N_6316,N_6075,N_6059);
xor U6317 (N_6317,N_6077,N_6079);
nand U6318 (N_6318,N_6197,N_6169);
nor U6319 (N_6319,N_6166,N_6116);
nand U6320 (N_6320,N_6004,N_6119);
or U6321 (N_6321,N_6166,N_6192);
and U6322 (N_6322,N_6149,N_6081);
xor U6323 (N_6323,N_6166,N_6186);
xnor U6324 (N_6324,N_6111,N_6126);
or U6325 (N_6325,N_6024,N_6103);
or U6326 (N_6326,N_6000,N_6074);
or U6327 (N_6327,N_6172,N_6071);
xor U6328 (N_6328,N_6196,N_6136);
xnor U6329 (N_6329,N_6084,N_6173);
or U6330 (N_6330,N_6148,N_6095);
nor U6331 (N_6331,N_6185,N_6120);
xor U6332 (N_6332,N_6030,N_6061);
nand U6333 (N_6333,N_6142,N_6191);
or U6334 (N_6334,N_6038,N_6109);
nor U6335 (N_6335,N_6121,N_6038);
xor U6336 (N_6336,N_6082,N_6080);
nand U6337 (N_6337,N_6174,N_6015);
nor U6338 (N_6338,N_6137,N_6077);
xor U6339 (N_6339,N_6140,N_6011);
and U6340 (N_6340,N_6179,N_6190);
nand U6341 (N_6341,N_6186,N_6077);
nand U6342 (N_6342,N_6075,N_6097);
xor U6343 (N_6343,N_6184,N_6089);
or U6344 (N_6344,N_6077,N_6029);
or U6345 (N_6345,N_6007,N_6038);
or U6346 (N_6346,N_6051,N_6199);
or U6347 (N_6347,N_6095,N_6054);
xor U6348 (N_6348,N_6171,N_6154);
xor U6349 (N_6349,N_6057,N_6018);
and U6350 (N_6350,N_6123,N_6173);
nand U6351 (N_6351,N_6149,N_6083);
nand U6352 (N_6352,N_6154,N_6038);
nor U6353 (N_6353,N_6102,N_6128);
nor U6354 (N_6354,N_6194,N_6015);
xnor U6355 (N_6355,N_6058,N_6189);
or U6356 (N_6356,N_6016,N_6117);
xnor U6357 (N_6357,N_6163,N_6167);
nand U6358 (N_6358,N_6147,N_6110);
and U6359 (N_6359,N_6197,N_6171);
nor U6360 (N_6360,N_6011,N_6122);
or U6361 (N_6361,N_6002,N_6005);
nor U6362 (N_6362,N_6142,N_6073);
nand U6363 (N_6363,N_6150,N_6192);
nor U6364 (N_6364,N_6176,N_6184);
nand U6365 (N_6365,N_6160,N_6175);
nor U6366 (N_6366,N_6131,N_6024);
nand U6367 (N_6367,N_6082,N_6104);
nand U6368 (N_6368,N_6155,N_6034);
or U6369 (N_6369,N_6158,N_6027);
xnor U6370 (N_6370,N_6043,N_6025);
nand U6371 (N_6371,N_6199,N_6020);
nand U6372 (N_6372,N_6137,N_6061);
or U6373 (N_6373,N_6152,N_6096);
xor U6374 (N_6374,N_6035,N_6133);
xnor U6375 (N_6375,N_6135,N_6112);
nor U6376 (N_6376,N_6011,N_6007);
or U6377 (N_6377,N_6131,N_6123);
nand U6378 (N_6378,N_6129,N_6082);
and U6379 (N_6379,N_6025,N_6014);
nor U6380 (N_6380,N_6035,N_6180);
nand U6381 (N_6381,N_6093,N_6062);
and U6382 (N_6382,N_6038,N_6059);
or U6383 (N_6383,N_6125,N_6089);
and U6384 (N_6384,N_6092,N_6100);
and U6385 (N_6385,N_6081,N_6003);
nand U6386 (N_6386,N_6110,N_6040);
and U6387 (N_6387,N_6069,N_6152);
and U6388 (N_6388,N_6135,N_6157);
nor U6389 (N_6389,N_6193,N_6097);
nand U6390 (N_6390,N_6183,N_6137);
xor U6391 (N_6391,N_6002,N_6191);
nand U6392 (N_6392,N_6075,N_6104);
and U6393 (N_6393,N_6047,N_6075);
and U6394 (N_6394,N_6037,N_6165);
or U6395 (N_6395,N_6158,N_6029);
or U6396 (N_6396,N_6039,N_6088);
nor U6397 (N_6397,N_6015,N_6009);
and U6398 (N_6398,N_6014,N_6071);
and U6399 (N_6399,N_6083,N_6012);
xnor U6400 (N_6400,N_6368,N_6278);
nor U6401 (N_6401,N_6299,N_6381);
nand U6402 (N_6402,N_6246,N_6307);
xor U6403 (N_6403,N_6280,N_6203);
and U6404 (N_6404,N_6377,N_6383);
xnor U6405 (N_6405,N_6320,N_6201);
xnor U6406 (N_6406,N_6347,N_6264);
and U6407 (N_6407,N_6217,N_6267);
nor U6408 (N_6408,N_6221,N_6250);
and U6409 (N_6409,N_6392,N_6310);
and U6410 (N_6410,N_6214,N_6272);
and U6411 (N_6411,N_6371,N_6372);
nor U6412 (N_6412,N_6385,N_6211);
nand U6413 (N_6413,N_6229,N_6205);
and U6414 (N_6414,N_6233,N_6399);
nand U6415 (N_6415,N_6282,N_6319);
and U6416 (N_6416,N_6329,N_6380);
nor U6417 (N_6417,N_6232,N_6312);
or U6418 (N_6418,N_6348,N_6294);
and U6419 (N_6419,N_6345,N_6353);
nor U6420 (N_6420,N_6226,N_6387);
and U6421 (N_6421,N_6367,N_6364);
or U6422 (N_6422,N_6216,N_6340);
nand U6423 (N_6423,N_6296,N_6209);
nand U6424 (N_6424,N_6281,N_6324);
nor U6425 (N_6425,N_6341,N_6379);
nand U6426 (N_6426,N_6289,N_6235);
nand U6427 (N_6427,N_6369,N_6208);
or U6428 (N_6428,N_6298,N_6395);
or U6429 (N_6429,N_6207,N_6394);
and U6430 (N_6430,N_6276,N_6332);
xnor U6431 (N_6431,N_6318,N_6228);
nand U6432 (N_6432,N_6331,N_6277);
nor U6433 (N_6433,N_6352,N_6382);
or U6434 (N_6434,N_6206,N_6397);
xnor U6435 (N_6435,N_6355,N_6265);
nand U6436 (N_6436,N_6252,N_6279);
nor U6437 (N_6437,N_6316,N_6315);
or U6438 (N_6438,N_6223,N_6251);
nand U6439 (N_6439,N_6247,N_6231);
xor U6440 (N_6440,N_6334,N_6269);
nand U6441 (N_6441,N_6327,N_6244);
nand U6442 (N_6442,N_6204,N_6378);
or U6443 (N_6443,N_6323,N_6255);
and U6444 (N_6444,N_6300,N_6257);
and U6445 (N_6445,N_6202,N_6225);
xnor U6446 (N_6446,N_6356,N_6230);
nor U6447 (N_6447,N_6236,N_6259);
xor U6448 (N_6448,N_6311,N_6303);
or U6449 (N_6449,N_6218,N_6262);
nand U6450 (N_6450,N_6391,N_6354);
xor U6451 (N_6451,N_6322,N_6238);
or U6452 (N_6452,N_6263,N_6239);
or U6453 (N_6453,N_6393,N_6346);
and U6454 (N_6454,N_6274,N_6330);
and U6455 (N_6455,N_6386,N_6291);
and U6456 (N_6456,N_6313,N_6240);
nor U6457 (N_6457,N_6254,N_6285);
or U6458 (N_6458,N_6237,N_6245);
and U6459 (N_6459,N_6212,N_6390);
nand U6460 (N_6460,N_6398,N_6325);
and U6461 (N_6461,N_6304,N_6219);
nor U6462 (N_6462,N_6362,N_6290);
nand U6463 (N_6463,N_6363,N_6295);
or U6464 (N_6464,N_6241,N_6375);
nand U6465 (N_6465,N_6342,N_6338);
xor U6466 (N_6466,N_6305,N_6365);
nand U6467 (N_6467,N_6336,N_6286);
nand U6468 (N_6468,N_6370,N_6308);
nand U6469 (N_6469,N_6256,N_6361);
xnor U6470 (N_6470,N_6261,N_6227);
or U6471 (N_6471,N_6302,N_6224);
nand U6472 (N_6472,N_6248,N_6349);
nand U6473 (N_6473,N_6213,N_6283);
or U6474 (N_6474,N_6249,N_6301);
nor U6475 (N_6475,N_6359,N_6374);
and U6476 (N_6476,N_6396,N_6388);
nor U6477 (N_6477,N_6321,N_6317);
or U6478 (N_6478,N_6288,N_6333);
xor U6479 (N_6479,N_6360,N_6215);
and U6480 (N_6480,N_6389,N_6366);
nand U6481 (N_6481,N_6234,N_6335);
and U6482 (N_6482,N_6376,N_6200);
nand U6483 (N_6483,N_6242,N_6260);
xor U6484 (N_6484,N_6326,N_6210);
nand U6485 (N_6485,N_6293,N_6306);
nor U6486 (N_6486,N_6273,N_6292);
xor U6487 (N_6487,N_6284,N_6275);
and U6488 (N_6488,N_6373,N_6287);
nor U6489 (N_6489,N_6358,N_6266);
and U6490 (N_6490,N_6268,N_6309);
and U6491 (N_6491,N_6271,N_6350);
and U6492 (N_6492,N_6339,N_6253);
nand U6493 (N_6493,N_6384,N_6351);
or U6494 (N_6494,N_6243,N_6258);
xor U6495 (N_6495,N_6297,N_6270);
and U6496 (N_6496,N_6220,N_6357);
nand U6497 (N_6497,N_6337,N_6328);
nor U6498 (N_6498,N_6343,N_6314);
xor U6499 (N_6499,N_6222,N_6344);
xnor U6500 (N_6500,N_6250,N_6204);
or U6501 (N_6501,N_6371,N_6275);
nor U6502 (N_6502,N_6244,N_6251);
and U6503 (N_6503,N_6361,N_6348);
nor U6504 (N_6504,N_6368,N_6238);
or U6505 (N_6505,N_6314,N_6279);
nand U6506 (N_6506,N_6368,N_6274);
or U6507 (N_6507,N_6386,N_6339);
and U6508 (N_6508,N_6238,N_6289);
and U6509 (N_6509,N_6223,N_6391);
xor U6510 (N_6510,N_6248,N_6313);
and U6511 (N_6511,N_6217,N_6386);
nor U6512 (N_6512,N_6245,N_6338);
nor U6513 (N_6513,N_6226,N_6374);
and U6514 (N_6514,N_6397,N_6393);
nand U6515 (N_6515,N_6303,N_6308);
or U6516 (N_6516,N_6308,N_6296);
nand U6517 (N_6517,N_6291,N_6383);
nor U6518 (N_6518,N_6219,N_6200);
xor U6519 (N_6519,N_6252,N_6211);
xor U6520 (N_6520,N_6350,N_6359);
nand U6521 (N_6521,N_6207,N_6328);
or U6522 (N_6522,N_6216,N_6259);
or U6523 (N_6523,N_6265,N_6337);
xnor U6524 (N_6524,N_6227,N_6215);
and U6525 (N_6525,N_6345,N_6373);
nand U6526 (N_6526,N_6394,N_6308);
xnor U6527 (N_6527,N_6205,N_6347);
nor U6528 (N_6528,N_6204,N_6224);
xor U6529 (N_6529,N_6252,N_6360);
and U6530 (N_6530,N_6328,N_6220);
xor U6531 (N_6531,N_6357,N_6218);
or U6532 (N_6532,N_6313,N_6243);
xor U6533 (N_6533,N_6364,N_6253);
nand U6534 (N_6534,N_6376,N_6261);
xnor U6535 (N_6535,N_6284,N_6212);
nand U6536 (N_6536,N_6363,N_6322);
nand U6537 (N_6537,N_6387,N_6217);
and U6538 (N_6538,N_6356,N_6369);
or U6539 (N_6539,N_6338,N_6284);
nand U6540 (N_6540,N_6332,N_6203);
nor U6541 (N_6541,N_6302,N_6355);
nand U6542 (N_6542,N_6233,N_6334);
nand U6543 (N_6543,N_6340,N_6200);
or U6544 (N_6544,N_6286,N_6236);
nor U6545 (N_6545,N_6245,N_6278);
nand U6546 (N_6546,N_6323,N_6251);
nor U6547 (N_6547,N_6322,N_6202);
and U6548 (N_6548,N_6296,N_6398);
nor U6549 (N_6549,N_6262,N_6254);
nor U6550 (N_6550,N_6354,N_6267);
or U6551 (N_6551,N_6278,N_6275);
and U6552 (N_6552,N_6396,N_6295);
xor U6553 (N_6553,N_6388,N_6281);
and U6554 (N_6554,N_6268,N_6214);
nand U6555 (N_6555,N_6347,N_6274);
xnor U6556 (N_6556,N_6213,N_6260);
or U6557 (N_6557,N_6299,N_6228);
and U6558 (N_6558,N_6375,N_6326);
and U6559 (N_6559,N_6212,N_6380);
or U6560 (N_6560,N_6308,N_6241);
or U6561 (N_6561,N_6328,N_6359);
nor U6562 (N_6562,N_6223,N_6213);
or U6563 (N_6563,N_6326,N_6233);
nand U6564 (N_6564,N_6256,N_6210);
xnor U6565 (N_6565,N_6357,N_6274);
nor U6566 (N_6566,N_6276,N_6252);
or U6567 (N_6567,N_6341,N_6364);
nand U6568 (N_6568,N_6348,N_6253);
and U6569 (N_6569,N_6309,N_6278);
nor U6570 (N_6570,N_6329,N_6353);
nor U6571 (N_6571,N_6296,N_6229);
xor U6572 (N_6572,N_6376,N_6391);
xor U6573 (N_6573,N_6237,N_6236);
xnor U6574 (N_6574,N_6275,N_6249);
or U6575 (N_6575,N_6378,N_6222);
nand U6576 (N_6576,N_6206,N_6267);
nand U6577 (N_6577,N_6349,N_6385);
and U6578 (N_6578,N_6247,N_6257);
xor U6579 (N_6579,N_6310,N_6325);
or U6580 (N_6580,N_6200,N_6278);
and U6581 (N_6581,N_6258,N_6366);
nand U6582 (N_6582,N_6283,N_6248);
xnor U6583 (N_6583,N_6272,N_6318);
and U6584 (N_6584,N_6294,N_6339);
nor U6585 (N_6585,N_6348,N_6214);
nor U6586 (N_6586,N_6250,N_6341);
nor U6587 (N_6587,N_6282,N_6273);
and U6588 (N_6588,N_6393,N_6348);
nand U6589 (N_6589,N_6367,N_6214);
or U6590 (N_6590,N_6343,N_6216);
nor U6591 (N_6591,N_6297,N_6267);
and U6592 (N_6592,N_6368,N_6276);
or U6593 (N_6593,N_6237,N_6258);
xnor U6594 (N_6594,N_6284,N_6293);
xnor U6595 (N_6595,N_6311,N_6362);
nor U6596 (N_6596,N_6218,N_6361);
or U6597 (N_6597,N_6237,N_6260);
and U6598 (N_6598,N_6378,N_6216);
nor U6599 (N_6599,N_6392,N_6321);
or U6600 (N_6600,N_6553,N_6401);
or U6601 (N_6601,N_6423,N_6531);
nor U6602 (N_6602,N_6432,N_6441);
nor U6603 (N_6603,N_6546,N_6521);
nand U6604 (N_6604,N_6417,N_6422);
nand U6605 (N_6605,N_6576,N_6438);
nor U6606 (N_6606,N_6545,N_6475);
or U6607 (N_6607,N_6437,N_6523);
or U6608 (N_6608,N_6565,N_6416);
or U6609 (N_6609,N_6492,N_6402);
and U6610 (N_6610,N_6486,N_6427);
nand U6611 (N_6611,N_6506,N_6453);
nor U6612 (N_6612,N_6561,N_6590);
xor U6613 (N_6613,N_6493,N_6562);
xor U6614 (N_6614,N_6413,N_6483);
nor U6615 (N_6615,N_6579,N_6444);
and U6616 (N_6616,N_6518,N_6514);
or U6617 (N_6617,N_6405,N_6505);
nand U6618 (N_6618,N_6460,N_6587);
and U6619 (N_6619,N_6508,N_6522);
nor U6620 (N_6620,N_6410,N_6425);
xnor U6621 (N_6621,N_6429,N_6472);
xnor U6622 (N_6622,N_6498,N_6554);
or U6623 (N_6623,N_6501,N_6516);
and U6624 (N_6624,N_6428,N_6591);
nor U6625 (N_6625,N_6434,N_6465);
xnor U6626 (N_6626,N_6584,N_6491);
xor U6627 (N_6627,N_6448,N_6536);
and U6628 (N_6628,N_6489,N_6552);
nor U6629 (N_6629,N_6527,N_6400);
or U6630 (N_6630,N_6403,N_6462);
xor U6631 (N_6631,N_6577,N_6412);
and U6632 (N_6632,N_6459,N_6450);
xor U6633 (N_6633,N_6513,N_6586);
nor U6634 (N_6634,N_6494,N_6535);
or U6635 (N_6635,N_6469,N_6511);
or U6636 (N_6636,N_6481,N_6426);
nor U6637 (N_6637,N_6502,N_6454);
nand U6638 (N_6638,N_6558,N_6446);
xnor U6639 (N_6639,N_6408,N_6443);
and U6640 (N_6640,N_6431,N_6592);
and U6641 (N_6641,N_6588,N_6497);
or U6642 (N_6642,N_6598,N_6550);
or U6643 (N_6643,N_6537,N_6542);
and U6644 (N_6644,N_6524,N_6510);
xnor U6645 (N_6645,N_6503,N_6596);
nor U6646 (N_6646,N_6525,N_6530);
nor U6647 (N_6647,N_6539,N_6420);
or U6648 (N_6648,N_6534,N_6452);
xor U6649 (N_6649,N_6570,N_6582);
nor U6650 (N_6650,N_6575,N_6589);
nand U6651 (N_6651,N_6415,N_6580);
or U6652 (N_6652,N_6517,N_6433);
or U6653 (N_6653,N_6519,N_6419);
nand U6654 (N_6654,N_6543,N_6585);
and U6655 (N_6655,N_6477,N_6457);
nor U6656 (N_6656,N_6512,N_6468);
and U6657 (N_6657,N_6541,N_6532);
xor U6658 (N_6658,N_6440,N_6476);
xor U6659 (N_6659,N_6424,N_6557);
nor U6660 (N_6660,N_6466,N_6567);
nand U6661 (N_6661,N_6583,N_6571);
and U6662 (N_6662,N_6555,N_6464);
and U6663 (N_6663,N_6436,N_6411);
nand U6664 (N_6664,N_6574,N_6406);
nand U6665 (N_6665,N_6495,N_6509);
xor U6666 (N_6666,N_6533,N_6445);
and U6667 (N_6667,N_6463,N_6487);
nor U6668 (N_6668,N_6479,N_6549);
nor U6669 (N_6669,N_6482,N_6520);
and U6670 (N_6670,N_6409,N_6488);
nand U6671 (N_6671,N_6581,N_6439);
and U6672 (N_6672,N_6451,N_6594);
or U6673 (N_6673,N_6499,N_6507);
and U6674 (N_6674,N_6564,N_6544);
xnor U6675 (N_6675,N_6490,N_6430);
or U6676 (N_6676,N_6559,N_6461);
or U6677 (N_6677,N_6421,N_6560);
xor U6678 (N_6678,N_6458,N_6569);
or U6679 (N_6679,N_6547,N_6485);
or U6680 (N_6680,N_6526,N_6528);
xor U6681 (N_6681,N_6566,N_6573);
xnor U6682 (N_6682,N_6414,N_6504);
or U6683 (N_6683,N_6470,N_6540);
and U6684 (N_6684,N_6404,N_6456);
or U6685 (N_6685,N_6480,N_6529);
and U6686 (N_6686,N_6474,N_6551);
xnor U6687 (N_6687,N_6548,N_6449);
nand U6688 (N_6688,N_6478,N_6563);
nor U6689 (N_6689,N_6407,N_6435);
or U6690 (N_6690,N_6572,N_6442);
or U6691 (N_6691,N_6500,N_6595);
nand U6692 (N_6692,N_6568,N_6515);
or U6693 (N_6693,N_6538,N_6484);
xor U6694 (N_6694,N_6455,N_6473);
or U6695 (N_6695,N_6599,N_6471);
nand U6696 (N_6696,N_6447,N_6578);
or U6697 (N_6697,N_6418,N_6467);
xor U6698 (N_6698,N_6593,N_6496);
and U6699 (N_6699,N_6597,N_6556);
nand U6700 (N_6700,N_6445,N_6454);
and U6701 (N_6701,N_6585,N_6547);
or U6702 (N_6702,N_6508,N_6575);
or U6703 (N_6703,N_6442,N_6430);
or U6704 (N_6704,N_6513,N_6512);
xor U6705 (N_6705,N_6538,N_6592);
nor U6706 (N_6706,N_6474,N_6564);
nor U6707 (N_6707,N_6591,N_6518);
or U6708 (N_6708,N_6563,N_6499);
nand U6709 (N_6709,N_6448,N_6417);
or U6710 (N_6710,N_6497,N_6453);
nor U6711 (N_6711,N_6469,N_6422);
nand U6712 (N_6712,N_6542,N_6516);
and U6713 (N_6713,N_6521,N_6501);
and U6714 (N_6714,N_6565,N_6507);
nor U6715 (N_6715,N_6407,N_6527);
or U6716 (N_6716,N_6472,N_6590);
nor U6717 (N_6717,N_6589,N_6418);
and U6718 (N_6718,N_6427,N_6537);
nand U6719 (N_6719,N_6455,N_6490);
and U6720 (N_6720,N_6572,N_6594);
or U6721 (N_6721,N_6447,N_6567);
nand U6722 (N_6722,N_6557,N_6515);
xnor U6723 (N_6723,N_6494,N_6577);
nand U6724 (N_6724,N_6541,N_6408);
xnor U6725 (N_6725,N_6416,N_6505);
nor U6726 (N_6726,N_6576,N_6440);
and U6727 (N_6727,N_6535,N_6520);
xor U6728 (N_6728,N_6579,N_6598);
xnor U6729 (N_6729,N_6594,N_6437);
nor U6730 (N_6730,N_6515,N_6549);
or U6731 (N_6731,N_6412,N_6576);
xor U6732 (N_6732,N_6490,N_6575);
and U6733 (N_6733,N_6423,N_6488);
xnor U6734 (N_6734,N_6493,N_6570);
nand U6735 (N_6735,N_6417,N_6509);
xnor U6736 (N_6736,N_6558,N_6426);
or U6737 (N_6737,N_6410,N_6511);
xor U6738 (N_6738,N_6418,N_6578);
nand U6739 (N_6739,N_6584,N_6524);
or U6740 (N_6740,N_6482,N_6483);
or U6741 (N_6741,N_6509,N_6546);
nor U6742 (N_6742,N_6419,N_6579);
and U6743 (N_6743,N_6415,N_6460);
and U6744 (N_6744,N_6511,N_6445);
and U6745 (N_6745,N_6510,N_6489);
or U6746 (N_6746,N_6540,N_6477);
nand U6747 (N_6747,N_6598,N_6462);
or U6748 (N_6748,N_6426,N_6422);
or U6749 (N_6749,N_6584,N_6438);
xnor U6750 (N_6750,N_6559,N_6417);
and U6751 (N_6751,N_6444,N_6470);
and U6752 (N_6752,N_6417,N_6542);
xnor U6753 (N_6753,N_6515,N_6421);
or U6754 (N_6754,N_6506,N_6560);
xnor U6755 (N_6755,N_6540,N_6400);
and U6756 (N_6756,N_6437,N_6441);
nand U6757 (N_6757,N_6523,N_6552);
nor U6758 (N_6758,N_6414,N_6527);
and U6759 (N_6759,N_6465,N_6420);
or U6760 (N_6760,N_6551,N_6562);
and U6761 (N_6761,N_6440,N_6466);
xnor U6762 (N_6762,N_6465,N_6477);
or U6763 (N_6763,N_6437,N_6402);
and U6764 (N_6764,N_6542,N_6408);
xnor U6765 (N_6765,N_6454,N_6477);
nor U6766 (N_6766,N_6566,N_6577);
or U6767 (N_6767,N_6558,N_6519);
or U6768 (N_6768,N_6560,N_6460);
nand U6769 (N_6769,N_6595,N_6466);
nor U6770 (N_6770,N_6444,N_6467);
xnor U6771 (N_6771,N_6454,N_6564);
and U6772 (N_6772,N_6551,N_6505);
and U6773 (N_6773,N_6599,N_6499);
nand U6774 (N_6774,N_6433,N_6481);
nor U6775 (N_6775,N_6404,N_6443);
and U6776 (N_6776,N_6529,N_6472);
xnor U6777 (N_6777,N_6474,N_6585);
nand U6778 (N_6778,N_6550,N_6485);
xor U6779 (N_6779,N_6457,N_6493);
xor U6780 (N_6780,N_6443,N_6516);
nand U6781 (N_6781,N_6556,N_6599);
xor U6782 (N_6782,N_6482,N_6491);
xor U6783 (N_6783,N_6586,N_6414);
xnor U6784 (N_6784,N_6539,N_6541);
and U6785 (N_6785,N_6416,N_6515);
nand U6786 (N_6786,N_6511,N_6454);
nand U6787 (N_6787,N_6518,N_6545);
xnor U6788 (N_6788,N_6544,N_6407);
xor U6789 (N_6789,N_6578,N_6570);
or U6790 (N_6790,N_6418,N_6574);
nor U6791 (N_6791,N_6462,N_6448);
nand U6792 (N_6792,N_6501,N_6528);
nand U6793 (N_6793,N_6486,N_6435);
nor U6794 (N_6794,N_6410,N_6576);
xor U6795 (N_6795,N_6542,N_6584);
or U6796 (N_6796,N_6401,N_6435);
xnor U6797 (N_6797,N_6451,N_6446);
nor U6798 (N_6798,N_6410,N_6518);
and U6799 (N_6799,N_6566,N_6518);
and U6800 (N_6800,N_6639,N_6775);
or U6801 (N_6801,N_6787,N_6681);
and U6802 (N_6802,N_6718,N_6600);
nand U6803 (N_6803,N_6697,N_6715);
nand U6804 (N_6804,N_6657,N_6680);
or U6805 (N_6805,N_6632,N_6741);
nand U6806 (N_6806,N_6769,N_6722);
or U6807 (N_6807,N_6702,N_6654);
and U6808 (N_6808,N_6713,N_6719);
and U6809 (N_6809,N_6730,N_6773);
nor U6810 (N_6810,N_6735,N_6695);
nand U6811 (N_6811,N_6688,N_6667);
or U6812 (N_6812,N_6686,N_6704);
or U6813 (N_6813,N_6646,N_6720);
nand U6814 (N_6814,N_6757,N_6669);
xnor U6815 (N_6815,N_6737,N_6601);
nand U6816 (N_6816,N_6708,N_6739);
nand U6817 (N_6817,N_6785,N_6711);
or U6818 (N_6818,N_6647,N_6649);
nand U6819 (N_6819,N_6609,N_6700);
xor U6820 (N_6820,N_6628,N_6640);
nand U6821 (N_6821,N_6738,N_6682);
nor U6822 (N_6822,N_6795,N_6659);
xnor U6823 (N_6823,N_6622,N_6666);
and U6824 (N_6824,N_6623,N_6749);
and U6825 (N_6825,N_6699,N_6652);
and U6826 (N_6826,N_6677,N_6616);
nand U6827 (N_6827,N_6793,N_6763);
and U6828 (N_6828,N_6693,N_6692);
nand U6829 (N_6829,N_6774,N_6764);
nor U6830 (N_6830,N_6798,N_6664);
xor U6831 (N_6831,N_6712,N_6629);
nand U6832 (N_6832,N_6759,N_6690);
xnor U6833 (N_6833,N_6608,N_6748);
xnor U6834 (N_6834,N_6671,N_6675);
xor U6835 (N_6835,N_6779,N_6771);
xor U6836 (N_6836,N_6750,N_6687);
and U6837 (N_6837,N_6602,N_6754);
and U6838 (N_6838,N_6613,N_6770);
nand U6839 (N_6839,N_6607,N_6625);
xnor U6840 (N_6840,N_6651,N_6620);
nand U6841 (N_6841,N_6645,N_6777);
or U6842 (N_6842,N_6752,N_6617);
or U6843 (N_6843,N_6781,N_6635);
xor U6844 (N_6844,N_6672,N_6746);
and U6845 (N_6845,N_6665,N_6604);
nand U6846 (N_6846,N_6612,N_6706);
and U6847 (N_6847,N_6791,N_6727);
xor U6848 (N_6848,N_6716,N_6728);
and U6849 (N_6849,N_6776,N_6606);
xor U6850 (N_6850,N_6734,N_6743);
nor U6851 (N_6851,N_6631,N_6627);
xnor U6852 (N_6852,N_6778,N_6767);
nor U6853 (N_6853,N_6758,N_6696);
and U6854 (N_6854,N_6709,N_6610);
nor U6855 (N_6855,N_6789,N_6618);
nor U6856 (N_6856,N_6745,N_6674);
nand U6857 (N_6857,N_6691,N_6655);
and U6858 (N_6858,N_6633,N_6661);
and U6859 (N_6859,N_6755,N_6637);
nand U6860 (N_6860,N_6783,N_6630);
xor U6861 (N_6861,N_6796,N_6685);
and U6862 (N_6862,N_6799,N_6698);
nor U6863 (N_6863,N_6644,N_6642);
xnor U6864 (N_6864,N_6772,N_6723);
nand U6865 (N_6865,N_6615,N_6760);
and U6866 (N_6866,N_6694,N_6673);
or U6867 (N_6867,N_6721,N_6753);
or U6868 (N_6868,N_6683,N_6689);
or U6869 (N_6869,N_6786,N_6624);
nand U6870 (N_6870,N_6762,N_6705);
nor U6871 (N_6871,N_6648,N_6614);
xnor U6872 (N_6872,N_6756,N_6660);
nor U6873 (N_6873,N_6643,N_6788);
nand U6874 (N_6874,N_6679,N_6792);
nand U6875 (N_6875,N_6794,N_6658);
and U6876 (N_6876,N_6668,N_6650);
nand U6877 (N_6877,N_6780,N_6731);
xnor U6878 (N_6878,N_6670,N_6656);
xor U6879 (N_6879,N_6747,N_6605);
nand U6880 (N_6880,N_6678,N_6736);
xnor U6881 (N_6881,N_6765,N_6684);
and U6882 (N_6882,N_6790,N_6611);
or U6883 (N_6883,N_6663,N_6751);
nor U6884 (N_6884,N_6621,N_6724);
nand U6885 (N_6885,N_6634,N_6784);
nor U6886 (N_6886,N_6703,N_6729);
xnor U6887 (N_6887,N_6768,N_6714);
or U6888 (N_6888,N_6653,N_6732);
nand U6889 (N_6889,N_6707,N_6726);
nand U6890 (N_6890,N_6638,N_6797);
xor U6891 (N_6891,N_6744,N_6742);
xnor U6892 (N_6892,N_6636,N_6662);
or U6893 (N_6893,N_6710,N_6626);
nand U6894 (N_6894,N_6725,N_6766);
and U6895 (N_6895,N_6782,N_6740);
or U6896 (N_6896,N_6619,N_6761);
nand U6897 (N_6897,N_6717,N_6733);
nand U6898 (N_6898,N_6641,N_6701);
or U6899 (N_6899,N_6603,N_6676);
and U6900 (N_6900,N_6605,N_6628);
nor U6901 (N_6901,N_6663,N_6792);
xor U6902 (N_6902,N_6666,N_6687);
or U6903 (N_6903,N_6792,N_6754);
nor U6904 (N_6904,N_6761,N_6748);
nand U6905 (N_6905,N_6658,N_6673);
or U6906 (N_6906,N_6676,N_6766);
nor U6907 (N_6907,N_6741,N_6776);
and U6908 (N_6908,N_6661,N_6788);
and U6909 (N_6909,N_6627,N_6633);
or U6910 (N_6910,N_6791,N_6709);
and U6911 (N_6911,N_6769,N_6703);
xnor U6912 (N_6912,N_6753,N_6637);
and U6913 (N_6913,N_6795,N_6663);
or U6914 (N_6914,N_6657,N_6638);
xor U6915 (N_6915,N_6791,N_6666);
nor U6916 (N_6916,N_6652,N_6736);
xnor U6917 (N_6917,N_6689,N_6785);
nand U6918 (N_6918,N_6609,N_6725);
nor U6919 (N_6919,N_6675,N_6655);
or U6920 (N_6920,N_6635,N_6710);
xnor U6921 (N_6921,N_6775,N_6604);
or U6922 (N_6922,N_6760,N_6748);
nand U6923 (N_6923,N_6690,N_6720);
or U6924 (N_6924,N_6735,N_6625);
xnor U6925 (N_6925,N_6757,N_6622);
and U6926 (N_6926,N_6665,N_6721);
nor U6927 (N_6927,N_6727,N_6709);
xor U6928 (N_6928,N_6722,N_6620);
and U6929 (N_6929,N_6738,N_6705);
nor U6930 (N_6930,N_6668,N_6712);
nor U6931 (N_6931,N_6601,N_6627);
and U6932 (N_6932,N_6664,N_6625);
nand U6933 (N_6933,N_6700,N_6706);
and U6934 (N_6934,N_6658,N_6785);
nor U6935 (N_6935,N_6714,N_6653);
or U6936 (N_6936,N_6680,N_6769);
or U6937 (N_6937,N_6605,N_6743);
and U6938 (N_6938,N_6751,N_6672);
or U6939 (N_6939,N_6631,N_6622);
nand U6940 (N_6940,N_6648,N_6788);
xor U6941 (N_6941,N_6653,N_6665);
xnor U6942 (N_6942,N_6607,N_6792);
and U6943 (N_6943,N_6751,N_6616);
and U6944 (N_6944,N_6627,N_6771);
and U6945 (N_6945,N_6750,N_6786);
and U6946 (N_6946,N_6627,N_6630);
or U6947 (N_6947,N_6606,N_6631);
nand U6948 (N_6948,N_6709,N_6638);
xor U6949 (N_6949,N_6671,N_6693);
nor U6950 (N_6950,N_6757,N_6793);
nor U6951 (N_6951,N_6621,N_6654);
or U6952 (N_6952,N_6617,N_6600);
nor U6953 (N_6953,N_6689,N_6730);
nand U6954 (N_6954,N_6728,N_6665);
nor U6955 (N_6955,N_6623,N_6767);
nand U6956 (N_6956,N_6631,N_6725);
nor U6957 (N_6957,N_6619,N_6744);
or U6958 (N_6958,N_6775,N_6621);
xnor U6959 (N_6959,N_6761,N_6692);
and U6960 (N_6960,N_6732,N_6613);
and U6961 (N_6961,N_6639,N_6681);
xnor U6962 (N_6962,N_6611,N_6704);
or U6963 (N_6963,N_6641,N_6736);
or U6964 (N_6964,N_6614,N_6735);
nor U6965 (N_6965,N_6663,N_6693);
nor U6966 (N_6966,N_6782,N_6724);
xnor U6967 (N_6967,N_6774,N_6716);
xor U6968 (N_6968,N_6689,N_6663);
nor U6969 (N_6969,N_6600,N_6723);
and U6970 (N_6970,N_6723,N_6742);
xor U6971 (N_6971,N_6635,N_6715);
nand U6972 (N_6972,N_6712,N_6660);
and U6973 (N_6973,N_6776,N_6674);
xnor U6974 (N_6974,N_6740,N_6771);
and U6975 (N_6975,N_6685,N_6629);
xor U6976 (N_6976,N_6798,N_6715);
and U6977 (N_6977,N_6768,N_6639);
and U6978 (N_6978,N_6628,N_6657);
nand U6979 (N_6979,N_6726,N_6656);
nor U6980 (N_6980,N_6738,N_6715);
nor U6981 (N_6981,N_6701,N_6728);
xnor U6982 (N_6982,N_6714,N_6799);
nor U6983 (N_6983,N_6677,N_6718);
and U6984 (N_6984,N_6661,N_6699);
xor U6985 (N_6985,N_6699,N_6768);
or U6986 (N_6986,N_6732,N_6769);
xnor U6987 (N_6987,N_6769,N_6767);
nand U6988 (N_6988,N_6616,N_6716);
nor U6989 (N_6989,N_6735,N_6731);
and U6990 (N_6990,N_6727,N_6641);
or U6991 (N_6991,N_6723,N_6765);
nor U6992 (N_6992,N_6611,N_6771);
and U6993 (N_6993,N_6664,N_6648);
and U6994 (N_6994,N_6753,N_6715);
nor U6995 (N_6995,N_6608,N_6756);
and U6996 (N_6996,N_6771,N_6767);
nand U6997 (N_6997,N_6672,N_6645);
xor U6998 (N_6998,N_6607,N_6618);
and U6999 (N_6999,N_6675,N_6742);
and U7000 (N_7000,N_6988,N_6834);
or U7001 (N_7001,N_6958,N_6804);
xor U7002 (N_7002,N_6817,N_6816);
nor U7003 (N_7003,N_6904,N_6927);
nand U7004 (N_7004,N_6897,N_6812);
xor U7005 (N_7005,N_6819,N_6860);
xnor U7006 (N_7006,N_6990,N_6872);
or U7007 (N_7007,N_6923,N_6846);
nand U7008 (N_7008,N_6915,N_6828);
nand U7009 (N_7009,N_6801,N_6971);
or U7010 (N_7010,N_6924,N_6840);
or U7011 (N_7011,N_6826,N_6864);
and U7012 (N_7012,N_6965,N_6818);
and U7013 (N_7013,N_6913,N_6909);
xor U7014 (N_7014,N_6926,N_6903);
and U7015 (N_7015,N_6972,N_6942);
nand U7016 (N_7016,N_6966,N_6961);
nor U7017 (N_7017,N_6914,N_6922);
and U7018 (N_7018,N_6892,N_6833);
nand U7019 (N_7019,N_6813,N_6898);
nand U7020 (N_7020,N_6824,N_6959);
xor U7021 (N_7021,N_6889,N_6825);
and U7022 (N_7022,N_6882,N_6838);
or U7023 (N_7023,N_6934,N_6861);
and U7024 (N_7024,N_6820,N_6932);
and U7025 (N_7025,N_6970,N_6830);
nand U7026 (N_7026,N_6953,N_6930);
or U7027 (N_7027,N_6806,N_6983);
and U7028 (N_7028,N_6906,N_6876);
and U7029 (N_7029,N_6852,N_6854);
nand U7030 (N_7030,N_6979,N_6902);
or U7031 (N_7031,N_6803,N_6884);
and U7032 (N_7032,N_6935,N_6885);
nand U7033 (N_7033,N_6862,N_6811);
nor U7034 (N_7034,N_6880,N_6982);
nand U7035 (N_7035,N_6821,N_6920);
xnor U7036 (N_7036,N_6807,N_6955);
nor U7037 (N_7037,N_6916,N_6857);
nand U7038 (N_7038,N_6962,N_6814);
nand U7039 (N_7039,N_6877,N_6874);
nand U7040 (N_7040,N_6900,N_6928);
nand U7041 (N_7041,N_6985,N_6967);
or U7042 (N_7042,N_6951,N_6858);
xnor U7043 (N_7043,N_6946,N_6894);
nor U7044 (N_7044,N_6978,N_6919);
xor U7045 (N_7045,N_6866,N_6936);
or U7046 (N_7046,N_6869,N_6856);
and U7047 (N_7047,N_6998,N_6851);
and U7048 (N_7048,N_6981,N_6855);
nor U7049 (N_7049,N_6917,N_6865);
xor U7050 (N_7050,N_6954,N_6957);
nor U7051 (N_7051,N_6960,N_6837);
nand U7052 (N_7052,N_6938,N_6950);
nor U7053 (N_7053,N_6994,N_6890);
or U7054 (N_7054,N_6879,N_6931);
xnor U7055 (N_7055,N_6996,N_6829);
nand U7056 (N_7056,N_6963,N_6842);
nor U7057 (N_7057,N_6991,N_6808);
and U7058 (N_7058,N_6964,N_6883);
or U7059 (N_7059,N_6896,N_6943);
nor U7060 (N_7060,N_6873,N_6997);
xnor U7061 (N_7061,N_6831,N_6944);
xnor U7062 (N_7062,N_6845,N_6976);
xnor U7063 (N_7063,N_6918,N_6952);
and U7064 (N_7064,N_6929,N_6867);
nand U7065 (N_7065,N_6899,N_6989);
xnor U7066 (N_7066,N_6868,N_6878);
nor U7067 (N_7067,N_6800,N_6945);
nor U7068 (N_7068,N_6980,N_6937);
or U7069 (N_7069,N_6810,N_6893);
xnor U7070 (N_7070,N_6901,N_6939);
nor U7071 (N_7071,N_6984,N_6999);
nand U7072 (N_7072,N_6948,N_6870);
or U7073 (N_7073,N_6847,N_6925);
nand U7074 (N_7074,N_6891,N_6908);
or U7075 (N_7075,N_6895,N_6859);
nand U7076 (N_7076,N_6836,N_6987);
xor U7077 (N_7077,N_6995,N_6905);
or U7078 (N_7078,N_6827,N_6968);
nor U7079 (N_7079,N_6823,N_6841);
nor U7080 (N_7080,N_6956,N_6992);
nand U7081 (N_7081,N_6853,N_6940);
and U7082 (N_7082,N_6973,N_6993);
and U7083 (N_7083,N_6912,N_6977);
or U7084 (N_7084,N_6822,N_6875);
nand U7085 (N_7085,N_6907,N_6911);
or U7086 (N_7086,N_6835,N_6832);
nor U7087 (N_7087,N_6815,N_6933);
nand U7088 (N_7088,N_6941,N_6843);
and U7089 (N_7089,N_6809,N_6850);
nor U7090 (N_7090,N_6986,N_6844);
or U7091 (N_7091,N_6805,N_6921);
xnor U7092 (N_7092,N_6975,N_6871);
or U7093 (N_7093,N_6887,N_6881);
nand U7094 (N_7094,N_6969,N_6863);
xor U7095 (N_7095,N_6839,N_6910);
nor U7096 (N_7096,N_6886,N_6974);
or U7097 (N_7097,N_6949,N_6888);
xor U7098 (N_7098,N_6802,N_6848);
nor U7099 (N_7099,N_6849,N_6947);
or U7100 (N_7100,N_6881,N_6950);
nor U7101 (N_7101,N_6904,N_6995);
xnor U7102 (N_7102,N_6959,N_6843);
nand U7103 (N_7103,N_6872,N_6993);
or U7104 (N_7104,N_6841,N_6992);
nor U7105 (N_7105,N_6920,N_6940);
nand U7106 (N_7106,N_6867,N_6950);
and U7107 (N_7107,N_6870,N_6803);
nand U7108 (N_7108,N_6930,N_6815);
or U7109 (N_7109,N_6805,N_6909);
nor U7110 (N_7110,N_6810,N_6827);
and U7111 (N_7111,N_6858,N_6888);
nand U7112 (N_7112,N_6830,N_6938);
xnor U7113 (N_7113,N_6897,N_6880);
and U7114 (N_7114,N_6821,N_6989);
nand U7115 (N_7115,N_6884,N_6909);
nand U7116 (N_7116,N_6860,N_6861);
nand U7117 (N_7117,N_6841,N_6910);
xnor U7118 (N_7118,N_6931,N_6952);
nand U7119 (N_7119,N_6999,N_6839);
and U7120 (N_7120,N_6984,N_6986);
and U7121 (N_7121,N_6836,N_6924);
xnor U7122 (N_7122,N_6873,N_6944);
nand U7123 (N_7123,N_6990,N_6800);
nand U7124 (N_7124,N_6845,N_6811);
nor U7125 (N_7125,N_6981,N_6873);
xor U7126 (N_7126,N_6993,N_6986);
nor U7127 (N_7127,N_6993,N_6867);
and U7128 (N_7128,N_6817,N_6928);
nor U7129 (N_7129,N_6875,N_6836);
and U7130 (N_7130,N_6808,N_6996);
nand U7131 (N_7131,N_6863,N_6899);
xnor U7132 (N_7132,N_6927,N_6928);
xor U7133 (N_7133,N_6903,N_6938);
nor U7134 (N_7134,N_6996,N_6948);
nand U7135 (N_7135,N_6831,N_6858);
nand U7136 (N_7136,N_6892,N_6949);
and U7137 (N_7137,N_6886,N_6986);
or U7138 (N_7138,N_6999,N_6838);
nand U7139 (N_7139,N_6835,N_6913);
nand U7140 (N_7140,N_6974,N_6968);
xor U7141 (N_7141,N_6919,N_6990);
and U7142 (N_7142,N_6880,N_6875);
nor U7143 (N_7143,N_6801,N_6992);
nor U7144 (N_7144,N_6977,N_6816);
or U7145 (N_7145,N_6892,N_6845);
nor U7146 (N_7146,N_6974,N_6955);
nand U7147 (N_7147,N_6993,N_6802);
nor U7148 (N_7148,N_6902,N_6930);
xor U7149 (N_7149,N_6882,N_6808);
and U7150 (N_7150,N_6954,N_6900);
nor U7151 (N_7151,N_6944,N_6940);
and U7152 (N_7152,N_6866,N_6855);
or U7153 (N_7153,N_6901,N_6921);
nor U7154 (N_7154,N_6920,N_6859);
and U7155 (N_7155,N_6926,N_6806);
or U7156 (N_7156,N_6863,N_6904);
nor U7157 (N_7157,N_6841,N_6869);
or U7158 (N_7158,N_6936,N_6880);
nand U7159 (N_7159,N_6918,N_6925);
nand U7160 (N_7160,N_6854,N_6824);
xor U7161 (N_7161,N_6922,N_6982);
or U7162 (N_7162,N_6977,N_6902);
nor U7163 (N_7163,N_6901,N_6883);
or U7164 (N_7164,N_6994,N_6842);
nor U7165 (N_7165,N_6959,N_6857);
xor U7166 (N_7166,N_6958,N_6982);
nor U7167 (N_7167,N_6973,N_6953);
nor U7168 (N_7168,N_6983,N_6951);
and U7169 (N_7169,N_6980,N_6929);
or U7170 (N_7170,N_6929,N_6936);
nor U7171 (N_7171,N_6831,N_6974);
nor U7172 (N_7172,N_6802,N_6849);
nand U7173 (N_7173,N_6860,N_6879);
nand U7174 (N_7174,N_6809,N_6937);
nand U7175 (N_7175,N_6963,N_6979);
xnor U7176 (N_7176,N_6922,N_6843);
or U7177 (N_7177,N_6852,N_6897);
nand U7178 (N_7178,N_6904,N_6854);
and U7179 (N_7179,N_6947,N_6884);
nand U7180 (N_7180,N_6875,N_6971);
and U7181 (N_7181,N_6859,N_6886);
nor U7182 (N_7182,N_6902,N_6990);
or U7183 (N_7183,N_6992,N_6888);
or U7184 (N_7184,N_6873,N_6850);
nor U7185 (N_7185,N_6809,N_6888);
or U7186 (N_7186,N_6953,N_6830);
nor U7187 (N_7187,N_6883,N_6993);
nand U7188 (N_7188,N_6999,N_6965);
xor U7189 (N_7189,N_6946,N_6925);
nand U7190 (N_7190,N_6979,N_6921);
nand U7191 (N_7191,N_6968,N_6858);
nor U7192 (N_7192,N_6995,N_6816);
nor U7193 (N_7193,N_6899,N_6957);
xor U7194 (N_7194,N_6930,N_6841);
and U7195 (N_7195,N_6976,N_6888);
or U7196 (N_7196,N_6848,N_6973);
xor U7197 (N_7197,N_6839,N_6835);
and U7198 (N_7198,N_6969,N_6914);
nor U7199 (N_7199,N_6916,N_6840);
nand U7200 (N_7200,N_7121,N_7046);
xor U7201 (N_7201,N_7105,N_7045);
or U7202 (N_7202,N_7119,N_7107);
and U7203 (N_7203,N_7135,N_7021);
or U7204 (N_7204,N_7130,N_7096);
or U7205 (N_7205,N_7133,N_7132);
nor U7206 (N_7206,N_7145,N_7093);
nand U7207 (N_7207,N_7103,N_7089);
nor U7208 (N_7208,N_7175,N_7193);
nor U7209 (N_7209,N_7012,N_7087);
nor U7210 (N_7210,N_7056,N_7188);
or U7211 (N_7211,N_7165,N_7110);
nor U7212 (N_7212,N_7034,N_7125);
nand U7213 (N_7213,N_7051,N_7078);
nand U7214 (N_7214,N_7083,N_7088);
and U7215 (N_7215,N_7134,N_7163);
nand U7216 (N_7216,N_7049,N_7111);
xor U7217 (N_7217,N_7167,N_7147);
nor U7218 (N_7218,N_7116,N_7137);
or U7219 (N_7219,N_7194,N_7108);
or U7220 (N_7220,N_7024,N_7029);
nand U7221 (N_7221,N_7126,N_7003);
or U7222 (N_7222,N_7198,N_7037);
nor U7223 (N_7223,N_7157,N_7118);
xnor U7224 (N_7224,N_7138,N_7004);
or U7225 (N_7225,N_7187,N_7054);
nand U7226 (N_7226,N_7176,N_7074);
nand U7227 (N_7227,N_7086,N_7191);
xnor U7228 (N_7228,N_7057,N_7189);
and U7229 (N_7229,N_7031,N_7178);
xnor U7230 (N_7230,N_7166,N_7060);
xor U7231 (N_7231,N_7052,N_7000);
nand U7232 (N_7232,N_7018,N_7156);
and U7233 (N_7233,N_7101,N_7035);
and U7234 (N_7234,N_7186,N_7079);
and U7235 (N_7235,N_7028,N_7128);
nor U7236 (N_7236,N_7124,N_7162);
nand U7237 (N_7237,N_7122,N_7113);
nor U7238 (N_7238,N_7071,N_7141);
or U7239 (N_7239,N_7170,N_7183);
or U7240 (N_7240,N_7005,N_7123);
and U7241 (N_7241,N_7195,N_7177);
and U7242 (N_7242,N_7050,N_7097);
xor U7243 (N_7243,N_7104,N_7181);
or U7244 (N_7244,N_7025,N_7013);
nand U7245 (N_7245,N_7055,N_7064);
nand U7246 (N_7246,N_7047,N_7171);
xnor U7247 (N_7247,N_7069,N_7102);
nor U7248 (N_7248,N_7146,N_7072);
xor U7249 (N_7249,N_7155,N_7148);
nand U7250 (N_7250,N_7094,N_7184);
nand U7251 (N_7251,N_7042,N_7112);
and U7252 (N_7252,N_7150,N_7010);
or U7253 (N_7253,N_7182,N_7164);
and U7254 (N_7254,N_7076,N_7061);
and U7255 (N_7255,N_7041,N_7063);
and U7256 (N_7256,N_7048,N_7023);
or U7257 (N_7257,N_7196,N_7077);
xnor U7258 (N_7258,N_7019,N_7039);
nand U7259 (N_7259,N_7106,N_7082);
nand U7260 (N_7260,N_7115,N_7142);
and U7261 (N_7261,N_7179,N_7009);
nor U7262 (N_7262,N_7090,N_7006);
or U7263 (N_7263,N_7015,N_7199);
nor U7264 (N_7264,N_7100,N_7151);
or U7265 (N_7265,N_7016,N_7131);
and U7266 (N_7266,N_7030,N_7085);
nand U7267 (N_7267,N_7092,N_7068);
or U7268 (N_7268,N_7169,N_7058);
nor U7269 (N_7269,N_7185,N_7020);
and U7270 (N_7270,N_7190,N_7140);
and U7271 (N_7271,N_7008,N_7152);
nor U7272 (N_7272,N_7027,N_7053);
or U7273 (N_7273,N_7109,N_7129);
xor U7274 (N_7274,N_7014,N_7043);
or U7275 (N_7275,N_7059,N_7022);
xnor U7276 (N_7276,N_7066,N_7036);
and U7277 (N_7277,N_7011,N_7172);
nor U7278 (N_7278,N_7174,N_7007);
nand U7279 (N_7279,N_7192,N_7091);
nand U7280 (N_7280,N_7017,N_7026);
nand U7281 (N_7281,N_7197,N_7154);
and U7282 (N_7282,N_7099,N_7158);
xor U7283 (N_7283,N_7001,N_7065);
xnor U7284 (N_7284,N_7084,N_7002);
and U7285 (N_7285,N_7161,N_7139);
and U7286 (N_7286,N_7143,N_7044);
nand U7287 (N_7287,N_7038,N_7160);
or U7288 (N_7288,N_7098,N_7127);
xor U7289 (N_7289,N_7153,N_7062);
xnor U7290 (N_7290,N_7180,N_7073);
and U7291 (N_7291,N_7032,N_7159);
or U7292 (N_7292,N_7075,N_7033);
nand U7293 (N_7293,N_7040,N_7120);
and U7294 (N_7294,N_7117,N_7136);
and U7295 (N_7295,N_7114,N_7080);
and U7296 (N_7296,N_7067,N_7144);
xnor U7297 (N_7297,N_7081,N_7070);
or U7298 (N_7298,N_7173,N_7168);
nand U7299 (N_7299,N_7149,N_7095);
nand U7300 (N_7300,N_7081,N_7026);
xnor U7301 (N_7301,N_7010,N_7160);
nand U7302 (N_7302,N_7054,N_7089);
nor U7303 (N_7303,N_7073,N_7129);
or U7304 (N_7304,N_7065,N_7105);
and U7305 (N_7305,N_7157,N_7043);
xnor U7306 (N_7306,N_7049,N_7195);
and U7307 (N_7307,N_7059,N_7026);
or U7308 (N_7308,N_7147,N_7045);
xor U7309 (N_7309,N_7034,N_7102);
xnor U7310 (N_7310,N_7021,N_7140);
or U7311 (N_7311,N_7043,N_7171);
and U7312 (N_7312,N_7166,N_7044);
nor U7313 (N_7313,N_7055,N_7114);
nor U7314 (N_7314,N_7074,N_7160);
xor U7315 (N_7315,N_7178,N_7174);
and U7316 (N_7316,N_7028,N_7041);
nor U7317 (N_7317,N_7071,N_7119);
and U7318 (N_7318,N_7114,N_7189);
xnor U7319 (N_7319,N_7187,N_7024);
or U7320 (N_7320,N_7132,N_7084);
nand U7321 (N_7321,N_7158,N_7169);
nor U7322 (N_7322,N_7161,N_7107);
nor U7323 (N_7323,N_7198,N_7081);
nor U7324 (N_7324,N_7049,N_7157);
nand U7325 (N_7325,N_7104,N_7057);
and U7326 (N_7326,N_7017,N_7149);
xnor U7327 (N_7327,N_7165,N_7075);
nand U7328 (N_7328,N_7110,N_7072);
and U7329 (N_7329,N_7127,N_7173);
or U7330 (N_7330,N_7012,N_7199);
nor U7331 (N_7331,N_7102,N_7014);
or U7332 (N_7332,N_7187,N_7059);
and U7333 (N_7333,N_7156,N_7080);
nor U7334 (N_7334,N_7031,N_7198);
xor U7335 (N_7335,N_7188,N_7103);
xnor U7336 (N_7336,N_7117,N_7077);
nand U7337 (N_7337,N_7139,N_7166);
nand U7338 (N_7338,N_7026,N_7148);
and U7339 (N_7339,N_7150,N_7104);
and U7340 (N_7340,N_7191,N_7048);
nand U7341 (N_7341,N_7016,N_7021);
nand U7342 (N_7342,N_7122,N_7179);
nor U7343 (N_7343,N_7179,N_7056);
nand U7344 (N_7344,N_7191,N_7097);
and U7345 (N_7345,N_7116,N_7068);
nor U7346 (N_7346,N_7116,N_7060);
nor U7347 (N_7347,N_7170,N_7031);
xor U7348 (N_7348,N_7040,N_7145);
and U7349 (N_7349,N_7177,N_7182);
xnor U7350 (N_7350,N_7011,N_7085);
and U7351 (N_7351,N_7045,N_7053);
nor U7352 (N_7352,N_7045,N_7082);
nand U7353 (N_7353,N_7090,N_7092);
nand U7354 (N_7354,N_7119,N_7095);
nor U7355 (N_7355,N_7173,N_7181);
nor U7356 (N_7356,N_7003,N_7018);
nor U7357 (N_7357,N_7198,N_7118);
or U7358 (N_7358,N_7023,N_7173);
and U7359 (N_7359,N_7167,N_7133);
or U7360 (N_7360,N_7095,N_7072);
or U7361 (N_7361,N_7164,N_7157);
or U7362 (N_7362,N_7183,N_7132);
nor U7363 (N_7363,N_7012,N_7194);
xor U7364 (N_7364,N_7150,N_7094);
nor U7365 (N_7365,N_7130,N_7154);
and U7366 (N_7366,N_7157,N_7171);
nor U7367 (N_7367,N_7182,N_7093);
or U7368 (N_7368,N_7103,N_7105);
nor U7369 (N_7369,N_7144,N_7145);
xnor U7370 (N_7370,N_7140,N_7029);
or U7371 (N_7371,N_7102,N_7039);
or U7372 (N_7372,N_7111,N_7155);
or U7373 (N_7373,N_7027,N_7112);
or U7374 (N_7374,N_7196,N_7041);
and U7375 (N_7375,N_7041,N_7113);
nor U7376 (N_7376,N_7118,N_7025);
or U7377 (N_7377,N_7139,N_7098);
xor U7378 (N_7378,N_7162,N_7067);
or U7379 (N_7379,N_7117,N_7019);
xor U7380 (N_7380,N_7189,N_7165);
nand U7381 (N_7381,N_7134,N_7164);
nand U7382 (N_7382,N_7027,N_7116);
nor U7383 (N_7383,N_7198,N_7107);
nor U7384 (N_7384,N_7143,N_7010);
nor U7385 (N_7385,N_7040,N_7007);
nor U7386 (N_7386,N_7063,N_7154);
and U7387 (N_7387,N_7125,N_7168);
or U7388 (N_7388,N_7151,N_7197);
xnor U7389 (N_7389,N_7001,N_7130);
nand U7390 (N_7390,N_7101,N_7043);
nand U7391 (N_7391,N_7124,N_7161);
xnor U7392 (N_7392,N_7032,N_7134);
nor U7393 (N_7393,N_7126,N_7067);
xor U7394 (N_7394,N_7101,N_7139);
or U7395 (N_7395,N_7199,N_7056);
nand U7396 (N_7396,N_7087,N_7122);
or U7397 (N_7397,N_7146,N_7086);
or U7398 (N_7398,N_7009,N_7101);
xnor U7399 (N_7399,N_7133,N_7036);
or U7400 (N_7400,N_7245,N_7259);
xor U7401 (N_7401,N_7224,N_7211);
and U7402 (N_7402,N_7253,N_7237);
or U7403 (N_7403,N_7317,N_7299);
or U7404 (N_7404,N_7239,N_7229);
and U7405 (N_7405,N_7208,N_7212);
nand U7406 (N_7406,N_7355,N_7391);
nand U7407 (N_7407,N_7303,N_7236);
or U7408 (N_7408,N_7261,N_7289);
and U7409 (N_7409,N_7282,N_7241);
and U7410 (N_7410,N_7354,N_7395);
nand U7411 (N_7411,N_7337,N_7288);
nand U7412 (N_7412,N_7295,N_7364);
nor U7413 (N_7413,N_7382,N_7207);
xor U7414 (N_7414,N_7221,N_7379);
nand U7415 (N_7415,N_7359,N_7389);
nor U7416 (N_7416,N_7386,N_7269);
or U7417 (N_7417,N_7396,N_7320);
and U7418 (N_7418,N_7277,N_7248);
or U7419 (N_7419,N_7281,N_7321);
nor U7420 (N_7420,N_7352,N_7315);
or U7421 (N_7421,N_7394,N_7250);
or U7422 (N_7422,N_7305,N_7361);
xnor U7423 (N_7423,N_7216,N_7378);
and U7424 (N_7424,N_7383,N_7214);
or U7425 (N_7425,N_7209,N_7326);
nand U7426 (N_7426,N_7292,N_7205);
nand U7427 (N_7427,N_7343,N_7341);
and U7428 (N_7428,N_7369,N_7275);
and U7429 (N_7429,N_7257,N_7206);
nand U7430 (N_7430,N_7256,N_7344);
nor U7431 (N_7431,N_7234,N_7384);
nor U7432 (N_7432,N_7370,N_7294);
and U7433 (N_7433,N_7274,N_7203);
or U7434 (N_7434,N_7246,N_7254);
or U7435 (N_7435,N_7372,N_7264);
nand U7436 (N_7436,N_7346,N_7351);
or U7437 (N_7437,N_7244,N_7327);
xor U7438 (N_7438,N_7318,N_7204);
nor U7439 (N_7439,N_7243,N_7371);
xnor U7440 (N_7440,N_7381,N_7302);
nand U7441 (N_7441,N_7331,N_7278);
and U7442 (N_7442,N_7312,N_7242);
nor U7443 (N_7443,N_7251,N_7265);
xnor U7444 (N_7444,N_7268,N_7210);
or U7445 (N_7445,N_7215,N_7373);
xnor U7446 (N_7446,N_7309,N_7358);
or U7447 (N_7447,N_7388,N_7357);
nor U7448 (N_7448,N_7335,N_7376);
nand U7449 (N_7449,N_7367,N_7290);
or U7450 (N_7450,N_7284,N_7232);
xor U7451 (N_7451,N_7385,N_7200);
nand U7452 (N_7452,N_7324,N_7231);
nand U7453 (N_7453,N_7339,N_7298);
and U7454 (N_7454,N_7306,N_7249);
xnor U7455 (N_7455,N_7347,N_7398);
nor U7456 (N_7456,N_7262,N_7226);
and U7457 (N_7457,N_7283,N_7368);
nor U7458 (N_7458,N_7316,N_7301);
and U7459 (N_7459,N_7330,N_7338);
nor U7460 (N_7460,N_7310,N_7363);
or U7461 (N_7461,N_7322,N_7349);
or U7462 (N_7462,N_7300,N_7360);
and U7463 (N_7463,N_7220,N_7366);
or U7464 (N_7464,N_7266,N_7260);
and U7465 (N_7465,N_7213,N_7336);
or U7466 (N_7466,N_7225,N_7255);
xor U7467 (N_7467,N_7319,N_7293);
nand U7468 (N_7468,N_7296,N_7240);
or U7469 (N_7469,N_7285,N_7267);
nor U7470 (N_7470,N_7323,N_7247);
or U7471 (N_7471,N_7333,N_7238);
nand U7472 (N_7472,N_7202,N_7287);
xor U7473 (N_7473,N_7345,N_7365);
xnor U7474 (N_7474,N_7276,N_7392);
nand U7475 (N_7475,N_7286,N_7356);
and U7476 (N_7476,N_7328,N_7217);
nor U7477 (N_7477,N_7399,N_7227);
and U7478 (N_7478,N_7311,N_7329);
xnor U7479 (N_7479,N_7314,N_7222);
xor U7480 (N_7480,N_7334,N_7258);
nand U7481 (N_7481,N_7279,N_7350);
nor U7482 (N_7482,N_7377,N_7233);
and U7483 (N_7483,N_7397,N_7270);
nand U7484 (N_7484,N_7307,N_7228);
and U7485 (N_7485,N_7223,N_7325);
or U7486 (N_7486,N_7340,N_7374);
nand U7487 (N_7487,N_7362,N_7263);
nand U7488 (N_7488,N_7332,N_7280);
or U7489 (N_7489,N_7271,N_7218);
and U7490 (N_7490,N_7353,N_7342);
and U7491 (N_7491,N_7348,N_7230);
nor U7492 (N_7492,N_7387,N_7375);
xnor U7493 (N_7493,N_7252,N_7304);
and U7494 (N_7494,N_7291,N_7390);
xor U7495 (N_7495,N_7297,N_7235);
nor U7496 (N_7496,N_7201,N_7380);
xnor U7497 (N_7497,N_7272,N_7219);
nand U7498 (N_7498,N_7313,N_7393);
nand U7499 (N_7499,N_7308,N_7273);
or U7500 (N_7500,N_7227,N_7376);
xor U7501 (N_7501,N_7283,N_7208);
nor U7502 (N_7502,N_7332,N_7322);
or U7503 (N_7503,N_7301,N_7232);
nand U7504 (N_7504,N_7393,N_7319);
or U7505 (N_7505,N_7356,N_7208);
and U7506 (N_7506,N_7342,N_7374);
and U7507 (N_7507,N_7304,N_7371);
xnor U7508 (N_7508,N_7332,N_7350);
or U7509 (N_7509,N_7235,N_7334);
xnor U7510 (N_7510,N_7229,N_7335);
or U7511 (N_7511,N_7258,N_7221);
nand U7512 (N_7512,N_7391,N_7231);
xnor U7513 (N_7513,N_7349,N_7357);
xnor U7514 (N_7514,N_7387,N_7354);
xnor U7515 (N_7515,N_7326,N_7381);
nand U7516 (N_7516,N_7361,N_7353);
xnor U7517 (N_7517,N_7306,N_7226);
nand U7518 (N_7518,N_7283,N_7274);
and U7519 (N_7519,N_7334,N_7394);
nor U7520 (N_7520,N_7390,N_7336);
or U7521 (N_7521,N_7356,N_7370);
and U7522 (N_7522,N_7204,N_7281);
nor U7523 (N_7523,N_7379,N_7273);
or U7524 (N_7524,N_7302,N_7257);
nor U7525 (N_7525,N_7295,N_7243);
nor U7526 (N_7526,N_7281,N_7369);
and U7527 (N_7527,N_7327,N_7375);
xor U7528 (N_7528,N_7361,N_7234);
and U7529 (N_7529,N_7388,N_7224);
nand U7530 (N_7530,N_7218,N_7246);
nor U7531 (N_7531,N_7228,N_7215);
and U7532 (N_7532,N_7263,N_7389);
nor U7533 (N_7533,N_7364,N_7241);
nor U7534 (N_7534,N_7389,N_7268);
or U7535 (N_7535,N_7307,N_7352);
or U7536 (N_7536,N_7259,N_7367);
or U7537 (N_7537,N_7308,N_7327);
and U7538 (N_7538,N_7354,N_7264);
or U7539 (N_7539,N_7382,N_7251);
and U7540 (N_7540,N_7347,N_7379);
nor U7541 (N_7541,N_7369,N_7256);
nor U7542 (N_7542,N_7318,N_7392);
nor U7543 (N_7543,N_7233,N_7399);
or U7544 (N_7544,N_7357,N_7220);
nand U7545 (N_7545,N_7315,N_7218);
and U7546 (N_7546,N_7281,N_7314);
or U7547 (N_7547,N_7316,N_7318);
and U7548 (N_7548,N_7292,N_7246);
nor U7549 (N_7549,N_7373,N_7283);
and U7550 (N_7550,N_7218,N_7236);
xnor U7551 (N_7551,N_7298,N_7296);
xnor U7552 (N_7552,N_7397,N_7347);
or U7553 (N_7553,N_7200,N_7284);
xor U7554 (N_7554,N_7339,N_7376);
and U7555 (N_7555,N_7395,N_7371);
and U7556 (N_7556,N_7340,N_7376);
nand U7557 (N_7557,N_7303,N_7269);
or U7558 (N_7558,N_7314,N_7288);
and U7559 (N_7559,N_7304,N_7339);
and U7560 (N_7560,N_7285,N_7225);
nor U7561 (N_7561,N_7250,N_7265);
nand U7562 (N_7562,N_7230,N_7291);
or U7563 (N_7563,N_7264,N_7324);
nor U7564 (N_7564,N_7243,N_7396);
nand U7565 (N_7565,N_7277,N_7309);
and U7566 (N_7566,N_7347,N_7287);
nand U7567 (N_7567,N_7209,N_7337);
or U7568 (N_7568,N_7218,N_7329);
xnor U7569 (N_7569,N_7290,N_7364);
nor U7570 (N_7570,N_7231,N_7202);
and U7571 (N_7571,N_7297,N_7368);
xnor U7572 (N_7572,N_7222,N_7226);
and U7573 (N_7573,N_7209,N_7297);
or U7574 (N_7574,N_7395,N_7363);
nand U7575 (N_7575,N_7206,N_7255);
nor U7576 (N_7576,N_7277,N_7296);
nand U7577 (N_7577,N_7328,N_7263);
nand U7578 (N_7578,N_7375,N_7229);
nor U7579 (N_7579,N_7268,N_7331);
nor U7580 (N_7580,N_7355,N_7250);
or U7581 (N_7581,N_7256,N_7232);
nor U7582 (N_7582,N_7387,N_7293);
xnor U7583 (N_7583,N_7395,N_7233);
or U7584 (N_7584,N_7339,N_7333);
and U7585 (N_7585,N_7231,N_7355);
xor U7586 (N_7586,N_7239,N_7320);
nand U7587 (N_7587,N_7352,N_7234);
nand U7588 (N_7588,N_7236,N_7345);
or U7589 (N_7589,N_7377,N_7273);
xor U7590 (N_7590,N_7302,N_7359);
xnor U7591 (N_7591,N_7345,N_7387);
xor U7592 (N_7592,N_7339,N_7208);
or U7593 (N_7593,N_7214,N_7344);
nand U7594 (N_7594,N_7294,N_7332);
xnor U7595 (N_7595,N_7295,N_7220);
nor U7596 (N_7596,N_7368,N_7375);
and U7597 (N_7597,N_7211,N_7352);
and U7598 (N_7598,N_7216,N_7339);
nand U7599 (N_7599,N_7204,N_7289);
nand U7600 (N_7600,N_7419,N_7477);
nor U7601 (N_7601,N_7566,N_7480);
and U7602 (N_7602,N_7444,N_7511);
or U7603 (N_7603,N_7462,N_7473);
nand U7604 (N_7604,N_7502,N_7548);
and U7605 (N_7605,N_7586,N_7488);
nor U7606 (N_7606,N_7506,N_7534);
nor U7607 (N_7607,N_7490,N_7539);
nor U7608 (N_7608,N_7595,N_7430);
or U7609 (N_7609,N_7496,N_7449);
and U7610 (N_7610,N_7493,N_7457);
nand U7611 (N_7611,N_7581,N_7483);
nand U7612 (N_7612,N_7459,N_7499);
and U7613 (N_7613,N_7479,N_7536);
xnor U7614 (N_7614,N_7554,N_7558);
or U7615 (N_7615,N_7423,N_7471);
and U7616 (N_7616,N_7470,N_7446);
xor U7617 (N_7617,N_7579,N_7561);
and U7618 (N_7618,N_7575,N_7532);
nand U7619 (N_7619,N_7522,N_7552);
and U7620 (N_7620,N_7460,N_7448);
xnor U7621 (N_7621,N_7508,N_7465);
or U7622 (N_7622,N_7414,N_7438);
and U7623 (N_7623,N_7464,N_7463);
and U7624 (N_7624,N_7596,N_7450);
xor U7625 (N_7625,N_7467,N_7518);
or U7626 (N_7626,N_7408,N_7478);
xor U7627 (N_7627,N_7571,N_7469);
and U7628 (N_7628,N_7402,N_7501);
nand U7629 (N_7629,N_7435,N_7409);
xor U7630 (N_7630,N_7598,N_7486);
nand U7631 (N_7631,N_7431,N_7434);
xor U7632 (N_7632,N_7489,N_7422);
nand U7633 (N_7633,N_7497,N_7553);
xnor U7634 (N_7634,N_7527,N_7513);
nand U7635 (N_7635,N_7474,N_7545);
nand U7636 (N_7636,N_7482,N_7599);
xnor U7637 (N_7637,N_7542,N_7447);
or U7638 (N_7638,N_7556,N_7546);
nand U7639 (N_7639,N_7559,N_7578);
and U7640 (N_7640,N_7413,N_7427);
xnor U7641 (N_7641,N_7588,N_7411);
nand U7642 (N_7642,N_7523,N_7436);
xnor U7643 (N_7643,N_7485,N_7439);
or U7644 (N_7644,N_7537,N_7452);
nor U7645 (N_7645,N_7594,N_7541);
xnor U7646 (N_7646,N_7582,N_7416);
nand U7647 (N_7647,N_7455,N_7557);
xor U7648 (N_7648,N_7504,N_7425);
xnor U7649 (N_7649,N_7570,N_7503);
or U7650 (N_7650,N_7475,N_7555);
nor U7651 (N_7651,N_7500,N_7583);
and U7652 (N_7652,N_7535,N_7573);
nand U7653 (N_7653,N_7404,N_7550);
xnor U7654 (N_7654,N_7544,N_7401);
or U7655 (N_7655,N_7529,N_7481);
nand U7656 (N_7656,N_7564,N_7517);
and U7657 (N_7657,N_7453,N_7420);
nor U7658 (N_7658,N_7562,N_7472);
xor U7659 (N_7659,N_7484,N_7424);
xnor U7660 (N_7660,N_7592,N_7567);
nand U7661 (N_7661,N_7412,N_7528);
or U7662 (N_7662,N_7533,N_7428);
nand U7663 (N_7663,N_7445,N_7543);
or U7664 (N_7664,N_7525,N_7591);
nand U7665 (N_7665,N_7405,N_7495);
or U7666 (N_7666,N_7589,N_7429);
nand U7667 (N_7667,N_7510,N_7432);
nor U7668 (N_7668,N_7530,N_7443);
nand U7669 (N_7669,N_7491,N_7584);
nand U7670 (N_7670,N_7512,N_7565);
nor U7671 (N_7671,N_7505,N_7587);
nor U7672 (N_7672,N_7476,N_7406);
nor U7673 (N_7673,N_7577,N_7442);
and U7674 (N_7674,N_7454,N_7593);
nand U7675 (N_7675,N_7520,N_7458);
nand U7676 (N_7676,N_7585,N_7487);
or U7677 (N_7677,N_7492,N_7433);
nand U7678 (N_7678,N_7466,N_7494);
nand U7679 (N_7679,N_7540,N_7597);
xor U7680 (N_7680,N_7572,N_7547);
or U7681 (N_7681,N_7515,N_7417);
xnor U7682 (N_7682,N_7451,N_7516);
or U7683 (N_7683,N_7407,N_7538);
nor U7684 (N_7684,N_7441,N_7569);
nand U7685 (N_7685,N_7551,N_7468);
or U7686 (N_7686,N_7426,N_7524);
xor U7687 (N_7687,N_7568,N_7440);
and U7688 (N_7688,N_7590,N_7519);
or U7689 (N_7689,N_7498,N_7531);
or U7690 (N_7690,N_7421,N_7410);
nand U7691 (N_7691,N_7437,N_7521);
nand U7692 (N_7692,N_7576,N_7507);
nor U7693 (N_7693,N_7456,N_7514);
xnor U7694 (N_7694,N_7418,N_7560);
nand U7695 (N_7695,N_7415,N_7461);
or U7696 (N_7696,N_7574,N_7580);
nand U7697 (N_7697,N_7509,N_7563);
nand U7698 (N_7698,N_7403,N_7526);
and U7699 (N_7699,N_7400,N_7549);
nor U7700 (N_7700,N_7485,N_7496);
xor U7701 (N_7701,N_7494,N_7426);
or U7702 (N_7702,N_7499,N_7535);
xnor U7703 (N_7703,N_7521,N_7493);
xor U7704 (N_7704,N_7427,N_7556);
xnor U7705 (N_7705,N_7483,N_7430);
and U7706 (N_7706,N_7550,N_7505);
nor U7707 (N_7707,N_7494,N_7581);
and U7708 (N_7708,N_7524,N_7481);
and U7709 (N_7709,N_7461,N_7594);
or U7710 (N_7710,N_7410,N_7455);
xnor U7711 (N_7711,N_7550,N_7518);
and U7712 (N_7712,N_7593,N_7435);
nand U7713 (N_7713,N_7421,N_7564);
xor U7714 (N_7714,N_7474,N_7544);
nor U7715 (N_7715,N_7475,N_7595);
nor U7716 (N_7716,N_7532,N_7432);
xnor U7717 (N_7717,N_7526,N_7502);
or U7718 (N_7718,N_7479,N_7481);
or U7719 (N_7719,N_7493,N_7509);
nand U7720 (N_7720,N_7476,N_7447);
xor U7721 (N_7721,N_7570,N_7434);
nand U7722 (N_7722,N_7562,N_7503);
or U7723 (N_7723,N_7524,N_7459);
xnor U7724 (N_7724,N_7514,N_7531);
nor U7725 (N_7725,N_7477,N_7575);
nor U7726 (N_7726,N_7549,N_7517);
or U7727 (N_7727,N_7462,N_7563);
xor U7728 (N_7728,N_7544,N_7596);
nand U7729 (N_7729,N_7568,N_7451);
nor U7730 (N_7730,N_7458,N_7459);
or U7731 (N_7731,N_7414,N_7412);
nor U7732 (N_7732,N_7528,N_7442);
and U7733 (N_7733,N_7400,N_7486);
xnor U7734 (N_7734,N_7555,N_7526);
nor U7735 (N_7735,N_7530,N_7570);
xnor U7736 (N_7736,N_7440,N_7426);
or U7737 (N_7737,N_7462,N_7429);
nand U7738 (N_7738,N_7505,N_7525);
nand U7739 (N_7739,N_7522,N_7455);
or U7740 (N_7740,N_7464,N_7466);
and U7741 (N_7741,N_7402,N_7586);
xnor U7742 (N_7742,N_7401,N_7525);
nor U7743 (N_7743,N_7475,N_7419);
nand U7744 (N_7744,N_7471,N_7520);
or U7745 (N_7745,N_7571,N_7552);
xnor U7746 (N_7746,N_7551,N_7548);
nand U7747 (N_7747,N_7469,N_7558);
and U7748 (N_7748,N_7432,N_7576);
and U7749 (N_7749,N_7483,N_7418);
xnor U7750 (N_7750,N_7456,N_7450);
xnor U7751 (N_7751,N_7521,N_7571);
nor U7752 (N_7752,N_7464,N_7435);
nor U7753 (N_7753,N_7463,N_7538);
nand U7754 (N_7754,N_7408,N_7549);
nand U7755 (N_7755,N_7474,N_7423);
nor U7756 (N_7756,N_7506,N_7554);
nor U7757 (N_7757,N_7484,N_7411);
nor U7758 (N_7758,N_7490,N_7415);
nor U7759 (N_7759,N_7432,N_7500);
or U7760 (N_7760,N_7575,N_7466);
xor U7761 (N_7761,N_7471,N_7432);
or U7762 (N_7762,N_7595,N_7575);
nor U7763 (N_7763,N_7573,N_7413);
or U7764 (N_7764,N_7568,N_7416);
or U7765 (N_7765,N_7598,N_7514);
and U7766 (N_7766,N_7496,N_7526);
and U7767 (N_7767,N_7513,N_7575);
xor U7768 (N_7768,N_7599,N_7540);
and U7769 (N_7769,N_7490,N_7420);
or U7770 (N_7770,N_7521,N_7464);
xor U7771 (N_7771,N_7427,N_7433);
or U7772 (N_7772,N_7547,N_7561);
and U7773 (N_7773,N_7429,N_7456);
or U7774 (N_7774,N_7484,N_7482);
nor U7775 (N_7775,N_7506,N_7599);
xor U7776 (N_7776,N_7417,N_7516);
and U7777 (N_7777,N_7452,N_7460);
xnor U7778 (N_7778,N_7589,N_7401);
nor U7779 (N_7779,N_7520,N_7518);
xor U7780 (N_7780,N_7431,N_7593);
nor U7781 (N_7781,N_7427,N_7431);
or U7782 (N_7782,N_7495,N_7490);
xor U7783 (N_7783,N_7407,N_7475);
and U7784 (N_7784,N_7563,N_7569);
nand U7785 (N_7785,N_7425,N_7406);
nand U7786 (N_7786,N_7407,N_7557);
and U7787 (N_7787,N_7438,N_7455);
xnor U7788 (N_7788,N_7452,N_7455);
and U7789 (N_7789,N_7536,N_7594);
xor U7790 (N_7790,N_7445,N_7458);
xor U7791 (N_7791,N_7542,N_7454);
or U7792 (N_7792,N_7592,N_7596);
nand U7793 (N_7793,N_7447,N_7483);
or U7794 (N_7794,N_7449,N_7417);
nor U7795 (N_7795,N_7451,N_7533);
xor U7796 (N_7796,N_7520,N_7473);
or U7797 (N_7797,N_7532,N_7475);
or U7798 (N_7798,N_7491,N_7464);
nor U7799 (N_7799,N_7435,N_7584);
xnor U7800 (N_7800,N_7793,N_7730);
and U7801 (N_7801,N_7675,N_7651);
nor U7802 (N_7802,N_7613,N_7690);
or U7803 (N_7803,N_7628,N_7668);
or U7804 (N_7804,N_7605,N_7641);
and U7805 (N_7805,N_7778,N_7799);
nand U7806 (N_7806,N_7643,N_7636);
or U7807 (N_7807,N_7685,N_7714);
or U7808 (N_7808,N_7633,N_7781);
nor U7809 (N_7809,N_7733,N_7602);
xnor U7810 (N_7810,N_7672,N_7657);
nor U7811 (N_7811,N_7742,N_7718);
nand U7812 (N_7812,N_7688,N_7782);
or U7813 (N_7813,N_7784,N_7796);
xor U7814 (N_7814,N_7728,N_7607);
nor U7815 (N_7815,N_7795,N_7755);
or U7816 (N_7816,N_7615,N_7756);
and U7817 (N_7817,N_7658,N_7706);
and U7818 (N_7818,N_7671,N_7725);
nand U7819 (N_7819,N_7779,N_7780);
or U7820 (N_7820,N_7773,N_7732);
xnor U7821 (N_7821,N_7749,N_7746);
nor U7822 (N_7822,N_7634,N_7786);
nor U7823 (N_7823,N_7741,N_7701);
or U7824 (N_7824,N_7712,N_7740);
and U7825 (N_7825,N_7702,N_7758);
nor U7826 (N_7826,N_7770,N_7600);
nor U7827 (N_7827,N_7709,N_7686);
nor U7828 (N_7828,N_7679,N_7654);
and U7829 (N_7829,N_7640,N_7724);
or U7830 (N_7830,N_7642,N_7644);
xor U7831 (N_7831,N_7700,N_7776);
xnor U7832 (N_7832,N_7699,N_7669);
nand U7833 (N_7833,N_7705,N_7797);
nand U7834 (N_7834,N_7715,N_7630);
or U7835 (N_7835,N_7761,N_7736);
nor U7836 (N_7836,N_7774,N_7622);
and U7837 (N_7837,N_7631,N_7635);
and U7838 (N_7838,N_7763,N_7610);
nand U7839 (N_7839,N_7771,N_7684);
and U7840 (N_7840,N_7754,N_7619);
or U7841 (N_7841,N_7789,N_7787);
nand U7842 (N_7842,N_7720,N_7738);
nor U7843 (N_7843,N_7665,N_7762);
and U7844 (N_7844,N_7767,N_7659);
or U7845 (N_7845,N_7663,N_7650);
and U7846 (N_7846,N_7670,N_7677);
nand U7847 (N_7847,N_7772,N_7608);
nand U7848 (N_7848,N_7783,N_7612);
or U7849 (N_7849,N_7618,N_7711);
or U7850 (N_7850,N_7614,N_7703);
nand U7851 (N_7851,N_7661,N_7707);
or U7852 (N_7852,N_7674,N_7710);
nor U7853 (N_7853,N_7791,N_7737);
and U7854 (N_7854,N_7768,N_7645);
xnor U7855 (N_7855,N_7673,N_7750);
and U7856 (N_7856,N_7683,N_7611);
or U7857 (N_7857,N_7693,N_7723);
and U7858 (N_7858,N_7639,N_7751);
xor U7859 (N_7859,N_7624,N_7626);
nand U7860 (N_7860,N_7759,N_7694);
nand U7861 (N_7861,N_7698,N_7721);
or U7862 (N_7862,N_7652,N_7726);
or U7863 (N_7863,N_7729,N_7760);
or U7864 (N_7864,N_7691,N_7646);
xor U7865 (N_7865,N_7716,N_7696);
nand U7866 (N_7866,N_7648,N_7743);
xor U7867 (N_7867,N_7689,N_7692);
or U7868 (N_7868,N_7617,N_7798);
or U7869 (N_7869,N_7719,N_7695);
nand U7870 (N_7870,N_7623,N_7734);
nand U7871 (N_7871,N_7731,N_7788);
and U7872 (N_7872,N_7747,N_7660);
nor U7873 (N_7873,N_7792,N_7704);
xor U7874 (N_7874,N_7748,N_7625);
nand U7875 (N_7875,N_7621,N_7777);
xor U7876 (N_7876,N_7653,N_7627);
or U7877 (N_7877,N_7735,N_7616);
xor U7878 (N_7878,N_7629,N_7676);
xnor U7879 (N_7879,N_7722,N_7757);
and U7880 (N_7880,N_7662,N_7766);
nor U7881 (N_7881,N_7794,N_7649);
nor U7882 (N_7882,N_7632,N_7667);
nor U7883 (N_7883,N_7769,N_7713);
and U7884 (N_7884,N_7764,N_7682);
and U7885 (N_7885,N_7601,N_7603);
nand U7886 (N_7886,N_7697,N_7620);
nor U7887 (N_7887,N_7664,N_7647);
or U7888 (N_7888,N_7609,N_7785);
nand U7889 (N_7889,N_7687,N_7727);
or U7890 (N_7890,N_7681,N_7604);
nor U7891 (N_7891,N_7637,N_7717);
nand U7892 (N_7892,N_7680,N_7744);
or U7893 (N_7893,N_7745,N_7739);
and U7894 (N_7894,N_7656,N_7666);
nand U7895 (N_7895,N_7765,N_7752);
xor U7896 (N_7896,N_7638,N_7655);
xor U7897 (N_7897,N_7775,N_7678);
or U7898 (N_7898,N_7790,N_7753);
xor U7899 (N_7899,N_7708,N_7606);
and U7900 (N_7900,N_7744,N_7675);
nor U7901 (N_7901,N_7762,N_7697);
and U7902 (N_7902,N_7747,N_7757);
nand U7903 (N_7903,N_7628,N_7624);
nand U7904 (N_7904,N_7675,N_7688);
or U7905 (N_7905,N_7765,N_7718);
or U7906 (N_7906,N_7738,N_7670);
nor U7907 (N_7907,N_7687,N_7602);
nand U7908 (N_7908,N_7661,N_7710);
nor U7909 (N_7909,N_7618,N_7678);
or U7910 (N_7910,N_7756,N_7701);
nor U7911 (N_7911,N_7775,N_7622);
nand U7912 (N_7912,N_7687,N_7722);
nand U7913 (N_7913,N_7761,N_7608);
and U7914 (N_7914,N_7753,N_7648);
nand U7915 (N_7915,N_7708,N_7699);
and U7916 (N_7916,N_7642,N_7703);
xor U7917 (N_7917,N_7778,N_7787);
xor U7918 (N_7918,N_7734,N_7774);
and U7919 (N_7919,N_7771,N_7784);
or U7920 (N_7920,N_7705,N_7626);
or U7921 (N_7921,N_7798,N_7687);
xor U7922 (N_7922,N_7656,N_7648);
nor U7923 (N_7923,N_7635,N_7607);
xnor U7924 (N_7924,N_7767,N_7742);
nand U7925 (N_7925,N_7634,N_7657);
and U7926 (N_7926,N_7615,N_7773);
or U7927 (N_7927,N_7623,N_7603);
nor U7928 (N_7928,N_7605,N_7679);
or U7929 (N_7929,N_7749,N_7775);
xnor U7930 (N_7930,N_7608,N_7660);
nand U7931 (N_7931,N_7741,N_7769);
or U7932 (N_7932,N_7709,N_7616);
and U7933 (N_7933,N_7788,N_7769);
xnor U7934 (N_7934,N_7773,N_7695);
nor U7935 (N_7935,N_7611,N_7676);
and U7936 (N_7936,N_7777,N_7678);
or U7937 (N_7937,N_7771,N_7776);
nor U7938 (N_7938,N_7655,N_7623);
nand U7939 (N_7939,N_7631,N_7739);
nand U7940 (N_7940,N_7617,N_7682);
or U7941 (N_7941,N_7697,N_7690);
xnor U7942 (N_7942,N_7703,N_7666);
and U7943 (N_7943,N_7715,N_7665);
or U7944 (N_7944,N_7621,N_7657);
nand U7945 (N_7945,N_7786,N_7658);
xor U7946 (N_7946,N_7731,N_7644);
nand U7947 (N_7947,N_7720,N_7632);
nor U7948 (N_7948,N_7601,N_7619);
or U7949 (N_7949,N_7613,N_7709);
nand U7950 (N_7950,N_7652,N_7793);
nand U7951 (N_7951,N_7781,N_7732);
nor U7952 (N_7952,N_7746,N_7600);
nand U7953 (N_7953,N_7768,N_7788);
nand U7954 (N_7954,N_7769,N_7717);
xor U7955 (N_7955,N_7684,N_7746);
or U7956 (N_7956,N_7642,N_7672);
nand U7957 (N_7957,N_7661,N_7605);
xor U7958 (N_7958,N_7749,N_7737);
and U7959 (N_7959,N_7689,N_7671);
nand U7960 (N_7960,N_7791,N_7670);
nor U7961 (N_7961,N_7682,N_7660);
nand U7962 (N_7962,N_7765,N_7660);
and U7963 (N_7963,N_7781,N_7753);
nor U7964 (N_7964,N_7671,N_7677);
or U7965 (N_7965,N_7642,N_7686);
and U7966 (N_7966,N_7775,N_7777);
or U7967 (N_7967,N_7650,N_7771);
nand U7968 (N_7968,N_7695,N_7711);
and U7969 (N_7969,N_7759,N_7776);
xnor U7970 (N_7970,N_7626,N_7795);
xor U7971 (N_7971,N_7787,N_7667);
or U7972 (N_7972,N_7738,N_7724);
xnor U7973 (N_7973,N_7742,N_7684);
and U7974 (N_7974,N_7701,N_7720);
nand U7975 (N_7975,N_7688,N_7696);
nor U7976 (N_7976,N_7737,N_7675);
xor U7977 (N_7977,N_7749,N_7638);
nand U7978 (N_7978,N_7773,N_7753);
and U7979 (N_7979,N_7790,N_7712);
xnor U7980 (N_7980,N_7741,N_7702);
nand U7981 (N_7981,N_7697,N_7615);
xor U7982 (N_7982,N_7730,N_7721);
and U7983 (N_7983,N_7719,N_7744);
xnor U7984 (N_7984,N_7728,N_7736);
nor U7985 (N_7985,N_7783,N_7792);
and U7986 (N_7986,N_7653,N_7771);
xnor U7987 (N_7987,N_7748,N_7603);
and U7988 (N_7988,N_7755,N_7716);
nor U7989 (N_7989,N_7728,N_7763);
nor U7990 (N_7990,N_7682,N_7700);
nand U7991 (N_7991,N_7725,N_7771);
or U7992 (N_7992,N_7712,N_7626);
nor U7993 (N_7993,N_7714,N_7759);
nand U7994 (N_7994,N_7765,N_7701);
or U7995 (N_7995,N_7655,N_7751);
and U7996 (N_7996,N_7745,N_7639);
xnor U7997 (N_7997,N_7620,N_7601);
nor U7998 (N_7998,N_7700,N_7723);
and U7999 (N_7999,N_7759,N_7754);
and U8000 (N_8000,N_7885,N_7819);
xor U8001 (N_8001,N_7945,N_7961);
or U8002 (N_8002,N_7997,N_7804);
nand U8003 (N_8003,N_7873,N_7979);
nor U8004 (N_8004,N_7848,N_7907);
nand U8005 (N_8005,N_7850,N_7881);
or U8006 (N_8006,N_7957,N_7944);
and U8007 (N_8007,N_7942,N_7946);
and U8008 (N_8008,N_7947,N_7840);
and U8009 (N_8009,N_7887,N_7967);
and U8010 (N_8010,N_7954,N_7878);
xnor U8011 (N_8011,N_7855,N_7884);
nand U8012 (N_8012,N_7914,N_7926);
or U8013 (N_8013,N_7801,N_7815);
xnor U8014 (N_8014,N_7920,N_7831);
or U8015 (N_8015,N_7998,N_7906);
nand U8016 (N_8016,N_7864,N_7928);
or U8017 (N_8017,N_7817,N_7976);
or U8018 (N_8018,N_7823,N_7843);
nand U8019 (N_8019,N_7988,N_7839);
and U8020 (N_8020,N_7844,N_7834);
or U8021 (N_8021,N_7821,N_7968);
or U8022 (N_8022,N_7975,N_7913);
nor U8023 (N_8023,N_7965,N_7858);
nor U8024 (N_8024,N_7836,N_7852);
or U8025 (N_8025,N_7974,N_7809);
and U8026 (N_8026,N_7985,N_7922);
xnor U8027 (N_8027,N_7832,N_7959);
nand U8028 (N_8028,N_7837,N_7802);
and U8029 (N_8029,N_7863,N_7956);
nor U8030 (N_8030,N_7896,N_7966);
and U8031 (N_8031,N_7842,N_7986);
nand U8032 (N_8032,N_7862,N_7962);
nor U8033 (N_8033,N_7814,N_7828);
and U8034 (N_8034,N_7847,N_7854);
or U8035 (N_8035,N_7857,N_7875);
nand U8036 (N_8036,N_7841,N_7808);
nor U8037 (N_8037,N_7827,N_7853);
nand U8038 (N_8038,N_7800,N_7856);
nor U8039 (N_8039,N_7903,N_7900);
nand U8040 (N_8040,N_7893,N_7989);
or U8041 (N_8041,N_7894,N_7937);
xor U8042 (N_8042,N_7803,N_7970);
xnor U8043 (N_8043,N_7950,N_7929);
and U8044 (N_8044,N_7870,N_7918);
nand U8045 (N_8045,N_7899,N_7867);
xor U8046 (N_8046,N_7934,N_7888);
or U8047 (N_8047,N_7830,N_7822);
nor U8048 (N_8048,N_7910,N_7943);
and U8049 (N_8049,N_7811,N_7851);
nor U8050 (N_8050,N_7995,N_7911);
xnor U8051 (N_8051,N_7935,N_7940);
nand U8052 (N_8052,N_7973,N_7820);
nand U8053 (N_8053,N_7931,N_7936);
nor U8054 (N_8054,N_7883,N_7845);
or U8055 (N_8055,N_7955,N_7859);
or U8056 (N_8056,N_7824,N_7912);
or U8057 (N_8057,N_7890,N_7939);
and U8058 (N_8058,N_7825,N_7813);
nor U8059 (N_8059,N_7952,N_7905);
nand U8060 (N_8060,N_7941,N_7807);
and U8061 (N_8061,N_7898,N_7932);
nand U8062 (N_8062,N_7958,N_7990);
or U8063 (N_8063,N_7818,N_7953);
or U8064 (N_8064,N_7964,N_7999);
nand U8065 (N_8065,N_7978,N_7904);
or U8066 (N_8066,N_7849,N_7917);
xor U8067 (N_8067,N_7933,N_7816);
xor U8068 (N_8068,N_7806,N_7984);
or U8069 (N_8069,N_7895,N_7861);
xor U8070 (N_8070,N_7951,N_7902);
nand U8071 (N_8071,N_7835,N_7865);
nor U8072 (N_8072,N_7860,N_7938);
xor U8073 (N_8073,N_7872,N_7919);
or U8074 (N_8074,N_7915,N_7874);
and U8075 (N_8075,N_7880,N_7996);
nand U8076 (N_8076,N_7921,N_7991);
xor U8077 (N_8077,N_7829,N_7924);
xnor U8078 (N_8078,N_7866,N_7908);
and U8079 (N_8079,N_7977,N_7876);
nand U8080 (N_8080,N_7960,N_7993);
and U8081 (N_8081,N_7869,N_7882);
nor U8082 (N_8082,N_7871,N_7805);
nand U8083 (N_8083,N_7886,N_7868);
nor U8084 (N_8084,N_7838,N_7901);
nand U8085 (N_8085,N_7897,N_7889);
xor U8086 (N_8086,N_7879,N_7909);
and U8087 (N_8087,N_7892,N_7812);
nor U8088 (N_8088,N_7987,N_7930);
nand U8089 (N_8089,N_7981,N_7826);
and U8090 (N_8090,N_7925,N_7983);
nor U8091 (N_8091,N_7992,N_7972);
and U8092 (N_8092,N_7948,N_7982);
nand U8093 (N_8093,N_7963,N_7969);
nor U8094 (N_8094,N_7927,N_7833);
nor U8095 (N_8095,N_7923,N_7891);
xnor U8096 (N_8096,N_7971,N_7846);
or U8097 (N_8097,N_7980,N_7877);
nand U8098 (N_8098,N_7994,N_7949);
or U8099 (N_8099,N_7916,N_7810);
nand U8100 (N_8100,N_7953,N_7963);
nor U8101 (N_8101,N_7988,N_7975);
nor U8102 (N_8102,N_7968,N_7879);
and U8103 (N_8103,N_7991,N_7846);
or U8104 (N_8104,N_7825,N_7902);
nor U8105 (N_8105,N_7861,N_7979);
xor U8106 (N_8106,N_7924,N_7910);
xor U8107 (N_8107,N_7815,N_7865);
nand U8108 (N_8108,N_7902,N_7987);
xor U8109 (N_8109,N_7951,N_7889);
xor U8110 (N_8110,N_7973,N_7929);
or U8111 (N_8111,N_7804,N_7879);
or U8112 (N_8112,N_7815,N_7854);
nor U8113 (N_8113,N_7849,N_7948);
or U8114 (N_8114,N_7818,N_7890);
nand U8115 (N_8115,N_7888,N_7968);
xor U8116 (N_8116,N_7806,N_7934);
nand U8117 (N_8117,N_7907,N_7802);
xnor U8118 (N_8118,N_7834,N_7827);
nor U8119 (N_8119,N_7863,N_7835);
nor U8120 (N_8120,N_7901,N_7979);
and U8121 (N_8121,N_7931,N_7935);
nand U8122 (N_8122,N_7982,N_7829);
or U8123 (N_8123,N_7851,N_7869);
nand U8124 (N_8124,N_7971,N_7874);
and U8125 (N_8125,N_7883,N_7891);
nor U8126 (N_8126,N_7977,N_7874);
or U8127 (N_8127,N_7958,N_7924);
nor U8128 (N_8128,N_7978,N_7997);
nor U8129 (N_8129,N_7816,N_7833);
and U8130 (N_8130,N_7948,N_7934);
or U8131 (N_8131,N_7973,N_7861);
nand U8132 (N_8132,N_7854,N_7919);
nor U8133 (N_8133,N_7882,N_7898);
and U8134 (N_8134,N_7923,N_7876);
nand U8135 (N_8135,N_7962,N_7945);
xnor U8136 (N_8136,N_7983,N_7839);
and U8137 (N_8137,N_7818,N_7896);
and U8138 (N_8138,N_7946,N_7913);
xnor U8139 (N_8139,N_7929,N_7990);
nand U8140 (N_8140,N_7935,N_7832);
nand U8141 (N_8141,N_7882,N_7814);
or U8142 (N_8142,N_7848,N_7804);
and U8143 (N_8143,N_7990,N_7994);
nand U8144 (N_8144,N_7969,N_7964);
nand U8145 (N_8145,N_7903,N_7892);
nand U8146 (N_8146,N_7976,N_7939);
xor U8147 (N_8147,N_7887,N_7923);
or U8148 (N_8148,N_7946,N_7841);
or U8149 (N_8149,N_7983,N_7815);
xnor U8150 (N_8150,N_7863,N_7836);
nand U8151 (N_8151,N_7832,N_7954);
nor U8152 (N_8152,N_7805,N_7862);
xnor U8153 (N_8153,N_7884,N_7815);
nor U8154 (N_8154,N_7966,N_7980);
xor U8155 (N_8155,N_7896,N_7949);
nor U8156 (N_8156,N_7977,N_7864);
nor U8157 (N_8157,N_7965,N_7952);
nand U8158 (N_8158,N_7934,N_7861);
or U8159 (N_8159,N_7943,N_7960);
nor U8160 (N_8160,N_7980,N_7999);
nor U8161 (N_8161,N_7924,N_7993);
nand U8162 (N_8162,N_7869,N_7840);
xor U8163 (N_8163,N_7890,N_7832);
nand U8164 (N_8164,N_7998,N_7888);
nor U8165 (N_8165,N_7807,N_7884);
nand U8166 (N_8166,N_7998,N_7870);
or U8167 (N_8167,N_7835,N_7997);
and U8168 (N_8168,N_7876,N_7886);
nand U8169 (N_8169,N_7824,N_7822);
xor U8170 (N_8170,N_7930,N_7808);
and U8171 (N_8171,N_7857,N_7945);
xnor U8172 (N_8172,N_7917,N_7858);
nor U8173 (N_8173,N_7899,N_7869);
nor U8174 (N_8174,N_7950,N_7908);
xnor U8175 (N_8175,N_7943,N_7818);
and U8176 (N_8176,N_7818,N_7927);
or U8177 (N_8177,N_7958,N_7839);
or U8178 (N_8178,N_7855,N_7893);
nand U8179 (N_8179,N_7839,N_7929);
nor U8180 (N_8180,N_7964,N_7898);
and U8181 (N_8181,N_7875,N_7861);
nor U8182 (N_8182,N_7812,N_7876);
or U8183 (N_8183,N_7833,N_7890);
and U8184 (N_8184,N_7833,N_7972);
or U8185 (N_8185,N_7985,N_7857);
nand U8186 (N_8186,N_7868,N_7961);
nand U8187 (N_8187,N_7984,N_7861);
or U8188 (N_8188,N_7872,N_7810);
and U8189 (N_8189,N_7855,N_7844);
xor U8190 (N_8190,N_7900,N_7808);
nand U8191 (N_8191,N_7855,N_7995);
or U8192 (N_8192,N_7875,N_7932);
and U8193 (N_8193,N_7836,N_7951);
nand U8194 (N_8194,N_7997,N_7954);
nor U8195 (N_8195,N_7941,N_7928);
or U8196 (N_8196,N_7898,N_7935);
and U8197 (N_8197,N_7885,N_7913);
nor U8198 (N_8198,N_7865,N_7838);
or U8199 (N_8199,N_7914,N_7932);
and U8200 (N_8200,N_8178,N_8185);
nor U8201 (N_8201,N_8054,N_8064);
and U8202 (N_8202,N_8000,N_8188);
and U8203 (N_8203,N_8171,N_8189);
nor U8204 (N_8204,N_8034,N_8088);
nand U8205 (N_8205,N_8150,N_8126);
nor U8206 (N_8206,N_8026,N_8163);
xor U8207 (N_8207,N_8193,N_8136);
and U8208 (N_8208,N_8035,N_8024);
and U8209 (N_8209,N_8104,N_8131);
nand U8210 (N_8210,N_8099,N_8084);
xor U8211 (N_8211,N_8111,N_8108);
and U8212 (N_8212,N_8128,N_8098);
nand U8213 (N_8213,N_8162,N_8165);
nand U8214 (N_8214,N_8044,N_8120);
xnor U8215 (N_8215,N_8109,N_8007);
or U8216 (N_8216,N_8018,N_8168);
and U8217 (N_8217,N_8187,N_8052);
and U8218 (N_8218,N_8135,N_8183);
nor U8219 (N_8219,N_8090,N_8115);
or U8220 (N_8220,N_8102,N_8137);
and U8221 (N_8221,N_8025,N_8086);
xor U8222 (N_8222,N_8033,N_8020);
nor U8223 (N_8223,N_8196,N_8145);
xor U8224 (N_8224,N_8029,N_8056);
nor U8225 (N_8225,N_8154,N_8057);
nand U8226 (N_8226,N_8142,N_8010);
nand U8227 (N_8227,N_8119,N_8148);
or U8228 (N_8228,N_8197,N_8139);
nor U8229 (N_8229,N_8008,N_8133);
nand U8230 (N_8230,N_8078,N_8093);
nor U8231 (N_8231,N_8181,N_8155);
and U8232 (N_8232,N_8005,N_8022);
and U8233 (N_8233,N_8070,N_8199);
nor U8234 (N_8234,N_8124,N_8149);
or U8235 (N_8235,N_8166,N_8031);
and U8236 (N_8236,N_8101,N_8058);
and U8237 (N_8237,N_8037,N_8112);
nor U8238 (N_8238,N_8055,N_8097);
nor U8239 (N_8239,N_8177,N_8184);
or U8240 (N_8240,N_8161,N_8114);
nand U8241 (N_8241,N_8105,N_8174);
xor U8242 (N_8242,N_8083,N_8127);
xnor U8243 (N_8243,N_8152,N_8074);
nor U8244 (N_8244,N_8110,N_8143);
nor U8245 (N_8245,N_8016,N_8063);
or U8246 (N_8246,N_8009,N_8125);
nand U8247 (N_8247,N_8118,N_8141);
and U8248 (N_8248,N_8198,N_8049);
or U8249 (N_8249,N_8032,N_8048);
nand U8250 (N_8250,N_8069,N_8076);
or U8251 (N_8251,N_8028,N_8151);
nor U8252 (N_8252,N_8147,N_8087);
or U8253 (N_8253,N_8053,N_8027);
xor U8254 (N_8254,N_8011,N_8144);
nor U8255 (N_8255,N_8030,N_8179);
and U8256 (N_8256,N_8158,N_8103);
nor U8257 (N_8257,N_8004,N_8160);
nand U8258 (N_8258,N_8012,N_8050);
and U8259 (N_8259,N_8191,N_8041);
nor U8260 (N_8260,N_8001,N_8067);
nand U8261 (N_8261,N_8023,N_8036);
nor U8262 (N_8262,N_8085,N_8095);
nor U8263 (N_8263,N_8073,N_8146);
nand U8264 (N_8264,N_8122,N_8182);
or U8265 (N_8265,N_8077,N_8042);
or U8266 (N_8266,N_8047,N_8106);
nor U8267 (N_8267,N_8172,N_8176);
nand U8268 (N_8268,N_8038,N_8003);
or U8269 (N_8269,N_8062,N_8089);
xnor U8270 (N_8270,N_8186,N_8117);
nand U8271 (N_8271,N_8173,N_8157);
xor U8272 (N_8272,N_8080,N_8092);
and U8273 (N_8273,N_8129,N_8094);
and U8274 (N_8274,N_8091,N_8071);
nand U8275 (N_8275,N_8153,N_8081);
or U8276 (N_8276,N_8045,N_8082);
nor U8277 (N_8277,N_8164,N_8194);
or U8278 (N_8278,N_8043,N_8156);
or U8279 (N_8279,N_8140,N_8061);
and U8280 (N_8280,N_8116,N_8017);
nand U8281 (N_8281,N_8014,N_8013);
xor U8282 (N_8282,N_8019,N_8134);
xor U8283 (N_8283,N_8046,N_8051);
nor U8284 (N_8284,N_8159,N_8167);
and U8285 (N_8285,N_8079,N_8123);
xor U8286 (N_8286,N_8175,N_8059);
xor U8287 (N_8287,N_8113,N_8075);
nor U8288 (N_8288,N_8100,N_8107);
xor U8289 (N_8289,N_8130,N_8066);
nor U8290 (N_8290,N_8132,N_8192);
nand U8291 (N_8291,N_8170,N_8040);
nor U8292 (N_8292,N_8096,N_8169);
nand U8293 (N_8293,N_8195,N_8006);
nor U8294 (N_8294,N_8002,N_8065);
nor U8295 (N_8295,N_8180,N_8060);
or U8296 (N_8296,N_8138,N_8015);
xor U8297 (N_8297,N_8068,N_8072);
and U8298 (N_8298,N_8190,N_8039);
xnor U8299 (N_8299,N_8121,N_8021);
and U8300 (N_8300,N_8011,N_8132);
xnor U8301 (N_8301,N_8198,N_8164);
nor U8302 (N_8302,N_8189,N_8178);
or U8303 (N_8303,N_8157,N_8092);
nor U8304 (N_8304,N_8096,N_8186);
nand U8305 (N_8305,N_8011,N_8101);
xnor U8306 (N_8306,N_8163,N_8161);
or U8307 (N_8307,N_8112,N_8180);
nor U8308 (N_8308,N_8014,N_8049);
and U8309 (N_8309,N_8058,N_8190);
xnor U8310 (N_8310,N_8043,N_8079);
nor U8311 (N_8311,N_8153,N_8143);
xor U8312 (N_8312,N_8040,N_8137);
nand U8313 (N_8313,N_8109,N_8132);
and U8314 (N_8314,N_8185,N_8033);
nand U8315 (N_8315,N_8022,N_8098);
or U8316 (N_8316,N_8029,N_8124);
xor U8317 (N_8317,N_8167,N_8137);
nor U8318 (N_8318,N_8124,N_8148);
or U8319 (N_8319,N_8139,N_8029);
xor U8320 (N_8320,N_8194,N_8156);
xor U8321 (N_8321,N_8016,N_8140);
or U8322 (N_8322,N_8062,N_8035);
nand U8323 (N_8323,N_8171,N_8133);
and U8324 (N_8324,N_8087,N_8113);
xor U8325 (N_8325,N_8003,N_8116);
nor U8326 (N_8326,N_8062,N_8178);
and U8327 (N_8327,N_8032,N_8118);
or U8328 (N_8328,N_8026,N_8142);
nor U8329 (N_8329,N_8129,N_8174);
nand U8330 (N_8330,N_8190,N_8107);
nand U8331 (N_8331,N_8073,N_8149);
nor U8332 (N_8332,N_8170,N_8045);
xnor U8333 (N_8333,N_8191,N_8084);
xnor U8334 (N_8334,N_8188,N_8058);
nor U8335 (N_8335,N_8193,N_8022);
and U8336 (N_8336,N_8145,N_8088);
nor U8337 (N_8337,N_8038,N_8013);
nor U8338 (N_8338,N_8001,N_8138);
xnor U8339 (N_8339,N_8112,N_8139);
nand U8340 (N_8340,N_8004,N_8102);
xnor U8341 (N_8341,N_8148,N_8070);
nand U8342 (N_8342,N_8077,N_8096);
nor U8343 (N_8343,N_8084,N_8133);
and U8344 (N_8344,N_8157,N_8052);
and U8345 (N_8345,N_8149,N_8074);
and U8346 (N_8346,N_8062,N_8015);
nand U8347 (N_8347,N_8170,N_8191);
or U8348 (N_8348,N_8184,N_8153);
nor U8349 (N_8349,N_8155,N_8141);
nor U8350 (N_8350,N_8045,N_8055);
nor U8351 (N_8351,N_8051,N_8087);
nor U8352 (N_8352,N_8069,N_8174);
xnor U8353 (N_8353,N_8022,N_8130);
nor U8354 (N_8354,N_8064,N_8193);
nand U8355 (N_8355,N_8132,N_8197);
or U8356 (N_8356,N_8122,N_8163);
nand U8357 (N_8357,N_8047,N_8121);
nand U8358 (N_8358,N_8092,N_8011);
xor U8359 (N_8359,N_8041,N_8110);
xor U8360 (N_8360,N_8004,N_8182);
xnor U8361 (N_8361,N_8038,N_8079);
or U8362 (N_8362,N_8028,N_8185);
nor U8363 (N_8363,N_8154,N_8176);
xor U8364 (N_8364,N_8049,N_8197);
nor U8365 (N_8365,N_8129,N_8025);
or U8366 (N_8366,N_8091,N_8015);
xor U8367 (N_8367,N_8157,N_8194);
nand U8368 (N_8368,N_8017,N_8016);
or U8369 (N_8369,N_8096,N_8177);
nand U8370 (N_8370,N_8007,N_8041);
nor U8371 (N_8371,N_8131,N_8129);
nand U8372 (N_8372,N_8126,N_8092);
or U8373 (N_8373,N_8029,N_8022);
nand U8374 (N_8374,N_8056,N_8128);
nor U8375 (N_8375,N_8108,N_8037);
nand U8376 (N_8376,N_8106,N_8128);
xor U8377 (N_8377,N_8046,N_8145);
and U8378 (N_8378,N_8026,N_8019);
or U8379 (N_8379,N_8090,N_8006);
and U8380 (N_8380,N_8116,N_8112);
xor U8381 (N_8381,N_8080,N_8165);
or U8382 (N_8382,N_8058,N_8129);
nor U8383 (N_8383,N_8045,N_8068);
nand U8384 (N_8384,N_8117,N_8014);
and U8385 (N_8385,N_8090,N_8058);
or U8386 (N_8386,N_8103,N_8005);
xor U8387 (N_8387,N_8166,N_8064);
xnor U8388 (N_8388,N_8001,N_8103);
xnor U8389 (N_8389,N_8146,N_8168);
or U8390 (N_8390,N_8193,N_8034);
or U8391 (N_8391,N_8001,N_8080);
nand U8392 (N_8392,N_8191,N_8093);
and U8393 (N_8393,N_8079,N_8019);
or U8394 (N_8394,N_8141,N_8058);
xnor U8395 (N_8395,N_8080,N_8121);
nand U8396 (N_8396,N_8065,N_8006);
nor U8397 (N_8397,N_8009,N_8088);
or U8398 (N_8398,N_8168,N_8006);
xor U8399 (N_8399,N_8130,N_8143);
and U8400 (N_8400,N_8280,N_8393);
nor U8401 (N_8401,N_8335,N_8321);
nor U8402 (N_8402,N_8270,N_8314);
nand U8403 (N_8403,N_8399,N_8392);
xnor U8404 (N_8404,N_8318,N_8397);
xnor U8405 (N_8405,N_8359,N_8217);
nand U8406 (N_8406,N_8291,N_8306);
or U8407 (N_8407,N_8281,N_8348);
nand U8408 (N_8408,N_8350,N_8374);
xnor U8409 (N_8409,N_8239,N_8279);
and U8410 (N_8410,N_8372,N_8282);
or U8411 (N_8411,N_8386,N_8349);
nand U8412 (N_8412,N_8228,N_8337);
nand U8413 (N_8413,N_8237,N_8304);
nand U8414 (N_8414,N_8285,N_8352);
and U8415 (N_8415,N_8251,N_8357);
xor U8416 (N_8416,N_8387,N_8278);
xnor U8417 (N_8417,N_8346,N_8389);
nor U8418 (N_8418,N_8264,N_8286);
or U8419 (N_8419,N_8311,N_8275);
or U8420 (N_8420,N_8269,N_8261);
xnor U8421 (N_8421,N_8378,N_8223);
and U8422 (N_8422,N_8302,N_8300);
xnor U8423 (N_8423,N_8292,N_8299);
nand U8424 (N_8424,N_8356,N_8385);
nor U8425 (N_8425,N_8289,N_8222);
xnor U8426 (N_8426,N_8255,N_8267);
nand U8427 (N_8427,N_8229,N_8277);
nand U8428 (N_8428,N_8268,N_8273);
nand U8429 (N_8429,N_8253,N_8344);
or U8430 (N_8430,N_8214,N_8340);
nand U8431 (N_8431,N_8295,N_8391);
nand U8432 (N_8432,N_8358,N_8259);
and U8433 (N_8433,N_8317,N_8218);
nand U8434 (N_8434,N_8327,N_8388);
xor U8435 (N_8435,N_8245,N_8343);
nand U8436 (N_8436,N_8227,N_8309);
nor U8437 (N_8437,N_8220,N_8342);
xor U8438 (N_8438,N_8398,N_8336);
nand U8439 (N_8439,N_8394,N_8246);
or U8440 (N_8440,N_8230,N_8363);
nor U8441 (N_8441,N_8206,N_8233);
nor U8442 (N_8442,N_8211,N_8215);
or U8443 (N_8443,N_8354,N_8303);
and U8444 (N_8444,N_8339,N_8276);
nor U8445 (N_8445,N_8226,N_8200);
or U8446 (N_8446,N_8351,N_8288);
or U8447 (N_8447,N_8345,N_8316);
and U8448 (N_8448,N_8274,N_8390);
nand U8449 (N_8449,N_8247,N_8293);
or U8450 (N_8450,N_8333,N_8312);
nand U8451 (N_8451,N_8373,N_8262);
and U8452 (N_8452,N_8257,N_8294);
nor U8453 (N_8453,N_8395,N_8263);
xor U8454 (N_8454,N_8371,N_8208);
xor U8455 (N_8455,N_8224,N_8361);
nor U8456 (N_8456,N_8322,N_8360);
or U8457 (N_8457,N_8201,N_8234);
xnor U8458 (N_8458,N_8382,N_8380);
xnor U8459 (N_8459,N_8250,N_8205);
nand U8460 (N_8460,N_8331,N_8383);
nor U8461 (N_8461,N_8203,N_8243);
nor U8462 (N_8462,N_8362,N_8396);
or U8463 (N_8463,N_8365,N_8265);
nand U8464 (N_8464,N_8235,N_8231);
and U8465 (N_8465,N_8315,N_8369);
nand U8466 (N_8466,N_8329,N_8313);
nor U8467 (N_8467,N_8326,N_8290);
nor U8468 (N_8468,N_8271,N_8225);
and U8469 (N_8469,N_8216,N_8284);
and U8470 (N_8470,N_8254,N_8308);
nor U8471 (N_8471,N_8377,N_8272);
or U8472 (N_8472,N_8320,N_8355);
nand U8473 (N_8473,N_8297,N_8301);
nor U8474 (N_8474,N_8375,N_8325);
nor U8475 (N_8475,N_8338,N_8283);
xnor U8476 (N_8476,N_8242,N_8332);
nand U8477 (N_8477,N_8323,N_8240);
or U8478 (N_8478,N_8370,N_8258);
xor U8479 (N_8479,N_8244,N_8256);
xnor U8480 (N_8480,N_8334,N_8307);
xor U8481 (N_8481,N_8384,N_8241);
and U8482 (N_8482,N_8368,N_8238);
or U8483 (N_8483,N_8367,N_8379);
xnor U8484 (N_8484,N_8236,N_8249);
nor U8485 (N_8485,N_8376,N_8366);
nand U8486 (N_8486,N_8209,N_8305);
nand U8487 (N_8487,N_8381,N_8260);
or U8488 (N_8488,N_8202,N_8207);
nor U8489 (N_8489,N_8328,N_8221);
nand U8490 (N_8490,N_8310,N_8266);
or U8491 (N_8491,N_8364,N_8248);
xnor U8492 (N_8492,N_8347,N_8330);
xnor U8493 (N_8493,N_8341,N_8319);
nand U8494 (N_8494,N_8210,N_8287);
nand U8495 (N_8495,N_8212,N_8252);
xnor U8496 (N_8496,N_8296,N_8353);
or U8497 (N_8497,N_8324,N_8298);
nor U8498 (N_8498,N_8219,N_8213);
and U8499 (N_8499,N_8232,N_8204);
nand U8500 (N_8500,N_8353,N_8284);
nand U8501 (N_8501,N_8321,N_8319);
or U8502 (N_8502,N_8315,N_8297);
and U8503 (N_8503,N_8288,N_8371);
nand U8504 (N_8504,N_8216,N_8363);
nand U8505 (N_8505,N_8381,N_8315);
nor U8506 (N_8506,N_8370,N_8315);
nand U8507 (N_8507,N_8297,N_8336);
or U8508 (N_8508,N_8386,N_8227);
and U8509 (N_8509,N_8246,N_8205);
or U8510 (N_8510,N_8304,N_8213);
nand U8511 (N_8511,N_8275,N_8262);
xnor U8512 (N_8512,N_8281,N_8395);
nand U8513 (N_8513,N_8357,N_8223);
nor U8514 (N_8514,N_8381,N_8263);
xnor U8515 (N_8515,N_8212,N_8369);
and U8516 (N_8516,N_8252,N_8318);
and U8517 (N_8517,N_8383,N_8358);
xor U8518 (N_8518,N_8215,N_8231);
or U8519 (N_8519,N_8288,N_8223);
and U8520 (N_8520,N_8363,N_8311);
nand U8521 (N_8521,N_8393,N_8285);
nand U8522 (N_8522,N_8314,N_8376);
or U8523 (N_8523,N_8260,N_8347);
and U8524 (N_8524,N_8312,N_8231);
or U8525 (N_8525,N_8370,N_8391);
or U8526 (N_8526,N_8228,N_8346);
nor U8527 (N_8527,N_8358,N_8287);
nor U8528 (N_8528,N_8363,N_8314);
xor U8529 (N_8529,N_8228,N_8286);
nor U8530 (N_8530,N_8350,N_8219);
or U8531 (N_8531,N_8217,N_8250);
nor U8532 (N_8532,N_8297,N_8248);
nor U8533 (N_8533,N_8351,N_8309);
nand U8534 (N_8534,N_8252,N_8247);
nor U8535 (N_8535,N_8227,N_8316);
and U8536 (N_8536,N_8264,N_8395);
nand U8537 (N_8537,N_8386,N_8219);
and U8538 (N_8538,N_8321,N_8260);
xor U8539 (N_8539,N_8302,N_8254);
and U8540 (N_8540,N_8346,N_8326);
or U8541 (N_8541,N_8295,N_8288);
nor U8542 (N_8542,N_8373,N_8308);
xnor U8543 (N_8543,N_8371,N_8283);
or U8544 (N_8544,N_8232,N_8315);
nand U8545 (N_8545,N_8245,N_8261);
or U8546 (N_8546,N_8241,N_8224);
and U8547 (N_8547,N_8330,N_8336);
and U8548 (N_8548,N_8357,N_8213);
xnor U8549 (N_8549,N_8255,N_8243);
nor U8550 (N_8550,N_8399,N_8304);
nand U8551 (N_8551,N_8219,N_8308);
and U8552 (N_8552,N_8238,N_8294);
xor U8553 (N_8553,N_8313,N_8358);
nor U8554 (N_8554,N_8212,N_8285);
xor U8555 (N_8555,N_8319,N_8218);
xnor U8556 (N_8556,N_8211,N_8230);
nand U8557 (N_8557,N_8203,N_8304);
nor U8558 (N_8558,N_8339,N_8254);
and U8559 (N_8559,N_8399,N_8374);
and U8560 (N_8560,N_8281,N_8234);
nor U8561 (N_8561,N_8258,N_8357);
nand U8562 (N_8562,N_8359,N_8288);
xor U8563 (N_8563,N_8262,N_8260);
xnor U8564 (N_8564,N_8263,N_8251);
nor U8565 (N_8565,N_8211,N_8292);
xnor U8566 (N_8566,N_8228,N_8218);
nand U8567 (N_8567,N_8210,N_8352);
xor U8568 (N_8568,N_8261,N_8328);
nor U8569 (N_8569,N_8368,N_8258);
nand U8570 (N_8570,N_8321,N_8259);
or U8571 (N_8571,N_8208,N_8281);
nor U8572 (N_8572,N_8285,N_8227);
or U8573 (N_8573,N_8247,N_8280);
and U8574 (N_8574,N_8397,N_8335);
and U8575 (N_8575,N_8275,N_8361);
xor U8576 (N_8576,N_8352,N_8321);
or U8577 (N_8577,N_8295,N_8373);
and U8578 (N_8578,N_8249,N_8374);
or U8579 (N_8579,N_8278,N_8254);
or U8580 (N_8580,N_8337,N_8387);
xnor U8581 (N_8581,N_8333,N_8391);
xnor U8582 (N_8582,N_8287,N_8253);
nor U8583 (N_8583,N_8229,N_8294);
nor U8584 (N_8584,N_8213,N_8271);
and U8585 (N_8585,N_8261,N_8208);
or U8586 (N_8586,N_8327,N_8234);
xor U8587 (N_8587,N_8379,N_8343);
nor U8588 (N_8588,N_8290,N_8356);
or U8589 (N_8589,N_8372,N_8225);
and U8590 (N_8590,N_8221,N_8222);
or U8591 (N_8591,N_8380,N_8354);
or U8592 (N_8592,N_8284,N_8303);
nor U8593 (N_8593,N_8273,N_8252);
and U8594 (N_8594,N_8364,N_8392);
or U8595 (N_8595,N_8254,N_8344);
or U8596 (N_8596,N_8228,N_8353);
or U8597 (N_8597,N_8284,N_8275);
and U8598 (N_8598,N_8280,N_8288);
nor U8599 (N_8599,N_8274,N_8397);
and U8600 (N_8600,N_8516,N_8517);
nand U8601 (N_8601,N_8580,N_8443);
nand U8602 (N_8602,N_8412,N_8575);
and U8603 (N_8603,N_8579,N_8413);
or U8604 (N_8604,N_8556,N_8467);
and U8605 (N_8605,N_8424,N_8460);
and U8606 (N_8606,N_8403,N_8567);
nor U8607 (N_8607,N_8593,N_8493);
nand U8608 (N_8608,N_8594,N_8474);
nand U8609 (N_8609,N_8465,N_8511);
and U8610 (N_8610,N_8546,N_8523);
nand U8611 (N_8611,N_8566,N_8598);
nand U8612 (N_8612,N_8586,N_8491);
and U8613 (N_8613,N_8433,N_8436);
xor U8614 (N_8614,N_8439,N_8535);
xnor U8615 (N_8615,N_8525,N_8448);
or U8616 (N_8616,N_8539,N_8519);
xnor U8617 (N_8617,N_8574,N_8479);
xor U8618 (N_8618,N_8522,N_8464);
and U8619 (N_8619,N_8520,N_8422);
nand U8620 (N_8620,N_8502,N_8428);
nor U8621 (N_8621,N_8489,N_8563);
or U8622 (N_8622,N_8402,N_8447);
xnor U8623 (N_8623,N_8527,N_8559);
nand U8624 (N_8624,N_8568,N_8503);
and U8625 (N_8625,N_8507,N_8496);
nand U8626 (N_8626,N_8531,N_8417);
and U8627 (N_8627,N_8584,N_8437);
nand U8628 (N_8628,N_8440,N_8442);
xor U8629 (N_8629,N_8453,N_8435);
xnor U8630 (N_8630,N_8501,N_8459);
xor U8631 (N_8631,N_8547,N_8513);
xor U8632 (N_8632,N_8452,N_8557);
and U8633 (N_8633,N_8476,N_8540);
nor U8634 (N_8634,N_8521,N_8405);
or U8635 (N_8635,N_8423,N_8581);
nand U8636 (N_8636,N_8471,N_8562);
nor U8637 (N_8637,N_8429,N_8466);
nand U8638 (N_8638,N_8419,N_8401);
or U8639 (N_8639,N_8532,N_8404);
and U8640 (N_8640,N_8414,N_8461);
or U8641 (N_8641,N_8478,N_8542);
and U8642 (N_8642,N_8510,N_8400);
xnor U8643 (N_8643,N_8455,N_8427);
or U8644 (N_8644,N_8578,N_8583);
or U8645 (N_8645,N_8481,N_8449);
or U8646 (N_8646,N_8468,N_8537);
nor U8647 (N_8647,N_8569,N_8490);
and U8648 (N_8648,N_8444,N_8555);
or U8649 (N_8649,N_8446,N_8571);
xnor U8650 (N_8650,N_8530,N_8512);
and U8651 (N_8651,N_8500,N_8469);
nor U8652 (N_8652,N_8420,N_8504);
or U8653 (N_8653,N_8497,N_8484);
nand U8654 (N_8654,N_8554,N_8411);
or U8655 (N_8655,N_8591,N_8408);
xor U8656 (N_8656,N_8548,N_8473);
and U8657 (N_8657,N_8553,N_8552);
nand U8658 (N_8658,N_8544,N_8434);
nor U8659 (N_8659,N_8589,N_8426);
or U8660 (N_8660,N_8470,N_8592);
xor U8661 (N_8661,N_8432,N_8526);
nor U8662 (N_8662,N_8475,N_8488);
or U8663 (N_8663,N_8518,N_8529);
and U8664 (N_8664,N_8450,N_8458);
xnor U8665 (N_8665,N_8498,N_8438);
and U8666 (N_8666,N_8538,N_8406);
nor U8667 (N_8667,N_8409,N_8418);
and U8668 (N_8668,N_8585,N_8590);
or U8669 (N_8669,N_8456,N_8508);
xor U8670 (N_8670,N_8445,N_8582);
xor U8671 (N_8671,N_8536,N_8492);
xnor U8672 (N_8672,N_8560,N_8485);
nor U8673 (N_8673,N_8499,N_8477);
xor U8674 (N_8674,N_8577,N_8543);
xor U8675 (N_8675,N_8587,N_8416);
nor U8676 (N_8676,N_8573,N_8533);
nand U8677 (N_8677,N_8483,N_8597);
and U8678 (N_8678,N_8482,N_8415);
and U8679 (N_8679,N_8451,N_8421);
nor U8680 (N_8680,N_8551,N_8425);
or U8681 (N_8681,N_8514,N_8549);
and U8682 (N_8682,N_8524,N_8430);
and U8683 (N_8683,N_8599,N_8528);
nand U8684 (N_8684,N_8565,N_8595);
xnor U8685 (N_8685,N_8407,N_8457);
or U8686 (N_8686,N_8486,N_8495);
nor U8687 (N_8687,N_8509,N_8441);
nor U8688 (N_8688,N_8494,N_8410);
and U8689 (N_8689,N_8454,N_8515);
or U8690 (N_8690,N_8534,N_8463);
xnor U8691 (N_8691,N_8505,N_8558);
and U8692 (N_8692,N_8541,N_8545);
nand U8693 (N_8693,N_8472,N_8572);
xor U8694 (N_8694,N_8561,N_8550);
or U8695 (N_8695,N_8576,N_8506);
nor U8696 (N_8696,N_8596,N_8564);
nor U8697 (N_8697,N_8588,N_8480);
nor U8698 (N_8698,N_8462,N_8431);
or U8699 (N_8699,N_8487,N_8570);
or U8700 (N_8700,N_8588,N_8432);
and U8701 (N_8701,N_8402,N_8544);
nor U8702 (N_8702,N_8460,N_8561);
or U8703 (N_8703,N_8525,N_8418);
or U8704 (N_8704,N_8438,N_8418);
nand U8705 (N_8705,N_8421,N_8437);
or U8706 (N_8706,N_8443,N_8464);
xor U8707 (N_8707,N_8442,N_8480);
nor U8708 (N_8708,N_8592,N_8545);
nand U8709 (N_8709,N_8528,N_8554);
and U8710 (N_8710,N_8568,N_8491);
nor U8711 (N_8711,N_8452,N_8462);
nor U8712 (N_8712,N_8517,N_8436);
or U8713 (N_8713,N_8424,N_8444);
nor U8714 (N_8714,N_8462,N_8406);
or U8715 (N_8715,N_8518,N_8521);
and U8716 (N_8716,N_8424,N_8401);
or U8717 (N_8717,N_8434,N_8548);
and U8718 (N_8718,N_8583,N_8515);
and U8719 (N_8719,N_8422,N_8544);
xor U8720 (N_8720,N_8568,N_8463);
xnor U8721 (N_8721,N_8564,N_8406);
xor U8722 (N_8722,N_8410,N_8503);
or U8723 (N_8723,N_8547,N_8586);
nor U8724 (N_8724,N_8495,N_8548);
nand U8725 (N_8725,N_8436,N_8534);
nand U8726 (N_8726,N_8573,N_8591);
xnor U8727 (N_8727,N_8538,N_8533);
nor U8728 (N_8728,N_8501,N_8451);
nand U8729 (N_8729,N_8412,N_8563);
and U8730 (N_8730,N_8488,N_8514);
nand U8731 (N_8731,N_8510,N_8478);
xor U8732 (N_8732,N_8442,N_8438);
nor U8733 (N_8733,N_8551,N_8404);
nor U8734 (N_8734,N_8445,N_8553);
xnor U8735 (N_8735,N_8573,N_8439);
xnor U8736 (N_8736,N_8430,N_8487);
and U8737 (N_8737,N_8502,N_8511);
nand U8738 (N_8738,N_8460,N_8448);
nand U8739 (N_8739,N_8405,N_8524);
nor U8740 (N_8740,N_8427,N_8493);
nor U8741 (N_8741,N_8536,N_8430);
nand U8742 (N_8742,N_8596,N_8584);
nor U8743 (N_8743,N_8537,N_8504);
or U8744 (N_8744,N_8538,N_8410);
nand U8745 (N_8745,N_8531,N_8533);
and U8746 (N_8746,N_8551,N_8586);
nand U8747 (N_8747,N_8443,N_8537);
or U8748 (N_8748,N_8577,N_8582);
or U8749 (N_8749,N_8403,N_8526);
xor U8750 (N_8750,N_8470,N_8436);
nand U8751 (N_8751,N_8409,N_8476);
or U8752 (N_8752,N_8586,N_8533);
xnor U8753 (N_8753,N_8490,N_8458);
xor U8754 (N_8754,N_8430,N_8550);
xor U8755 (N_8755,N_8417,N_8542);
nor U8756 (N_8756,N_8546,N_8562);
or U8757 (N_8757,N_8520,N_8586);
and U8758 (N_8758,N_8494,N_8422);
nor U8759 (N_8759,N_8553,N_8598);
and U8760 (N_8760,N_8544,N_8464);
and U8761 (N_8761,N_8422,N_8517);
and U8762 (N_8762,N_8534,N_8487);
and U8763 (N_8763,N_8452,N_8564);
nand U8764 (N_8764,N_8410,N_8509);
and U8765 (N_8765,N_8569,N_8501);
nand U8766 (N_8766,N_8505,N_8584);
nor U8767 (N_8767,N_8422,N_8442);
or U8768 (N_8768,N_8576,N_8502);
or U8769 (N_8769,N_8574,N_8495);
and U8770 (N_8770,N_8562,N_8534);
xnor U8771 (N_8771,N_8527,N_8488);
or U8772 (N_8772,N_8496,N_8443);
or U8773 (N_8773,N_8403,N_8487);
xor U8774 (N_8774,N_8501,N_8449);
and U8775 (N_8775,N_8529,N_8510);
nor U8776 (N_8776,N_8562,N_8470);
nand U8777 (N_8777,N_8566,N_8498);
nand U8778 (N_8778,N_8444,N_8594);
xor U8779 (N_8779,N_8404,N_8568);
or U8780 (N_8780,N_8463,N_8512);
and U8781 (N_8781,N_8443,N_8531);
nor U8782 (N_8782,N_8540,N_8517);
or U8783 (N_8783,N_8459,N_8576);
xnor U8784 (N_8784,N_8464,N_8453);
nor U8785 (N_8785,N_8445,N_8436);
or U8786 (N_8786,N_8555,N_8500);
or U8787 (N_8787,N_8427,N_8483);
nand U8788 (N_8788,N_8554,N_8579);
or U8789 (N_8789,N_8566,N_8564);
nand U8790 (N_8790,N_8542,N_8419);
nand U8791 (N_8791,N_8524,N_8492);
nor U8792 (N_8792,N_8499,N_8484);
xor U8793 (N_8793,N_8593,N_8437);
and U8794 (N_8794,N_8460,N_8523);
or U8795 (N_8795,N_8467,N_8511);
nand U8796 (N_8796,N_8506,N_8465);
nand U8797 (N_8797,N_8474,N_8572);
nor U8798 (N_8798,N_8506,N_8521);
nand U8799 (N_8799,N_8549,N_8577);
nor U8800 (N_8800,N_8609,N_8704);
xor U8801 (N_8801,N_8781,N_8710);
and U8802 (N_8802,N_8799,N_8721);
nand U8803 (N_8803,N_8771,N_8720);
xor U8804 (N_8804,N_8715,N_8755);
xor U8805 (N_8805,N_8770,N_8775);
nand U8806 (N_8806,N_8631,N_8675);
and U8807 (N_8807,N_8669,N_8772);
or U8808 (N_8808,N_8688,N_8727);
and U8809 (N_8809,N_8757,N_8694);
xnor U8810 (N_8810,N_8706,N_8790);
nor U8811 (N_8811,N_8712,N_8789);
nor U8812 (N_8812,N_8606,N_8700);
and U8813 (N_8813,N_8782,N_8634);
nor U8814 (N_8814,N_8645,N_8760);
nand U8815 (N_8815,N_8768,N_8730);
nor U8816 (N_8816,N_8797,N_8649);
nand U8817 (N_8817,N_8708,N_8713);
nand U8818 (N_8818,N_8640,N_8732);
xnor U8819 (N_8819,N_8660,N_8601);
nand U8820 (N_8820,N_8679,N_8671);
and U8821 (N_8821,N_8641,N_8703);
xnor U8822 (N_8822,N_8729,N_8756);
nor U8823 (N_8823,N_8745,N_8627);
or U8824 (N_8824,N_8636,N_8743);
nor U8825 (N_8825,N_8600,N_8655);
nand U8826 (N_8826,N_8659,N_8728);
nand U8827 (N_8827,N_8750,N_8615);
nor U8828 (N_8828,N_8722,N_8748);
xor U8829 (N_8829,N_8714,N_8647);
and U8830 (N_8830,N_8698,N_8709);
or U8831 (N_8831,N_8644,N_8736);
nor U8832 (N_8832,N_8603,N_8677);
and U8833 (N_8833,N_8765,N_8749);
nand U8834 (N_8834,N_8784,N_8666);
and U8835 (N_8835,N_8786,N_8758);
and U8836 (N_8836,N_8608,N_8651);
and U8837 (N_8837,N_8739,N_8624);
xnor U8838 (N_8838,N_8718,N_8761);
or U8839 (N_8839,N_8779,N_8637);
nor U8840 (N_8840,N_8658,N_8733);
nand U8841 (N_8841,N_8662,N_8629);
nor U8842 (N_8842,N_8726,N_8780);
nor U8843 (N_8843,N_8602,N_8626);
xor U8844 (N_8844,N_8687,N_8740);
or U8845 (N_8845,N_8751,N_8796);
and U8846 (N_8846,N_8793,N_8696);
nor U8847 (N_8847,N_8676,N_8664);
nand U8848 (N_8848,N_8791,N_8723);
nand U8849 (N_8849,N_8734,N_8635);
and U8850 (N_8850,N_8663,N_8693);
nor U8851 (N_8851,N_8737,N_8621);
xnor U8852 (N_8852,N_8618,N_8652);
nand U8853 (N_8853,N_8762,N_8678);
nand U8854 (N_8854,N_8668,N_8691);
and U8855 (N_8855,N_8632,N_8616);
nand U8856 (N_8856,N_8656,N_8628);
and U8857 (N_8857,N_8605,N_8759);
or U8858 (N_8858,N_8633,N_8686);
xor U8859 (N_8859,N_8744,N_8643);
and U8860 (N_8860,N_8735,N_8705);
nand U8861 (N_8861,N_8701,N_8612);
and U8862 (N_8862,N_8672,N_8648);
nor U8863 (N_8863,N_8630,N_8763);
nand U8864 (N_8864,N_8683,N_8690);
or U8865 (N_8865,N_8638,N_8613);
nand U8866 (N_8866,N_8753,N_8766);
xor U8867 (N_8867,N_8680,N_8661);
and U8868 (N_8868,N_8610,N_8724);
nand U8869 (N_8869,N_8699,N_8716);
or U8870 (N_8870,N_8769,N_8614);
nand U8871 (N_8871,N_8767,N_8682);
and U8872 (N_8872,N_8795,N_8695);
and U8873 (N_8873,N_8673,N_8692);
nand U8874 (N_8874,N_8717,N_8617);
nand U8875 (N_8875,N_8741,N_8667);
nor U8876 (N_8876,N_8697,N_8611);
xor U8877 (N_8877,N_8738,N_8702);
or U8878 (N_8878,N_8689,N_8774);
or U8879 (N_8879,N_8776,N_8747);
nand U8880 (N_8880,N_8711,N_8646);
nor U8881 (N_8881,N_8639,N_8681);
nor U8882 (N_8882,N_8719,N_8625);
nand U8883 (N_8883,N_8684,N_8783);
nand U8884 (N_8884,N_8764,N_8731);
nor U8885 (N_8885,N_8607,N_8707);
or U8886 (N_8886,N_8754,N_8650);
nor U8887 (N_8887,N_8623,N_8794);
nor U8888 (N_8888,N_8665,N_8798);
and U8889 (N_8889,N_8773,N_8792);
nand U8890 (N_8890,N_8619,N_8657);
nand U8891 (N_8891,N_8653,N_8604);
or U8892 (N_8892,N_8620,N_8654);
xnor U8893 (N_8893,N_8642,N_8778);
and U8894 (N_8894,N_8622,N_8725);
and U8895 (N_8895,N_8787,N_8777);
xor U8896 (N_8896,N_8785,N_8742);
nor U8897 (N_8897,N_8674,N_8670);
nand U8898 (N_8898,N_8788,N_8752);
and U8899 (N_8899,N_8685,N_8746);
and U8900 (N_8900,N_8714,N_8791);
and U8901 (N_8901,N_8600,N_8634);
nand U8902 (N_8902,N_8744,N_8665);
nor U8903 (N_8903,N_8700,N_8638);
or U8904 (N_8904,N_8664,N_8691);
or U8905 (N_8905,N_8660,N_8728);
nand U8906 (N_8906,N_8704,N_8676);
and U8907 (N_8907,N_8612,N_8726);
or U8908 (N_8908,N_8607,N_8649);
nand U8909 (N_8909,N_8700,N_8678);
xnor U8910 (N_8910,N_8767,N_8607);
xnor U8911 (N_8911,N_8764,N_8664);
or U8912 (N_8912,N_8705,N_8611);
and U8913 (N_8913,N_8610,N_8692);
nand U8914 (N_8914,N_8686,N_8707);
xnor U8915 (N_8915,N_8669,N_8703);
nand U8916 (N_8916,N_8654,N_8739);
or U8917 (N_8917,N_8759,N_8703);
and U8918 (N_8918,N_8751,N_8719);
nand U8919 (N_8919,N_8627,N_8749);
or U8920 (N_8920,N_8636,N_8662);
nand U8921 (N_8921,N_8610,N_8710);
and U8922 (N_8922,N_8766,N_8609);
xnor U8923 (N_8923,N_8675,N_8764);
nand U8924 (N_8924,N_8749,N_8735);
nor U8925 (N_8925,N_8675,N_8611);
nand U8926 (N_8926,N_8733,N_8774);
nand U8927 (N_8927,N_8607,N_8712);
xor U8928 (N_8928,N_8710,N_8620);
nor U8929 (N_8929,N_8764,N_8613);
or U8930 (N_8930,N_8650,N_8605);
xnor U8931 (N_8931,N_8665,N_8713);
xor U8932 (N_8932,N_8773,N_8649);
xor U8933 (N_8933,N_8738,N_8637);
and U8934 (N_8934,N_8704,N_8610);
nand U8935 (N_8935,N_8755,N_8683);
and U8936 (N_8936,N_8616,N_8714);
or U8937 (N_8937,N_8620,N_8633);
xnor U8938 (N_8938,N_8764,N_8676);
and U8939 (N_8939,N_8759,N_8607);
and U8940 (N_8940,N_8745,N_8668);
nor U8941 (N_8941,N_8794,N_8778);
nand U8942 (N_8942,N_8631,N_8671);
and U8943 (N_8943,N_8799,N_8715);
and U8944 (N_8944,N_8710,N_8611);
xor U8945 (N_8945,N_8664,N_8681);
nor U8946 (N_8946,N_8710,N_8798);
nand U8947 (N_8947,N_8649,N_8618);
nor U8948 (N_8948,N_8628,N_8676);
and U8949 (N_8949,N_8689,N_8602);
nor U8950 (N_8950,N_8656,N_8610);
nor U8951 (N_8951,N_8741,N_8660);
or U8952 (N_8952,N_8720,N_8750);
xnor U8953 (N_8953,N_8630,N_8783);
nor U8954 (N_8954,N_8627,N_8707);
or U8955 (N_8955,N_8777,N_8732);
or U8956 (N_8956,N_8625,N_8702);
nand U8957 (N_8957,N_8766,N_8788);
nor U8958 (N_8958,N_8696,N_8748);
xor U8959 (N_8959,N_8748,N_8612);
and U8960 (N_8960,N_8655,N_8649);
or U8961 (N_8961,N_8738,N_8765);
or U8962 (N_8962,N_8734,N_8755);
or U8963 (N_8963,N_8678,N_8775);
nand U8964 (N_8964,N_8654,N_8601);
nor U8965 (N_8965,N_8688,N_8767);
xnor U8966 (N_8966,N_8737,N_8691);
xnor U8967 (N_8967,N_8667,N_8796);
xnor U8968 (N_8968,N_8776,N_8628);
or U8969 (N_8969,N_8741,N_8677);
or U8970 (N_8970,N_8755,N_8623);
nand U8971 (N_8971,N_8716,N_8600);
or U8972 (N_8972,N_8717,N_8719);
nand U8973 (N_8973,N_8766,N_8656);
or U8974 (N_8974,N_8600,N_8787);
or U8975 (N_8975,N_8748,N_8618);
xor U8976 (N_8976,N_8787,N_8682);
nor U8977 (N_8977,N_8738,N_8655);
nor U8978 (N_8978,N_8637,N_8619);
nor U8979 (N_8979,N_8697,N_8729);
or U8980 (N_8980,N_8610,N_8737);
nand U8981 (N_8981,N_8607,N_8736);
xnor U8982 (N_8982,N_8787,N_8684);
or U8983 (N_8983,N_8705,N_8762);
and U8984 (N_8984,N_8655,N_8739);
or U8985 (N_8985,N_8616,N_8718);
or U8986 (N_8986,N_8706,N_8679);
nand U8987 (N_8987,N_8612,N_8624);
or U8988 (N_8988,N_8676,N_8654);
nand U8989 (N_8989,N_8619,N_8734);
nor U8990 (N_8990,N_8645,N_8750);
or U8991 (N_8991,N_8661,N_8767);
and U8992 (N_8992,N_8799,N_8684);
nor U8993 (N_8993,N_8761,N_8679);
or U8994 (N_8994,N_8791,N_8670);
nand U8995 (N_8995,N_8735,N_8704);
or U8996 (N_8996,N_8775,N_8604);
or U8997 (N_8997,N_8654,N_8779);
nor U8998 (N_8998,N_8638,N_8761);
or U8999 (N_8999,N_8635,N_8623);
or U9000 (N_9000,N_8852,N_8900);
nor U9001 (N_9001,N_8965,N_8804);
xor U9002 (N_9002,N_8979,N_8993);
or U9003 (N_9003,N_8917,N_8801);
nor U9004 (N_9004,N_8836,N_8942);
xor U9005 (N_9005,N_8894,N_8991);
or U9006 (N_9006,N_8937,N_8901);
nand U9007 (N_9007,N_8858,N_8998);
and U9008 (N_9008,N_8975,N_8859);
nand U9009 (N_9009,N_8841,N_8924);
nand U9010 (N_9010,N_8983,N_8995);
nor U9011 (N_9011,N_8854,N_8954);
or U9012 (N_9012,N_8881,N_8961);
or U9013 (N_9013,N_8839,N_8985);
nor U9014 (N_9014,N_8948,N_8892);
or U9015 (N_9015,N_8884,N_8811);
xor U9016 (N_9016,N_8989,N_8887);
xnor U9017 (N_9017,N_8981,N_8889);
or U9018 (N_9018,N_8963,N_8909);
xnor U9019 (N_9019,N_8997,N_8810);
and U9020 (N_9020,N_8941,N_8912);
nor U9021 (N_9021,N_8932,N_8972);
nor U9022 (N_9022,N_8971,N_8931);
and U9023 (N_9023,N_8980,N_8960);
nor U9024 (N_9024,N_8815,N_8830);
or U9025 (N_9025,N_8949,N_8896);
and U9026 (N_9026,N_8822,N_8809);
or U9027 (N_9027,N_8862,N_8976);
nor U9028 (N_9028,N_8846,N_8853);
nand U9029 (N_9029,N_8819,N_8844);
or U9030 (N_9030,N_8927,N_8869);
nand U9031 (N_9031,N_8977,N_8920);
or U9032 (N_9032,N_8842,N_8870);
and U9033 (N_9033,N_8899,N_8866);
xnor U9034 (N_9034,N_8848,N_8970);
or U9035 (N_9035,N_8969,N_8863);
xor U9036 (N_9036,N_8888,N_8933);
or U9037 (N_9037,N_8945,N_8918);
xor U9038 (N_9038,N_8802,N_8906);
xor U9039 (N_9039,N_8907,N_8902);
and U9040 (N_9040,N_8895,N_8905);
and U9041 (N_9041,N_8818,N_8856);
nor U9042 (N_9042,N_8925,N_8832);
nand U9043 (N_9043,N_8956,N_8807);
or U9044 (N_9044,N_8908,N_8934);
nand U9045 (N_9045,N_8929,N_8939);
nor U9046 (N_9046,N_8915,N_8879);
and U9047 (N_9047,N_8827,N_8868);
or U9048 (N_9048,N_8872,N_8957);
nand U9049 (N_9049,N_8845,N_8861);
xnor U9050 (N_9050,N_8871,N_8978);
and U9051 (N_9051,N_8875,N_8886);
nand U9052 (N_9052,N_8880,N_8820);
xnor U9053 (N_9053,N_8851,N_8834);
or U9054 (N_9054,N_8926,N_8883);
or U9055 (N_9055,N_8816,N_8930);
or U9056 (N_9056,N_8857,N_8999);
or U9057 (N_9057,N_8953,N_8951);
or U9058 (N_9058,N_8987,N_8946);
xor U9059 (N_9059,N_8921,N_8885);
or U9060 (N_9060,N_8964,N_8877);
xor U9061 (N_9061,N_8867,N_8800);
and U9062 (N_9062,N_8911,N_8966);
nor U9063 (N_9063,N_8855,N_8805);
nand U9064 (N_9064,N_8974,N_8882);
nor U9065 (N_9065,N_8944,N_8916);
nand U9066 (N_9066,N_8840,N_8829);
or U9067 (N_9067,N_8984,N_8943);
nand U9068 (N_9068,N_8837,N_8986);
nor U9069 (N_9069,N_8824,N_8996);
nor U9070 (N_9070,N_8923,N_8847);
and U9071 (N_9071,N_8982,N_8950);
or U9072 (N_9072,N_8865,N_8828);
xnor U9073 (N_9073,N_8903,N_8947);
and U9074 (N_9074,N_8973,N_8878);
and U9075 (N_9075,N_8940,N_8919);
xor U9076 (N_9076,N_8835,N_8860);
and U9077 (N_9077,N_8914,N_8922);
and U9078 (N_9078,N_8833,N_8959);
nand U9079 (N_9079,N_8817,N_8814);
and U9080 (N_9080,N_8967,N_8803);
xnor U9081 (N_9081,N_8890,N_8808);
nor U9082 (N_9082,N_8994,N_8864);
nor U9083 (N_9083,N_8893,N_8988);
and U9084 (N_9084,N_8813,N_8938);
nor U9085 (N_9085,N_8850,N_8891);
xor U9086 (N_9086,N_8936,N_8806);
and U9087 (N_9087,N_8955,N_8873);
nand U9088 (N_9088,N_8874,N_8910);
or U9089 (N_9089,N_8904,N_8962);
xnor U9090 (N_9090,N_8935,N_8823);
or U9091 (N_9091,N_8849,N_8952);
or U9092 (N_9092,N_8897,N_8821);
or U9093 (N_9093,N_8843,N_8990);
nand U9094 (N_9094,N_8913,N_8826);
or U9095 (N_9095,N_8928,N_8825);
and U9096 (N_9096,N_8876,N_8958);
nand U9097 (N_9097,N_8992,N_8812);
nand U9098 (N_9098,N_8838,N_8898);
xor U9099 (N_9099,N_8831,N_8968);
xor U9100 (N_9100,N_8895,N_8965);
nor U9101 (N_9101,N_8889,N_8946);
and U9102 (N_9102,N_8825,N_8916);
or U9103 (N_9103,N_8825,N_8866);
nand U9104 (N_9104,N_8923,N_8948);
nand U9105 (N_9105,N_8934,N_8917);
or U9106 (N_9106,N_8854,N_8858);
nand U9107 (N_9107,N_8816,N_8810);
xor U9108 (N_9108,N_8929,N_8971);
and U9109 (N_9109,N_8927,N_8917);
and U9110 (N_9110,N_8854,N_8902);
nand U9111 (N_9111,N_8825,N_8914);
xor U9112 (N_9112,N_8905,N_8913);
or U9113 (N_9113,N_8940,N_8992);
or U9114 (N_9114,N_8830,N_8979);
or U9115 (N_9115,N_8907,N_8820);
and U9116 (N_9116,N_8961,N_8937);
or U9117 (N_9117,N_8842,N_8921);
xor U9118 (N_9118,N_8846,N_8816);
nor U9119 (N_9119,N_8813,N_8979);
or U9120 (N_9120,N_8936,N_8940);
nand U9121 (N_9121,N_8918,N_8831);
nor U9122 (N_9122,N_8920,N_8826);
xnor U9123 (N_9123,N_8833,N_8907);
and U9124 (N_9124,N_8957,N_8802);
nand U9125 (N_9125,N_8872,N_8981);
xnor U9126 (N_9126,N_8883,N_8845);
nor U9127 (N_9127,N_8979,N_8917);
or U9128 (N_9128,N_8919,N_8996);
nand U9129 (N_9129,N_8906,N_8826);
or U9130 (N_9130,N_8943,N_8965);
and U9131 (N_9131,N_8889,N_8956);
or U9132 (N_9132,N_8996,N_8822);
or U9133 (N_9133,N_8888,N_8844);
and U9134 (N_9134,N_8964,N_8979);
or U9135 (N_9135,N_8832,N_8807);
or U9136 (N_9136,N_8995,N_8828);
nand U9137 (N_9137,N_8838,N_8881);
nand U9138 (N_9138,N_8850,N_8846);
xnor U9139 (N_9139,N_8975,N_8947);
and U9140 (N_9140,N_8826,N_8982);
and U9141 (N_9141,N_8978,N_8955);
or U9142 (N_9142,N_8860,N_8824);
nand U9143 (N_9143,N_8931,N_8843);
nand U9144 (N_9144,N_8970,N_8855);
nor U9145 (N_9145,N_8992,N_8934);
and U9146 (N_9146,N_8955,N_8849);
and U9147 (N_9147,N_8845,N_8855);
or U9148 (N_9148,N_8964,N_8842);
nor U9149 (N_9149,N_8882,N_8903);
nand U9150 (N_9150,N_8924,N_8874);
nand U9151 (N_9151,N_8962,N_8913);
nand U9152 (N_9152,N_8980,N_8827);
or U9153 (N_9153,N_8878,N_8979);
nand U9154 (N_9154,N_8853,N_8859);
nor U9155 (N_9155,N_8847,N_8808);
nor U9156 (N_9156,N_8978,N_8891);
nor U9157 (N_9157,N_8982,N_8917);
nor U9158 (N_9158,N_8868,N_8801);
nor U9159 (N_9159,N_8960,N_8902);
nand U9160 (N_9160,N_8968,N_8816);
nand U9161 (N_9161,N_8898,N_8897);
or U9162 (N_9162,N_8980,N_8987);
nor U9163 (N_9163,N_8952,N_8807);
nor U9164 (N_9164,N_8899,N_8816);
nor U9165 (N_9165,N_8997,N_8963);
or U9166 (N_9166,N_8955,N_8801);
or U9167 (N_9167,N_8849,N_8940);
nor U9168 (N_9168,N_8827,N_8822);
nor U9169 (N_9169,N_8916,N_8950);
xnor U9170 (N_9170,N_8873,N_8878);
nand U9171 (N_9171,N_8984,N_8976);
nand U9172 (N_9172,N_8850,N_8937);
xnor U9173 (N_9173,N_8831,N_8875);
xnor U9174 (N_9174,N_8896,N_8824);
xor U9175 (N_9175,N_8924,N_8870);
or U9176 (N_9176,N_8985,N_8929);
nor U9177 (N_9177,N_8873,N_8862);
xor U9178 (N_9178,N_8995,N_8851);
xnor U9179 (N_9179,N_8815,N_8932);
nor U9180 (N_9180,N_8998,N_8956);
xnor U9181 (N_9181,N_8863,N_8802);
nand U9182 (N_9182,N_8958,N_8832);
nor U9183 (N_9183,N_8845,N_8998);
nand U9184 (N_9184,N_8967,N_8895);
and U9185 (N_9185,N_8945,N_8922);
nor U9186 (N_9186,N_8864,N_8827);
nand U9187 (N_9187,N_8998,N_8800);
and U9188 (N_9188,N_8836,N_8971);
xnor U9189 (N_9189,N_8953,N_8968);
nor U9190 (N_9190,N_8901,N_8913);
xnor U9191 (N_9191,N_8949,N_8899);
or U9192 (N_9192,N_8929,N_8926);
and U9193 (N_9193,N_8828,N_8918);
xnor U9194 (N_9194,N_8818,N_8965);
xor U9195 (N_9195,N_8824,N_8989);
nor U9196 (N_9196,N_8910,N_8869);
nand U9197 (N_9197,N_8919,N_8838);
nand U9198 (N_9198,N_8837,N_8999);
and U9199 (N_9199,N_8951,N_8808);
nand U9200 (N_9200,N_9050,N_9082);
or U9201 (N_9201,N_9181,N_9143);
nand U9202 (N_9202,N_9100,N_9025);
or U9203 (N_9203,N_9095,N_9020);
or U9204 (N_9204,N_9006,N_9156);
or U9205 (N_9205,N_9047,N_9105);
xnor U9206 (N_9206,N_9071,N_9176);
nand U9207 (N_9207,N_9014,N_9033);
xor U9208 (N_9208,N_9118,N_9192);
xnor U9209 (N_9209,N_9193,N_9116);
nor U9210 (N_9210,N_9067,N_9174);
nor U9211 (N_9211,N_9115,N_9180);
and U9212 (N_9212,N_9102,N_9128);
or U9213 (N_9213,N_9109,N_9088);
xor U9214 (N_9214,N_9195,N_9114);
xor U9215 (N_9215,N_9106,N_9149);
and U9216 (N_9216,N_9093,N_9089);
xnor U9217 (N_9217,N_9189,N_9055);
xor U9218 (N_9218,N_9157,N_9019);
or U9219 (N_9219,N_9043,N_9096);
or U9220 (N_9220,N_9099,N_9085);
xnor U9221 (N_9221,N_9135,N_9015);
nand U9222 (N_9222,N_9173,N_9198);
nor U9223 (N_9223,N_9162,N_9197);
and U9224 (N_9224,N_9098,N_9112);
or U9225 (N_9225,N_9134,N_9130);
or U9226 (N_9226,N_9132,N_9147);
or U9227 (N_9227,N_9002,N_9107);
xor U9228 (N_9228,N_9026,N_9196);
xnor U9229 (N_9229,N_9138,N_9178);
or U9230 (N_9230,N_9078,N_9042);
nor U9231 (N_9231,N_9150,N_9171);
nor U9232 (N_9232,N_9104,N_9139);
and U9233 (N_9233,N_9076,N_9090);
nor U9234 (N_9234,N_9072,N_9077);
nor U9235 (N_9235,N_9080,N_9123);
or U9236 (N_9236,N_9191,N_9040);
nand U9237 (N_9237,N_9003,N_9053);
or U9238 (N_9238,N_9068,N_9008);
and U9239 (N_9239,N_9166,N_9129);
nand U9240 (N_9240,N_9169,N_9185);
xnor U9241 (N_9241,N_9187,N_9190);
nor U9242 (N_9242,N_9137,N_9086);
nor U9243 (N_9243,N_9029,N_9092);
xnor U9244 (N_9244,N_9152,N_9167);
or U9245 (N_9245,N_9126,N_9108);
xnor U9246 (N_9246,N_9037,N_9060);
nand U9247 (N_9247,N_9151,N_9188);
and U9248 (N_9248,N_9079,N_9016);
or U9249 (N_9249,N_9087,N_9120);
nor U9250 (N_9250,N_9165,N_9124);
nor U9251 (N_9251,N_9061,N_9034);
xnor U9252 (N_9252,N_9035,N_9127);
nor U9253 (N_9253,N_9010,N_9009);
nor U9254 (N_9254,N_9011,N_9119);
and U9255 (N_9255,N_9172,N_9063);
or U9256 (N_9256,N_9199,N_9094);
xor U9257 (N_9257,N_9057,N_9177);
nand U9258 (N_9258,N_9121,N_9031);
or U9259 (N_9259,N_9027,N_9039);
nand U9260 (N_9260,N_9045,N_9044);
and U9261 (N_9261,N_9141,N_9160);
nor U9262 (N_9262,N_9184,N_9021);
nand U9263 (N_9263,N_9049,N_9194);
or U9264 (N_9264,N_9164,N_9070);
nor U9265 (N_9265,N_9113,N_9153);
or U9266 (N_9266,N_9030,N_9133);
nand U9267 (N_9267,N_9065,N_9028);
or U9268 (N_9268,N_9110,N_9144);
or U9269 (N_9269,N_9001,N_9125);
or U9270 (N_9270,N_9073,N_9154);
xor U9271 (N_9271,N_9148,N_9056);
nor U9272 (N_9272,N_9117,N_9101);
xnor U9273 (N_9273,N_9179,N_9059);
and U9274 (N_9274,N_9022,N_9048);
nor U9275 (N_9275,N_9159,N_9182);
nor U9276 (N_9276,N_9066,N_9024);
nand U9277 (N_9277,N_9052,N_9142);
nor U9278 (N_9278,N_9032,N_9136);
and U9279 (N_9279,N_9081,N_9005);
or U9280 (N_9280,N_9122,N_9062);
nand U9281 (N_9281,N_9097,N_9064);
nor U9282 (N_9282,N_9038,N_9023);
and U9283 (N_9283,N_9007,N_9046);
nor U9284 (N_9284,N_9013,N_9004);
xnor U9285 (N_9285,N_9069,N_9054);
and U9286 (N_9286,N_9018,N_9170);
xor U9287 (N_9287,N_9161,N_9146);
and U9288 (N_9288,N_9186,N_9163);
xor U9289 (N_9289,N_9091,N_9084);
nor U9290 (N_9290,N_9075,N_9058);
nor U9291 (N_9291,N_9155,N_9168);
nor U9292 (N_9292,N_9158,N_9103);
nand U9293 (N_9293,N_9012,N_9017);
and U9294 (N_9294,N_9041,N_9036);
nand U9295 (N_9295,N_9083,N_9140);
and U9296 (N_9296,N_9175,N_9051);
and U9297 (N_9297,N_9131,N_9111);
nor U9298 (N_9298,N_9183,N_9000);
nor U9299 (N_9299,N_9074,N_9145);
and U9300 (N_9300,N_9018,N_9027);
xor U9301 (N_9301,N_9189,N_9069);
nor U9302 (N_9302,N_9196,N_9122);
or U9303 (N_9303,N_9074,N_9041);
or U9304 (N_9304,N_9183,N_9119);
xnor U9305 (N_9305,N_9024,N_9061);
xnor U9306 (N_9306,N_9192,N_9000);
nor U9307 (N_9307,N_9062,N_9113);
or U9308 (N_9308,N_9061,N_9177);
and U9309 (N_9309,N_9033,N_9025);
xnor U9310 (N_9310,N_9105,N_9016);
and U9311 (N_9311,N_9021,N_9140);
nor U9312 (N_9312,N_9110,N_9018);
or U9313 (N_9313,N_9191,N_9070);
nor U9314 (N_9314,N_9136,N_9055);
nand U9315 (N_9315,N_9173,N_9037);
nand U9316 (N_9316,N_9195,N_9028);
or U9317 (N_9317,N_9036,N_9061);
xor U9318 (N_9318,N_9162,N_9154);
xor U9319 (N_9319,N_9020,N_9097);
and U9320 (N_9320,N_9137,N_9198);
and U9321 (N_9321,N_9145,N_9016);
or U9322 (N_9322,N_9039,N_9190);
xnor U9323 (N_9323,N_9012,N_9122);
xor U9324 (N_9324,N_9058,N_9192);
and U9325 (N_9325,N_9002,N_9164);
nand U9326 (N_9326,N_9144,N_9027);
or U9327 (N_9327,N_9188,N_9127);
nor U9328 (N_9328,N_9006,N_9163);
xor U9329 (N_9329,N_9059,N_9041);
or U9330 (N_9330,N_9027,N_9109);
nor U9331 (N_9331,N_9121,N_9114);
and U9332 (N_9332,N_9007,N_9030);
xor U9333 (N_9333,N_9096,N_9120);
nand U9334 (N_9334,N_9002,N_9086);
xnor U9335 (N_9335,N_9197,N_9121);
xor U9336 (N_9336,N_9060,N_9131);
and U9337 (N_9337,N_9156,N_9025);
xor U9338 (N_9338,N_9030,N_9004);
nor U9339 (N_9339,N_9054,N_9178);
nor U9340 (N_9340,N_9156,N_9029);
nand U9341 (N_9341,N_9107,N_9008);
nor U9342 (N_9342,N_9186,N_9130);
nand U9343 (N_9343,N_9056,N_9176);
xnor U9344 (N_9344,N_9003,N_9186);
nor U9345 (N_9345,N_9023,N_9166);
xnor U9346 (N_9346,N_9121,N_9030);
and U9347 (N_9347,N_9038,N_9098);
xor U9348 (N_9348,N_9195,N_9135);
and U9349 (N_9349,N_9002,N_9134);
nand U9350 (N_9350,N_9050,N_9106);
and U9351 (N_9351,N_9161,N_9025);
nand U9352 (N_9352,N_9095,N_9128);
and U9353 (N_9353,N_9054,N_9160);
or U9354 (N_9354,N_9161,N_9089);
nor U9355 (N_9355,N_9081,N_9175);
xor U9356 (N_9356,N_9110,N_9120);
xor U9357 (N_9357,N_9176,N_9066);
xnor U9358 (N_9358,N_9020,N_9105);
nand U9359 (N_9359,N_9042,N_9158);
xor U9360 (N_9360,N_9197,N_9182);
xor U9361 (N_9361,N_9040,N_9187);
or U9362 (N_9362,N_9018,N_9041);
or U9363 (N_9363,N_9078,N_9053);
xor U9364 (N_9364,N_9090,N_9192);
xor U9365 (N_9365,N_9031,N_9068);
nand U9366 (N_9366,N_9113,N_9154);
xor U9367 (N_9367,N_9141,N_9134);
nand U9368 (N_9368,N_9071,N_9154);
and U9369 (N_9369,N_9105,N_9072);
nor U9370 (N_9370,N_9155,N_9121);
or U9371 (N_9371,N_9007,N_9075);
nand U9372 (N_9372,N_9070,N_9112);
nor U9373 (N_9373,N_9066,N_9057);
xnor U9374 (N_9374,N_9032,N_9033);
and U9375 (N_9375,N_9094,N_9102);
nand U9376 (N_9376,N_9151,N_9034);
xnor U9377 (N_9377,N_9131,N_9078);
or U9378 (N_9378,N_9068,N_9162);
and U9379 (N_9379,N_9093,N_9011);
nand U9380 (N_9380,N_9098,N_9179);
nor U9381 (N_9381,N_9124,N_9097);
xor U9382 (N_9382,N_9167,N_9116);
or U9383 (N_9383,N_9113,N_9158);
or U9384 (N_9384,N_9063,N_9153);
xor U9385 (N_9385,N_9150,N_9159);
nand U9386 (N_9386,N_9098,N_9197);
and U9387 (N_9387,N_9008,N_9051);
nor U9388 (N_9388,N_9172,N_9039);
and U9389 (N_9389,N_9067,N_9192);
or U9390 (N_9390,N_9158,N_9011);
or U9391 (N_9391,N_9159,N_9167);
nor U9392 (N_9392,N_9157,N_9161);
and U9393 (N_9393,N_9032,N_9098);
xor U9394 (N_9394,N_9156,N_9160);
xor U9395 (N_9395,N_9016,N_9097);
or U9396 (N_9396,N_9101,N_9115);
nor U9397 (N_9397,N_9167,N_9031);
xnor U9398 (N_9398,N_9198,N_9079);
or U9399 (N_9399,N_9104,N_9186);
or U9400 (N_9400,N_9285,N_9373);
nand U9401 (N_9401,N_9335,N_9225);
or U9402 (N_9402,N_9256,N_9207);
xor U9403 (N_9403,N_9346,N_9269);
and U9404 (N_9404,N_9265,N_9280);
and U9405 (N_9405,N_9267,N_9314);
nor U9406 (N_9406,N_9291,N_9200);
or U9407 (N_9407,N_9251,N_9388);
nand U9408 (N_9408,N_9220,N_9208);
or U9409 (N_9409,N_9254,N_9253);
nor U9410 (N_9410,N_9232,N_9309);
or U9411 (N_9411,N_9336,N_9294);
or U9412 (N_9412,N_9320,N_9264);
xnor U9413 (N_9413,N_9355,N_9352);
and U9414 (N_9414,N_9237,N_9293);
or U9415 (N_9415,N_9261,N_9268);
nor U9416 (N_9416,N_9382,N_9387);
nand U9417 (N_9417,N_9215,N_9378);
or U9418 (N_9418,N_9363,N_9283);
and U9419 (N_9419,N_9235,N_9218);
and U9420 (N_9420,N_9216,N_9273);
or U9421 (N_9421,N_9376,N_9340);
or U9422 (N_9422,N_9255,N_9386);
and U9423 (N_9423,N_9205,N_9379);
xnor U9424 (N_9424,N_9206,N_9296);
nand U9425 (N_9425,N_9368,N_9371);
nand U9426 (N_9426,N_9375,N_9324);
and U9427 (N_9427,N_9372,N_9203);
xnor U9428 (N_9428,N_9311,N_9334);
and U9429 (N_9429,N_9213,N_9303);
and U9430 (N_9430,N_9211,N_9305);
and U9431 (N_9431,N_9377,N_9343);
and U9432 (N_9432,N_9222,N_9279);
nand U9433 (N_9433,N_9330,N_9250);
or U9434 (N_9434,N_9361,N_9332);
nor U9435 (N_9435,N_9395,N_9300);
xnor U9436 (N_9436,N_9366,N_9327);
nor U9437 (N_9437,N_9323,N_9317);
and U9438 (N_9438,N_9307,N_9274);
and U9439 (N_9439,N_9230,N_9337);
xor U9440 (N_9440,N_9374,N_9289);
nand U9441 (N_9441,N_9282,N_9201);
xnor U9442 (N_9442,N_9292,N_9262);
and U9443 (N_9443,N_9369,N_9301);
and U9444 (N_9444,N_9266,N_9329);
xnor U9445 (N_9445,N_9272,N_9241);
nand U9446 (N_9446,N_9242,N_9257);
and U9447 (N_9447,N_9316,N_9302);
and U9448 (N_9448,N_9246,N_9362);
xor U9449 (N_9449,N_9227,N_9217);
xnor U9450 (N_9450,N_9306,N_9381);
or U9451 (N_9451,N_9202,N_9350);
nor U9452 (N_9452,N_9319,N_9214);
nor U9453 (N_9453,N_9312,N_9259);
nor U9454 (N_9454,N_9252,N_9299);
nand U9455 (N_9455,N_9276,N_9263);
xor U9456 (N_9456,N_9318,N_9397);
xor U9457 (N_9457,N_9236,N_9271);
or U9458 (N_9458,N_9351,N_9353);
or U9459 (N_9459,N_9228,N_9275);
or U9460 (N_9460,N_9231,N_9290);
and U9461 (N_9461,N_9287,N_9224);
nand U9462 (N_9462,N_9380,N_9365);
and U9463 (N_9463,N_9249,N_9219);
nor U9464 (N_9464,N_9244,N_9308);
or U9465 (N_9465,N_9229,N_9357);
nor U9466 (N_9466,N_9295,N_9243);
nand U9467 (N_9467,N_9248,N_9389);
nand U9468 (N_9468,N_9358,N_9245);
and U9469 (N_9469,N_9325,N_9281);
nor U9470 (N_9470,N_9394,N_9284);
xnor U9471 (N_9471,N_9321,N_9328);
or U9472 (N_9472,N_9278,N_9247);
or U9473 (N_9473,N_9383,N_9399);
or U9474 (N_9474,N_9349,N_9298);
nor U9475 (N_9475,N_9364,N_9367);
nand U9476 (N_9476,N_9370,N_9304);
or U9477 (N_9477,N_9209,N_9348);
nor U9478 (N_9478,N_9391,N_9359);
or U9479 (N_9479,N_9338,N_9210);
xnor U9480 (N_9480,N_9322,N_9221);
nor U9481 (N_9481,N_9260,N_9270);
and U9482 (N_9482,N_9342,N_9233);
nor U9483 (N_9483,N_9258,N_9288);
nand U9484 (N_9484,N_9277,N_9212);
and U9485 (N_9485,N_9313,N_9297);
xor U9486 (N_9486,N_9344,N_9360);
and U9487 (N_9487,N_9234,N_9396);
nor U9488 (N_9488,N_9204,N_9341);
xnor U9489 (N_9489,N_9239,N_9333);
nand U9490 (N_9490,N_9326,N_9240);
xor U9491 (N_9491,N_9226,N_9398);
nand U9492 (N_9492,N_9354,N_9331);
nand U9493 (N_9493,N_9339,N_9223);
xnor U9494 (N_9494,N_9384,N_9286);
or U9495 (N_9495,N_9238,N_9356);
xor U9496 (N_9496,N_9385,N_9315);
nand U9497 (N_9497,N_9310,N_9345);
and U9498 (N_9498,N_9390,N_9393);
nor U9499 (N_9499,N_9347,N_9392);
and U9500 (N_9500,N_9264,N_9235);
nor U9501 (N_9501,N_9320,N_9372);
nand U9502 (N_9502,N_9325,N_9250);
nor U9503 (N_9503,N_9260,N_9207);
or U9504 (N_9504,N_9394,N_9249);
nor U9505 (N_9505,N_9308,N_9360);
nor U9506 (N_9506,N_9324,N_9217);
nor U9507 (N_9507,N_9317,N_9377);
nand U9508 (N_9508,N_9315,N_9209);
xnor U9509 (N_9509,N_9295,N_9244);
or U9510 (N_9510,N_9391,N_9207);
nand U9511 (N_9511,N_9370,N_9306);
or U9512 (N_9512,N_9298,N_9364);
and U9513 (N_9513,N_9371,N_9290);
and U9514 (N_9514,N_9222,N_9269);
xor U9515 (N_9515,N_9221,N_9262);
nand U9516 (N_9516,N_9302,N_9285);
xnor U9517 (N_9517,N_9331,N_9270);
nand U9518 (N_9518,N_9320,N_9395);
or U9519 (N_9519,N_9217,N_9355);
nand U9520 (N_9520,N_9379,N_9323);
and U9521 (N_9521,N_9330,N_9298);
or U9522 (N_9522,N_9343,N_9385);
nor U9523 (N_9523,N_9387,N_9257);
or U9524 (N_9524,N_9204,N_9237);
nand U9525 (N_9525,N_9362,N_9351);
or U9526 (N_9526,N_9366,N_9251);
or U9527 (N_9527,N_9340,N_9294);
xnor U9528 (N_9528,N_9260,N_9370);
nand U9529 (N_9529,N_9291,N_9394);
nor U9530 (N_9530,N_9350,N_9368);
or U9531 (N_9531,N_9302,N_9260);
nand U9532 (N_9532,N_9332,N_9222);
and U9533 (N_9533,N_9304,N_9254);
nor U9534 (N_9534,N_9390,N_9335);
nand U9535 (N_9535,N_9223,N_9267);
and U9536 (N_9536,N_9351,N_9229);
nand U9537 (N_9537,N_9256,N_9232);
xor U9538 (N_9538,N_9303,N_9350);
xnor U9539 (N_9539,N_9290,N_9237);
xnor U9540 (N_9540,N_9220,N_9324);
nand U9541 (N_9541,N_9223,N_9329);
nand U9542 (N_9542,N_9225,N_9298);
and U9543 (N_9543,N_9213,N_9297);
nand U9544 (N_9544,N_9221,N_9305);
xnor U9545 (N_9545,N_9344,N_9374);
and U9546 (N_9546,N_9328,N_9226);
nor U9547 (N_9547,N_9208,N_9375);
and U9548 (N_9548,N_9277,N_9347);
nor U9549 (N_9549,N_9395,N_9240);
nand U9550 (N_9550,N_9341,N_9346);
nor U9551 (N_9551,N_9397,N_9377);
xnor U9552 (N_9552,N_9218,N_9356);
or U9553 (N_9553,N_9352,N_9378);
nor U9554 (N_9554,N_9248,N_9215);
and U9555 (N_9555,N_9230,N_9362);
or U9556 (N_9556,N_9259,N_9214);
nand U9557 (N_9557,N_9399,N_9201);
nand U9558 (N_9558,N_9233,N_9232);
and U9559 (N_9559,N_9260,N_9327);
nand U9560 (N_9560,N_9307,N_9326);
nor U9561 (N_9561,N_9329,N_9365);
nand U9562 (N_9562,N_9350,N_9292);
nor U9563 (N_9563,N_9262,N_9350);
xor U9564 (N_9564,N_9236,N_9299);
and U9565 (N_9565,N_9246,N_9347);
or U9566 (N_9566,N_9226,N_9220);
nand U9567 (N_9567,N_9215,N_9263);
nor U9568 (N_9568,N_9203,N_9209);
xor U9569 (N_9569,N_9345,N_9237);
xnor U9570 (N_9570,N_9282,N_9216);
or U9571 (N_9571,N_9324,N_9382);
and U9572 (N_9572,N_9380,N_9242);
nand U9573 (N_9573,N_9207,N_9303);
or U9574 (N_9574,N_9284,N_9249);
nand U9575 (N_9575,N_9388,N_9213);
or U9576 (N_9576,N_9244,N_9282);
nor U9577 (N_9577,N_9293,N_9294);
nor U9578 (N_9578,N_9284,N_9288);
or U9579 (N_9579,N_9232,N_9252);
and U9580 (N_9580,N_9292,N_9264);
nand U9581 (N_9581,N_9204,N_9366);
and U9582 (N_9582,N_9206,N_9225);
nor U9583 (N_9583,N_9334,N_9350);
or U9584 (N_9584,N_9377,N_9258);
or U9585 (N_9585,N_9364,N_9252);
xor U9586 (N_9586,N_9215,N_9318);
nor U9587 (N_9587,N_9280,N_9206);
xor U9588 (N_9588,N_9306,N_9392);
or U9589 (N_9589,N_9267,N_9323);
or U9590 (N_9590,N_9345,N_9388);
nand U9591 (N_9591,N_9259,N_9325);
and U9592 (N_9592,N_9342,N_9323);
nor U9593 (N_9593,N_9215,N_9254);
xnor U9594 (N_9594,N_9356,N_9273);
nand U9595 (N_9595,N_9287,N_9382);
nand U9596 (N_9596,N_9387,N_9233);
nor U9597 (N_9597,N_9264,N_9380);
xnor U9598 (N_9598,N_9293,N_9249);
or U9599 (N_9599,N_9213,N_9394);
xor U9600 (N_9600,N_9444,N_9421);
xnor U9601 (N_9601,N_9595,N_9540);
nor U9602 (N_9602,N_9585,N_9452);
or U9603 (N_9603,N_9410,N_9538);
xor U9604 (N_9604,N_9493,N_9434);
or U9605 (N_9605,N_9520,N_9537);
nor U9606 (N_9606,N_9532,N_9415);
and U9607 (N_9607,N_9462,N_9599);
nor U9608 (N_9608,N_9594,N_9589);
or U9609 (N_9609,N_9424,N_9571);
xor U9610 (N_9610,N_9572,N_9474);
or U9611 (N_9611,N_9411,N_9484);
or U9612 (N_9612,N_9560,N_9563);
and U9613 (N_9613,N_9522,N_9443);
and U9614 (N_9614,N_9466,N_9527);
or U9615 (N_9615,N_9500,N_9497);
and U9616 (N_9616,N_9551,N_9561);
nand U9617 (N_9617,N_9596,N_9549);
xnor U9618 (N_9618,N_9582,N_9584);
or U9619 (N_9619,N_9554,N_9543);
nor U9620 (N_9620,N_9591,N_9420);
or U9621 (N_9621,N_9499,N_9529);
xnor U9622 (N_9622,N_9573,N_9469);
nand U9623 (N_9623,N_9491,N_9478);
nand U9624 (N_9624,N_9578,N_9505);
or U9625 (N_9625,N_9577,N_9400);
xnor U9626 (N_9626,N_9464,N_9545);
nand U9627 (N_9627,N_9473,N_9442);
nor U9628 (N_9628,N_9558,N_9559);
nand U9629 (N_9629,N_9453,N_9472);
nor U9630 (N_9630,N_9502,N_9450);
xor U9631 (N_9631,N_9583,N_9459);
xnor U9632 (N_9632,N_9509,N_9440);
and U9633 (N_9633,N_9508,N_9542);
xor U9634 (N_9634,N_9438,N_9516);
xnor U9635 (N_9635,N_9448,N_9486);
nand U9636 (N_9636,N_9564,N_9492);
nand U9637 (N_9637,N_9514,N_9477);
or U9638 (N_9638,N_9433,N_9455);
or U9639 (N_9639,N_9557,N_9562);
nand U9640 (N_9640,N_9405,N_9428);
nor U9641 (N_9641,N_9510,N_9429);
or U9642 (N_9642,N_9457,N_9533);
xnor U9643 (N_9643,N_9460,N_9446);
nand U9644 (N_9644,N_9586,N_9550);
xor U9645 (N_9645,N_9476,N_9461);
nand U9646 (N_9646,N_9467,N_9521);
and U9647 (N_9647,N_9528,N_9547);
or U9648 (N_9648,N_9437,N_9430);
xor U9649 (N_9649,N_9471,N_9436);
and U9650 (N_9650,N_9414,N_9506);
nand U9651 (N_9651,N_9413,N_9402);
or U9652 (N_9652,N_9470,N_9489);
and U9653 (N_9653,N_9555,N_9458);
nand U9654 (N_9654,N_9512,N_9552);
xor U9655 (N_9655,N_9412,N_9518);
and U9656 (N_9656,N_9556,N_9495);
nor U9657 (N_9657,N_9567,N_9581);
and U9658 (N_9658,N_9449,N_9511);
xnor U9659 (N_9659,N_9468,N_9524);
nor U9660 (N_9660,N_9485,N_9546);
xnor U9661 (N_9661,N_9530,N_9513);
or U9662 (N_9662,N_9479,N_9481);
xnor U9663 (N_9663,N_9487,N_9423);
or U9664 (N_9664,N_9465,N_9566);
nand U9665 (N_9665,N_9544,N_9575);
nand U9666 (N_9666,N_9419,N_9406);
and U9667 (N_9667,N_9503,N_9531);
and U9668 (N_9668,N_9570,N_9409);
xnor U9669 (N_9669,N_9569,N_9403);
and U9670 (N_9670,N_9574,N_9507);
and U9671 (N_9671,N_9579,N_9590);
and U9672 (N_9672,N_9535,N_9408);
xnor U9673 (N_9673,N_9536,N_9587);
nand U9674 (N_9674,N_9425,N_9498);
and U9675 (N_9675,N_9501,N_9565);
or U9676 (N_9676,N_9496,N_9475);
nand U9677 (N_9677,N_9580,N_9456);
nor U9678 (N_9678,N_9488,N_9525);
and U9679 (N_9679,N_9598,N_9463);
xor U9680 (N_9680,N_9431,N_9490);
or U9681 (N_9681,N_9407,N_9548);
nor U9682 (N_9682,N_9480,N_9427);
and U9683 (N_9683,N_9597,N_9534);
and U9684 (N_9684,N_9426,N_9482);
or U9685 (N_9685,N_9401,N_9515);
nor U9686 (N_9686,N_9494,N_9441);
xnor U9687 (N_9687,N_9553,N_9588);
nor U9688 (N_9688,N_9593,N_9422);
and U9689 (N_9689,N_9447,N_9517);
or U9690 (N_9690,N_9435,N_9445);
and U9691 (N_9691,N_9418,N_9451);
or U9692 (N_9692,N_9483,N_9404);
or U9693 (N_9693,N_9439,N_9432);
nor U9694 (N_9694,N_9504,N_9523);
xor U9695 (N_9695,N_9454,N_9519);
nor U9696 (N_9696,N_9526,N_9592);
nand U9697 (N_9697,N_9576,N_9539);
nor U9698 (N_9698,N_9541,N_9568);
or U9699 (N_9699,N_9416,N_9417);
or U9700 (N_9700,N_9549,N_9529);
xor U9701 (N_9701,N_9437,N_9484);
xor U9702 (N_9702,N_9435,N_9412);
xor U9703 (N_9703,N_9417,N_9536);
or U9704 (N_9704,N_9461,N_9538);
nor U9705 (N_9705,N_9565,N_9410);
xnor U9706 (N_9706,N_9415,N_9438);
nand U9707 (N_9707,N_9526,N_9560);
xor U9708 (N_9708,N_9426,N_9528);
nand U9709 (N_9709,N_9536,N_9444);
and U9710 (N_9710,N_9511,N_9530);
and U9711 (N_9711,N_9469,N_9430);
and U9712 (N_9712,N_9544,N_9483);
nand U9713 (N_9713,N_9480,N_9423);
nand U9714 (N_9714,N_9474,N_9588);
and U9715 (N_9715,N_9478,N_9404);
xnor U9716 (N_9716,N_9520,N_9579);
nand U9717 (N_9717,N_9414,N_9453);
or U9718 (N_9718,N_9415,N_9400);
nand U9719 (N_9719,N_9586,N_9540);
nor U9720 (N_9720,N_9463,N_9427);
nand U9721 (N_9721,N_9542,N_9454);
or U9722 (N_9722,N_9548,N_9546);
or U9723 (N_9723,N_9400,N_9463);
and U9724 (N_9724,N_9554,N_9552);
nand U9725 (N_9725,N_9415,N_9594);
or U9726 (N_9726,N_9467,N_9529);
or U9727 (N_9727,N_9410,N_9566);
or U9728 (N_9728,N_9430,N_9506);
nor U9729 (N_9729,N_9560,N_9515);
xor U9730 (N_9730,N_9400,N_9494);
xnor U9731 (N_9731,N_9450,N_9426);
xnor U9732 (N_9732,N_9514,N_9471);
nand U9733 (N_9733,N_9593,N_9408);
and U9734 (N_9734,N_9406,N_9529);
or U9735 (N_9735,N_9491,N_9494);
nand U9736 (N_9736,N_9540,N_9566);
or U9737 (N_9737,N_9527,N_9516);
and U9738 (N_9738,N_9596,N_9598);
or U9739 (N_9739,N_9438,N_9496);
xnor U9740 (N_9740,N_9473,N_9580);
and U9741 (N_9741,N_9419,N_9495);
or U9742 (N_9742,N_9405,N_9472);
or U9743 (N_9743,N_9584,N_9467);
or U9744 (N_9744,N_9492,N_9571);
xnor U9745 (N_9745,N_9404,N_9581);
and U9746 (N_9746,N_9456,N_9490);
nand U9747 (N_9747,N_9436,N_9473);
or U9748 (N_9748,N_9435,N_9599);
xnor U9749 (N_9749,N_9575,N_9430);
and U9750 (N_9750,N_9497,N_9505);
and U9751 (N_9751,N_9437,N_9525);
and U9752 (N_9752,N_9570,N_9411);
and U9753 (N_9753,N_9525,N_9400);
xor U9754 (N_9754,N_9527,N_9561);
nor U9755 (N_9755,N_9594,N_9559);
nor U9756 (N_9756,N_9547,N_9451);
and U9757 (N_9757,N_9545,N_9508);
xor U9758 (N_9758,N_9433,N_9578);
nand U9759 (N_9759,N_9456,N_9529);
xnor U9760 (N_9760,N_9596,N_9532);
xor U9761 (N_9761,N_9531,N_9437);
or U9762 (N_9762,N_9567,N_9414);
or U9763 (N_9763,N_9426,N_9431);
nor U9764 (N_9764,N_9593,N_9429);
or U9765 (N_9765,N_9541,N_9526);
nand U9766 (N_9766,N_9590,N_9589);
nor U9767 (N_9767,N_9429,N_9413);
nand U9768 (N_9768,N_9443,N_9551);
and U9769 (N_9769,N_9534,N_9560);
xor U9770 (N_9770,N_9545,N_9537);
or U9771 (N_9771,N_9566,N_9496);
nand U9772 (N_9772,N_9447,N_9436);
nor U9773 (N_9773,N_9454,N_9572);
xor U9774 (N_9774,N_9512,N_9567);
xor U9775 (N_9775,N_9452,N_9409);
or U9776 (N_9776,N_9463,N_9522);
and U9777 (N_9777,N_9536,N_9408);
xor U9778 (N_9778,N_9513,N_9408);
or U9779 (N_9779,N_9522,N_9406);
and U9780 (N_9780,N_9527,N_9441);
xnor U9781 (N_9781,N_9416,N_9558);
or U9782 (N_9782,N_9536,N_9413);
nor U9783 (N_9783,N_9424,N_9425);
xor U9784 (N_9784,N_9504,N_9422);
xor U9785 (N_9785,N_9460,N_9442);
nand U9786 (N_9786,N_9508,N_9433);
and U9787 (N_9787,N_9435,N_9456);
and U9788 (N_9788,N_9509,N_9489);
nor U9789 (N_9789,N_9472,N_9467);
nor U9790 (N_9790,N_9521,N_9485);
nand U9791 (N_9791,N_9512,N_9559);
nor U9792 (N_9792,N_9434,N_9595);
nand U9793 (N_9793,N_9563,N_9575);
nand U9794 (N_9794,N_9523,N_9562);
or U9795 (N_9795,N_9526,N_9480);
nand U9796 (N_9796,N_9403,N_9591);
xor U9797 (N_9797,N_9512,N_9451);
or U9798 (N_9798,N_9441,N_9510);
nand U9799 (N_9799,N_9401,N_9444);
or U9800 (N_9800,N_9697,N_9681);
or U9801 (N_9801,N_9738,N_9602);
nand U9802 (N_9802,N_9643,N_9795);
nor U9803 (N_9803,N_9688,N_9601);
and U9804 (N_9804,N_9605,N_9661);
and U9805 (N_9805,N_9788,N_9674);
and U9806 (N_9806,N_9737,N_9623);
xnor U9807 (N_9807,N_9687,N_9778);
xnor U9808 (N_9808,N_9609,N_9761);
nand U9809 (N_9809,N_9678,N_9696);
and U9810 (N_9810,N_9743,N_9786);
nand U9811 (N_9811,N_9727,N_9797);
xor U9812 (N_9812,N_9620,N_9693);
nor U9813 (N_9813,N_9704,N_9637);
or U9814 (N_9814,N_9732,N_9621);
xor U9815 (N_9815,N_9691,N_9703);
or U9816 (N_9816,N_9783,N_9610);
nor U9817 (N_9817,N_9717,N_9714);
or U9818 (N_9818,N_9769,N_9614);
nand U9819 (N_9819,N_9731,N_9771);
and U9820 (N_9820,N_9646,N_9702);
nand U9821 (N_9821,N_9709,N_9730);
nor U9822 (N_9822,N_9745,N_9612);
nand U9823 (N_9823,N_9728,N_9622);
nand U9824 (N_9824,N_9753,N_9790);
and U9825 (N_9825,N_9652,N_9660);
xor U9826 (N_9826,N_9784,N_9644);
nor U9827 (N_9827,N_9711,N_9664);
nor U9828 (N_9828,N_9757,N_9780);
nor U9829 (N_9829,N_9650,N_9774);
xnor U9830 (N_9830,N_9735,N_9680);
xor U9831 (N_9831,N_9626,N_9789);
nand U9832 (N_9832,N_9754,N_9690);
xnor U9833 (N_9833,N_9669,N_9642);
or U9834 (N_9834,N_9663,N_9751);
or U9835 (N_9835,N_9740,N_9755);
nand U9836 (N_9836,N_9679,N_9676);
nand U9837 (N_9837,N_9758,N_9766);
and U9838 (N_9838,N_9686,N_9793);
nand U9839 (N_9839,N_9775,N_9734);
nor U9840 (N_9840,N_9628,N_9630);
xnor U9841 (N_9841,N_9746,N_9645);
nand U9842 (N_9842,N_9787,N_9773);
nand U9843 (N_9843,N_9694,N_9712);
nor U9844 (N_9844,N_9635,N_9724);
and U9845 (N_9845,N_9750,N_9736);
xor U9846 (N_9846,N_9762,N_9729);
and U9847 (N_9847,N_9744,N_9776);
xnor U9848 (N_9848,N_9782,N_9716);
or U9849 (N_9849,N_9673,N_9632);
or U9850 (N_9850,N_9682,N_9792);
or U9851 (N_9851,N_9647,N_9685);
or U9852 (N_9852,N_9600,N_9653);
xor U9853 (N_9853,N_9699,N_9684);
or U9854 (N_9854,N_9659,N_9760);
nand U9855 (N_9855,N_9617,N_9768);
nand U9856 (N_9856,N_9700,N_9733);
or U9857 (N_9857,N_9627,N_9631);
nor U9858 (N_9858,N_9655,N_9747);
and U9859 (N_9859,N_9634,N_9668);
nand U9860 (N_9860,N_9794,N_9779);
and U9861 (N_9861,N_9765,N_9624);
xor U9862 (N_9862,N_9657,N_9796);
and U9863 (N_9863,N_9723,N_9648);
nor U9864 (N_9864,N_9639,N_9695);
xor U9865 (N_9865,N_9615,N_9756);
nand U9866 (N_9866,N_9633,N_9689);
xnor U9867 (N_9867,N_9798,N_9662);
xor U9868 (N_9868,N_9748,N_9777);
and U9869 (N_9869,N_9741,N_9772);
or U9870 (N_9870,N_9708,N_9677);
xor U9871 (N_9871,N_9770,N_9715);
and U9872 (N_9872,N_9619,N_9705);
xor U9873 (N_9873,N_9701,N_9706);
and U9874 (N_9874,N_9742,N_9656);
and U9875 (N_9875,N_9618,N_9613);
nand U9876 (N_9876,N_9667,N_9654);
or U9877 (N_9877,N_9785,N_9608);
and U9878 (N_9878,N_9799,N_9791);
nand U9879 (N_9879,N_9651,N_9604);
and U9880 (N_9880,N_9752,N_9665);
nand U9881 (N_9881,N_9641,N_9616);
and U9882 (N_9882,N_9739,N_9636);
nor U9883 (N_9883,N_9607,N_9720);
nor U9884 (N_9884,N_9658,N_9719);
and U9885 (N_9885,N_9670,N_9764);
or U9886 (N_9886,N_9625,N_9722);
xnor U9887 (N_9887,N_9759,N_9675);
and U9888 (N_9888,N_9606,N_9726);
nand U9889 (N_9889,N_9713,N_9603);
nand U9890 (N_9890,N_9629,N_9725);
xnor U9891 (N_9891,N_9672,N_9749);
or U9892 (N_9892,N_9692,N_9721);
and U9893 (N_9893,N_9649,N_9781);
and U9894 (N_9894,N_9638,N_9683);
xor U9895 (N_9895,N_9698,N_9640);
and U9896 (N_9896,N_9671,N_9767);
nor U9897 (N_9897,N_9611,N_9763);
and U9898 (N_9898,N_9710,N_9707);
and U9899 (N_9899,N_9718,N_9666);
xor U9900 (N_9900,N_9652,N_9736);
nand U9901 (N_9901,N_9711,N_9773);
xor U9902 (N_9902,N_9799,N_9654);
nand U9903 (N_9903,N_9769,N_9615);
or U9904 (N_9904,N_9664,N_9744);
nand U9905 (N_9905,N_9648,N_9710);
nand U9906 (N_9906,N_9601,N_9721);
or U9907 (N_9907,N_9632,N_9762);
nand U9908 (N_9908,N_9602,N_9684);
or U9909 (N_9909,N_9646,N_9666);
or U9910 (N_9910,N_9621,N_9601);
nand U9911 (N_9911,N_9794,N_9672);
nand U9912 (N_9912,N_9687,N_9707);
or U9913 (N_9913,N_9789,N_9708);
or U9914 (N_9914,N_9723,N_9724);
or U9915 (N_9915,N_9696,N_9660);
or U9916 (N_9916,N_9731,N_9655);
nor U9917 (N_9917,N_9700,N_9673);
nand U9918 (N_9918,N_9616,N_9648);
nand U9919 (N_9919,N_9647,N_9763);
nor U9920 (N_9920,N_9785,N_9708);
or U9921 (N_9921,N_9762,N_9750);
and U9922 (N_9922,N_9643,N_9683);
and U9923 (N_9923,N_9754,N_9606);
nor U9924 (N_9924,N_9753,N_9747);
and U9925 (N_9925,N_9612,N_9781);
xnor U9926 (N_9926,N_9661,N_9651);
nor U9927 (N_9927,N_9644,N_9752);
nor U9928 (N_9928,N_9626,N_9618);
nand U9929 (N_9929,N_9745,N_9704);
and U9930 (N_9930,N_9613,N_9652);
and U9931 (N_9931,N_9668,N_9728);
nor U9932 (N_9932,N_9695,N_9676);
and U9933 (N_9933,N_9757,N_9631);
nor U9934 (N_9934,N_9619,N_9780);
nand U9935 (N_9935,N_9733,N_9695);
xor U9936 (N_9936,N_9630,N_9633);
nor U9937 (N_9937,N_9729,N_9704);
nor U9938 (N_9938,N_9710,N_9638);
and U9939 (N_9939,N_9792,N_9735);
xor U9940 (N_9940,N_9652,N_9615);
nor U9941 (N_9941,N_9790,N_9780);
or U9942 (N_9942,N_9629,N_9641);
or U9943 (N_9943,N_9789,N_9624);
and U9944 (N_9944,N_9770,N_9681);
or U9945 (N_9945,N_9637,N_9674);
xnor U9946 (N_9946,N_9707,N_9745);
xnor U9947 (N_9947,N_9674,N_9638);
nor U9948 (N_9948,N_9679,N_9696);
xor U9949 (N_9949,N_9732,N_9771);
nand U9950 (N_9950,N_9662,N_9633);
xor U9951 (N_9951,N_9663,N_9606);
or U9952 (N_9952,N_9765,N_9617);
and U9953 (N_9953,N_9663,N_9783);
or U9954 (N_9954,N_9746,N_9749);
xor U9955 (N_9955,N_9628,N_9645);
or U9956 (N_9956,N_9601,N_9794);
nor U9957 (N_9957,N_9791,N_9647);
nand U9958 (N_9958,N_9786,N_9754);
or U9959 (N_9959,N_9701,N_9697);
nor U9960 (N_9960,N_9725,N_9633);
and U9961 (N_9961,N_9749,N_9724);
and U9962 (N_9962,N_9787,N_9713);
and U9963 (N_9963,N_9698,N_9731);
or U9964 (N_9964,N_9793,N_9663);
or U9965 (N_9965,N_9673,N_9721);
nand U9966 (N_9966,N_9665,N_9622);
or U9967 (N_9967,N_9693,N_9643);
nand U9968 (N_9968,N_9766,N_9781);
nor U9969 (N_9969,N_9709,N_9688);
nand U9970 (N_9970,N_9780,N_9705);
nor U9971 (N_9971,N_9779,N_9741);
xnor U9972 (N_9972,N_9776,N_9771);
nor U9973 (N_9973,N_9715,N_9609);
or U9974 (N_9974,N_9645,N_9658);
nand U9975 (N_9975,N_9702,N_9748);
and U9976 (N_9976,N_9644,N_9712);
nor U9977 (N_9977,N_9783,N_9698);
xnor U9978 (N_9978,N_9744,N_9746);
xnor U9979 (N_9979,N_9760,N_9651);
nand U9980 (N_9980,N_9728,N_9718);
xnor U9981 (N_9981,N_9738,N_9789);
nor U9982 (N_9982,N_9671,N_9774);
xnor U9983 (N_9983,N_9650,N_9676);
and U9984 (N_9984,N_9746,N_9652);
nor U9985 (N_9985,N_9671,N_9778);
nor U9986 (N_9986,N_9705,N_9712);
xor U9987 (N_9987,N_9780,N_9674);
nor U9988 (N_9988,N_9684,N_9697);
nor U9989 (N_9989,N_9640,N_9733);
nand U9990 (N_9990,N_9737,N_9741);
xor U9991 (N_9991,N_9784,N_9652);
xnor U9992 (N_9992,N_9739,N_9698);
nor U9993 (N_9993,N_9670,N_9615);
nor U9994 (N_9994,N_9692,N_9753);
nor U9995 (N_9995,N_9793,N_9764);
xnor U9996 (N_9996,N_9626,N_9770);
and U9997 (N_9997,N_9685,N_9755);
nor U9998 (N_9998,N_9609,N_9744);
nor U9999 (N_9999,N_9649,N_9638);
xnor U10000 (N_10000,N_9980,N_9955);
nor U10001 (N_10001,N_9828,N_9863);
nor U10002 (N_10002,N_9855,N_9897);
nor U10003 (N_10003,N_9882,N_9886);
and U10004 (N_10004,N_9989,N_9909);
xor U10005 (N_10005,N_9858,N_9829);
nor U10006 (N_10006,N_9842,N_9912);
and U10007 (N_10007,N_9803,N_9987);
and U10008 (N_10008,N_9946,N_9936);
nand U10009 (N_10009,N_9973,N_9969);
nor U10010 (N_10010,N_9937,N_9919);
nand U10011 (N_10011,N_9885,N_9899);
or U10012 (N_10012,N_9983,N_9970);
nand U10013 (N_10013,N_9875,N_9822);
or U10014 (N_10014,N_9949,N_9952);
nor U10015 (N_10015,N_9836,N_9893);
nor U10016 (N_10016,N_9956,N_9824);
or U10017 (N_10017,N_9877,N_9881);
and U10018 (N_10018,N_9979,N_9941);
nor U10019 (N_10019,N_9923,N_9975);
nor U10020 (N_10020,N_9994,N_9808);
nand U10021 (N_10021,N_9837,N_9958);
and U10022 (N_10022,N_9910,N_9845);
nand U10023 (N_10023,N_9966,N_9962);
or U10024 (N_10024,N_9904,N_9894);
and U10025 (N_10025,N_9876,N_9898);
nor U10026 (N_10026,N_9818,N_9986);
nand U10027 (N_10027,N_9996,N_9874);
or U10028 (N_10028,N_9891,N_9879);
xnor U10029 (N_10029,N_9963,N_9888);
or U10030 (N_10030,N_9957,N_9843);
or U10031 (N_10031,N_9947,N_9853);
or U10032 (N_10032,N_9985,N_9981);
nand U10033 (N_10033,N_9943,N_9911);
xor U10034 (N_10034,N_9872,N_9817);
nor U10035 (N_10035,N_9951,N_9964);
and U10036 (N_10036,N_9913,N_9988);
nand U10037 (N_10037,N_9926,N_9925);
and U10038 (N_10038,N_9868,N_9826);
nor U10039 (N_10039,N_9895,N_9800);
or U10040 (N_10040,N_9892,N_9961);
or U10041 (N_10041,N_9922,N_9960);
xor U10042 (N_10042,N_9862,N_9838);
xor U10043 (N_10043,N_9977,N_9915);
nand U10044 (N_10044,N_9993,N_9861);
nand U10045 (N_10045,N_9825,N_9802);
nand U10046 (N_10046,N_9851,N_9865);
and U10047 (N_10047,N_9814,N_9847);
nand U10048 (N_10048,N_9849,N_9850);
xor U10049 (N_10049,N_9990,N_9972);
or U10050 (N_10050,N_9827,N_9942);
xnor U10051 (N_10051,N_9860,N_9991);
nand U10052 (N_10052,N_9917,N_9992);
xor U10053 (N_10053,N_9965,N_9953);
nand U10054 (N_10054,N_9869,N_9916);
nand U10055 (N_10055,N_9920,N_9906);
xor U10056 (N_10056,N_9889,N_9831);
or U10057 (N_10057,N_9830,N_9998);
xnor U10058 (N_10058,N_9927,N_9834);
xnor U10059 (N_10059,N_9968,N_9978);
or U10060 (N_10060,N_9806,N_9867);
and U10061 (N_10061,N_9852,N_9866);
nand U10062 (N_10062,N_9908,N_9984);
or U10063 (N_10063,N_9940,N_9809);
nor U10064 (N_10064,N_9887,N_9832);
or U10065 (N_10065,N_9902,N_9854);
xor U10066 (N_10066,N_9921,N_9859);
and U10067 (N_10067,N_9846,N_9821);
or U10068 (N_10068,N_9907,N_9924);
nand U10069 (N_10069,N_9959,N_9878);
and U10070 (N_10070,N_9930,N_9950);
nor U10071 (N_10071,N_9835,N_9905);
and U10072 (N_10072,N_9804,N_9856);
or U10073 (N_10073,N_9807,N_9820);
xor U10074 (N_10074,N_9967,N_9857);
nand U10075 (N_10075,N_9801,N_9945);
nand U10076 (N_10076,N_9934,N_9840);
nor U10077 (N_10077,N_9971,N_9813);
xnor U10078 (N_10078,N_9812,N_9954);
and U10079 (N_10079,N_9914,N_9982);
nand U10080 (N_10080,N_9816,N_9864);
nor U10081 (N_10081,N_9805,N_9884);
xor U10082 (N_10082,N_9997,N_9810);
or U10083 (N_10083,N_9841,N_9839);
xor U10084 (N_10084,N_9890,N_9931);
nor U10085 (N_10085,N_9999,N_9918);
xor U10086 (N_10086,N_9901,N_9819);
and U10087 (N_10087,N_9933,N_9844);
nor U10088 (N_10088,N_9848,N_9976);
xnor U10089 (N_10089,N_9938,N_9944);
xor U10090 (N_10090,N_9823,N_9900);
nor U10091 (N_10091,N_9935,N_9896);
nand U10092 (N_10092,N_9815,N_9974);
or U10093 (N_10093,N_9811,N_9883);
or U10094 (N_10094,N_9932,N_9873);
and U10095 (N_10095,N_9928,N_9995);
nor U10096 (N_10096,N_9870,N_9929);
nand U10097 (N_10097,N_9948,N_9903);
and U10098 (N_10098,N_9871,N_9880);
or U10099 (N_10099,N_9833,N_9939);
nor U10100 (N_10100,N_9803,N_9897);
and U10101 (N_10101,N_9826,N_9907);
and U10102 (N_10102,N_9978,N_9979);
or U10103 (N_10103,N_9919,N_9828);
nand U10104 (N_10104,N_9846,N_9834);
nor U10105 (N_10105,N_9979,N_9852);
or U10106 (N_10106,N_9890,N_9995);
or U10107 (N_10107,N_9816,N_9821);
nand U10108 (N_10108,N_9896,N_9942);
or U10109 (N_10109,N_9965,N_9984);
xor U10110 (N_10110,N_9897,N_9887);
nand U10111 (N_10111,N_9932,N_9883);
nor U10112 (N_10112,N_9953,N_9998);
nand U10113 (N_10113,N_9881,N_9913);
nand U10114 (N_10114,N_9827,N_9944);
nor U10115 (N_10115,N_9884,N_9854);
and U10116 (N_10116,N_9821,N_9879);
or U10117 (N_10117,N_9999,N_9980);
or U10118 (N_10118,N_9888,N_9958);
nand U10119 (N_10119,N_9838,N_9850);
xor U10120 (N_10120,N_9900,N_9996);
and U10121 (N_10121,N_9801,N_9964);
xor U10122 (N_10122,N_9950,N_9871);
or U10123 (N_10123,N_9846,N_9939);
and U10124 (N_10124,N_9922,N_9901);
and U10125 (N_10125,N_9850,N_9992);
or U10126 (N_10126,N_9806,N_9830);
or U10127 (N_10127,N_9829,N_9827);
or U10128 (N_10128,N_9990,N_9914);
and U10129 (N_10129,N_9903,N_9960);
and U10130 (N_10130,N_9816,N_9804);
and U10131 (N_10131,N_9999,N_9859);
and U10132 (N_10132,N_9898,N_9930);
or U10133 (N_10133,N_9834,N_9848);
or U10134 (N_10134,N_9830,N_9800);
nor U10135 (N_10135,N_9931,N_9881);
and U10136 (N_10136,N_9855,N_9905);
xor U10137 (N_10137,N_9855,N_9808);
xnor U10138 (N_10138,N_9987,N_9826);
xor U10139 (N_10139,N_9943,N_9813);
and U10140 (N_10140,N_9987,N_9836);
nand U10141 (N_10141,N_9978,N_9918);
or U10142 (N_10142,N_9980,N_9936);
nor U10143 (N_10143,N_9867,N_9809);
nor U10144 (N_10144,N_9866,N_9826);
nand U10145 (N_10145,N_9888,N_9883);
nor U10146 (N_10146,N_9849,N_9942);
nor U10147 (N_10147,N_9853,N_9816);
or U10148 (N_10148,N_9964,N_9928);
nand U10149 (N_10149,N_9927,N_9803);
nor U10150 (N_10150,N_9939,N_9831);
nand U10151 (N_10151,N_9929,N_9953);
nor U10152 (N_10152,N_9992,N_9932);
or U10153 (N_10153,N_9986,N_9867);
xnor U10154 (N_10154,N_9868,N_9955);
and U10155 (N_10155,N_9806,N_9927);
nand U10156 (N_10156,N_9850,N_9828);
xnor U10157 (N_10157,N_9969,N_9863);
nand U10158 (N_10158,N_9868,N_9932);
xor U10159 (N_10159,N_9813,N_9898);
and U10160 (N_10160,N_9892,N_9948);
nand U10161 (N_10161,N_9899,N_9862);
and U10162 (N_10162,N_9979,N_9866);
or U10163 (N_10163,N_9866,N_9967);
nand U10164 (N_10164,N_9806,N_9819);
nor U10165 (N_10165,N_9840,N_9918);
xor U10166 (N_10166,N_9829,N_9814);
nor U10167 (N_10167,N_9900,N_9985);
xor U10168 (N_10168,N_9949,N_9941);
xnor U10169 (N_10169,N_9924,N_9887);
nand U10170 (N_10170,N_9971,N_9829);
or U10171 (N_10171,N_9834,N_9926);
xor U10172 (N_10172,N_9802,N_9943);
xor U10173 (N_10173,N_9953,N_9961);
and U10174 (N_10174,N_9860,N_9953);
nand U10175 (N_10175,N_9845,N_9870);
or U10176 (N_10176,N_9903,N_9983);
and U10177 (N_10177,N_9853,N_9875);
xnor U10178 (N_10178,N_9913,N_9933);
and U10179 (N_10179,N_9969,N_9836);
nand U10180 (N_10180,N_9807,N_9939);
nand U10181 (N_10181,N_9881,N_9906);
and U10182 (N_10182,N_9814,N_9990);
or U10183 (N_10183,N_9974,N_9867);
nor U10184 (N_10184,N_9813,N_9839);
nand U10185 (N_10185,N_9869,N_9932);
nand U10186 (N_10186,N_9941,N_9895);
xor U10187 (N_10187,N_9919,N_9953);
nand U10188 (N_10188,N_9926,N_9970);
or U10189 (N_10189,N_9941,N_9824);
and U10190 (N_10190,N_9835,N_9958);
nand U10191 (N_10191,N_9862,N_9918);
or U10192 (N_10192,N_9962,N_9900);
nor U10193 (N_10193,N_9978,N_9987);
and U10194 (N_10194,N_9975,N_9955);
nor U10195 (N_10195,N_9865,N_9843);
xor U10196 (N_10196,N_9920,N_9848);
and U10197 (N_10197,N_9813,N_9820);
nor U10198 (N_10198,N_9856,N_9833);
xor U10199 (N_10199,N_9940,N_9956);
nand U10200 (N_10200,N_10164,N_10032);
nand U10201 (N_10201,N_10117,N_10144);
or U10202 (N_10202,N_10149,N_10073);
or U10203 (N_10203,N_10155,N_10014);
xnor U10204 (N_10204,N_10006,N_10038);
xnor U10205 (N_10205,N_10180,N_10054);
xor U10206 (N_10206,N_10145,N_10085);
or U10207 (N_10207,N_10047,N_10178);
xnor U10208 (N_10208,N_10005,N_10094);
nand U10209 (N_10209,N_10165,N_10170);
nand U10210 (N_10210,N_10010,N_10099);
xnor U10211 (N_10211,N_10160,N_10098);
and U10212 (N_10212,N_10007,N_10041);
nor U10213 (N_10213,N_10028,N_10030);
and U10214 (N_10214,N_10056,N_10096);
or U10215 (N_10215,N_10091,N_10045);
nor U10216 (N_10216,N_10163,N_10008);
and U10217 (N_10217,N_10040,N_10179);
nor U10218 (N_10218,N_10115,N_10132);
xnor U10219 (N_10219,N_10123,N_10001);
xnor U10220 (N_10220,N_10183,N_10020);
nor U10221 (N_10221,N_10184,N_10078);
xnor U10222 (N_10222,N_10104,N_10093);
and U10223 (N_10223,N_10072,N_10173);
xnor U10224 (N_10224,N_10012,N_10147);
or U10225 (N_10225,N_10055,N_10036);
or U10226 (N_10226,N_10022,N_10166);
nand U10227 (N_10227,N_10171,N_10189);
and U10228 (N_10228,N_10168,N_10157);
and U10229 (N_10229,N_10074,N_10172);
xnor U10230 (N_10230,N_10049,N_10043);
nand U10231 (N_10231,N_10097,N_10197);
or U10232 (N_10232,N_10086,N_10159);
nand U10233 (N_10233,N_10194,N_10196);
nand U10234 (N_10234,N_10000,N_10103);
xnor U10235 (N_10235,N_10191,N_10017);
nand U10236 (N_10236,N_10199,N_10037);
and U10237 (N_10237,N_10065,N_10102);
and U10238 (N_10238,N_10119,N_10044);
nor U10239 (N_10239,N_10161,N_10081);
xor U10240 (N_10240,N_10108,N_10193);
and U10241 (N_10241,N_10127,N_10029);
nor U10242 (N_10242,N_10152,N_10080);
xor U10243 (N_10243,N_10198,N_10068);
nor U10244 (N_10244,N_10105,N_10134);
or U10245 (N_10245,N_10142,N_10111);
and U10246 (N_10246,N_10181,N_10060);
or U10247 (N_10247,N_10138,N_10195);
and U10248 (N_10248,N_10109,N_10087);
nor U10249 (N_10249,N_10024,N_10046);
nand U10250 (N_10250,N_10083,N_10063);
xnor U10251 (N_10251,N_10131,N_10069);
xnor U10252 (N_10252,N_10021,N_10016);
or U10253 (N_10253,N_10084,N_10025);
nand U10254 (N_10254,N_10059,N_10133);
nand U10255 (N_10255,N_10071,N_10141);
or U10256 (N_10256,N_10015,N_10034);
xor U10257 (N_10257,N_10092,N_10100);
xnor U10258 (N_10258,N_10050,N_10107);
and U10259 (N_10259,N_10140,N_10129);
nor U10260 (N_10260,N_10130,N_10192);
or U10261 (N_10261,N_10167,N_10070);
and U10262 (N_10262,N_10148,N_10075);
xnor U10263 (N_10263,N_10057,N_10002);
and U10264 (N_10264,N_10095,N_10048);
or U10265 (N_10265,N_10088,N_10110);
xnor U10266 (N_10266,N_10176,N_10018);
nand U10267 (N_10267,N_10188,N_10150);
nand U10268 (N_10268,N_10162,N_10122);
or U10269 (N_10269,N_10136,N_10064);
and U10270 (N_10270,N_10120,N_10053);
nor U10271 (N_10271,N_10175,N_10077);
xnor U10272 (N_10272,N_10039,N_10187);
and U10273 (N_10273,N_10079,N_10076);
nand U10274 (N_10274,N_10019,N_10190);
nand U10275 (N_10275,N_10082,N_10052);
nand U10276 (N_10276,N_10158,N_10058);
or U10277 (N_10277,N_10143,N_10169);
xor U10278 (N_10278,N_10061,N_10013);
xor U10279 (N_10279,N_10177,N_10023);
nor U10280 (N_10280,N_10114,N_10186);
xor U10281 (N_10281,N_10116,N_10033);
or U10282 (N_10282,N_10066,N_10042);
nand U10283 (N_10283,N_10124,N_10135);
nor U10284 (N_10284,N_10027,N_10156);
nand U10285 (N_10285,N_10113,N_10035);
xnor U10286 (N_10286,N_10101,N_10003);
nand U10287 (N_10287,N_10153,N_10026);
nand U10288 (N_10288,N_10139,N_10151);
xnor U10289 (N_10289,N_10031,N_10009);
nand U10290 (N_10290,N_10154,N_10118);
nand U10291 (N_10291,N_10121,N_10137);
nor U10292 (N_10292,N_10146,N_10112);
and U10293 (N_10293,N_10089,N_10004);
and U10294 (N_10294,N_10051,N_10090);
or U10295 (N_10295,N_10185,N_10011);
xnor U10296 (N_10296,N_10062,N_10126);
nor U10297 (N_10297,N_10106,N_10128);
nand U10298 (N_10298,N_10125,N_10174);
nand U10299 (N_10299,N_10182,N_10067);
nand U10300 (N_10300,N_10016,N_10121);
nand U10301 (N_10301,N_10053,N_10096);
xnor U10302 (N_10302,N_10154,N_10143);
xor U10303 (N_10303,N_10085,N_10115);
or U10304 (N_10304,N_10066,N_10165);
or U10305 (N_10305,N_10027,N_10076);
xnor U10306 (N_10306,N_10188,N_10120);
xnor U10307 (N_10307,N_10139,N_10071);
or U10308 (N_10308,N_10052,N_10150);
nor U10309 (N_10309,N_10080,N_10056);
nor U10310 (N_10310,N_10163,N_10027);
or U10311 (N_10311,N_10163,N_10176);
nand U10312 (N_10312,N_10090,N_10010);
xnor U10313 (N_10313,N_10190,N_10152);
nor U10314 (N_10314,N_10138,N_10167);
and U10315 (N_10315,N_10062,N_10004);
xnor U10316 (N_10316,N_10163,N_10180);
nor U10317 (N_10317,N_10034,N_10126);
xnor U10318 (N_10318,N_10173,N_10092);
xnor U10319 (N_10319,N_10033,N_10139);
xor U10320 (N_10320,N_10025,N_10184);
and U10321 (N_10321,N_10006,N_10097);
and U10322 (N_10322,N_10041,N_10036);
nor U10323 (N_10323,N_10017,N_10122);
nor U10324 (N_10324,N_10164,N_10161);
xnor U10325 (N_10325,N_10136,N_10023);
and U10326 (N_10326,N_10060,N_10184);
and U10327 (N_10327,N_10022,N_10078);
nand U10328 (N_10328,N_10188,N_10040);
xnor U10329 (N_10329,N_10198,N_10095);
nor U10330 (N_10330,N_10170,N_10162);
nand U10331 (N_10331,N_10002,N_10028);
nor U10332 (N_10332,N_10107,N_10047);
and U10333 (N_10333,N_10034,N_10140);
nor U10334 (N_10334,N_10000,N_10077);
and U10335 (N_10335,N_10172,N_10111);
or U10336 (N_10336,N_10068,N_10101);
nand U10337 (N_10337,N_10193,N_10094);
or U10338 (N_10338,N_10013,N_10072);
or U10339 (N_10339,N_10043,N_10148);
or U10340 (N_10340,N_10140,N_10146);
nand U10341 (N_10341,N_10072,N_10086);
and U10342 (N_10342,N_10019,N_10153);
and U10343 (N_10343,N_10135,N_10138);
and U10344 (N_10344,N_10190,N_10073);
or U10345 (N_10345,N_10133,N_10051);
or U10346 (N_10346,N_10127,N_10180);
nor U10347 (N_10347,N_10010,N_10151);
nor U10348 (N_10348,N_10018,N_10076);
and U10349 (N_10349,N_10014,N_10116);
nor U10350 (N_10350,N_10174,N_10057);
xnor U10351 (N_10351,N_10121,N_10147);
nor U10352 (N_10352,N_10061,N_10101);
nand U10353 (N_10353,N_10062,N_10152);
or U10354 (N_10354,N_10193,N_10130);
and U10355 (N_10355,N_10004,N_10168);
or U10356 (N_10356,N_10021,N_10191);
nand U10357 (N_10357,N_10108,N_10122);
nor U10358 (N_10358,N_10108,N_10086);
nor U10359 (N_10359,N_10134,N_10136);
and U10360 (N_10360,N_10063,N_10158);
xor U10361 (N_10361,N_10121,N_10190);
nand U10362 (N_10362,N_10035,N_10038);
or U10363 (N_10363,N_10175,N_10140);
xnor U10364 (N_10364,N_10105,N_10185);
nor U10365 (N_10365,N_10129,N_10029);
xnor U10366 (N_10366,N_10107,N_10153);
nor U10367 (N_10367,N_10013,N_10122);
nand U10368 (N_10368,N_10116,N_10155);
nand U10369 (N_10369,N_10094,N_10085);
nand U10370 (N_10370,N_10082,N_10143);
nand U10371 (N_10371,N_10184,N_10153);
nand U10372 (N_10372,N_10177,N_10165);
xor U10373 (N_10373,N_10122,N_10195);
xnor U10374 (N_10374,N_10194,N_10126);
xor U10375 (N_10375,N_10104,N_10049);
and U10376 (N_10376,N_10069,N_10087);
xor U10377 (N_10377,N_10113,N_10052);
xnor U10378 (N_10378,N_10102,N_10069);
and U10379 (N_10379,N_10149,N_10046);
and U10380 (N_10380,N_10115,N_10105);
nand U10381 (N_10381,N_10077,N_10114);
and U10382 (N_10382,N_10014,N_10102);
xnor U10383 (N_10383,N_10054,N_10097);
nand U10384 (N_10384,N_10197,N_10049);
nand U10385 (N_10385,N_10102,N_10125);
nand U10386 (N_10386,N_10089,N_10052);
or U10387 (N_10387,N_10057,N_10058);
and U10388 (N_10388,N_10155,N_10080);
xnor U10389 (N_10389,N_10177,N_10118);
nand U10390 (N_10390,N_10049,N_10009);
and U10391 (N_10391,N_10194,N_10151);
and U10392 (N_10392,N_10115,N_10142);
nor U10393 (N_10393,N_10020,N_10084);
nor U10394 (N_10394,N_10113,N_10189);
and U10395 (N_10395,N_10193,N_10024);
or U10396 (N_10396,N_10076,N_10071);
and U10397 (N_10397,N_10021,N_10056);
and U10398 (N_10398,N_10008,N_10031);
and U10399 (N_10399,N_10195,N_10056);
nand U10400 (N_10400,N_10329,N_10226);
nor U10401 (N_10401,N_10299,N_10383);
or U10402 (N_10402,N_10375,N_10271);
nor U10403 (N_10403,N_10302,N_10265);
or U10404 (N_10404,N_10394,N_10392);
nor U10405 (N_10405,N_10266,N_10246);
or U10406 (N_10406,N_10211,N_10393);
nor U10407 (N_10407,N_10335,N_10376);
nor U10408 (N_10408,N_10336,N_10253);
and U10409 (N_10409,N_10256,N_10239);
or U10410 (N_10410,N_10233,N_10369);
or U10411 (N_10411,N_10309,N_10210);
xnor U10412 (N_10412,N_10371,N_10349);
and U10413 (N_10413,N_10292,N_10387);
and U10414 (N_10414,N_10379,N_10240);
and U10415 (N_10415,N_10305,N_10268);
and U10416 (N_10416,N_10347,N_10352);
nor U10417 (N_10417,N_10332,N_10202);
or U10418 (N_10418,N_10304,N_10370);
nor U10419 (N_10419,N_10356,N_10326);
nand U10420 (N_10420,N_10200,N_10251);
xnor U10421 (N_10421,N_10362,N_10348);
and U10422 (N_10422,N_10346,N_10244);
nand U10423 (N_10423,N_10390,N_10212);
nand U10424 (N_10424,N_10248,N_10290);
nor U10425 (N_10425,N_10337,N_10238);
xnor U10426 (N_10426,N_10365,N_10316);
or U10427 (N_10427,N_10355,N_10245);
nor U10428 (N_10428,N_10317,N_10338);
xnor U10429 (N_10429,N_10324,N_10223);
and U10430 (N_10430,N_10220,N_10327);
nand U10431 (N_10431,N_10330,N_10322);
or U10432 (N_10432,N_10391,N_10232);
or U10433 (N_10433,N_10333,N_10366);
or U10434 (N_10434,N_10209,N_10255);
xnor U10435 (N_10435,N_10217,N_10206);
nor U10436 (N_10436,N_10364,N_10272);
xor U10437 (N_10437,N_10275,N_10307);
xnor U10438 (N_10438,N_10397,N_10399);
nand U10439 (N_10439,N_10353,N_10306);
and U10440 (N_10440,N_10247,N_10205);
nor U10441 (N_10441,N_10368,N_10341);
or U10442 (N_10442,N_10310,N_10340);
or U10443 (N_10443,N_10320,N_10385);
nand U10444 (N_10444,N_10313,N_10361);
or U10445 (N_10445,N_10285,N_10208);
and U10446 (N_10446,N_10230,N_10331);
xor U10447 (N_10447,N_10389,N_10325);
or U10448 (N_10448,N_10345,N_10237);
nor U10449 (N_10449,N_10300,N_10288);
nor U10450 (N_10450,N_10374,N_10204);
and U10451 (N_10451,N_10207,N_10225);
xnor U10452 (N_10452,N_10314,N_10295);
and U10453 (N_10453,N_10203,N_10218);
or U10454 (N_10454,N_10201,N_10318);
and U10455 (N_10455,N_10339,N_10367);
nor U10456 (N_10456,N_10291,N_10278);
and U10457 (N_10457,N_10298,N_10270);
and U10458 (N_10458,N_10283,N_10372);
and U10459 (N_10459,N_10213,N_10274);
nand U10460 (N_10460,N_10334,N_10219);
or U10461 (N_10461,N_10343,N_10377);
nor U10462 (N_10462,N_10354,N_10308);
xnor U10463 (N_10463,N_10235,N_10269);
or U10464 (N_10464,N_10328,N_10229);
nand U10465 (N_10465,N_10277,N_10294);
or U10466 (N_10466,N_10321,N_10359);
nand U10467 (N_10467,N_10351,N_10358);
xor U10468 (N_10468,N_10231,N_10243);
xnor U10469 (N_10469,N_10242,N_10344);
xnor U10470 (N_10470,N_10254,N_10357);
nor U10471 (N_10471,N_10216,N_10280);
nor U10472 (N_10472,N_10214,N_10315);
or U10473 (N_10473,N_10276,N_10279);
or U10474 (N_10474,N_10281,N_10384);
nor U10475 (N_10475,N_10222,N_10297);
nor U10476 (N_10476,N_10373,N_10282);
nand U10477 (N_10477,N_10311,N_10234);
or U10478 (N_10478,N_10250,N_10293);
and U10479 (N_10479,N_10342,N_10259);
nand U10480 (N_10480,N_10386,N_10264);
xor U10481 (N_10481,N_10323,N_10289);
nor U10482 (N_10482,N_10267,N_10252);
and U10483 (N_10483,N_10262,N_10360);
xnor U10484 (N_10484,N_10221,N_10363);
nand U10485 (N_10485,N_10378,N_10396);
nand U10486 (N_10486,N_10286,N_10312);
and U10487 (N_10487,N_10296,N_10301);
xnor U10488 (N_10488,N_10388,N_10303);
xor U10489 (N_10489,N_10273,N_10350);
xor U10490 (N_10490,N_10227,N_10382);
xnor U10491 (N_10491,N_10395,N_10241);
and U10492 (N_10492,N_10380,N_10257);
and U10493 (N_10493,N_10287,N_10381);
xnor U10494 (N_10494,N_10258,N_10249);
and U10495 (N_10495,N_10263,N_10260);
xnor U10496 (N_10496,N_10284,N_10236);
and U10497 (N_10497,N_10224,N_10319);
and U10498 (N_10498,N_10228,N_10261);
or U10499 (N_10499,N_10215,N_10398);
and U10500 (N_10500,N_10374,N_10348);
nor U10501 (N_10501,N_10399,N_10291);
xnor U10502 (N_10502,N_10389,N_10271);
nor U10503 (N_10503,N_10266,N_10249);
nand U10504 (N_10504,N_10255,N_10339);
and U10505 (N_10505,N_10278,N_10369);
nor U10506 (N_10506,N_10298,N_10375);
and U10507 (N_10507,N_10354,N_10358);
nor U10508 (N_10508,N_10380,N_10293);
or U10509 (N_10509,N_10245,N_10268);
and U10510 (N_10510,N_10321,N_10242);
nand U10511 (N_10511,N_10372,N_10224);
or U10512 (N_10512,N_10278,N_10266);
nor U10513 (N_10513,N_10215,N_10332);
nand U10514 (N_10514,N_10206,N_10274);
nand U10515 (N_10515,N_10333,N_10336);
nand U10516 (N_10516,N_10263,N_10212);
nand U10517 (N_10517,N_10228,N_10229);
nand U10518 (N_10518,N_10212,N_10265);
nand U10519 (N_10519,N_10355,N_10303);
nor U10520 (N_10520,N_10226,N_10377);
and U10521 (N_10521,N_10355,N_10281);
and U10522 (N_10522,N_10275,N_10370);
nand U10523 (N_10523,N_10373,N_10303);
or U10524 (N_10524,N_10270,N_10321);
nor U10525 (N_10525,N_10249,N_10375);
xor U10526 (N_10526,N_10388,N_10362);
nand U10527 (N_10527,N_10381,N_10321);
nor U10528 (N_10528,N_10372,N_10312);
nand U10529 (N_10529,N_10316,N_10231);
xnor U10530 (N_10530,N_10343,N_10349);
nand U10531 (N_10531,N_10302,N_10240);
or U10532 (N_10532,N_10280,N_10396);
nand U10533 (N_10533,N_10325,N_10245);
and U10534 (N_10534,N_10318,N_10243);
xnor U10535 (N_10535,N_10288,N_10261);
nand U10536 (N_10536,N_10363,N_10232);
nor U10537 (N_10537,N_10348,N_10278);
xor U10538 (N_10538,N_10300,N_10342);
xor U10539 (N_10539,N_10205,N_10220);
and U10540 (N_10540,N_10376,N_10369);
nor U10541 (N_10541,N_10268,N_10201);
xnor U10542 (N_10542,N_10240,N_10227);
nand U10543 (N_10543,N_10334,N_10321);
nor U10544 (N_10544,N_10301,N_10214);
and U10545 (N_10545,N_10304,N_10219);
xnor U10546 (N_10546,N_10341,N_10295);
xnor U10547 (N_10547,N_10329,N_10274);
nand U10548 (N_10548,N_10356,N_10241);
or U10549 (N_10549,N_10205,N_10388);
and U10550 (N_10550,N_10290,N_10373);
and U10551 (N_10551,N_10291,N_10363);
or U10552 (N_10552,N_10394,N_10233);
nor U10553 (N_10553,N_10213,N_10261);
and U10554 (N_10554,N_10258,N_10203);
nand U10555 (N_10555,N_10371,N_10387);
or U10556 (N_10556,N_10214,N_10224);
or U10557 (N_10557,N_10255,N_10354);
and U10558 (N_10558,N_10269,N_10296);
xor U10559 (N_10559,N_10354,N_10253);
nor U10560 (N_10560,N_10253,N_10217);
or U10561 (N_10561,N_10278,N_10328);
and U10562 (N_10562,N_10237,N_10351);
xnor U10563 (N_10563,N_10217,N_10378);
xnor U10564 (N_10564,N_10387,N_10308);
xor U10565 (N_10565,N_10386,N_10310);
or U10566 (N_10566,N_10246,N_10216);
or U10567 (N_10567,N_10259,N_10337);
xnor U10568 (N_10568,N_10291,N_10397);
nor U10569 (N_10569,N_10320,N_10288);
nand U10570 (N_10570,N_10337,N_10258);
or U10571 (N_10571,N_10217,N_10360);
or U10572 (N_10572,N_10301,N_10229);
and U10573 (N_10573,N_10359,N_10269);
xnor U10574 (N_10574,N_10364,N_10385);
or U10575 (N_10575,N_10250,N_10302);
nand U10576 (N_10576,N_10353,N_10259);
or U10577 (N_10577,N_10321,N_10210);
xnor U10578 (N_10578,N_10346,N_10315);
nor U10579 (N_10579,N_10324,N_10310);
nand U10580 (N_10580,N_10377,N_10238);
nand U10581 (N_10581,N_10224,N_10262);
xor U10582 (N_10582,N_10305,N_10378);
and U10583 (N_10583,N_10310,N_10211);
nand U10584 (N_10584,N_10348,N_10346);
xnor U10585 (N_10585,N_10390,N_10286);
xnor U10586 (N_10586,N_10234,N_10393);
xnor U10587 (N_10587,N_10272,N_10311);
and U10588 (N_10588,N_10272,N_10282);
xor U10589 (N_10589,N_10222,N_10225);
nor U10590 (N_10590,N_10223,N_10236);
xnor U10591 (N_10591,N_10278,N_10366);
nor U10592 (N_10592,N_10274,N_10341);
xor U10593 (N_10593,N_10291,N_10221);
and U10594 (N_10594,N_10251,N_10359);
nor U10595 (N_10595,N_10226,N_10331);
nand U10596 (N_10596,N_10354,N_10212);
xor U10597 (N_10597,N_10349,N_10339);
nor U10598 (N_10598,N_10384,N_10392);
or U10599 (N_10599,N_10286,N_10316);
xnor U10600 (N_10600,N_10447,N_10564);
and U10601 (N_10601,N_10426,N_10569);
or U10602 (N_10602,N_10599,N_10524);
nand U10603 (N_10603,N_10483,N_10450);
or U10604 (N_10604,N_10583,N_10449);
nor U10605 (N_10605,N_10441,N_10516);
and U10606 (N_10606,N_10493,N_10455);
xor U10607 (N_10607,N_10507,N_10579);
nor U10608 (N_10608,N_10578,N_10418);
nand U10609 (N_10609,N_10532,N_10557);
and U10610 (N_10610,N_10460,N_10407);
xor U10611 (N_10611,N_10434,N_10548);
xor U10612 (N_10612,N_10560,N_10463);
nand U10613 (N_10613,N_10526,N_10502);
xor U10614 (N_10614,N_10542,N_10475);
nor U10615 (N_10615,N_10503,N_10527);
nor U10616 (N_10616,N_10577,N_10458);
nor U10617 (N_10617,N_10467,N_10535);
and U10618 (N_10618,N_10432,N_10506);
or U10619 (N_10619,N_10427,N_10484);
or U10620 (N_10620,N_10570,N_10592);
or U10621 (N_10621,N_10496,N_10525);
or U10622 (N_10622,N_10466,N_10423);
and U10623 (N_10623,N_10480,N_10587);
nand U10624 (N_10624,N_10582,N_10487);
nor U10625 (N_10625,N_10454,N_10541);
xnor U10626 (N_10626,N_10485,N_10510);
nand U10627 (N_10627,N_10400,N_10430);
nor U10628 (N_10628,N_10531,N_10437);
nand U10629 (N_10629,N_10595,N_10433);
nor U10630 (N_10630,N_10438,N_10403);
xnor U10631 (N_10631,N_10537,N_10566);
nand U10632 (N_10632,N_10443,N_10546);
or U10633 (N_10633,N_10576,N_10405);
nor U10634 (N_10634,N_10580,N_10585);
nor U10635 (N_10635,N_10590,N_10513);
xor U10636 (N_10636,N_10536,N_10464);
xor U10637 (N_10637,N_10511,N_10422);
nand U10638 (N_10638,N_10482,N_10545);
and U10639 (N_10639,N_10440,N_10534);
or U10640 (N_10640,N_10494,N_10573);
nor U10641 (N_10641,N_10567,N_10591);
xor U10642 (N_10642,N_10508,N_10445);
or U10643 (N_10643,N_10406,N_10554);
nand U10644 (N_10644,N_10492,N_10490);
xor U10645 (N_10645,N_10424,N_10439);
nand U10646 (N_10646,N_10584,N_10498);
or U10647 (N_10647,N_10425,N_10529);
and U10648 (N_10648,N_10470,N_10465);
nor U10649 (N_10649,N_10509,N_10562);
or U10650 (N_10650,N_10409,N_10501);
nor U10651 (N_10651,N_10549,N_10551);
nor U10652 (N_10652,N_10597,N_10575);
nand U10653 (N_10653,N_10488,N_10408);
nand U10654 (N_10654,N_10481,N_10420);
nand U10655 (N_10655,N_10540,N_10572);
nand U10656 (N_10656,N_10435,N_10552);
or U10657 (N_10657,N_10495,N_10581);
xor U10658 (N_10658,N_10448,N_10412);
or U10659 (N_10659,N_10469,N_10456);
or U10660 (N_10660,N_10568,N_10512);
or U10661 (N_10661,N_10558,N_10431);
xnor U10662 (N_10662,N_10559,N_10574);
and U10663 (N_10663,N_10528,N_10596);
nor U10664 (N_10664,N_10411,N_10462);
nor U10665 (N_10665,N_10556,N_10533);
and U10666 (N_10666,N_10598,N_10586);
xor U10667 (N_10667,N_10518,N_10539);
or U10668 (N_10668,N_10404,N_10523);
or U10669 (N_10669,N_10515,N_10517);
nor U10670 (N_10670,N_10429,N_10413);
or U10671 (N_10671,N_10538,N_10442);
nand U10672 (N_10672,N_10474,N_10415);
or U10673 (N_10673,N_10504,N_10477);
nand U10674 (N_10674,N_10473,N_10410);
and U10675 (N_10675,N_10571,N_10519);
or U10676 (N_10676,N_10547,N_10436);
or U10677 (N_10677,N_10520,N_10553);
xor U10678 (N_10678,N_10461,N_10453);
nand U10679 (N_10679,N_10505,N_10491);
xor U10680 (N_10680,N_10446,N_10489);
or U10681 (N_10681,N_10402,N_10472);
xnor U10682 (N_10682,N_10452,N_10476);
nor U10683 (N_10683,N_10522,N_10544);
or U10684 (N_10684,N_10451,N_10594);
and U10685 (N_10685,N_10444,N_10555);
or U10686 (N_10686,N_10417,N_10428);
or U10687 (N_10687,N_10589,N_10478);
and U10688 (N_10688,N_10468,N_10550);
nand U10689 (N_10689,N_10514,N_10416);
or U10690 (N_10690,N_10479,N_10486);
or U10691 (N_10691,N_10530,N_10414);
and U10692 (N_10692,N_10521,N_10401);
xnor U10693 (N_10693,N_10561,N_10593);
nor U10694 (N_10694,N_10497,N_10471);
nor U10695 (N_10695,N_10500,N_10459);
nor U10696 (N_10696,N_10457,N_10543);
or U10697 (N_10697,N_10588,N_10419);
xnor U10698 (N_10698,N_10499,N_10565);
nand U10699 (N_10699,N_10421,N_10563);
xnor U10700 (N_10700,N_10419,N_10564);
nand U10701 (N_10701,N_10520,N_10430);
or U10702 (N_10702,N_10540,N_10519);
and U10703 (N_10703,N_10522,N_10449);
xnor U10704 (N_10704,N_10413,N_10557);
xor U10705 (N_10705,N_10540,N_10426);
nand U10706 (N_10706,N_10564,N_10408);
xor U10707 (N_10707,N_10405,N_10525);
or U10708 (N_10708,N_10531,N_10490);
and U10709 (N_10709,N_10437,N_10489);
or U10710 (N_10710,N_10520,N_10594);
xnor U10711 (N_10711,N_10589,N_10590);
or U10712 (N_10712,N_10462,N_10580);
xor U10713 (N_10713,N_10404,N_10517);
and U10714 (N_10714,N_10498,N_10555);
and U10715 (N_10715,N_10435,N_10433);
nor U10716 (N_10716,N_10482,N_10417);
nor U10717 (N_10717,N_10531,N_10445);
xor U10718 (N_10718,N_10435,N_10502);
and U10719 (N_10719,N_10417,N_10588);
and U10720 (N_10720,N_10407,N_10426);
nand U10721 (N_10721,N_10422,N_10474);
and U10722 (N_10722,N_10428,N_10565);
nor U10723 (N_10723,N_10521,N_10493);
nor U10724 (N_10724,N_10496,N_10503);
nor U10725 (N_10725,N_10419,N_10453);
or U10726 (N_10726,N_10503,N_10421);
and U10727 (N_10727,N_10513,N_10576);
or U10728 (N_10728,N_10464,N_10520);
and U10729 (N_10729,N_10504,N_10450);
nand U10730 (N_10730,N_10413,N_10428);
xor U10731 (N_10731,N_10526,N_10468);
or U10732 (N_10732,N_10407,N_10488);
xnor U10733 (N_10733,N_10523,N_10477);
or U10734 (N_10734,N_10553,N_10405);
or U10735 (N_10735,N_10409,N_10487);
xnor U10736 (N_10736,N_10524,N_10519);
nand U10737 (N_10737,N_10514,N_10462);
and U10738 (N_10738,N_10409,N_10470);
or U10739 (N_10739,N_10542,N_10431);
and U10740 (N_10740,N_10423,N_10524);
nand U10741 (N_10741,N_10457,N_10471);
or U10742 (N_10742,N_10444,N_10446);
xnor U10743 (N_10743,N_10408,N_10567);
nor U10744 (N_10744,N_10593,N_10590);
nor U10745 (N_10745,N_10599,N_10414);
nand U10746 (N_10746,N_10541,N_10455);
and U10747 (N_10747,N_10440,N_10437);
nor U10748 (N_10748,N_10483,N_10427);
nor U10749 (N_10749,N_10553,N_10473);
nand U10750 (N_10750,N_10469,N_10428);
and U10751 (N_10751,N_10585,N_10557);
and U10752 (N_10752,N_10479,N_10453);
nor U10753 (N_10753,N_10448,N_10503);
and U10754 (N_10754,N_10509,N_10569);
or U10755 (N_10755,N_10579,N_10508);
nand U10756 (N_10756,N_10597,N_10401);
nand U10757 (N_10757,N_10464,N_10586);
nor U10758 (N_10758,N_10573,N_10437);
or U10759 (N_10759,N_10423,N_10413);
nor U10760 (N_10760,N_10597,N_10413);
or U10761 (N_10761,N_10562,N_10495);
or U10762 (N_10762,N_10497,N_10440);
and U10763 (N_10763,N_10481,N_10476);
nand U10764 (N_10764,N_10400,N_10460);
and U10765 (N_10765,N_10546,N_10419);
or U10766 (N_10766,N_10597,N_10479);
or U10767 (N_10767,N_10516,N_10403);
nand U10768 (N_10768,N_10567,N_10491);
nand U10769 (N_10769,N_10418,N_10505);
xnor U10770 (N_10770,N_10434,N_10456);
or U10771 (N_10771,N_10443,N_10464);
and U10772 (N_10772,N_10450,N_10416);
xnor U10773 (N_10773,N_10400,N_10557);
and U10774 (N_10774,N_10506,N_10465);
or U10775 (N_10775,N_10543,N_10456);
xor U10776 (N_10776,N_10570,N_10587);
nand U10777 (N_10777,N_10505,N_10475);
nand U10778 (N_10778,N_10468,N_10536);
or U10779 (N_10779,N_10531,N_10444);
nor U10780 (N_10780,N_10492,N_10432);
xnor U10781 (N_10781,N_10461,N_10594);
xor U10782 (N_10782,N_10465,N_10554);
nor U10783 (N_10783,N_10413,N_10491);
or U10784 (N_10784,N_10406,N_10576);
nor U10785 (N_10785,N_10444,N_10400);
or U10786 (N_10786,N_10478,N_10564);
nor U10787 (N_10787,N_10513,N_10517);
or U10788 (N_10788,N_10511,N_10526);
nor U10789 (N_10789,N_10590,N_10599);
nor U10790 (N_10790,N_10438,N_10522);
xnor U10791 (N_10791,N_10466,N_10585);
nor U10792 (N_10792,N_10569,N_10429);
nor U10793 (N_10793,N_10411,N_10576);
nor U10794 (N_10794,N_10473,N_10433);
xnor U10795 (N_10795,N_10582,N_10457);
xor U10796 (N_10796,N_10519,N_10405);
nand U10797 (N_10797,N_10530,N_10596);
xor U10798 (N_10798,N_10559,N_10510);
or U10799 (N_10799,N_10599,N_10567);
and U10800 (N_10800,N_10687,N_10714);
nor U10801 (N_10801,N_10790,N_10672);
nor U10802 (N_10802,N_10622,N_10775);
nor U10803 (N_10803,N_10782,N_10638);
or U10804 (N_10804,N_10635,N_10716);
nor U10805 (N_10805,N_10666,N_10774);
nor U10806 (N_10806,N_10679,N_10670);
and U10807 (N_10807,N_10626,N_10603);
and U10808 (N_10808,N_10772,N_10715);
and U10809 (N_10809,N_10776,N_10700);
nand U10810 (N_10810,N_10769,N_10722);
nor U10811 (N_10811,N_10667,N_10606);
nor U10812 (N_10812,N_10657,N_10780);
nor U10813 (N_10813,N_10720,N_10758);
xnor U10814 (N_10814,N_10612,N_10711);
nor U10815 (N_10815,N_10724,N_10602);
and U10816 (N_10816,N_10784,N_10639);
or U10817 (N_10817,N_10773,N_10668);
nor U10818 (N_10818,N_10767,N_10743);
xor U10819 (N_10819,N_10727,N_10712);
or U10820 (N_10820,N_10601,N_10628);
nand U10821 (N_10821,N_10702,N_10740);
and U10822 (N_10822,N_10614,N_10731);
nand U10823 (N_10823,N_10631,N_10721);
nand U10824 (N_10824,N_10797,N_10733);
nand U10825 (N_10825,N_10704,N_10734);
nor U10826 (N_10826,N_10749,N_10744);
nand U10827 (N_10827,N_10732,N_10678);
nand U10828 (N_10828,N_10762,N_10786);
xnor U10829 (N_10829,N_10680,N_10699);
and U10830 (N_10830,N_10739,N_10696);
nand U10831 (N_10831,N_10779,N_10695);
or U10832 (N_10832,N_10761,N_10619);
nand U10833 (N_10833,N_10757,N_10755);
nand U10834 (N_10834,N_10798,N_10613);
nand U10835 (N_10835,N_10765,N_10600);
and U10836 (N_10836,N_10736,N_10634);
nand U10837 (N_10837,N_10741,N_10685);
nand U10838 (N_10838,N_10694,N_10609);
and U10839 (N_10839,N_10691,N_10725);
and U10840 (N_10840,N_10616,N_10728);
or U10841 (N_10841,N_10747,N_10750);
or U10842 (N_10842,N_10756,N_10665);
nor U10843 (N_10843,N_10697,N_10642);
nor U10844 (N_10844,N_10663,N_10726);
or U10845 (N_10845,N_10647,N_10682);
and U10846 (N_10846,N_10627,N_10701);
nor U10847 (N_10847,N_10783,N_10791);
and U10848 (N_10848,N_10737,N_10641);
nand U10849 (N_10849,N_10754,N_10763);
nand U10850 (N_10850,N_10677,N_10674);
xnor U10851 (N_10851,N_10708,N_10729);
nand U10852 (N_10852,N_10633,N_10673);
and U10853 (N_10853,N_10793,N_10766);
and U10854 (N_10854,N_10611,N_10751);
and U10855 (N_10855,N_10605,N_10799);
nor U10856 (N_10856,N_10618,N_10604);
nand U10857 (N_10857,N_10660,N_10698);
nor U10858 (N_10858,N_10764,N_10617);
or U10859 (N_10859,N_10796,N_10615);
and U10860 (N_10860,N_10640,N_10646);
xnor U10861 (N_10861,N_10686,N_10654);
xnor U10862 (N_10862,N_10636,N_10676);
or U10863 (N_10863,N_10620,N_10661);
or U10864 (N_10864,N_10649,N_10645);
or U10865 (N_10865,N_10794,N_10681);
xor U10866 (N_10866,N_10787,N_10759);
xnor U10867 (N_10867,N_10652,N_10777);
or U10868 (N_10868,N_10789,N_10662);
or U10869 (N_10869,N_10655,N_10738);
and U10870 (N_10870,N_10735,N_10753);
and U10871 (N_10871,N_10653,N_10643);
nor U10872 (N_10872,N_10656,N_10650);
nand U10873 (N_10873,N_10723,N_10709);
or U10874 (N_10874,N_10664,N_10717);
nor U10875 (N_10875,N_10692,N_10719);
nor U10876 (N_10876,N_10629,N_10671);
xor U10877 (N_10877,N_10689,N_10644);
nand U10878 (N_10878,N_10785,N_10637);
nand U10879 (N_10879,N_10745,N_10623);
xor U10880 (N_10880,N_10703,N_10770);
or U10881 (N_10881,N_10710,N_10705);
nor U10882 (N_10882,N_10706,N_10658);
or U10883 (N_10883,N_10788,N_10792);
and U10884 (N_10884,N_10693,N_10608);
or U10885 (N_10885,N_10621,N_10684);
nand U10886 (N_10886,N_10707,N_10768);
or U10887 (N_10887,N_10651,N_10659);
or U10888 (N_10888,N_10690,N_10781);
nor U10889 (N_10889,N_10632,N_10771);
xor U10890 (N_10890,N_10625,N_10610);
and U10891 (N_10891,N_10760,N_10752);
or U10892 (N_10892,N_10778,N_10742);
and U10893 (N_10893,N_10683,N_10669);
or U10894 (N_10894,N_10607,N_10718);
nand U10895 (N_10895,N_10748,N_10648);
nand U10896 (N_10896,N_10675,N_10795);
xnor U10897 (N_10897,N_10730,N_10630);
xnor U10898 (N_10898,N_10624,N_10713);
nor U10899 (N_10899,N_10688,N_10746);
nor U10900 (N_10900,N_10702,N_10750);
or U10901 (N_10901,N_10677,N_10725);
nor U10902 (N_10902,N_10707,N_10759);
nand U10903 (N_10903,N_10694,N_10651);
or U10904 (N_10904,N_10684,N_10751);
nor U10905 (N_10905,N_10621,N_10769);
and U10906 (N_10906,N_10625,N_10604);
xnor U10907 (N_10907,N_10613,N_10799);
nor U10908 (N_10908,N_10667,N_10797);
or U10909 (N_10909,N_10746,N_10608);
nand U10910 (N_10910,N_10765,N_10732);
or U10911 (N_10911,N_10702,N_10790);
xnor U10912 (N_10912,N_10669,N_10796);
xnor U10913 (N_10913,N_10615,N_10706);
xnor U10914 (N_10914,N_10744,N_10611);
xnor U10915 (N_10915,N_10761,N_10654);
or U10916 (N_10916,N_10600,N_10784);
nand U10917 (N_10917,N_10633,N_10695);
nor U10918 (N_10918,N_10719,N_10608);
or U10919 (N_10919,N_10690,N_10685);
xor U10920 (N_10920,N_10763,N_10782);
nor U10921 (N_10921,N_10655,N_10732);
nand U10922 (N_10922,N_10641,N_10632);
and U10923 (N_10923,N_10750,N_10631);
nor U10924 (N_10924,N_10679,N_10682);
nand U10925 (N_10925,N_10737,N_10720);
nor U10926 (N_10926,N_10677,N_10608);
nor U10927 (N_10927,N_10630,N_10657);
or U10928 (N_10928,N_10734,N_10741);
or U10929 (N_10929,N_10781,N_10631);
and U10930 (N_10930,N_10635,N_10712);
or U10931 (N_10931,N_10768,N_10727);
nor U10932 (N_10932,N_10696,N_10623);
nor U10933 (N_10933,N_10664,N_10676);
xor U10934 (N_10934,N_10654,N_10622);
and U10935 (N_10935,N_10676,N_10750);
nor U10936 (N_10936,N_10625,N_10622);
nand U10937 (N_10937,N_10701,N_10761);
or U10938 (N_10938,N_10775,N_10766);
or U10939 (N_10939,N_10736,N_10796);
xnor U10940 (N_10940,N_10711,N_10797);
and U10941 (N_10941,N_10785,N_10615);
or U10942 (N_10942,N_10617,N_10668);
xor U10943 (N_10943,N_10630,N_10629);
or U10944 (N_10944,N_10616,N_10621);
or U10945 (N_10945,N_10715,N_10625);
nor U10946 (N_10946,N_10788,N_10756);
and U10947 (N_10947,N_10666,N_10735);
nand U10948 (N_10948,N_10724,N_10645);
and U10949 (N_10949,N_10646,N_10674);
nor U10950 (N_10950,N_10603,N_10709);
and U10951 (N_10951,N_10774,N_10756);
nand U10952 (N_10952,N_10796,N_10641);
nand U10953 (N_10953,N_10696,N_10763);
or U10954 (N_10954,N_10746,N_10678);
nor U10955 (N_10955,N_10784,N_10721);
or U10956 (N_10956,N_10610,N_10620);
and U10957 (N_10957,N_10788,N_10661);
xnor U10958 (N_10958,N_10703,N_10631);
xor U10959 (N_10959,N_10624,N_10703);
and U10960 (N_10960,N_10735,N_10682);
xor U10961 (N_10961,N_10631,N_10611);
nand U10962 (N_10962,N_10700,N_10697);
nor U10963 (N_10963,N_10713,N_10621);
or U10964 (N_10964,N_10662,N_10762);
and U10965 (N_10965,N_10657,N_10623);
or U10966 (N_10966,N_10609,N_10637);
nand U10967 (N_10967,N_10679,N_10603);
nor U10968 (N_10968,N_10685,N_10644);
nor U10969 (N_10969,N_10698,N_10703);
nor U10970 (N_10970,N_10758,N_10726);
nand U10971 (N_10971,N_10715,N_10646);
nand U10972 (N_10972,N_10637,N_10762);
nor U10973 (N_10973,N_10692,N_10788);
nor U10974 (N_10974,N_10742,N_10671);
and U10975 (N_10975,N_10748,N_10797);
xnor U10976 (N_10976,N_10758,N_10649);
nor U10977 (N_10977,N_10699,N_10758);
xnor U10978 (N_10978,N_10611,N_10615);
nand U10979 (N_10979,N_10625,N_10635);
nor U10980 (N_10980,N_10674,N_10686);
nand U10981 (N_10981,N_10747,N_10787);
nand U10982 (N_10982,N_10667,N_10704);
and U10983 (N_10983,N_10792,N_10690);
or U10984 (N_10984,N_10728,N_10625);
nand U10985 (N_10985,N_10717,N_10706);
and U10986 (N_10986,N_10705,N_10761);
nand U10987 (N_10987,N_10731,N_10650);
nand U10988 (N_10988,N_10706,N_10757);
nor U10989 (N_10989,N_10711,N_10616);
nor U10990 (N_10990,N_10796,N_10688);
and U10991 (N_10991,N_10734,N_10746);
nand U10992 (N_10992,N_10730,N_10684);
nand U10993 (N_10993,N_10700,N_10744);
and U10994 (N_10994,N_10795,N_10628);
nor U10995 (N_10995,N_10603,N_10604);
nor U10996 (N_10996,N_10659,N_10698);
nand U10997 (N_10997,N_10789,N_10793);
and U10998 (N_10998,N_10673,N_10775);
nand U10999 (N_10999,N_10653,N_10796);
and U11000 (N_11000,N_10803,N_10947);
xnor U11001 (N_11001,N_10935,N_10960);
or U11002 (N_11002,N_10923,N_10823);
and U11003 (N_11003,N_10998,N_10824);
nand U11004 (N_11004,N_10847,N_10886);
nand U11005 (N_11005,N_10915,N_10927);
nand U11006 (N_11006,N_10995,N_10993);
or U11007 (N_11007,N_10811,N_10882);
nor U11008 (N_11008,N_10940,N_10950);
nand U11009 (N_11009,N_10958,N_10913);
or U11010 (N_11010,N_10836,N_10875);
nand U11011 (N_11011,N_10817,N_10837);
and U11012 (N_11012,N_10897,N_10980);
and U11013 (N_11013,N_10890,N_10864);
or U11014 (N_11014,N_10999,N_10968);
nor U11015 (N_11015,N_10894,N_10843);
and U11016 (N_11016,N_10848,N_10990);
and U11017 (N_11017,N_10978,N_10945);
nand U11018 (N_11018,N_10876,N_10939);
xnor U11019 (N_11019,N_10851,N_10802);
and U11020 (N_11020,N_10832,N_10926);
xnor U11021 (N_11021,N_10889,N_10867);
and U11022 (N_11022,N_10961,N_10825);
xor U11023 (N_11023,N_10933,N_10849);
nor U11024 (N_11024,N_10946,N_10911);
or U11025 (N_11025,N_10866,N_10975);
or U11026 (N_11026,N_10973,N_10878);
nor U11027 (N_11027,N_10887,N_10865);
nor U11028 (N_11028,N_10879,N_10903);
xor U11029 (N_11029,N_10841,N_10856);
nand U11030 (N_11030,N_10905,N_10810);
and U11031 (N_11031,N_10954,N_10839);
or U11032 (N_11032,N_10868,N_10800);
or U11033 (N_11033,N_10895,N_10853);
or U11034 (N_11034,N_10988,N_10969);
nor U11035 (N_11035,N_10924,N_10912);
and U11036 (N_11036,N_10914,N_10937);
xor U11037 (N_11037,N_10959,N_10970);
xor U11038 (N_11038,N_10992,N_10949);
and U11039 (N_11039,N_10925,N_10822);
and U11040 (N_11040,N_10852,N_10979);
nand U11041 (N_11041,N_10840,N_10909);
nor U11042 (N_11042,N_10854,N_10986);
and U11043 (N_11043,N_10870,N_10942);
xnor U11044 (N_11044,N_10902,N_10835);
nor U11045 (N_11045,N_10919,N_10855);
and U11046 (N_11046,N_10971,N_10953);
or U11047 (N_11047,N_10957,N_10918);
or U11048 (N_11048,N_10932,N_10842);
nand U11049 (N_11049,N_10908,N_10863);
nand U11050 (N_11050,N_10991,N_10891);
and U11051 (N_11051,N_10831,N_10828);
and U11052 (N_11052,N_10801,N_10815);
nand U11053 (N_11053,N_10858,N_10983);
or U11054 (N_11054,N_10936,N_10845);
xor U11055 (N_11055,N_10833,N_10859);
and U11056 (N_11056,N_10952,N_10907);
nor U11057 (N_11057,N_10910,N_10892);
or U11058 (N_11058,N_10928,N_10819);
xor U11059 (N_11059,N_10974,N_10981);
or U11060 (N_11060,N_10884,N_10846);
or U11061 (N_11061,N_10877,N_10938);
nand U11062 (N_11062,N_10898,N_10930);
nor U11063 (N_11063,N_10943,N_10885);
xor U11064 (N_11064,N_10873,N_10963);
or U11065 (N_11065,N_10955,N_10916);
nand U11066 (N_11066,N_10826,N_10862);
xnor U11067 (N_11067,N_10900,N_10857);
nand U11068 (N_11068,N_10921,N_10996);
or U11069 (N_11069,N_10965,N_10818);
or U11070 (N_11070,N_10964,N_10920);
xnor U11071 (N_11071,N_10929,N_10967);
nand U11072 (N_11072,N_10820,N_10888);
or U11073 (N_11073,N_10944,N_10809);
xor U11074 (N_11074,N_10893,N_10989);
nand U11075 (N_11075,N_10951,N_10880);
xnor U11076 (N_11076,N_10838,N_10994);
nor U11077 (N_11077,N_10816,N_10813);
nand U11078 (N_11078,N_10984,N_10966);
nor U11079 (N_11079,N_10807,N_10872);
nand U11080 (N_11080,N_10985,N_10805);
and U11081 (N_11081,N_10976,N_10899);
xnor U11082 (N_11082,N_10860,N_10901);
and U11083 (N_11083,N_10871,N_10861);
nor U11084 (N_11084,N_10931,N_10906);
nand U11085 (N_11085,N_10934,N_10962);
xnor U11086 (N_11086,N_10987,N_10869);
xnor U11087 (N_11087,N_10844,N_10977);
or U11088 (N_11088,N_10972,N_10814);
nor U11089 (N_11089,N_10904,N_10804);
or U11090 (N_11090,N_10982,N_10896);
nand U11091 (N_11091,N_10829,N_10806);
and U11092 (N_11092,N_10812,N_10850);
and U11093 (N_11093,N_10948,N_10881);
nand U11094 (N_11094,N_10997,N_10941);
or U11095 (N_11095,N_10883,N_10834);
nor U11096 (N_11096,N_10830,N_10874);
or U11097 (N_11097,N_10922,N_10821);
or U11098 (N_11098,N_10917,N_10808);
nor U11099 (N_11099,N_10827,N_10956);
or U11100 (N_11100,N_10829,N_10998);
nor U11101 (N_11101,N_10987,N_10932);
xnor U11102 (N_11102,N_10854,N_10840);
xor U11103 (N_11103,N_10925,N_10852);
nand U11104 (N_11104,N_10871,N_10800);
xor U11105 (N_11105,N_10902,N_10895);
xor U11106 (N_11106,N_10807,N_10985);
nor U11107 (N_11107,N_10813,N_10951);
nor U11108 (N_11108,N_10894,N_10823);
xnor U11109 (N_11109,N_10990,N_10950);
nand U11110 (N_11110,N_10913,N_10941);
or U11111 (N_11111,N_10822,N_10971);
and U11112 (N_11112,N_10907,N_10966);
and U11113 (N_11113,N_10919,N_10931);
xor U11114 (N_11114,N_10806,N_10889);
nand U11115 (N_11115,N_10861,N_10884);
and U11116 (N_11116,N_10880,N_10948);
and U11117 (N_11117,N_10984,N_10912);
nor U11118 (N_11118,N_10872,N_10825);
nor U11119 (N_11119,N_10812,N_10874);
nor U11120 (N_11120,N_10880,N_10844);
nor U11121 (N_11121,N_10818,N_10812);
and U11122 (N_11122,N_10832,N_10917);
nand U11123 (N_11123,N_10930,N_10901);
xor U11124 (N_11124,N_10984,N_10903);
and U11125 (N_11125,N_10851,N_10867);
or U11126 (N_11126,N_10909,N_10950);
or U11127 (N_11127,N_10903,N_10814);
nor U11128 (N_11128,N_10929,N_10842);
nand U11129 (N_11129,N_10923,N_10992);
xnor U11130 (N_11130,N_10989,N_10964);
or U11131 (N_11131,N_10852,N_10895);
nor U11132 (N_11132,N_10895,N_10959);
xnor U11133 (N_11133,N_10963,N_10849);
nand U11134 (N_11134,N_10883,N_10993);
nand U11135 (N_11135,N_10837,N_10971);
and U11136 (N_11136,N_10886,N_10874);
and U11137 (N_11137,N_10862,N_10995);
xor U11138 (N_11138,N_10976,N_10881);
nand U11139 (N_11139,N_10816,N_10865);
nand U11140 (N_11140,N_10828,N_10962);
or U11141 (N_11141,N_10949,N_10834);
and U11142 (N_11142,N_10981,N_10839);
or U11143 (N_11143,N_10939,N_10934);
and U11144 (N_11144,N_10950,N_10971);
or U11145 (N_11145,N_10892,N_10993);
nand U11146 (N_11146,N_10848,N_10859);
nor U11147 (N_11147,N_10930,N_10931);
nor U11148 (N_11148,N_10817,N_10900);
xnor U11149 (N_11149,N_10872,N_10808);
or U11150 (N_11150,N_10988,N_10849);
or U11151 (N_11151,N_10938,N_10940);
xnor U11152 (N_11152,N_10879,N_10866);
nand U11153 (N_11153,N_10895,N_10825);
or U11154 (N_11154,N_10825,N_10851);
nor U11155 (N_11155,N_10999,N_10958);
and U11156 (N_11156,N_10896,N_10839);
xnor U11157 (N_11157,N_10871,N_10905);
nand U11158 (N_11158,N_10888,N_10997);
or U11159 (N_11159,N_10952,N_10888);
or U11160 (N_11160,N_10860,N_10825);
nand U11161 (N_11161,N_10983,N_10943);
nor U11162 (N_11162,N_10878,N_10972);
and U11163 (N_11163,N_10963,N_10883);
nor U11164 (N_11164,N_10933,N_10972);
nor U11165 (N_11165,N_10894,N_10974);
nor U11166 (N_11166,N_10922,N_10941);
nand U11167 (N_11167,N_10884,N_10927);
or U11168 (N_11168,N_10820,N_10893);
nor U11169 (N_11169,N_10890,N_10952);
or U11170 (N_11170,N_10962,N_10918);
nor U11171 (N_11171,N_10855,N_10925);
xnor U11172 (N_11172,N_10836,N_10904);
or U11173 (N_11173,N_10996,N_10968);
xnor U11174 (N_11174,N_10985,N_10982);
nor U11175 (N_11175,N_10852,N_10975);
xor U11176 (N_11176,N_10965,N_10801);
nor U11177 (N_11177,N_10982,N_10857);
nor U11178 (N_11178,N_10994,N_10913);
or U11179 (N_11179,N_10832,N_10854);
nand U11180 (N_11180,N_10991,N_10853);
nand U11181 (N_11181,N_10806,N_10952);
and U11182 (N_11182,N_10803,N_10917);
nor U11183 (N_11183,N_10870,N_10872);
xnor U11184 (N_11184,N_10803,N_10885);
xor U11185 (N_11185,N_10835,N_10950);
xor U11186 (N_11186,N_10873,N_10965);
nand U11187 (N_11187,N_10926,N_10841);
xor U11188 (N_11188,N_10837,N_10862);
or U11189 (N_11189,N_10913,N_10931);
and U11190 (N_11190,N_10940,N_10930);
or U11191 (N_11191,N_10941,N_10990);
xnor U11192 (N_11192,N_10858,N_10889);
xor U11193 (N_11193,N_10833,N_10964);
or U11194 (N_11194,N_10910,N_10969);
nor U11195 (N_11195,N_10990,N_10882);
or U11196 (N_11196,N_10922,N_10926);
or U11197 (N_11197,N_10854,N_10868);
nand U11198 (N_11198,N_10870,N_10984);
nand U11199 (N_11199,N_10918,N_10852);
and U11200 (N_11200,N_11036,N_11092);
and U11201 (N_11201,N_11156,N_11031);
xnor U11202 (N_11202,N_11128,N_11091);
xor U11203 (N_11203,N_11097,N_11130);
and U11204 (N_11204,N_11023,N_11027);
nand U11205 (N_11205,N_11005,N_11154);
xor U11206 (N_11206,N_11009,N_11180);
and U11207 (N_11207,N_11077,N_11134);
or U11208 (N_11208,N_11033,N_11054);
xnor U11209 (N_11209,N_11153,N_11049);
and U11210 (N_11210,N_11021,N_11171);
nor U11211 (N_11211,N_11137,N_11120);
nor U11212 (N_11212,N_11022,N_11157);
nand U11213 (N_11213,N_11122,N_11047);
xnor U11214 (N_11214,N_11151,N_11170);
xnor U11215 (N_11215,N_11136,N_11155);
and U11216 (N_11216,N_11184,N_11085);
nor U11217 (N_11217,N_11191,N_11145);
and U11218 (N_11218,N_11080,N_11198);
and U11219 (N_11219,N_11032,N_11175);
xor U11220 (N_11220,N_11006,N_11041);
nand U11221 (N_11221,N_11152,N_11182);
nand U11222 (N_11222,N_11161,N_11076);
nor U11223 (N_11223,N_11042,N_11095);
and U11224 (N_11224,N_11146,N_11017);
or U11225 (N_11225,N_11039,N_11040);
nand U11226 (N_11226,N_11125,N_11002);
nor U11227 (N_11227,N_11069,N_11075);
and U11228 (N_11228,N_11149,N_11070);
xnor U11229 (N_11229,N_11107,N_11147);
nor U11230 (N_11230,N_11043,N_11016);
nor U11231 (N_11231,N_11018,N_11074);
xor U11232 (N_11232,N_11189,N_11081);
xor U11233 (N_11233,N_11139,N_11104);
and U11234 (N_11234,N_11164,N_11094);
nand U11235 (N_11235,N_11179,N_11056);
or U11236 (N_11236,N_11173,N_11133);
or U11237 (N_11237,N_11186,N_11062);
xor U11238 (N_11238,N_11068,N_11132);
nor U11239 (N_11239,N_11096,N_11112);
xnor U11240 (N_11240,N_11116,N_11083);
nor U11241 (N_11241,N_11008,N_11088);
and U11242 (N_11242,N_11163,N_11127);
and U11243 (N_11243,N_11020,N_11007);
or U11244 (N_11244,N_11129,N_11144);
nor U11245 (N_11245,N_11141,N_11121);
and U11246 (N_11246,N_11183,N_11038);
xor U11247 (N_11247,N_11113,N_11061);
nand U11248 (N_11248,N_11194,N_11168);
nor U11249 (N_11249,N_11174,N_11188);
or U11250 (N_11250,N_11162,N_11098);
nor U11251 (N_11251,N_11108,N_11148);
or U11252 (N_11252,N_11046,N_11159);
nor U11253 (N_11253,N_11037,N_11115);
or U11254 (N_11254,N_11169,N_11195);
xnor U11255 (N_11255,N_11109,N_11078);
nor U11256 (N_11256,N_11167,N_11196);
and U11257 (N_11257,N_11187,N_11052);
nor U11258 (N_11258,N_11138,N_11048);
nor U11259 (N_11259,N_11193,N_11012);
or U11260 (N_11260,N_11131,N_11067);
xnor U11261 (N_11261,N_11025,N_11126);
nor U11262 (N_11262,N_11089,N_11100);
nor U11263 (N_11263,N_11026,N_11172);
or U11264 (N_11264,N_11190,N_11051);
nand U11265 (N_11265,N_11199,N_11057);
xor U11266 (N_11266,N_11071,N_11044);
nand U11267 (N_11267,N_11066,N_11181);
or U11268 (N_11268,N_11101,N_11178);
or U11269 (N_11269,N_11103,N_11053);
and U11270 (N_11270,N_11063,N_11087);
nor U11271 (N_11271,N_11035,N_11019);
xor U11272 (N_11272,N_11014,N_11197);
nand U11273 (N_11273,N_11000,N_11015);
and U11274 (N_11274,N_11045,N_11105);
xnor U11275 (N_11275,N_11065,N_11124);
xnor U11276 (N_11276,N_11106,N_11084);
nor U11277 (N_11277,N_11142,N_11114);
and U11278 (N_11278,N_11177,N_11117);
or U11279 (N_11279,N_11086,N_11111);
nor U11280 (N_11280,N_11011,N_11055);
and U11281 (N_11281,N_11140,N_11185);
xor U11282 (N_11282,N_11143,N_11118);
xnor U11283 (N_11283,N_11059,N_11165);
and U11284 (N_11284,N_11034,N_11010);
nand U11285 (N_11285,N_11079,N_11004);
nand U11286 (N_11286,N_11003,N_11028);
and U11287 (N_11287,N_11123,N_11093);
and U11288 (N_11288,N_11030,N_11013);
and U11289 (N_11289,N_11192,N_11072);
xor U11290 (N_11290,N_11119,N_11176);
nor U11291 (N_11291,N_11050,N_11024);
nor U11292 (N_11292,N_11090,N_11060);
and U11293 (N_11293,N_11150,N_11082);
nor U11294 (N_11294,N_11058,N_11102);
xnor U11295 (N_11295,N_11099,N_11064);
or U11296 (N_11296,N_11166,N_11135);
nor U11297 (N_11297,N_11001,N_11073);
nand U11298 (N_11298,N_11158,N_11160);
nand U11299 (N_11299,N_11029,N_11110);
nand U11300 (N_11300,N_11122,N_11014);
or U11301 (N_11301,N_11005,N_11031);
or U11302 (N_11302,N_11062,N_11069);
or U11303 (N_11303,N_11134,N_11009);
nand U11304 (N_11304,N_11038,N_11027);
xor U11305 (N_11305,N_11049,N_11130);
xnor U11306 (N_11306,N_11061,N_11078);
nand U11307 (N_11307,N_11039,N_11180);
or U11308 (N_11308,N_11178,N_11059);
xor U11309 (N_11309,N_11131,N_11154);
or U11310 (N_11310,N_11021,N_11105);
nor U11311 (N_11311,N_11113,N_11069);
nor U11312 (N_11312,N_11074,N_11162);
nor U11313 (N_11313,N_11125,N_11000);
xor U11314 (N_11314,N_11185,N_11037);
xnor U11315 (N_11315,N_11083,N_11160);
or U11316 (N_11316,N_11149,N_11102);
nand U11317 (N_11317,N_11094,N_11138);
xnor U11318 (N_11318,N_11157,N_11072);
xnor U11319 (N_11319,N_11136,N_11123);
nor U11320 (N_11320,N_11039,N_11044);
or U11321 (N_11321,N_11073,N_11135);
nor U11322 (N_11322,N_11050,N_11135);
and U11323 (N_11323,N_11185,N_11079);
and U11324 (N_11324,N_11021,N_11145);
and U11325 (N_11325,N_11119,N_11118);
or U11326 (N_11326,N_11149,N_11074);
nand U11327 (N_11327,N_11059,N_11154);
xnor U11328 (N_11328,N_11096,N_11006);
or U11329 (N_11329,N_11170,N_11165);
or U11330 (N_11330,N_11005,N_11179);
xor U11331 (N_11331,N_11135,N_11029);
nand U11332 (N_11332,N_11126,N_11153);
xnor U11333 (N_11333,N_11026,N_11111);
xnor U11334 (N_11334,N_11056,N_11107);
or U11335 (N_11335,N_11112,N_11028);
or U11336 (N_11336,N_11159,N_11095);
xor U11337 (N_11337,N_11123,N_11113);
and U11338 (N_11338,N_11123,N_11121);
or U11339 (N_11339,N_11194,N_11116);
xor U11340 (N_11340,N_11167,N_11042);
or U11341 (N_11341,N_11047,N_11172);
xor U11342 (N_11342,N_11019,N_11098);
nand U11343 (N_11343,N_11190,N_11021);
or U11344 (N_11344,N_11020,N_11147);
xor U11345 (N_11345,N_11068,N_11056);
and U11346 (N_11346,N_11179,N_11021);
nand U11347 (N_11347,N_11068,N_11125);
xor U11348 (N_11348,N_11133,N_11155);
or U11349 (N_11349,N_11198,N_11038);
and U11350 (N_11350,N_11133,N_11179);
nand U11351 (N_11351,N_11141,N_11147);
nand U11352 (N_11352,N_11119,N_11141);
nand U11353 (N_11353,N_11005,N_11118);
nand U11354 (N_11354,N_11073,N_11120);
and U11355 (N_11355,N_11150,N_11164);
and U11356 (N_11356,N_11040,N_11074);
xor U11357 (N_11357,N_11037,N_11110);
nor U11358 (N_11358,N_11058,N_11018);
xnor U11359 (N_11359,N_11199,N_11093);
and U11360 (N_11360,N_11011,N_11082);
nand U11361 (N_11361,N_11092,N_11139);
nand U11362 (N_11362,N_11109,N_11126);
nor U11363 (N_11363,N_11130,N_11132);
xnor U11364 (N_11364,N_11113,N_11125);
xnor U11365 (N_11365,N_11150,N_11171);
nand U11366 (N_11366,N_11026,N_11184);
or U11367 (N_11367,N_11003,N_11032);
or U11368 (N_11368,N_11128,N_11009);
xor U11369 (N_11369,N_11093,N_11033);
or U11370 (N_11370,N_11079,N_11038);
nand U11371 (N_11371,N_11179,N_11046);
nand U11372 (N_11372,N_11177,N_11137);
nor U11373 (N_11373,N_11115,N_11150);
nor U11374 (N_11374,N_11015,N_11175);
nor U11375 (N_11375,N_11025,N_11061);
or U11376 (N_11376,N_11081,N_11070);
nor U11377 (N_11377,N_11065,N_11197);
and U11378 (N_11378,N_11055,N_11045);
xor U11379 (N_11379,N_11007,N_11085);
xnor U11380 (N_11380,N_11160,N_11082);
nor U11381 (N_11381,N_11043,N_11081);
nand U11382 (N_11382,N_11133,N_11110);
xor U11383 (N_11383,N_11111,N_11177);
nand U11384 (N_11384,N_11154,N_11057);
and U11385 (N_11385,N_11124,N_11170);
nor U11386 (N_11386,N_11156,N_11166);
or U11387 (N_11387,N_11000,N_11020);
nor U11388 (N_11388,N_11168,N_11012);
nand U11389 (N_11389,N_11101,N_11065);
xor U11390 (N_11390,N_11152,N_11141);
xor U11391 (N_11391,N_11192,N_11009);
or U11392 (N_11392,N_11115,N_11009);
xor U11393 (N_11393,N_11194,N_11005);
nor U11394 (N_11394,N_11042,N_11127);
nor U11395 (N_11395,N_11138,N_11135);
nor U11396 (N_11396,N_11166,N_11064);
nand U11397 (N_11397,N_11029,N_11146);
nand U11398 (N_11398,N_11174,N_11182);
nor U11399 (N_11399,N_11074,N_11067);
or U11400 (N_11400,N_11398,N_11399);
nand U11401 (N_11401,N_11302,N_11312);
nand U11402 (N_11402,N_11205,N_11392);
nand U11403 (N_11403,N_11325,N_11318);
nand U11404 (N_11404,N_11344,N_11244);
xnor U11405 (N_11405,N_11267,N_11270);
and U11406 (N_11406,N_11394,N_11339);
xor U11407 (N_11407,N_11276,N_11364);
xor U11408 (N_11408,N_11215,N_11360);
nor U11409 (N_11409,N_11251,N_11211);
nand U11410 (N_11410,N_11261,N_11236);
xor U11411 (N_11411,N_11308,N_11338);
xor U11412 (N_11412,N_11369,N_11390);
nor U11413 (N_11413,N_11271,N_11388);
xor U11414 (N_11414,N_11377,N_11375);
xnor U11415 (N_11415,N_11291,N_11387);
xor U11416 (N_11416,N_11201,N_11333);
and U11417 (N_11417,N_11239,N_11385);
or U11418 (N_11418,N_11245,N_11395);
xor U11419 (N_11419,N_11252,N_11268);
nor U11420 (N_11420,N_11259,N_11289);
xor U11421 (N_11421,N_11393,N_11351);
or U11422 (N_11422,N_11356,N_11349);
and U11423 (N_11423,N_11342,N_11269);
xnor U11424 (N_11424,N_11224,N_11240);
nor U11425 (N_11425,N_11250,N_11214);
nand U11426 (N_11426,N_11223,N_11320);
xnor U11427 (N_11427,N_11335,N_11359);
xnor U11428 (N_11428,N_11346,N_11221);
xor U11429 (N_11429,N_11357,N_11226);
xor U11430 (N_11430,N_11371,N_11286);
nand U11431 (N_11431,N_11370,N_11274);
and U11432 (N_11432,N_11353,N_11336);
or U11433 (N_11433,N_11248,N_11258);
nor U11434 (N_11434,N_11292,N_11367);
nor U11435 (N_11435,N_11288,N_11262);
or U11436 (N_11436,N_11202,N_11212);
and U11437 (N_11437,N_11222,N_11343);
and U11438 (N_11438,N_11254,N_11311);
xor U11439 (N_11439,N_11210,N_11361);
nand U11440 (N_11440,N_11200,N_11229);
nand U11441 (N_11441,N_11378,N_11382);
or U11442 (N_11442,N_11303,N_11220);
xnor U11443 (N_11443,N_11260,N_11266);
nand U11444 (N_11444,N_11279,N_11397);
or U11445 (N_11445,N_11204,N_11323);
nor U11446 (N_11446,N_11310,N_11278);
or U11447 (N_11447,N_11256,N_11253);
xor U11448 (N_11448,N_11216,N_11368);
or U11449 (N_11449,N_11396,N_11362);
nand U11450 (N_11450,N_11281,N_11213);
nor U11451 (N_11451,N_11337,N_11321);
and U11452 (N_11452,N_11247,N_11317);
nand U11453 (N_11453,N_11206,N_11373);
xnor U11454 (N_11454,N_11294,N_11327);
and U11455 (N_11455,N_11386,N_11242);
nor U11456 (N_11456,N_11280,N_11227);
xor U11457 (N_11457,N_11263,N_11230);
or U11458 (N_11458,N_11307,N_11391);
xor U11459 (N_11459,N_11316,N_11299);
nor U11460 (N_11460,N_11319,N_11381);
nand U11461 (N_11461,N_11237,N_11301);
nor U11462 (N_11462,N_11284,N_11228);
and U11463 (N_11463,N_11293,N_11257);
or U11464 (N_11464,N_11374,N_11376);
nor U11465 (N_11465,N_11309,N_11383);
xnor U11466 (N_11466,N_11366,N_11314);
or U11467 (N_11467,N_11379,N_11352);
or U11468 (N_11468,N_11218,N_11207);
nor U11469 (N_11469,N_11322,N_11298);
or U11470 (N_11470,N_11241,N_11329);
or U11471 (N_11471,N_11255,N_11358);
nor U11472 (N_11472,N_11334,N_11290);
and U11473 (N_11473,N_11347,N_11354);
nand U11474 (N_11474,N_11348,N_11235);
nand U11475 (N_11475,N_11285,N_11306);
xor U11476 (N_11476,N_11372,N_11246);
and U11477 (N_11477,N_11272,N_11234);
xnor U11478 (N_11478,N_11225,N_11328);
nor U11479 (N_11479,N_11380,N_11389);
nand U11480 (N_11480,N_11384,N_11265);
nor U11481 (N_11481,N_11313,N_11283);
nand U11482 (N_11482,N_11264,N_11282);
or U11483 (N_11483,N_11277,N_11249);
xor U11484 (N_11484,N_11305,N_11238);
xor U11485 (N_11485,N_11330,N_11287);
nand U11486 (N_11486,N_11217,N_11243);
nor U11487 (N_11487,N_11340,N_11363);
xor U11488 (N_11488,N_11296,N_11203);
and U11489 (N_11489,N_11295,N_11345);
or U11490 (N_11490,N_11232,N_11208);
and U11491 (N_11491,N_11331,N_11209);
xnor U11492 (N_11492,N_11315,N_11300);
or U11493 (N_11493,N_11332,N_11341);
and U11494 (N_11494,N_11324,N_11233);
and U11495 (N_11495,N_11304,N_11326);
xor U11496 (N_11496,N_11275,N_11365);
nand U11497 (N_11497,N_11355,N_11231);
or U11498 (N_11498,N_11273,N_11219);
nand U11499 (N_11499,N_11297,N_11350);
and U11500 (N_11500,N_11367,N_11327);
xnor U11501 (N_11501,N_11248,N_11296);
and U11502 (N_11502,N_11367,N_11284);
xor U11503 (N_11503,N_11394,N_11312);
nand U11504 (N_11504,N_11285,N_11230);
xor U11505 (N_11505,N_11266,N_11378);
or U11506 (N_11506,N_11340,N_11367);
or U11507 (N_11507,N_11335,N_11203);
nor U11508 (N_11508,N_11224,N_11362);
nand U11509 (N_11509,N_11275,N_11321);
or U11510 (N_11510,N_11263,N_11312);
nand U11511 (N_11511,N_11314,N_11374);
nand U11512 (N_11512,N_11360,N_11372);
nor U11513 (N_11513,N_11204,N_11289);
nand U11514 (N_11514,N_11298,N_11201);
or U11515 (N_11515,N_11292,N_11364);
xnor U11516 (N_11516,N_11256,N_11272);
nand U11517 (N_11517,N_11379,N_11381);
and U11518 (N_11518,N_11223,N_11337);
xor U11519 (N_11519,N_11325,N_11235);
or U11520 (N_11520,N_11382,N_11328);
xor U11521 (N_11521,N_11342,N_11207);
xnor U11522 (N_11522,N_11259,N_11218);
or U11523 (N_11523,N_11334,N_11372);
nor U11524 (N_11524,N_11241,N_11348);
and U11525 (N_11525,N_11376,N_11288);
or U11526 (N_11526,N_11257,N_11227);
and U11527 (N_11527,N_11387,N_11331);
nand U11528 (N_11528,N_11244,N_11378);
and U11529 (N_11529,N_11257,N_11218);
nand U11530 (N_11530,N_11367,N_11222);
nor U11531 (N_11531,N_11298,N_11287);
nor U11532 (N_11532,N_11252,N_11288);
or U11533 (N_11533,N_11265,N_11303);
and U11534 (N_11534,N_11371,N_11226);
and U11535 (N_11535,N_11275,N_11208);
or U11536 (N_11536,N_11215,N_11304);
nand U11537 (N_11537,N_11376,N_11237);
nor U11538 (N_11538,N_11222,N_11244);
nand U11539 (N_11539,N_11222,N_11315);
or U11540 (N_11540,N_11378,N_11326);
or U11541 (N_11541,N_11238,N_11394);
xnor U11542 (N_11542,N_11268,N_11261);
nor U11543 (N_11543,N_11215,N_11234);
nand U11544 (N_11544,N_11257,N_11233);
and U11545 (N_11545,N_11233,N_11356);
and U11546 (N_11546,N_11210,N_11321);
nand U11547 (N_11547,N_11277,N_11225);
and U11548 (N_11548,N_11342,N_11244);
xor U11549 (N_11549,N_11261,N_11243);
xor U11550 (N_11550,N_11214,N_11385);
nand U11551 (N_11551,N_11281,N_11241);
and U11552 (N_11552,N_11332,N_11363);
nor U11553 (N_11553,N_11314,N_11326);
and U11554 (N_11554,N_11380,N_11395);
nor U11555 (N_11555,N_11320,N_11389);
xor U11556 (N_11556,N_11355,N_11224);
nor U11557 (N_11557,N_11232,N_11227);
or U11558 (N_11558,N_11343,N_11321);
or U11559 (N_11559,N_11226,N_11211);
nand U11560 (N_11560,N_11360,N_11358);
nor U11561 (N_11561,N_11286,N_11361);
or U11562 (N_11562,N_11302,N_11288);
and U11563 (N_11563,N_11225,N_11387);
or U11564 (N_11564,N_11246,N_11263);
xnor U11565 (N_11565,N_11342,N_11209);
xor U11566 (N_11566,N_11347,N_11353);
nand U11567 (N_11567,N_11260,N_11317);
or U11568 (N_11568,N_11378,N_11393);
nor U11569 (N_11569,N_11398,N_11359);
and U11570 (N_11570,N_11257,N_11391);
nand U11571 (N_11571,N_11344,N_11206);
nor U11572 (N_11572,N_11320,N_11203);
nor U11573 (N_11573,N_11287,N_11280);
nand U11574 (N_11574,N_11331,N_11358);
and U11575 (N_11575,N_11327,N_11233);
nand U11576 (N_11576,N_11344,N_11250);
or U11577 (N_11577,N_11332,N_11356);
xnor U11578 (N_11578,N_11361,N_11378);
nand U11579 (N_11579,N_11343,N_11208);
or U11580 (N_11580,N_11303,N_11338);
and U11581 (N_11581,N_11318,N_11368);
or U11582 (N_11582,N_11245,N_11358);
xor U11583 (N_11583,N_11365,N_11376);
xnor U11584 (N_11584,N_11220,N_11376);
or U11585 (N_11585,N_11204,N_11372);
xor U11586 (N_11586,N_11358,N_11357);
and U11587 (N_11587,N_11364,N_11255);
nand U11588 (N_11588,N_11311,N_11309);
or U11589 (N_11589,N_11234,N_11380);
and U11590 (N_11590,N_11333,N_11365);
nor U11591 (N_11591,N_11373,N_11294);
and U11592 (N_11592,N_11211,N_11276);
nor U11593 (N_11593,N_11366,N_11361);
nor U11594 (N_11594,N_11204,N_11290);
and U11595 (N_11595,N_11236,N_11367);
or U11596 (N_11596,N_11399,N_11330);
and U11597 (N_11597,N_11315,N_11288);
and U11598 (N_11598,N_11280,N_11266);
nand U11599 (N_11599,N_11252,N_11222);
or U11600 (N_11600,N_11558,N_11586);
xnor U11601 (N_11601,N_11555,N_11531);
nand U11602 (N_11602,N_11526,N_11585);
xor U11603 (N_11603,N_11493,N_11520);
nand U11604 (N_11604,N_11412,N_11424);
xor U11605 (N_11605,N_11487,N_11500);
or U11606 (N_11606,N_11496,N_11402);
nand U11607 (N_11607,N_11430,N_11518);
xor U11608 (N_11608,N_11588,N_11401);
xnor U11609 (N_11609,N_11449,N_11599);
xor U11610 (N_11610,N_11543,N_11525);
nor U11611 (N_11611,N_11418,N_11409);
nand U11612 (N_11612,N_11565,N_11407);
xnor U11613 (N_11613,N_11420,N_11521);
and U11614 (N_11614,N_11499,N_11421);
and U11615 (N_11615,N_11538,N_11497);
or U11616 (N_11616,N_11523,N_11471);
xnor U11617 (N_11617,N_11484,N_11447);
nor U11618 (N_11618,N_11463,N_11466);
xnor U11619 (N_11619,N_11508,N_11587);
nand U11620 (N_11620,N_11436,N_11580);
or U11621 (N_11621,N_11476,N_11549);
nand U11622 (N_11622,N_11514,N_11417);
nand U11623 (N_11623,N_11532,N_11485);
xnor U11624 (N_11624,N_11503,N_11512);
xor U11625 (N_11625,N_11426,N_11429);
and U11626 (N_11626,N_11576,N_11589);
xnor U11627 (N_11627,N_11438,N_11489);
nor U11628 (N_11628,N_11492,N_11416);
or U11629 (N_11629,N_11579,N_11477);
and U11630 (N_11630,N_11551,N_11529);
xor U11631 (N_11631,N_11460,N_11459);
and U11632 (N_11632,N_11536,N_11535);
xnor U11633 (N_11633,N_11486,N_11482);
xnor U11634 (N_11634,N_11583,N_11440);
nor U11635 (N_11635,N_11572,N_11578);
nor U11636 (N_11636,N_11427,N_11480);
xnor U11637 (N_11637,N_11504,N_11542);
or U11638 (N_11638,N_11524,N_11509);
nand U11639 (N_11639,N_11511,N_11577);
nor U11640 (N_11640,N_11422,N_11465);
xnor U11641 (N_11641,N_11574,N_11554);
xnor U11642 (N_11642,N_11425,N_11562);
nand U11643 (N_11643,N_11570,N_11468);
or U11644 (N_11644,N_11483,N_11410);
xor U11645 (N_11645,N_11462,N_11419);
or U11646 (N_11646,N_11563,N_11534);
nor U11647 (N_11647,N_11550,N_11404);
xor U11648 (N_11648,N_11561,N_11467);
and U11649 (N_11649,N_11584,N_11594);
and U11650 (N_11650,N_11569,N_11461);
nand U11651 (N_11651,N_11495,N_11453);
nor U11652 (N_11652,N_11546,N_11552);
nand U11653 (N_11653,N_11411,N_11457);
or U11654 (N_11654,N_11522,N_11433);
and U11655 (N_11655,N_11544,N_11510);
nor U11656 (N_11656,N_11435,N_11590);
or U11657 (N_11657,N_11539,N_11559);
nand U11658 (N_11658,N_11553,N_11414);
nor U11659 (N_11659,N_11517,N_11481);
nor U11660 (N_11660,N_11506,N_11479);
nor U11661 (N_11661,N_11441,N_11446);
and U11662 (N_11662,N_11498,N_11519);
and U11663 (N_11663,N_11455,N_11450);
or U11664 (N_11664,N_11437,N_11456);
and U11665 (N_11665,N_11494,N_11575);
nand U11666 (N_11666,N_11557,N_11405);
nor U11667 (N_11667,N_11581,N_11595);
xor U11668 (N_11668,N_11406,N_11488);
or U11669 (N_11669,N_11458,N_11472);
nand U11670 (N_11670,N_11448,N_11431);
and U11671 (N_11671,N_11475,N_11507);
nor U11672 (N_11672,N_11582,N_11528);
and U11673 (N_11673,N_11444,N_11560);
and U11674 (N_11674,N_11478,N_11415);
or U11675 (N_11675,N_11474,N_11469);
xnor U11676 (N_11676,N_11505,N_11571);
and U11677 (N_11677,N_11464,N_11540);
or U11678 (N_11678,N_11573,N_11423);
nand U11679 (N_11679,N_11564,N_11502);
nor U11680 (N_11680,N_11439,N_11452);
xnor U11681 (N_11681,N_11547,N_11413);
or U11682 (N_11682,N_11530,N_11516);
nor U11683 (N_11683,N_11545,N_11501);
xor U11684 (N_11684,N_11533,N_11556);
nor U11685 (N_11685,N_11445,N_11596);
or U11686 (N_11686,N_11591,N_11451);
nand U11687 (N_11687,N_11548,N_11432);
and U11688 (N_11688,N_11566,N_11593);
nand U11689 (N_11689,N_11598,N_11428);
and U11690 (N_11690,N_11597,N_11434);
nor U11691 (N_11691,N_11513,N_11515);
and U11692 (N_11692,N_11491,N_11454);
nand U11693 (N_11693,N_11400,N_11568);
and U11694 (N_11694,N_11541,N_11470);
or U11695 (N_11695,N_11443,N_11490);
nand U11696 (N_11696,N_11473,N_11408);
nor U11697 (N_11697,N_11567,N_11403);
nor U11698 (N_11698,N_11592,N_11537);
xnor U11699 (N_11699,N_11442,N_11527);
nor U11700 (N_11700,N_11432,N_11421);
xnor U11701 (N_11701,N_11579,N_11584);
and U11702 (N_11702,N_11570,N_11539);
or U11703 (N_11703,N_11487,N_11506);
or U11704 (N_11704,N_11497,N_11468);
xor U11705 (N_11705,N_11467,N_11444);
and U11706 (N_11706,N_11571,N_11547);
xnor U11707 (N_11707,N_11412,N_11404);
nor U11708 (N_11708,N_11566,N_11534);
or U11709 (N_11709,N_11528,N_11447);
nor U11710 (N_11710,N_11409,N_11424);
and U11711 (N_11711,N_11403,N_11594);
or U11712 (N_11712,N_11457,N_11577);
nor U11713 (N_11713,N_11510,N_11529);
xnor U11714 (N_11714,N_11584,N_11511);
or U11715 (N_11715,N_11415,N_11404);
and U11716 (N_11716,N_11538,N_11448);
or U11717 (N_11717,N_11400,N_11442);
nor U11718 (N_11718,N_11547,N_11418);
nor U11719 (N_11719,N_11551,N_11409);
and U11720 (N_11720,N_11518,N_11508);
and U11721 (N_11721,N_11522,N_11476);
or U11722 (N_11722,N_11485,N_11479);
and U11723 (N_11723,N_11482,N_11441);
nor U11724 (N_11724,N_11426,N_11458);
and U11725 (N_11725,N_11532,N_11476);
xor U11726 (N_11726,N_11533,N_11531);
and U11727 (N_11727,N_11446,N_11428);
and U11728 (N_11728,N_11598,N_11532);
or U11729 (N_11729,N_11435,N_11400);
xor U11730 (N_11730,N_11462,N_11478);
nor U11731 (N_11731,N_11495,N_11406);
or U11732 (N_11732,N_11409,N_11530);
nor U11733 (N_11733,N_11455,N_11511);
and U11734 (N_11734,N_11517,N_11465);
or U11735 (N_11735,N_11420,N_11576);
nand U11736 (N_11736,N_11509,N_11593);
and U11737 (N_11737,N_11430,N_11460);
nand U11738 (N_11738,N_11565,N_11459);
nand U11739 (N_11739,N_11503,N_11490);
xnor U11740 (N_11740,N_11540,N_11476);
and U11741 (N_11741,N_11550,N_11493);
nand U11742 (N_11742,N_11473,N_11418);
xor U11743 (N_11743,N_11538,N_11436);
nor U11744 (N_11744,N_11422,N_11490);
nand U11745 (N_11745,N_11500,N_11474);
or U11746 (N_11746,N_11410,N_11524);
nor U11747 (N_11747,N_11583,N_11520);
nand U11748 (N_11748,N_11467,N_11469);
nand U11749 (N_11749,N_11519,N_11499);
xor U11750 (N_11750,N_11445,N_11428);
xnor U11751 (N_11751,N_11524,N_11473);
or U11752 (N_11752,N_11518,N_11515);
and U11753 (N_11753,N_11458,N_11445);
and U11754 (N_11754,N_11591,N_11507);
or U11755 (N_11755,N_11468,N_11591);
or U11756 (N_11756,N_11479,N_11445);
nor U11757 (N_11757,N_11402,N_11512);
nand U11758 (N_11758,N_11502,N_11417);
xnor U11759 (N_11759,N_11581,N_11503);
and U11760 (N_11760,N_11485,N_11517);
or U11761 (N_11761,N_11536,N_11515);
or U11762 (N_11762,N_11437,N_11597);
and U11763 (N_11763,N_11559,N_11499);
xnor U11764 (N_11764,N_11451,N_11542);
nand U11765 (N_11765,N_11447,N_11545);
nor U11766 (N_11766,N_11504,N_11587);
nand U11767 (N_11767,N_11434,N_11463);
nor U11768 (N_11768,N_11549,N_11567);
and U11769 (N_11769,N_11489,N_11538);
or U11770 (N_11770,N_11401,N_11478);
xor U11771 (N_11771,N_11448,N_11521);
nand U11772 (N_11772,N_11513,N_11416);
or U11773 (N_11773,N_11547,N_11593);
xnor U11774 (N_11774,N_11469,N_11458);
and U11775 (N_11775,N_11563,N_11452);
nand U11776 (N_11776,N_11515,N_11512);
nand U11777 (N_11777,N_11415,N_11567);
nor U11778 (N_11778,N_11515,N_11457);
xnor U11779 (N_11779,N_11561,N_11508);
nor U11780 (N_11780,N_11461,N_11412);
nor U11781 (N_11781,N_11561,N_11411);
nand U11782 (N_11782,N_11516,N_11563);
and U11783 (N_11783,N_11571,N_11479);
nand U11784 (N_11784,N_11443,N_11497);
or U11785 (N_11785,N_11514,N_11511);
nand U11786 (N_11786,N_11460,N_11466);
or U11787 (N_11787,N_11511,N_11573);
nor U11788 (N_11788,N_11472,N_11511);
nor U11789 (N_11789,N_11575,N_11469);
xnor U11790 (N_11790,N_11461,N_11527);
xnor U11791 (N_11791,N_11507,N_11447);
or U11792 (N_11792,N_11543,N_11589);
xor U11793 (N_11793,N_11596,N_11556);
xor U11794 (N_11794,N_11597,N_11491);
nor U11795 (N_11795,N_11524,N_11443);
or U11796 (N_11796,N_11533,N_11558);
nand U11797 (N_11797,N_11580,N_11589);
nand U11798 (N_11798,N_11420,N_11435);
xor U11799 (N_11799,N_11552,N_11574);
nand U11800 (N_11800,N_11731,N_11660);
nor U11801 (N_11801,N_11714,N_11648);
xor U11802 (N_11802,N_11680,N_11737);
and U11803 (N_11803,N_11676,N_11705);
nor U11804 (N_11804,N_11709,N_11695);
or U11805 (N_11805,N_11798,N_11713);
nor U11806 (N_11806,N_11744,N_11618);
nor U11807 (N_11807,N_11781,N_11613);
and U11808 (N_11808,N_11673,N_11639);
or U11809 (N_11809,N_11703,N_11726);
and U11810 (N_11810,N_11759,N_11644);
xor U11811 (N_11811,N_11698,N_11780);
nand U11812 (N_11812,N_11720,N_11752);
xor U11813 (N_11813,N_11716,N_11617);
or U11814 (N_11814,N_11769,N_11643);
nor U11815 (N_11815,N_11730,N_11692);
nand U11816 (N_11816,N_11758,N_11640);
and U11817 (N_11817,N_11756,N_11763);
nor U11818 (N_11818,N_11792,N_11665);
xnor U11819 (N_11819,N_11637,N_11717);
nand U11820 (N_11820,N_11670,N_11658);
or U11821 (N_11821,N_11710,N_11719);
nand U11822 (N_11822,N_11605,N_11642);
nor U11823 (N_11823,N_11600,N_11693);
and U11824 (N_11824,N_11632,N_11602);
or U11825 (N_11825,N_11782,N_11741);
nand U11826 (N_11826,N_11690,N_11646);
xor U11827 (N_11827,N_11764,N_11702);
and U11828 (N_11828,N_11668,N_11754);
nand U11829 (N_11829,N_11604,N_11651);
or U11830 (N_11830,N_11706,N_11649);
or U11831 (N_11831,N_11748,N_11608);
and U11832 (N_11832,N_11625,N_11610);
xor U11833 (N_11833,N_11657,N_11789);
nand U11834 (N_11834,N_11662,N_11691);
nor U11835 (N_11835,N_11677,N_11607);
xnor U11836 (N_11836,N_11689,N_11761);
xor U11837 (N_11837,N_11794,N_11772);
xor U11838 (N_11838,N_11749,N_11675);
and U11839 (N_11839,N_11628,N_11795);
and U11840 (N_11840,N_11715,N_11739);
or U11841 (N_11841,N_11738,N_11788);
nand U11842 (N_11842,N_11653,N_11609);
nand U11843 (N_11843,N_11757,N_11686);
xnor U11844 (N_11844,N_11740,N_11770);
or U11845 (N_11845,N_11614,N_11626);
xnor U11846 (N_11846,N_11685,N_11656);
or U11847 (N_11847,N_11636,N_11783);
xor U11848 (N_11848,N_11633,N_11619);
or U11849 (N_11849,N_11683,N_11684);
nand U11850 (N_11850,N_11606,N_11760);
or U11851 (N_11851,N_11681,N_11616);
xnor U11852 (N_11852,N_11712,N_11700);
or U11853 (N_11853,N_11791,N_11655);
and U11854 (N_11854,N_11793,N_11638);
nand U11855 (N_11855,N_11736,N_11629);
nand U11856 (N_11856,N_11722,N_11745);
nor U11857 (N_11857,N_11697,N_11620);
nand U11858 (N_11858,N_11721,N_11679);
nor U11859 (N_11859,N_11615,N_11762);
or U11860 (N_11860,N_11678,N_11612);
xor U11861 (N_11861,N_11733,N_11775);
and U11862 (N_11862,N_11735,N_11696);
or U11863 (N_11863,N_11767,N_11611);
xnor U11864 (N_11864,N_11711,N_11797);
nand U11865 (N_11865,N_11799,N_11768);
and U11866 (N_11866,N_11641,N_11652);
xor U11867 (N_11867,N_11766,N_11663);
nor U11868 (N_11868,N_11645,N_11773);
or U11869 (N_11869,N_11661,N_11765);
or U11870 (N_11870,N_11630,N_11750);
nor U11871 (N_11871,N_11672,N_11627);
or U11872 (N_11872,N_11732,N_11659);
and U11873 (N_11873,N_11723,N_11687);
nand U11874 (N_11874,N_11669,N_11777);
and U11875 (N_11875,N_11755,N_11624);
nand U11876 (N_11876,N_11779,N_11694);
nand U11877 (N_11877,N_11724,N_11664);
and U11878 (N_11878,N_11746,N_11725);
and U11879 (N_11879,N_11776,N_11601);
nand U11880 (N_11880,N_11790,N_11634);
xor U11881 (N_11881,N_11603,N_11771);
nor U11882 (N_11882,N_11742,N_11753);
xor U11883 (N_11883,N_11784,N_11621);
nor U11884 (N_11884,N_11654,N_11623);
nor U11885 (N_11885,N_11747,N_11674);
nor U11886 (N_11886,N_11708,N_11729);
or U11887 (N_11887,N_11778,N_11728);
and U11888 (N_11888,N_11718,N_11707);
xor U11889 (N_11889,N_11786,N_11699);
nor U11890 (N_11890,N_11667,N_11701);
nor U11891 (N_11891,N_11734,N_11631);
nor U11892 (N_11892,N_11774,N_11751);
nand U11893 (N_11893,N_11635,N_11671);
and U11894 (N_11894,N_11650,N_11727);
and U11895 (N_11895,N_11666,N_11787);
nor U11896 (N_11896,N_11647,N_11743);
xor U11897 (N_11897,N_11796,N_11622);
nand U11898 (N_11898,N_11785,N_11688);
nand U11899 (N_11899,N_11704,N_11682);
nand U11900 (N_11900,N_11701,N_11684);
or U11901 (N_11901,N_11755,N_11616);
nand U11902 (N_11902,N_11731,N_11794);
xnor U11903 (N_11903,N_11669,N_11772);
xnor U11904 (N_11904,N_11749,N_11671);
nand U11905 (N_11905,N_11749,N_11676);
nand U11906 (N_11906,N_11639,N_11783);
nand U11907 (N_11907,N_11707,N_11605);
xnor U11908 (N_11908,N_11640,N_11691);
nand U11909 (N_11909,N_11665,N_11604);
nand U11910 (N_11910,N_11791,N_11708);
nand U11911 (N_11911,N_11675,N_11710);
or U11912 (N_11912,N_11648,N_11765);
or U11913 (N_11913,N_11623,N_11729);
nand U11914 (N_11914,N_11799,N_11666);
and U11915 (N_11915,N_11641,N_11610);
or U11916 (N_11916,N_11706,N_11773);
or U11917 (N_11917,N_11666,N_11625);
or U11918 (N_11918,N_11743,N_11616);
xnor U11919 (N_11919,N_11709,N_11751);
or U11920 (N_11920,N_11713,N_11680);
and U11921 (N_11921,N_11699,N_11707);
or U11922 (N_11922,N_11655,N_11677);
nand U11923 (N_11923,N_11706,N_11618);
nor U11924 (N_11924,N_11600,N_11613);
xnor U11925 (N_11925,N_11754,N_11627);
and U11926 (N_11926,N_11783,N_11732);
and U11927 (N_11927,N_11782,N_11796);
xnor U11928 (N_11928,N_11623,N_11700);
or U11929 (N_11929,N_11763,N_11603);
and U11930 (N_11930,N_11784,N_11633);
nand U11931 (N_11931,N_11693,N_11667);
nand U11932 (N_11932,N_11710,N_11608);
nor U11933 (N_11933,N_11647,N_11655);
and U11934 (N_11934,N_11624,N_11681);
nor U11935 (N_11935,N_11602,N_11683);
nor U11936 (N_11936,N_11693,N_11678);
nor U11937 (N_11937,N_11794,N_11757);
and U11938 (N_11938,N_11734,N_11707);
nand U11939 (N_11939,N_11794,N_11785);
xnor U11940 (N_11940,N_11729,N_11689);
nor U11941 (N_11941,N_11785,N_11777);
nor U11942 (N_11942,N_11750,N_11660);
xnor U11943 (N_11943,N_11646,N_11733);
nand U11944 (N_11944,N_11615,N_11792);
and U11945 (N_11945,N_11601,N_11669);
xnor U11946 (N_11946,N_11745,N_11738);
and U11947 (N_11947,N_11609,N_11605);
xnor U11948 (N_11948,N_11614,N_11642);
xor U11949 (N_11949,N_11651,N_11790);
nor U11950 (N_11950,N_11633,N_11604);
or U11951 (N_11951,N_11711,N_11758);
xor U11952 (N_11952,N_11764,N_11759);
and U11953 (N_11953,N_11630,N_11602);
nor U11954 (N_11954,N_11784,N_11615);
or U11955 (N_11955,N_11739,N_11797);
xor U11956 (N_11956,N_11632,N_11796);
nor U11957 (N_11957,N_11744,N_11643);
nor U11958 (N_11958,N_11743,N_11652);
and U11959 (N_11959,N_11767,N_11751);
nand U11960 (N_11960,N_11745,N_11733);
nor U11961 (N_11961,N_11673,N_11720);
nor U11962 (N_11962,N_11683,N_11664);
nor U11963 (N_11963,N_11787,N_11623);
nor U11964 (N_11964,N_11648,N_11726);
nor U11965 (N_11965,N_11740,N_11639);
nor U11966 (N_11966,N_11670,N_11797);
xor U11967 (N_11967,N_11710,N_11767);
nand U11968 (N_11968,N_11784,N_11608);
xnor U11969 (N_11969,N_11783,N_11713);
nor U11970 (N_11970,N_11755,N_11651);
or U11971 (N_11971,N_11671,N_11644);
nand U11972 (N_11972,N_11729,N_11793);
nor U11973 (N_11973,N_11713,N_11601);
xor U11974 (N_11974,N_11715,N_11600);
nand U11975 (N_11975,N_11699,N_11666);
xor U11976 (N_11976,N_11742,N_11625);
and U11977 (N_11977,N_11656,N_11668);
xnor U11978 (N_11978,N_11667,N_11603);
xnor U11979 (N_11979,N_11700,N_11750);
nand U11980 (N_11980,N_11626,N_11721);
nand U11981 (N_11981,N_11687,N_11787);
xor U11982 (N_11982,N_11724,N_11669);
xnor U11983 (N_11983,N_11725,N_11656);
nand U11984 (N_11984,N_11652,N_11776);
nor U11985 (N_11985,N_11735,N_11627);
nor U11986 (N_11986,N_11794,N_11667);
xnor U11987 (N_11987,N_11786,N_11716);
xor U11988 (N_11988,N_11653,N_11739);
xor U11989 (N_11989,N_11768,N_11642);
or U11990 (N_11990,N_11662,N_11763);
nand U11991 (N_11991,N_11601,N_11751);
or U11992 (N_11992,N_11665,N_11729);
and U11993 (N_11993,N_11677,N_11699);
and U11994 (N_11994,N_11707,N_11670);
and U11995 (N_11995,N_11756,N_11775);
nand U11996 (N_11996,N_11707,N_11640);
or U11997 (N_11997,N_11622,N_11763);
nor U11998 (N_11998,N_11754,N_11740);
or U11999 (N_11999,N_11757,N_11731);
xnor U12000 (N_12000,N_11867,N_11813);
nor U12001 (N_12001,N_11984,N_11839);
and U12002 (N_12002,N_11838,N_11983);
nand U12003 (N_12003,N_11951,N_11831);
nor U12004 (N_12004,N_11934,N_11835);
xor U12005 (N_12005,N_11965,N_11880);
xor U12006 (N_12006,N_11846,N_11808);
xnor U12007 (N_12007,N_11985,N_11950);
and U12008 (N_12008,N_11942,N_11829);
or U12009 (N_12009,N_11809,N_11865);
and U12010 (N_12010,N_11891,N_11817);
and U12011 (N_12011,N_11810,N_11890);
nand U12012 (N_12012,N_11894,N_11904);
xor U12013 (N_12013,N_11933,N_11971);
or U12014 (N_12014,N_11958,N_11992);
nand U12015 (N_12015,N_11820,N_11849);
and U12016 (N_12016,N_11818,N_11804);
xor U12017 (N_12017,N_11910,N_11889);
nand U12018 (N_12018,N_11929,N_11801);
nand U12019 (N_12019,N_11938,N_11981);
nand U12020 (N_12020,N_11932,N_11848);
or U12021 (N_12021,N_11979,N_11995);
and U12022 (N_12022,N_11896,N_11954);
xor U12023 (N_12023,N_11842,N_11960);
and U12024 (N_12024,N_11850,N_11953);
or U12025 (N_12025,N_11859,N_11967);
and U12026 (N_12026,N_11921,N_11861);
and U12027 (N_12027,N_11852,N_11897);
nor U12028 (N_12028,N_11991,N_11874);
or U12029 (N_12029,N_11819,N_11976);
xnor U12030 (N_12030,N_11858,N_11836);
and U12031 (N_12031,N_11925,N_11902);
nand U12032 (N_12032,N_11977,N_11847);
nand U12033 (N_12033,N_11968,N_11988);
and U12034 (N_12034,N_11827,N_11937);
nor U12035 (N_12035,N_11893,N_11828);
nand U12036 (N_12036,N_11906,N_11916);
xnor U12037 (N_12037,N_11803,N_11924);
xor U12038 (N_12038,N_11821,N_11966);
or U12039 (N_12039,N_11907,N_11993);
xnor U12040 (N_12040,N_11826,N_11879);
xnor U12041 (N_12041,N_11941,N_11935);
xor U12042 (N_12042,N_11816,N_11901);
nand U12043 (N_12043,N_11844,N_11898);
nand U12044 (N_12044,N_11961,N_11980);
nand U12045 (N_12045,N_11974,N_11882);
nand U12046 (N_12046,N_11918,N_11853);
or U12047 (N_12047,N_11870,N_11860);
or U12048 (N_12048,N_11866,N_11956);
nor U12049 (N_12049,N_11923,N_11973);
nand U12050 (N_12050,N_11963,N_11875);
nor U12051 (N_12051,N_11952,N_11903);
nor U12052 (N_12052,N_11917,N_11940);
and U12053 (N_12053,N_11946,N_11944);
nand U12054 (N_12054,N_11825,N_11845);
nor U12055 (N_12055,N_11999,N_11948);
or U12056 (N_12056,N_11883,N_11833);
or U12057 (N_12057,N_11877,N_11878);
nor U12058 (N_12058,N_11996,N_11943);
and U12059 (N_12059,N_11868,N_11851);
nand U12060 (N_12060,N_11911,N_11947);
xnor U12061 (N_12061,N_11945,N_11990);
nand U12062 (N_12062,N_11857,N_11823);
nor U12063 (N_12063,N_11872,N_11840);
xnor U12064 (N_12064,N_11997,N_11873);
and U12065 (N_12065,N_11869,N_11892);
nand U12066 (N_12066,N_11912,N_11915);
or U12067 (N_12067,N_11982,N_11811);
and U12068 (N_12068,N_11936,N_11928);
xor U12069 (N_12069,N_11855,N_11806);
xor U12070 (N_12070,N_11899,N_11909);
nor U12071 (N_12071,N_11824,N_11905);
nor U12072 (N_12072,N_11815,N_11962);
or U12073 (N_12073,N_11931,N_11871);
or U12074 (N_12074,N_11986,N_11989);
or U12075 (N_12075,N_11886,N_11888);
nand U12076 (N_12076,N_11884,N_11900);
xnor U12077 (N_12077,N_11919,N_11856);
or U12078 (N_12078,N_11805,N_11998);
and U12079 (N_12079,N_11895,N_11876);
nand U12080 (N_12080,N_11807,N_11920);
xnor U12081 (N_12081,N_11969,N_11930);
nand U12082 (N_12082,N_11927,N_11881);
and U12083 (N_12083,N_11939,N_11854);
or U12084 (N_12084,N_11863,N_11841);
nor U12085 (N_12085,N_11955,N_11970);
or U12086 (N_12086,N_11843,N_11800);
or U12087 (N_12087,N_11978,N_11802);
and U12088 (N_12088,N_11914,N_11864);
nor U12089 (N_12089,N_11814,N_11922);
or U12090 (N_12090,N_11812,N_11887);
and U12091 (N_12091,N_11913,N_11959);
xnor U12092 (N_12092,N_11822,N_11987);
or U12093 (N_12093,N_11837,N_11975);
nor U12094 (N_12094,N_11957,N_11964);
and U12095 (N_12095,N_11885,N_11908);
or U12096 (N_12096,N_11949,N_11926);
nand U12097 (N_12097,N_11832,N_11862);
nand U12098 (N_12098,N_11972,N_11834);
nand U12099 (N_12099,N_11830,N_11994);
xnor U12100 (N_12100,N_11952,N_11822);
nand U12101 (N_12101,N_11864,N_11867);
or U12102 (N_12102,N_11902,N_11837);
xor U12103 (N_12103,N_11859,N_11837);
nand U12104 (N_12104,N_11839,N_11980);
nand U12105 (N_12105,N_11987,N_11956);
or U12106 (N_12106,N_11876,N_11897);
and U12107 (N_12107,N_11852,N_11987);
or U12108 (N_12108,N_11936,N_11973);
and U12109 (N_12109,N_11887,N_11808);
xnor U12110 (N_12110,N_11840,N_11836);
or U12111 (N_12111,N_11881,N_11971);
and U12112 (N_12112,N_11801,N_11919);
or U12113 (N_12113,N_11814,N_11893);
xnor U12114 (N_12114,N_11956,N_11969);
and U12115 (N_12115,N_11826,N_11968);
and U12116 (N_12116,N_11843,N_11974);
nand U12117 (N_12117,N_11864,N_11860);
or U12118 (N_12118,N_11819,N_11895);
nor U12119 (N_12119,N_11931,N_11895);
xnor U12120 (N_12120,N_11973,N_11825);
nor U12121 (N_12121,N_11800,N_11914);
and U12122 (N_12122,N_11993,N_11845);
or U12123 (N_12123,N_11884,N_11870);
or U12124 (N_12124,N_11962,N_11836);
and U12125 (N_12125,N_11924,N_11842);
or U12126 (N_12126,N_11924,N_11860);
and U12127 (N_12127,N_11837,N_11805);
xor U12128 (N_12128,N_11862,N_11973);
and U12129 (N_12129,N_11808,N_11950);
xor U12130 (N_12130,N_11932,N_11945);
nor U12131 (N_12131,N_11884,N_11974);
nor U12132 (N_12132,N_11830,N_11905);
nand U12133 (N_12133,N_11951,N_11992);
xor U12134 (N_12134,N_11828,N_11904);
nand U12135 (N_12135,N_11985,N_11870);
or U12136 (N_12136,N_11927,N_11834);
xnor U12137 (N_12137,N_11831,N_11979);
nor U12138 (N_12138,N_11845,N_11849);
xnor U12139 (N_12139,N_11817,N_11987);
xnor U12140 (N_12140,N_11988,N_11924);
nor U12141 (N_12141,N_11867,N_11837);
or U12142 (N_12142,N_11909,N_11916);
nor U12143 (N_12143,N_11824,N_11995);
nor U12144 (N_12144,N_11801,N_11889);
xnor U12145 (N_12145,N_11980,N_11984);
xor U12146 (N_12146,N_11959,N_11802);
xor U12147 (N_12147,N_11865,N_11846);
xnor U12148 (N_12148,N_11846,N_11907);
nor U12149 (N_12149,N_11958,N_11988);
and U12150 (N_12150,N_11957,N_11907);
nand U12151 (N_12151,N_11823,N_11929);
or U12152 (N_12152,N_11886,N_11878);
nor U12153 (N_12153,N_11979,N_11871);
or U12154 (N_12154,N_11981,N_11902);
nor U12155 (N_12155,N_11933,N_11860);
or U12156 (N_12156,N_11994,N_11825);
or U12157 (N_12157,N_11944,N_11860);
or U12158 (N_12158,N_11816,N_11910);
or U12159 (N_12159,N_11975,N_11863);
xnor U12160 (N_12160,N_11843,N_11829);
xor U12161 (N_12161,N_11886,N_11961);
or U12162 (N_12162,N_11837,N_11830);
nand U12163 (N_12163,N_11882,N_11918);
and U12164 (N_12164,N_11838,N_11910);
nor U12165 (N_12165,N_11993,N_11886);
or U12166 (N_12166,N_11832,N_11833);
xor U12167 (N_12167,N_11990,N_11950);
and U12168 (N_12168,N_11834,N_11811);
nor U12169 (N_12169,N_11907,N_11868);
and U12170 (N_12170,N_11914,N_11984);
nor U12171 (N_12171,N_11821,N_11824);
xor U12172 (N_12172,N_11999,N_11868);
or U12173 (N_12173,N_11942,N_11805);
nand U12174 (N_12174,N_11919,N_11834);
nor U12175 (N_12175,N_11824,N_11877);
nand U12176 (N_12176,N_11991,N_11863);
nor U12177 (N_12177,N_11949,N_11842);
nor U12178 (N_12178,N_11896,N_11996);
xor U12179 (N_12179,N_11884,N_11831);
or U12180 (N_12180,N_11890,N_11984);
nor U12181 (N_12181,N_11870,N_11890);
and U12182 (N_12182,N_11817,N_11838);
xor U12183 (N_12183,N_11897,N_11921);
nand U12184 (N_12184,N_11831,N_11894);
nor U12185 (N_12185,N_11988,N_11935);
xor U12186 (N_12186,N_11981,N_11836);
nand U12187 (N_12187,N_11923,N_11846);
nor U12188 (N_12188,N_11900,N_11929);
xnor U12189 (N_12189,N_11925,N_11811);
or U12190 (N_12190,N_11972,N_11892);
nand U12191 (N_12191,N_11943,N_11849);
xor U12192 (N_12192,N_11963,N_11971);
nand U12193 (N_12193,N_11972,N_11821);
or U12194 (N_12194,N_11936,N_11984);
nor U12195 (N_12195,N_11871,N_11844);
nand U12196 (N_12196,N_11890,N_11850);
nand U12197 (N_12197,N_11833,N_11945);
nand U12198 (N_12198,N_11957,N_11908);
or U12199 (N_12199,N_11972,N_11929);
nor U12200 (N_12200,N_12052,N_12023);
nor U12201 (N_12201,N_12040,N_12104);
or U12202 (N_12202,N_12025,N_12181);
nor U12203 (N_12203,N_12072,N_12064);
nor U12204 (N_12204,N_12071,N_12082);
nor U12205 (N_12205,N_12192,N_12037);
nor U12206 (N_12206,N_12050,N_12122);
nor U12207 (N_12207,N_12036,N_12191);
nor U12208 (N_12208,N_12039,N_12041);
or U12209 (N_12209,N_12046,N_12070);
xor U12210 (N_12210,N_12068,N_12038);
or U12211 (N_12211,N_12076,N_12145);
nor U12212 (N_12212,N_12043,N_12093);
xor U12213 (N_12213,N_12148,N_12128);
nor U12214 (N_12214,N_12012,N_12097);
nor U12215 (N_12215,N_12024,N_12010);
nor U12216 (N_12216,N_12014,N_12144);
and U12217 (N_12217,N_12149,N_12141);
xor U12218 (N_12218,N_12170,N_12103);
nor U12219 (N_12219,N_12178,N_12047);
nor U12220 (N_12220,N_12188,N_12013);
nor U12221 (N_12221,N_12173,N_12008);
or U12222 (N_12222,N_12180,N_12094);
and U12223 (N_12223,N_12033,N_12101);
nor U12224 (N_12224,N_12183,N_12019);
or U12225 (N_12225,N_12140,N_12190);
nor U12226 (N_12226,N_12150,N_12127);
nor U12227 (N_12227,N_12078,N_12113);
nor U12228 (N_12228,N_12118,N_12098);
nand U12229 (N_12229,N_12117,N_12179);
and U12230 (N_12230,N_12116,N_12086);
xnor U12231 (N_12231,N_12137,N_12080);
xor U12232 (N_12232,N_12074,N_12184);
xor U12233 (N_12233,N_12091,N_12151);
or U12234 (N_12234,N_12139,N_12168);
or U12235 (N_12235,N_12108,N_12169);
xnor U12236 (N_12236,N_12085,N_12102);
nor U12237 (N_12237,N_12121,N_12146);
xnor U12238 (N_12238,N_12177,N_12032);
or U12239 (N_12239,N_12090,N_12026);
and U12240 (N_12240,N_12016,N_12042);
nor U12241 (N_12241,N_12194,N_12163);
xnor U12242 (N_12242,N_12199,N_12002);
or U12243 (N_12243,N_12197,N_12020);
nor U12244 (N_12244,N_12106,N_12028);
nor U12245 (N_12245,N_12054,N_12143);
and U12246 (N_12246,N_12182,N_12000);
xnor U12247 (N_12247,N_12115,N_12065);
nor U12248 (N_12248,N_12073,N_12147);
nand U12249 (N_12249,N_12011,N_12152);
or U12250 (N_12250,N_12089,N_12109);
nand U12251 (N_12251,N_12079,N_12027);
and U12252 (N_12252,N_12049,N_12165);
or U12253 (N_12253,N_12196,N_12006);
nand U12254 (N_12254,N_12135,N_12056);
and U12255 (N_12255,N_12001,N_12185);
or U12256 (N_12256,N_12095,N_12167);
nand U12257 (N_12257,N_12112,N_12132);
or U12258 (N_12258,N_12142,N_12100);
or U12259 (N_12259,N_12134,N_12017);
nand U12260 (N_12260,N_12081,N_12129);
nor U12261 (N_12261,N_12159,N_12105);
xnor U12262 (N_12262,N_12171,N_12058);
nor U12263 (N_12263,N_12030,N_12186);
nand U12264 (N_12264,N_12174,N_12005);
or U12265 (N_12265,N_12077,N_12031);
xor U12266 (N_12266,N_12075,N_12018);
nor U12267 (N_12267,N_12066,N_12069);
nor U12268 (N_12268,N_12045,N_12126);
xnor U12269 (N_12269,N_12034,N_12176);
and U12270 (N_12270,N_12189,N_12063);
nor U12271 (N_12271,N_12007,N_12138);
or U12272 (N_12272,N_12107,N_12004);
or U12273 (N_12273,N_12125,N_12029);
nor U12274 (N_12274,N_12021,N_12061);
nor U12275 (N_12275,N_12120,N_12124);
and U12276 (N_12276,N_12158,N_12133);
nand U12277 (N_12277,N_12160,N_12154);
nor U12278 (N_12278,N_12123,N_12156);
nor U12279 (N_12279,N_12164,N_12083);
nand U12280 (N_12280,N_12053,N_12048);
or U12281 (N_12281,N_12087,N_12111);
or U12282 (N_12282,N_12051,N_12015);
xnor U12283 (N_12283,N_12119,N_12009);
or U12284 (N_12284,N_12099,N_12062);
nand U12285 (N_12285,N_12059,N_12172);
nand U12286 (N_12286,N_12193,N_12088);
and U12287 (N_12287,N_12166,N_12084);
xor U12288 (N_12288,N_12057,N_12055);
and U12289 (N_12289,N_12130,N_12161);
xor U12290 (N_12290,N_12060,N_12035);
or U12291 (N_12291,N_12162,N_12131);
nand U12292 (N_12292,N_12003,N_12067);
nand U12293 (N_12293,N_12022,N_12044);
xnor U12294 (N_12294,N_12114,N_12195);
xor U12295 (N_12295,N_12155,N_12157);
or U12296 (N_12296,N_12187,N_12175);
and U12297 (N_12297,N_12198,N_12110);
nor U12298 (N_12298,N_12096,N_12136);
xnor U12299 (N_12299,N_12153,N_12092);
nand U12300 (N_12300,N_12093,N_12107);
xnor U12301 (N_12301,N_12018,N_12139);
xnor U12302 (N_12302,N_12188,N_12175);
nand U12303 (N_12303,N_12109,N_12152);
or U12304 (N_12304,N_12054,N_12018);
nor U12305 (N_12305,N_12093,N_12005);
xor U12306 (N_12306,N_12113,N_12056);
nand U12307 (N_12307,N_12151,N_12097);
and U12308 (N_12308,N_12008,N_12171);
xor U12309 (N_12309,N_12189,N_12076);
nand U12310 (N_12310,N_12020,N_12054);
nor U12311 (N_12311,N_12165,N_12008);
or U12312 (N_12312,N_12147,N_12195);
or U12313 (N_12313,N_12006,N_12021);
or U12314 (N_12314,N_12122,N_12103);
nor U12315 (N_12315,N_12090,N_12161);
nor U12316 (N_12316,N_12139,N_12086);
and U12317 (N_12317,N_12142,N_12073);
xor U12318 (N_12318,N_12109,N_12149);
nand U12319 (N_12319,N_12005,N_12064);
and U12320 (N_12320,N_12186,N_12077);
xnor U12321 (N_12321,N_12148,N_12086);
xor U12322 (N_12322,N_12169,N_12144);
nor U12323 (N_12323,N_12113,N_12082);
nor U12324 (N_12324,N_12022,N_12186);
nand U12325 (N_12325,N_12074,N_12032);
or U12326 (N_12326,N_12074,N_12102);
nand U12327 (N_12327,N_12105,N_12068);
nor U12328 (N_12328,N_12141,N_12098);
or U12329 (N_12329,N_12099,N_12106);
and U12330 (N_12330,N_12140,N_12058);
xnor U12331 (N_12331,N_12000,N_12072);
or U12332 (N_12332,N_12027,N_12115);
nand U12333 (N_12333,N_12128,N_12020);
and U12334 (N_12334,N_12097,N_12165);
and U12335 (N_12335,N_12193,N_12139);
nor U12336 (N_12336,N_12020,N_12146);
and U12337 (N_12337,N_12020,N_12059);
or U12338 (N_12338,N_12192,N_12159);
xor U12339 (N_12339,N_12054,N_12139);
nand U12340 (N_12340,N_12023,N_12123);
and U12341 (N_12341,N_12067,N_12041);
and U12342 (N_12342,N_12114,N_12058);
and U12343 (N_12343,N_12007,N_12020);
nand U12344 (N_12344,N_12122,N_12056);
and U12345 (N_12345,N_12031,N_12133);
xnor U12346 (N_12346,N_12181,N_12086);
nor U12347 (N_12347,N_12101,N_12079);
xnor U12348 (N_12348,N_12177,N_12178);
and U12349 (N_12349,N_12015,N_12175);
xnor U12350 (N_12350,N_12156,N_12049);
xor U12351 (N_12351,N_12191,N_12068);
nor U12352 (N_12352,N_12154,N_12167);
nand U12353 (N_12353,N_12008,N_12007);
or U12354 (N_12354,N_12077,N_12114);
nand U12355 (N_12355,N_12148,N_12151);
nand U12356 (N_12356,N_12014,N_12181);
xnor U12357 (N_12357,N_12089,N_12164);
and U12358 (N_12358,N_12060,N_12099);
and U12359 (N_12359,N_12151,N_12057);
and U12360 (N_12360,N_12060,N_12150);
xor U12361 (N_12361,N_12002,N_12120);
nand U12362 (N_12362,N_12128,N_12101);
and U12363 (N_12363,N_12180,N_12176);
xnor U12364 (N_12364,N_12190,N_12004);
xnor U12365 (N_12365,N_12087,N_12102);
nor U12366 (N_12366,N_12023,N_12042);
nand U12367 (N_12367,N_12001,N_12070);
and U12368 (N_12368,N_12132,N_12173);
and U12369 (N_12369,N_12157,N_12010);
xor U12370 (N_12370,N_12014,N_12123);
xnor U12371 (N_12371,N_12160,N_12058);
nand U12372 (N_12372,N_12115,N_12074);
or U12373 (N_12373,N_12046,N_12042);
xnor U12374 (N_12374,N_12116,N_12031);
and U12375 (N_12375,N_12082,N_12175);
nor U12376 (N_12376,N_12120,N_12147);
and U12377 (N_12377,N_12141,N_12128);
nand U12378 (N_12378,N_12052,N_12061);
nand U12379 (N_12379,N_12045,N_12087);
nand U12380 (N_12380,N_12081,N_12065);
xnor U12381 (N_12381,N_12084,N_12050);
or U12382 (N_12382,N_12143,N_12149);
nor U12383 (N_12383,N_12055,N_12095);
nand U12384 (N_12384,N_12176,N_12070);
xnor U12385 (N_12385,N_12024,N_12081);
nand U12386 (N_12386,N_12104,N_12138);
or U12387 (N_12387,N_12127,N_12101);
xnor U12388 (N_12388,N_12052,N_12097);
and U12389 (N_12389,N_12026,N_12023);
and U12390 (N_12390,N_12186,N_12123);
or U12391 (N_12391,N_12180,N_12190);
and U12392 (N_12392,N_12192,N_12169);
nand U12393 (N_12393,N_12036,N_12177);
nor U12394 (N_12394,N_12048,N_12062);
xor U12395 (N_12395,N_12139,N_12091);
and U12396 (N_12396,N_12095,N_12169);
or U12397 (N_12397,N_12007,N_12136);
or U12398 (N_12398,N_12181,N_12091);
or U12399 (N_12399,N_12067,N_12038);
nor U12400 (N_12400,N_12391,N_12285);
or U12401 (N_12401,N_12271,N_12304);
or U12402 (N_12402,N_12338,N_12233);
and U12403 (N_12403,N_12278,N_12242);
and U12404 (N_12404,N_12267,N_12337);
or U12405 (N_12405,N_12293,N_12254);
xnor U12406 (N_12406,N_12274,N_12286);
or U12407 (N_12407,N_12346,N_12394);
nor U12408 (N_12408,N_12206,N_12297);
and U12409 (N_12409,N_12247,N_12389);
nand U12410 (N_12410,N_12288,N_12224);
or U12411 (N_12411,N_12357,N_12273);
nand U12412 (N_12412,N_12317,N_12232);
or U12413 (N_12413,N_12381,N_12359);
xnor U12414 (N_12414,N_12301,N_12373);
nor U12415 (N_12415,N_12272,N_12200);
and U12416 (N_12416,N_12344,N_12318);
xnor U12417 (N_12417,N_12340,N_12253);
or U12418 (N_12418,N_12299,N_12269);
or U12419 (N_12419,N_12364,N_12398);
xor U12420 (N_12420,N_12214,N_12252);
nand U12421 (N_12421,N_12308,N_12343);
nor U12422 (N_12422,N_12323,N_12264);
and U12423 (N_12423,N_12202,N_12270);
nand U12424 (N_12424,N_12289,N_12309);
and U12425 (N_12425,N_12368,N_12372);
nand U12426 (N_12426,N_12383,N_12305);
nand U12427 (N_12427,N_12213,N_12259);
nor U12428 (N_12428,N_12386,N_12326);
and U12429 (N_12429,N_12203,N_12369);
xnor U12430 (N_12430,N_12234,N_12370);
nand U12431 (N_12431,N_12230,N_12324);
nand U12432 (N_12432,N_12312,N_12399);
and U12433 (N_12433,N_12260,N_12223);
or U12434 (N_12434,N_12333,N_12240);
xor U12435 (N_12435,N_12377,N_12235);
and U12436 (N_12436,N_12294,N_12282);
and U12437 (N_12437,N_12210,N_12284);
nand U12438 (N_12438,N_12315,N_12311);
or U12439 (N_12439,N_12397,N_12376);
nand U12440 (N_12440,N_12204,N_12392);
nor U12441 (N_12441,N_12212,N_12251);
nor U12442 (N_12442,N_12395,N_12291);
xnor U12443 (N_12443,N_12296,N_12246);
nand U12444 (N_12444,N_12355,N_12396);
or U12445 (N_12445,N_12275,N_12320);
nand U12446 (N_12446,N_12336,N_12290);
and U12447 (N_12447,N_12217,N_12295);
or U12448 (N_12448,N_12280,N_12390);
and U12449 (N_12449,N_12265,N_12255);
nor U12450 (N_12450,N_12365,N_12244);
and U12451 (N_12451,N_12287,N_12216);
and U12452 (N_12452,N_12302,N_12360);
and U12453 (N_12453,N_12358,N_12222);
xnor U12454 (N_12454,N_12292,N_12226);
nand U12455 (N_12455,N_12283,N_12227);
nand U12456 (N_12456,N_12387,N_12201);
xnor U12457 (N_12457,N_12374,N_12266);
nor U12458 (N_12458,N_12352,N_12319);
and U12459 (N_12459,N_12229,N_12325);
and U12460 (N_12460,N_12354,N_12361);
nand U12461 (N_12461,N_12379,N_12221);
and U12462 (N_12462,N_12277,N_12367);
or U12463 (N_12463,N_12219,N_12300);
nor U12464 (N_12464,N_12238,N_12329);
nand U12465 (N_12465,N_12393,N_12349);
or U12466 (N_12466,N_12347,N_12268);
xor U12467 (N_12467,N_12281,N_12225);
nor U12468 (N_12468,N_12362,N_12248);
xnor U12469 (N_12469,N_12384,N_12375);
or U12470 (N_12470,N_12261,N_12243);
or U12471 (N_12471,N_12388,N_12330);
and U12472 (N_12472,N_12339,N_12366);
xor U12473 (N_12473,N_12205,N_12316);
nand U12474 (N_12474,N_12237,N_12342);
and U12475 (N_12475,N_12332,N_12353);
and U12476 (N_12476,N_12371,N_12310);
and U12477 (N_12477,N_12279,N_12341);
and U12478 (N_12478,N_12356,N_12321);
or U12479 (N_12479,N_12350,N_12250);
xor U12480 (N_12480,N_12218,N_12215);
or U12481 (N_12481,N_12378,N_12327);
and U12482 (N_12482,N_12382,N_12298);
xor U12483 (N_12483,N_12328,N_12231);
nand U12484 (N_12484,N_12334,N_12306);
nor U12485 (N_12485,N_12241,N_12348);
or U12486 (N_12486,N_12276,N_12258);
xor U12487 (N_12487,N_12208,N_12335);
or U12488 (N_12488,N_12263,N_12303);
and U12489 (N_12489,N_12345,N_12262);
and U12490 (N_12490,N_12257,N_12228);
and U12491 (N_12491,N_12313,N_12307);
nand U12492 (N_12492,N_12314,N_12209);
nand U12493 (N_12493,N_12249,N_12236);
xnor U12494 (N_12494,N_12351,N_12331);
and U12495 (N_12495,N_12245,N_12380);
or U12496 (N_12496,N_12256,N_12363);
nor U12497 (N_12497,N_12239,N_12385);
nor U12498 (N_12498,N_12322,N_12211);
and U12499 (N_12499,N_12220,N_12207);
nand U12500 (N_12500,N_12383,N_12203);
and U12501 (N_12501,N_12294,N_12396);
or U12502 (N_12502,N_12305,N_12280);
nand U12503 (N_12503,N_12371,N_12228);
xor U12504 (N_12504,N_12228,N_12245);
xnor U12505 (N_12505,N_12305,N_12399);
nor U12506 (N_12506,N_12343,N_12282);
nor U12507 (N_12507,N_12375,N_12266);
xnor U12508 (N_12508,N_12330,N_12319);
nor U12509 (N_12509,N_12377,N_12220);
xor U12510 (N_12510,N_12301,N_12204);
or U12511 (N_12511,N_12317,N_12319);
nor U12512 (N_12512,N_12334,N_12239);
xnor U12513 (N_12513,N_12397,N_12271);
nor U12514 (N_12514,N_12258,N_12332);
xor U12515 (N_12515,N_12266,N_12382);
nand U12516 (N_12516,N_12275,N_12235);
nand U12517 (N_12517,N_12320,N_12230);
nand U12518 (N_12518,N_12342,N_12393);
or U12519 (N_12519,N_12325,N_12204);
nand U12520 (N_12520,N_12339,N_12336);
and U12521 (N_12521,N_12364,N_12270);
or U12522 (N_12522,N_12373,N_12219);
or U12523 (N_12523,N_12246,N_12273);
and U12524 (N_12524,N_12258,N_12268);
nand U12525 (N_12525,N_12201,N_12358);
and U12526 (N_12526,N_12329,N_12231);
and U12527 (N_12527,N_12360,N_12371);
nor U12528 (N_12528,N_12378,N_12242);
nor U12529 (N_12529,N_12345,N_12246);
xor U12530 (N_12530,N_12373,N_12276);
nand U12531 (N_12531,N_12207,N_12392);
nand U12532 (N_12532,N_12252,N_12353);
or U12533 (N_12533,N_12340,N_12232);
nor U12534 (N_12534,N_12220,N_12206);
nor U12535 (N_12535,N_12268,N_12270);
nand U12536 (N_12536,N_12310,N_12209);
nand U12537 (N_12537,N_12361,N_12228);
and U12538 (N_12538,N_12351,N_12231);
and U12539 (N_12539,N_12333,N_12382);
xnor U12540 (N_12540,N_12254,N_12329);
and U12541 (N_12541,N_12252,N_12222);
xnor U12542 (N_12542,N_12247,N_12309);
and U12543 (N_12543,N_12339,N_12310);
nand U12544 (N_12544,N_12213,N_12312);
and U12545 (N_12545,N_12241,N_12375);
nor U12546 (N_12546,N_12238,N_12243);
nand U12547 (N_12547,N_12274,N_12390);
and U12548 (N_12548,N_12230,N_12359);
and U12549 (N_12549,N_12298,N_12269);
or U12550 (N_12550,N_12230,N_12286);
nor U12551 (N_12551,N_12212,N_12340);
xor U12552 (N_12552,N_12242,N_12281);
xor U12553 (N_12553,N_12365,N_12302);
and U12554 (N_12554,N_12242,N_12325);
and U12555 (N_12555,N_12248,N_12201);
nand U12556 (N_12556,N_12357,N_12248);
nor U12557 (N_12557,N_12208,N_12368);
nor U12558 (N_12558,N_12358,N_12283);
xnor U12559 (N_12559,N_12259,N_12226);
and U12560 (N_12560,N_12264,N_12267);
and U12561 (N_12561,N_12335,N_12200);
xor U12562 (N_12562,N_12242,N_12322);
and U12563 (N_12563,N_12326,N_12294);
xor U12564 (N_12564,N_12371,N_12248);
nand U12565 (N_12565,N_12203,N_12371);
and U12566 (N_12566,N_12334,N_12216);
nor U12567 (N_12567,N_12252,N_12379);
nor U12568 (N_12568,N_12316,N_12218);
and U12569 (N_12569,N_12389,N_12204);
xor U12570 (N_12570,N_12250,N_12271);
and U12571 (N_12571,N_12343,N_12380);
or U12572 (N_12572,N_12310,N_12295);
and U12573 (N_12573,N_12298,N_12314);
xnor U12574 (N_12574,N_12382,N_12340);
and U12575 (N_12575,N_12368,N_12264);
nor U12576 (N_12576,N_12340,N_12388);
xnor U12577 (N_12577,N_12217,N_12377);
nand U12578 (N_12578,N_12276,N_12308);
xor U12579 (N_12579,N_12275,N_12363);
xor U12580 (N_12580,N_12377,N_12250);
nor U12581 (N_12581,N_12366,N_12320);
xor U12582 (N_12582,N_12316,N_12285);
nand U12583 (N_12583,N_12311,N_12224);
and U12584 (N_12584,N_12385,N_12363);
xor U12585 (N_12585,N_12387,N_12347);
nand U12586 (N_12586,N_12325,N_12368);
and U12587 (N_12587,N_12343,N_12366);
nand U12588 (N_12588,N_12330,N_12295);
and U12589 (N_12589,N_12333,N_12291);
xor U12590 (N_12590,N_12386,N_12272);
or U12591 (N_12591,N_12224,N_12237);
nand U12592 (N_12592,N_12310,N_12375);
or U12593 (N_12593,N_12264,N_12363);
nor U12594 (N_12594,N_12328,N_12324);
or U12595 (N_12595,N_12216,N_12300);
and U12596 (N_12596,N_12353,N_12242);
nor U12597 (N_12597,N_12273,N_12308);
and U12598 (N_12598,N_12381,N_12303);
and U12599 (N_12599,N_12372,N_12306);
nand U12600 (N_12600,N_12495,N_12417);
xor U12601 (N_12601,N_12589,N_12434);
or U12602 (N_12602,N_12583,N_12555);
xor U12603 (N_12603,N_12592,N_12453);
or U12604 (N_12604,N_12430,N_12446);
or U12605 (N_12605,N_12519,N_12467);
xor U12606 (N_12606,N_12455,N_12457);
nand U12607 (N_12607,N_12481,N_12549);
or U12608 (N_12608,N_12415,N_12503);
xnor U12609 (N_12609,N_12498,N_12512);
and U12610 (N_12610,N_12531,N_12480);
and U12611 (N_12611,N_12522,N_12536);
and U12612 (N_12612,N_12471,N_12586);
nor U12613 (N_12613,N_12587,N_12411);
nand U12614 (N_12614,N_12462,N_12575);
and U12615 (N_12615,N_12533,N_12454);
nand U12616 (N_12616,N_12576,N_12568);
nor U12617 (N_12617,N_12598,N_12582);
and U12618 (N_12618,N_12530,N_12410);
nand U12619 (N_12619,N_12593,N_12448);
xnor U12620 (N_12620,N_12511,N_12500);
nor U12621 (N_12621,N_12513,N_12594);
nand U12622 (N_12622,N_12477,N_12432);
or U12623 (N_12623,N_12579,N_12482);
nor U12624 (N_12624,N_12561,N_12558);
nand U12625 (N_12625,N_12479,N_12416);
nand U12626 (N_12626,N_12547,N_12445);
xnor U12627 (N_12627,N_12515,N_12517);
xnor U12628 (N_12628,N_12459,N_12567);
or U12629 (N_12629,N_12418,N_12532);
nand U12630 (N_12630,N_12505,N_12559);
xor U12631 (N_12631,N_12447,N_12550);
nand U12632 (N_12632,N_12553,N_12412);
nor U12633 (N_12633,N_12486,N_12565);
xnor U12634 (N_12634,N_12591,N_12490);
nor U12635 (N_12635,N_12494,N_12421);
or U12636 (N_12636,N_12590,N_12422);
nor U12637 (N_12637,N_12473,N_12507);
and U12638 (N_12638,N_12470,N_12560);
nand U12639 (N_12639,N_12406,N_12580);
or U12640 (N_12640,N_12525,N_12572);
nor U12641 (N_12641,N_12527,N_12543);
nand U12642 (N_12642,N_12508,N_12489);
xor U12643 (N_12643,N_12518,N_12574);
nor U12644 (N_12644,N_12521,N_12557);
nand U12645 (N_12645,N_12440,N_12509);
nor U12646 (N_12646,N_12444,N_12407);
nand U12647 (N_12647,N_12431,N_12595);
and U12648 (N_12648,N_12581,N_12597);
or U12649 (N_12649,N_12475,N_12524);
nor U12650 (N_12650,N_12537,N_12546);
xnor U12651 (N_12651,N_12499,N_12544);
nor U12652 (N_12652,N_12488,N_12469);
and U12653 (N_12653,N_12433,N_12427);
and U12654 (N_12654,N_12452,N_12578);
nand U12655 (N_12655,N_12556,N_12529);
or U12656 (N_12656,N_12449,N_12439);
nand U12657 (N_12657,N_12425,N_12435);
xor U12658 (N_12658,N_12487,N_12424);
or U12659 (N_12659,N_12501,N_12573);
nand U12660 (N_12660,N_12552,N_12483);
and U12661 (N_12661,N_12493,N_12400);
or U12662 (N_12662,N_12441,N_12577);
or U12663 (N_12663,N_12596,N_12484);
and U12664 (N_12664,N_12414,N_12456);
nand U12665 (N_12665,N_12563,N_12588);
nor U12666 (N_12666,N_12570,N_12538);
nand U12667 (N_12667,N_12516,N_12497);
or U12668 (N_12668,N_12485,N_12451);
and U12669 (N_12669,N_12554,N_12474);
and U12670 (N_12670,N_12491,N_12472);
xor U12671 (N_12671,N_12420,N_12535);
nand U12672 (N_12672,N_12403,N_12496);
and U12673 (N_12673,N_12569,N_12514);
nand U12674 (N_12674,N_12436,N_12465);
or U12675 (N_12675,N_12504,N_12478);
xor U12676 (N_12676,N_12426,N_12506);
or U12677 (N_12677,N_12523,N_12401);
nand U12678 (N_12678,N_12534,N_12442);
nand U12679 (N_12679,N_12492,N_12545);
and U12680 (N_12680,N_12409,N_12423);
and U12681 (N_12681,N_12464,N_12428);
or U12682 (N_12682,N_12429,N_12541);
nand U12683 (N_12683,N_12443,N_12461);
or U12684 (N_12684,N_12520,N_12404);
xor U12685 (N_12685,N_12566,N_12438);
nor U12686 (N_12686,N_12468,N_12458);
nor U12687 (N_12687,N_12413,N_12599);
or U12688 (N_12688,N_12510,N_12551);
nor U12689 (N_12689,N_12476,N_12526);
xor U12690 (N_12690,N_12528,N_12460);
xnor U12691 (N_12691,N_12402,N_12540);
xor U12692 (N_12692,N_12408,N_12539);
nand U12693 (N_12693,N_12584,N_12564);
or U12694 (N_12694,N_12405,N_12450);
or U12695 (N_12695,N_12548,N_12463);
and U12696 (N_12696,N_12437,N_12571);
nor U12697 (N_12697,N_12585,N_12502);
nor U12698 (N_12698,N_12419,N_12466);
xnor U12699 (N_12699,N_12542,N_12562);
and U12700 (N_12700,N_12446,N_12475);
nand U12701 (N_12701,N_12538,N_12403);
xnor U12702 (N_12702,N_12499,N_12529);
nand U12703 (N_12703,N_12424,N_12511);
xnor U12704 (N_12704,N_12405,N_12458);
xor U12705 (N_12705,N_12581,N_12589);
nand U12706 (N_12706,N_12525,N_12494);
and U12707 (N_12707,N_12572,N_12589);
nor U12708 (N_12708,N_12595,N_12487);
nand U12709 (N_12709,N_12426,N_12515);
nand U12710 (N_12710,N_12515,N_12585);
nor U12711 (N_12711,N_12511,N_12572);
nand U12712 (N_12712,N_12490,N_12442);
or U12713 (N_12713,N_12414,N_12598);
and U12714 (N_12714,N_12582,N_12443);
and U12715 (N_12715,N_12458,N_12587);
xnor U12716 (N_12716,N_12494,N_12404);
or U12717 (N_12717,N_12405,N_12515);
or U12718 (N_12718,N_12477,N_12574);
xnor U12719 (N_12719,N_12463,N_12542);
nor U12720 (N_12720,N_12538,N_12442);
xnor U12721 (N_12721,N_12593,N_12439);
and U12722 (N_12722,N_12479,N_12553);
and U12723 (N_12723,N_12439,N_12446);
and U12724 (N_12724,N_12509,N_12549);
or U12725 (N_12725,N_12580,N_12534);
xor U12726 (N_12726,N_12538,N_12585);
nand U12727 (N_12727,N_12525,N_12484);
nand U12728 (N_12728,N_12479,N_12411);
xnor U12729 (N_12729,N_12494,N_12532);
or U12730 (N_12730,N_12514,N_12477);
or U12731 (N_12731,N_12591,N_12580);
or U12732 (N_12732,N_12435,N_12499);
xor U12733 (N_12733,N_12445,N_12598);
nor U12734 (N_12734,N_12473,N_12555);
or U12735 (N_12735,N_12422,N_12547);
and U12736 (N_12736,N_12489,N_12456);
xnor U12737 (N_12737,N_12568,N_12400);
or U12738 (N_12738,N_12471,N_12584);
nand U12739 (N_12739,N_12562,N_12512);
and U12740 (N_12740,N_12491,N_12470);
and U12741 (N_12741,N_12524,N_12581);
xor U12742 (N_12742,N_12558,N_12568);
and U12743 (N_12743,N_12437,N_12453);
or U12744 (N_12744,N_12503,N_12437);
and U12745 (N_12745,N_12486,N_12488);
xnor U12746 (N_12746,N_12534,N_12500);
nor U12747 (N_12747,N_12554,N_12502);
and U12748 (N_12748,N_12525,N_12423);
and U12749 (N_12749,N_12575,N_12594);
or U12750 (N_12750,N_12481,N_12509);
and U12751 (N_12751,N_12476,N_12556);
xnor U12752 (N_12752,N_12493,N_12596);
xnor U12753 (N_12753,N_12508,N_12437);
and U12754 (N_12754,N_12533,N_12516);
or U12755 (N_12755,N_12484,N_12569);
and U12756 (N_12756,N_12478,N_12457);
nand U12757 (N_12757,N_12428,N_12570);
nand U12758 (N_12758,N_12494,N_12434);
and U12759 (N_12759,N_12537,N_12455);
or U12760 (N_12760,N_12554,N_12468);
nand U12761 (N_12761,N_12404,N_12469);
and U12762 (N_12762,N_12401,N_12450);
or U12763 (N_12763,N_12578,N_12598);
and U12764 (N_12764,N_12555,N_12411);
or U12765 (N_12765,N_12595,N_12503);
xor U12766 (N_12766,N_12505,N_12574);
and U12767 (N_12767,N_12586,N_12581);
or U12768 (N_12768,N_12522,N_12475);
nor U12769 (N_12769,N_12415,N_12573);
nand U12770 (N_12770,N_12571,N_12486);
and U12771 (N_12771,N_12409,N_12488);
and U12772 (N_12772,N_12474,N_12538);
or U12773 (N_12773,N_12585,N_12495);
and U12774 (N_12774,N_12537,N_12528);
xor U12775 (N_12775,N_12578,N_12402);
xor U12776 (N_12776,N_12416,N_12434);
nand U12777 (N_12777,N_12552,N_12479);
xnor U12778 (N_12778,N_12557,N_12569);
and U12779 (N_12779,N_12425,N_12415);
nand U12780 (N_12780,N_12479,N_12577);
and U12781 (N_12781,N_12565,N_12483);
nand U12782 (N_12782,N_12595,N_12401);
nand U12783 (N_12783,N_12406,N_12400);
nor U12784 (N_12784,N_12525,N_12476);
xnor U12785 (N_12785,N_12558,N_12450);
or U12786 (N_12786,N_12508,N_12507);
or U12787 (N_12787,N_12553,N_12428);
or U12788 (N_12788,N_12452,N_12588);
nand U12789 (N_12789,N_12585,N_12529);
and U12790 (N_12790,N_12520,N_12522);
nor U12791 (N_12791,N_12471,N_12514);
and U12792 (N_12792,N_12565,N_12480);
and U12793 (N_12793,N_12534,N_12493);
xor U12794 (N_12794,N_12551,N_12429);
nand U12795 (N_12795,N_12596,N_12579);
xor U12796 (N_12796,N_12598,N_12403);
or U12797 (N_12797,N_12429,N_12554);
xnor U12798 (N_12798,N_12425,N_12596);
nor U12799 (N_12799,N_12485,N_12548);
nand U12800 (N_12800,N_12623,N_12711);
xor U12801 (N_12801,N_12660,N_12608);
or U12802 (N_12802,N_12609,N_12702);
or U12803 (N_12803,N_12652,N_12676);
and U12804 (N_12804,N_12692,N_12651);
or U12805 (N_12805,N_12749,N_12686);
nor U12806 (N_12806,N_12671,N_12705);
nand U12807 (N_12807,N_12781,N_12699);
nand U12808 (N_12808,N_12739,N_12765);
and U12809 (N_12809,N_12618,N_12738);
nor U12810 (N_12810,N_12703,N_12675);
and U12811 (N_12811,N_12688,N_12669);
xor U12812 (N_12812,N_12714,N_12641);
and U12813 (N_12813,N_12610,N_12744);
nor U12814 (N_12814,N_12691,N_12696);
xnor U12815 (N_12815,N_12764,N_12659);
or U12816 (N_12816,N_12783,N_12758);
xnor U12817 (N_12817,N_12697,N_12681);
nor U12818 (N_12818,N_12616,N_12662);
or U12819 (N_12819,N_12720,N_12753);
nand U12820 (N_12820,N_12730,N_12638);
or U12821 (N_12821,N_12734,N_12663);
nor U12822 (N_12822,N_12726,N_12771);
and U12823 (N_12823,N_12630,N_12622);
nand U12824 (N_12824,N_12754,N_12786);
and U12825 (N_12825,N_12762,N_12644);
xor U12826 (N_12826,N_12679,N_12729);
nand U12827 (N_12827,N_12747,N_12621);
xor U12828 (N_12828,N_12633,N_12721);
xor U12829 (N_12829,N_12724,N_12643);
and U12830 (N_12830,N_12668,N_12784);
nand U12831 (N_12831,N_12656,N_12766);
xor U12832 (N_12832,N_12645,N_12606);
nand U12833 (N_12833,N_12787,N_12603);
or U12834 (N_12834,N_12667,N_12690);
or U12835 (N_12835,N_12627,N_12760);
nand U12836 (N_12836,N_12634,N_12752);
or U12837 (N_12837,N_12664,N_12712);
nor U12838 (N_12838,N_12773,N_12670);
nor U12839 (N_12839,N_12646,N_12731);
or U12840 (N_12840,N_12782,N_12661);
and U12841 (N_12841,N_12612,N_12768);
or U12842 (N_12842,N_12790,N_12629);
and U12843 (N_12843,N_12694,N_12673);
and U12844 (N_12844,N_12698,N_12665);
or U12845 (N_12845,N_12613,N_12789);
nor U12846 (N_12846,N_12687,N_12636);
nand U12847 (N_12847,N_12746,N_12732);
xor U12848 (N_12848,N_12718,N_12793);
or U12849 (N_12849,N_12788,N_12796);
nor U12850 (N_12850,N_12763,N_12683);
nand U12851 (N_12851,N_12778,N_12756);
nor U12852 (N_12852,N_12759,N_12795);
nand U12853 (N_12853,N_12799,N_12740);
and U12854 (N_12854,N_12631,N_12710);
xnor U12855 (N_12855,N_12736,N_12672);
xnor U12856 (N_12856,N_12727,N_12785);
or U12857 (N_12857,N_12625,N_12770);
nand U12858 (N_12858,N_12619,N_12617);
nor U12859 (N_12859,N_12713,N_12745);
nand U12860 (N_12860,N_12715,N_12605);
nor U12861 (N_12861,N_12695,N_12678);
nand U12862 (N_12862,N_12769,N_12742);
and U12863 (N_12863,N_12750,N_12716);
nand U12864 (N_12864,N_12761,N_12751);
xnor U12865 (N_12865,N_12626,N_12655);
xnor U12866 (N_12866,N_12743,N_12735);
nand U12867 (N_12867,N_12653,N_12684);
or U12868 (N_12868,N_12654,N_12658);
xnor U12869 (N_12869,N_12757,N_12649);
xor U12870 (N_12870,N_12722,N_12737);
nand U12871 (N_12871,N_12647,N_12741);
or U12872 (N_12872,N_12728,N_12682);
or U12873 (N_12873,N_12719,N_12704);
or U12874 (N_12874,N_12689,N_12725);
or U12875 (N_12875,N_12637,N_12639);
nor U12876 (N_12876,N_12604,N_12693);
or U12877 (N_12877,N_12642,N_12797);
nor U12878 (N_12878,N_12708,N_12680);
nand U12879 (N_12879,N_12707,N_12615);
nor U12880 (N_12880,N_12794,N_12772);
and U12881 (N_12881,N_12706,N_12709);
xnor U12882 (N_12882,N_12767,N_12776);
xnor U12883 (N_12883,N_12620,N_12777);
or U12884 (N_12884,N_12632,N_12601);
nand U12885 (N_12885,N_12780,N_12701);
nand U12886 (N_12886,N_12640,N_12685);
and U12887 (N_12887,N_12624,N_12628);
xnor U12888 (N_12888,N_12635,N_12733);
nor U12889 (N_12889,N_12674,N_12717);
xor U12890 (N_12890,N_12700,N_12607);
and U12891 (N_12891,N_12611,N_12779);
or U12892 (N_12892,N_12723,N_12748);
nand U12893 (N_12893,N_12775,N_12677);
nand U12894 (N_12894,N_12792,N_12798);
xor U12895 (N_12895,N_12614,N_12666);
or U12896 (N_12896,N_12755,N_12648);
nor U12897 (N_12897,N_12774,N_12602);
nand U12898 (N_12898,N_12600,N_12791);
and U12899 (N_12899,N_12650,N_12657);
nand U12900 (N_12900,N_12778,N_12624);
xnor U12901 (N_12901,N_12785,N_12678);
nand U12902 (N_12902,N_12706,N_12788);
nor U12903 (N_12903,N_12772,N_12651);
and U12904 (N_12904,N_12717,N_12629);
and U12905 (N_12905,N_12667,N_12701);
or U12906 (N_12906,N_12749,N_12766);
nand U12907 (N_12907,N_12787,N_12774);
nor U12908 (N_12908,N_12663,N_12646);
or U12909 (N_12909,N_12735,N_12625);
nand U12910 (N_12910,N_12752,N_12725);
nand U12911 (N_12911,N_12798,N_12610);
nand U12912 (N_12912,N_12705,N_12746);
xnor U12913 (N_12913,N_12610,N_12708);
and U12914 (N_12914,N_12796,N_12751);
or U12915 (N_12915,N_12645,N_12777);
and U12916 (N_12916,N_12751,N_12747);
and U12917 (N_12917,N_12686,N_12631);
xor U12918 (N_12918,N_12701,N_12651);
nor U12919 (N_12919,N_12747,N_12682);
and U12920 (N_12920,N_12668,N_12747);
and U12921 (N_12921,N_12716,N_12696);
nand U12922 (N_12922,N_12777,N_12785);
nand U12923 (N_12923,N_12722,N_12602);
or U12924 (N_12924,N_12780,N_12790);
xor U12925 (N_12925,N_12773,N_12647);
or U12926 (N_12926,N_12605,N_12690);
xor U12927 (N_12927,N_12720,N_12771);
and U12928 (N_12928,N_12694,N_12612);
xnor U12929 (N_12929,N_12766,N_12623);
nand U12930 (N_12930,N_12719,N_12610);
or U12931 (N_12931,N_12764,N_12634);
nor U12932 (N_12932,N_12646,N_12620);
xnor U12933 (N_12933,N_12785,N_12660);
xor U12934 (N_12934,N_12755,N_12638);
xnor U12935 (N_12935,N_12635,N_12688);
xnor U12936 (N_12936,N_12606,N_12760);
nand U12937 (N_12937,N_12672,N_12693);
nand U12938 (N_12938,N_12776,N_12651);
xor U12939 (N_12939,N_12735,N_12704);
or U12940 (N_12940,N_12691,N_12624);
and U12941 (N_12941,N_12769,N_12733);
or U12942 (N_12942,N_12727,N_12756);
nor U12943 (N_12943,N_12678,N_12697);
or U12944 (N_12944,N_12635,N_12780);
xnor U12945 (N_12945,N_12759,N_12753);
nor U12946 (N_12946,N_12735,N_12646);
xnor U12947 (N_12947,N_12617,N_12782);
or U12948 (N_12948,N_12734,N_12626);
or U12949 (N_12949,N_12788,N_12717);
nand U12950 (N_12950,N_12644,N_12648);
and U12951 (N_12951,N_12665,N_12756);
or U12952 (N_12952,N_12720,N_12743);
nand U12953 (N_12953,N_12684,N_12739);
or U12954 (N_12954,N_12742,N_12648);
and U12955 (N_12955,N_12692,N_12670);
xnor U12956 (N_12956,N_12612,N_12611);
and U12957 (N_12957,N_12781,N_12619);
xnor U12958 (N_12958,N_12610,N_12784);
nand U12959 (N_12959,N_12776,N_12744);
nand U12960 (N_12960,N_12700,N_12671);
nand U12961 (N_12961,N_12653,N_12654);
nor U12962 (N_12962,N_12764,N_12775);
nand U12963 (N_12963,N_12632,N_12664);
nor U12964 (N_12964,N_12698,N_12713);
nor U12965 (N_12965,N_12761,N_12727);
nor U12966 (N_12966,N_12737,N_12690);
or U12967 (N_12967,N_12735,N_12623);
or U12968 (N_12968,N_12714,N_12742);
or U12969 (N_12969,N_12784,N_12741);
nand U12970 (N_12970,N_12769,N_12653);
and U12971 (N_12971,N_12742,N_12726);
xor U12972 (N_12972,N_12716,N_12743);
nand U12973 (N_12973,N_12715,N_12613);
and U12974 (N_12974,N_12673,N_12665);
xnor U12975 (N_12975,N_12738,N_12619);
and U12976 (N_12976,N_12773,N_12649);
xnor U12977 (N_12977,N_12645,N_12770);
nand U12978 (N_12978,N_12791,N_12740);
and U12979 (N_12979,N_12670,N_12777);
nand U12980 (N_12980,N_12678,N_12659);
and U12981 (N_12981,N_12620,N_12763);
xor U12982 (N_12982,N_12635,N_12615);
nor U12983 (N_12983,N_12734,N_12792);
nor U12984 (N_12984,N_12786,N_12678);
and U12985 (N_12985,N_12635,N_12679);
and U12986 (N_12986,N_12797,N_12610);
nor U12987 (N_12987,N_12628,N_12724);
nor U12988 (N_12988,N_12722,N_12612);
or U12989 (N_12989,N_12600,N_12719);
xor U12990 (N_12990,N_12631,N_12717);
nor U12991 (N_12991,N_12630,N_12631);
and U12992 (N_12992,N_12751,N_12703);
and U12993 (N_12993,N_12774,N_12781);
nand U12994 (N_12994,N_12796,N_12724);
xor U12995 (N_12995,N_12695,N_12611);
nand U12996 (N_12996,N_12606,N_12799);
and U12997 (N_12997,N_12771,N_12609);
nand U12998 (N_12998,N_12613,N_12721);
nand U12999 (N_12999,N_12706,N_12732);
and U13000 (N_13000,N_12917,N_12934);
and U13001 (N_13001,N_12842,N_12984);
nor U13002 (N_13002,N_12849,N_12838);
xnor U13003 (N_13003,N_12806,N_12811);
nor U13004 (N_13004,N_12906,N_12879);
xor U13005 (N_13005,N_12922,N_12882);
nor U13006 (N_13006,N_12877,N_12981);
xnor U13007 (N_13007,N_12946,N_12897);
nor U13008 (N_13008,N_12825,N_12937);
and U13009 (N_13009,N_12830,N_12943);
and U13010 (N_13010,N_12927,N_12935);
nand U13011 (N_13011,N_12853,N_12965);
or U13012 (N_13012,N_12858,N_12973);
nand U13013 (N_13013,N_12878,N_12868);
and U13014 (N_13014,N_12862,N_12867);
nor U13015 (N_13015,N_12885,N_12861);
nor U13016 (N_13016,N_12963,N_12987);
nor U13017 (N_13017,N_12964,N_12971);
nor U13018 (N_13018,N_12813,N_12953);
and U13019 (N_13019,N_12938,N_12900);
or U13020 (N_13020,N_12968,N_12939);
or U13021 (N_13021,N_12857,N_12915);
nand U13022 (N_13022,N_12816,N_12910);
nor U13023 (N_13023,N_12911,N_12957);
xor U13024 (N_13024,N_12855,N_12810);
and U13025 (N_13025,N_12817,N_12818);
nor U13026 (N_13026,N_12933,N_12836);
or U13027 (N_13027,N_12977,N_12989);
or U13028 (N_13028,N_12932,N_12834);
or U13029 (N_13029,N_12902,N_12908);
xnor U13030 (N_13030,N_12936,N_12831);
and U13031 (N_13031,N_12876,N_12966);
and U13032 (N_13032,N_12873,N_12845);
nand U13033 (N_13033,N_12829,N_12851);
xor U13034 (N_13034,N_12999,N_12983);
nand U13035 (N_13035,N_12924,N_12837);
or U13036 (N_13036,N_12846,N_12998);
nor U13037 (N_13037,N_12950,N_12880);
xnor U13038 (N_13038,N_12992,N_12931);
xor U13039 (N_13039,N_12852,N_12928);
or U13040 (N_13040,N_12925,N_12930);
or U13041 (N_13041,N_12812,N_12870);
nor U13042 (N_13042,N_12832,N_12843);
and U13043 (N_13043,N_12912,N_12982);
xor U13044 (N_13044,N_12893,N_12823);
and U13045 (N_13045,N_12909,N_12800);
or U13046 (N_13046,N_12884,N_12828);
xor U13047 (N_13047,N_12865,N_12951);
xnor U13048 (N_13048,N_12920,N_12807);
xnor U13049 (N_13049,N_12821,N_12994);
or U13050 (N_13050,N_12955,N_12802);
xnor U13051 (N_13051,N_12926,N_12850);
xor U13052 (N_13052,N_12907,N_12972);
xor U13053 (N_13053,N_12859,N_12889);
or U13054 (N_13054,N_12975,N_12980);
or U13055 (N_13055,N_12803,N_12895);
or U13056 (N_13056,N_12919,N_12967);
nor U13057 (N_13057,N_12847,N_12904);
xnor U13058 (N_13058,N_12815,N_12929);
and U13059 (N_13059,N_12949,N_12947);
xnor U13060 (N_13060,N_12988,N_12854);
and U13061 (N_13061,N_12901,N_12974);
nand U13062 (N_13062,N_12962,N_12995);
xnor U13063 (N_13063,N_12945,N_12820);
nand U13064 (N_13064,N_12941,N_12986);
nand U13065 (N_13065,N_12991,N_12864);
nand U13066 (N_13066,N_12863,N_12819);
xor U13067 (N_13067,N_12990,N_12805);
and U13068 (N_13068,N_12948,N_12954);
nand U13069 (N_13069,N_12894,N_12886);
nand U13070 (N_13070,N_12916,N_12979);
or U13071 (N_13071,N_12905,N_12835);
nor U13072 (N_13072,N_12961,N_12942);
xor U13073 (N_13073,N_12869,N_12969);
or U13074 (N_13074,N_12860,N_12890);
xor U13075 (N_13075,N_12956,N_12918);
or U13076 (N_13076,N_12952,N_12898);
or U13077 (N_13077,N_12944,N_12826);
or U13078 (N_13078,N_12940,N_12913);
xnor U13079 (N_13079,N_12978,N_12814);
nand U13080 (N_13080,N_12899,N_12844);
or U13081 (N_13081,N_12833,N_12993);
nand U13082 (N_13082,N_12856,N_12887);
nand U13083 (N_13083,N_12839,N_12866);
or U13084 (N_13084,N_12801,N_12840);
and U13085 (N_13085,N_12914,N_12841);
or U13086 (N_13086,N_12921,N_12804);
nor U13087 (N_13087,N_12996,N_12960);
xnor U13088 (N_13088,N_12883,N_12923);
and U13089 (N_13089,N_12848,N_12891);
nor U13090 (N_13090,N_12872,N_12824);
nor U13091 (N_13091,N_12827,N_12896);
nand U13092 (N_13092,N_12985,N_12809);
and U13093 (N_13093,N_12958,N_12888);
nand U13094 (N_13094,N_12874,N_12808);
nand U13095 (N_13095,N_12997,N_12881);
xor U13096 (N_13096,N_12976,N_12822);
nand U13097 (N_13097,N_12970,N_12903);
nand U13098 (N_13098,N_12871,N_12875);
or U13099 (N_13099,N_12959,N_12892);
or U13100 (N_13100,N_12862,N_12991);
xor U13101 (N_13101,N_12828,N_12944);
and U13102 (N_13102,N_12950,N_12828);
xnor U13103 (N_13103,N_12952,N_12802);
and U13104 (N_13104,N_12951,N_12915);
xor U13105 (N_13105,N_12813,N_12902);
nor U13106 (N_13106,N_12825,N_12972);
nor U13107 (N_13107,N_12832,N_12862);
nand U13108 (N_13108,N_12962,N_12812);
and U13109 (N_13109,N_12978,N_12897);
nor U13110 (N_13110,N_12995,N_12985);
xor U13111 (N_13111,N_12910,N_12866);
or U13112 (N_13112,N_12999,N_12946);
nor U13113 (N_13113,N_12984,N_12854);
nor U13114 (N_13114,N_12885,N_12963);
xor U13115 (N_13115,N_12907,N_12911);
nand U13116 (N_13116,N_12986,N_12853);
or U13117 (N_13117,N_12810,N_12944);
nand U13118 (N_13118,N_12804,N_12910);
and U13119 (N_13119,N_12923,N_12965);
xor U13120 (N_13120,N_12923,N_12945);
xor U13121 (N_13121,N_12931,N_12878);
nand U13122 (N_13122,N_12861,N_12896);
nand U13123 (N_13123,N_12887,N_12820);
or U13124 (N_13124,N_12857,N_12886);
xnor U13125 (N_13125,N_12825,N_12836);
xor U13126 (N_13126,N_12959,N_12945);
nand U13127 (N_13127,N_12953,N_12965);
and U13128 (N_13128,N_12933,N_12893);
nor U13129 (N_13129,N_12969,N_12976);
and U13130 (N_13130,N_12969,N_12901);
nor U13131 (N_13131,N_12880,N_12970);
and U13132 (N_13132,N_12830,N_12855);
nor U13133 (N_13133,N_12960,N_12894);
nand U13134 (N_13134,N_12894,N_12904);
xnor U13135 (N_13135,N_12939,N_12812);
xor U13136 (N_13136,N_12969,N_12837);
or U13137 (N_13137,N_12823,N_12979);
nor U13138 (N_13138,N_12847,N_12976);
or U13139 (N_13139,N_12829,N_12813);
xnor U13140 (N_13140,N_12857,N_12948);
and U13141 (N_13141,N_12932,N_12808);
or U13142 (N_13142,N_12806,N_12961);
xor U13143 (N_13143,N_12818,N_12919);
and U13144 (N_13144,N_12823,N_12940);
and U13145 (N_13145,N_12993,N_12801);
xor U13146 (N_13146,N_12854,N_12941);
or U13147 (N_13147,N_12818,N_12987);
xnor U13148 (N_13148,N_12906,N_12825);
and U13149 (N_13149,N_12801,N_12988);
and U13150 (N_13150,N_12952,N_12970);
and U13151 (N_13151,N_12858,N_12835);
nand U13152 (N_13152,N_12840,N_12966);
xnor U13153 (N_13153,N_12963,N_12865);
nor U13154 (N_13154,N_12901,N_12817);
and U13155 (N_13155,N_12872,N_12840);
nor U13156 (N_13156,N_12948,N_12961);
nor U13157 (N_13157,N_12931,N_12999);
and U13158 (N_13158,N_12874,N_12883);
nor U13159 (N_13159,N_12982,N_12871);
xnor U13160 (N_13160,N_12827,N_12937);
and U13161 (N_13161,N_12977,N_12887);
or U13162 (N_13162,N_12869,N_12845);
nor U13163 (N_13163,N_12934,N_12945);
xnor U13164 (N_13164,N_12885,N_12933);
nor U13165 (N_13165,N_12882,N_12985);
and U13166 (N_13166,N_12874,N_12924);
nand U13167 (N_13167,N_12974,N_12903);
or U13168 (N_13168,N_12928,N_12870);
and U13169 (N_13169,N_12886,N_12929);
or U13170 (N_13170,N_12935,N_12863);
or U13171 (N_13171,N_12855,N_12864);
nand U13172 (N_13172,N_12821,N_12804);
and U13173 (N_13173,N_12971,N_12954);
xnor U13174 (N_13174,N_12932,N_12924);
nand U13175 (N_13175,N_12954,N_12950);
nor U13176 (N_13176,N_12918,N_12834);
nand U13177 (N_13177,N_12880,N_12951);
nor U13178 (N_13178,N_12855,N_12965);
nor U13179 (N_13179,N_12839,N_12816);
nand U13180 (N_13180,N_12922,N_12841);
xnor U13181 (N_13181,N_12969,N_12927);
or U13182 (N_13182,N_12870,N_12847);
nand U13183 (N_13183,N_12817,N_12826);
nand U13184 (N_13184,N_12848,N_12980);
xnor U13185 (N_13185,N_12857,N_12847);
nor U13186 (N_13186,N_12986,N_12887);
and U13187 (N_13187,N_12890,N_12855);
nand U13188 (N_13188,N_12950,N_12854);
or U13189 (N_13189,N_12850,N_12934);
nand U13190 (N_13190,N_12959,N_12987);
nand U13191 (N_13191,N_12800,N_12826);
xor U13192 (N_13192,N_12934,N_12860);
nor U13193 (N_13193,N_12903,N_12845);
nor U13194 (N_13194,N_12970,N_12979);
nand U13195 (N_13195,N_12809,N_12955);
or U13196 (N_13196,N_12990,N_12960);
or U13197 (N_13197,N_12911,N_12952);
nor U13198 (N_13198,N_12827,N_12872);
or U13199 (N_13199,N_12825,N_12993);
nor U13200 (N_13200,N_13174,N_13152);
nor U13201 (N_13201,N_13017,N_13082);
xor U13202 (N_13202,N_13184,N_13068);
and U13203 (N_13203,N_13144,N_13097);
nor U13204 (N_13204,N_13000,N_13065);
and U13205 (N_13205,N_13071,N_13064);
xor U13206 (N_13206,N_13126,N_13104);
and U13207 (N_13207,N_13128,N_13175);
nor U13208 (N_13208,N_13042,N_13046);
or U13209 (N_13209,N_13167,N_13086);
xor U13210 (N_13210,N_13194,N_13037);
or U13211 (N_13211,N_13093,N_13009);
nand U13212 (N_13212,N_13157,N_13185);
nand U13213 (N_13213,N_13051,N_13008);
xnor U13214 (N_13214,N_13183,N_13199);
nand U13215 (N_13215,N_13039,N_13127);
nor U13216 (N_13216,N_13111,N_13158);
or U13217 (N_13217,N_13117,N_13058);
nor U13218 (N_13218,N_13193,N_13196);
xor U13219 (N_13219,N_13024,N_13136);
and U13220 (N_13220,N_13055,N_13066);
or U13221 (N_13221,N_13029,N_13160);
xor U13222 (N_13222,N_13062,N_13176);
nand U13223 (N_13223,N_13163,N_13032);
xor U13224 (N_13224,N_13074,N_13133);
nand U13225 (N_13225,N_13145,N_13018);
xnor U13226 (N_13226,N_13069,N_13125);
and U13227 (N_13227,N_13143,N_13007);
nand U13228 (N_13228,N_13028,N_13181);
or U13229 (N_13229,N_13186,N_13169);
xnor U13230 (N_13230,N_13159,N_13070);
nand U13231 (N_13231,N_13197,N_13044);
or U13232 (N_13232,N_13122,N_13001);
nor U13233 (N_13233,N_13013,N_13146);
xor U13234 (N_13234,N_13166,N_13137);
or U13235 (N_13235,N_13049,N_13191);
xnor U13236 (N_13236,N_13002,N_13150);
and U13237 (N_13237,N_13130,N_13182);
or U13238 (N_13238,N_13105,N_13102);
nand U13239 (N_13239,N_13079,N_13112);
or U13240 (N_13240,N_13192,N_13005);
or U13241 (N_13241,N_13045,N_13020);
nor U13242 (N_13242,N_13003,N_13031);
nand U13243 (N_13243,N_13010,N_13121);
and U13244 (N_13244,N_13006,N_13048);
xnor U13245 (N_13245,N_13047,N_13161);
or U13246 (N_13246,N_13014,N_13187);
xor U13247 (N_13247,N_13188,N_13141);
and U13248 (N_13248,N_13153,N_13113);
xor U13249 (N_13249,N_13178,N_13059);
nand U13250 (N_13250,N_13078,N_13076);
and U13251 (N_13251,N_13073,N_13142);
nor U13252 (N_13252,N_13151,N_13107);
and U13253 (N_13253,N_13004,N_13131);
and U13254 (N_13254,N_13081,N_13095);
and U13255 (N_13255,N_13094,N_13114);
or U13256 (N_13256,N_13154,N_13057);
and U13257 (N_13257,N_13156,N_13147);
nor U13258 (N_13258,N_13092,N_13067);
or U13259 (N_13259,N_13036,N_13135);
or U13260 (N_13260,N_13180,N_13026);
xor U13261 (N_13261,N_13129,N_13019);
or U13262 (N_13262,N_13155,N_13162);
xor U13263 (N_13263,N_13021,N_13139);
nor U13264 (N_13264,N_13088,N_13172);
nor U13265 (N_13265,N_13030,N_13043);
or U13266 (N_13266,N_13116,N_13165);
xnor U13267 (N_13267,N_13179,N_13110);
nor U13268 (N_13268,N_13189,N_13138);
nand U13269 (N_13269,N_13011,N_13106);
and U13270 (N_13270,N_13164,N_13115);
or U13271 (N_13271,N_13089,N_13075);
or U13272 (N_13272,N_13050,N_13091);
nand U13273 (N_13273,N_13103,N_13099);
or U13274 (N_13274,N_13177,N_13118);
nor U13275 (N_13275,N_13173,N_13056);
nand U13276 (N_13276,N_13060,N_13038);
and U13277 (N_13277,N_13054,N_13134);
xnor U13278 (N_13278,N_13016,N_13080);
xnor U13279 (N_13279,N_13090,N_13084);
xnor U13280 (N_13280,N_13170,N_13072);
and U13281 (N_13281,N_13195,N_13101);
nor U13282 (N_13282,N_13040,N_13149);
nor U13283 (N_13283,N_13015,N_13140);
or U13284 (N_13284,N_13085,N_13096);
nand U13285 (N_13285,N_13063,N_13132);
nand U13286 (N_13286,N_13012,N_13022);
xor U13287 (N_13287,N_13198,N_13120);
or U13288 (N_13288,N_13190,N_13035);
and U13289 (N_13289,N_13171,N_13027);
xor U13290 (N_13290,N_13025,N_13168);
and U13291 (N_13291,N_13109,N_13100);
and U13292 (N_13292,N_13123,N_13098);
xor U13293 (N_13293,N_13053,N_13023);
nand U13294 (N_13294,N_13077,N_13124);
or U13295 (N_13295,N_13148,N_13041);
nand U13296 (N_13296,N_13061,N_13033);
xor U13297 (N_13297,N_13087,N_13052);
nand U13298 (N_13298,N_13083,N_13108);
or U13299 (N_13299,N_13034,N_13119);
nand U13300 (N_13300,N_13064,N_13123);
nand U13301 (N_13301,N_13103,N_13045);
nor U13302 (N_13302,N_13075,N_13170);
xnor U13303 (N_13303,N_13175,N_13033);
and U13304 (N_13304,N_13031,N_13153);
or U13305 (N_13305,N_13003,N_13113);
xor U13306 (N_13306,N_13151,N_13095);
xnor U13307 (N_13307,N_13128,N_13056);
nor U13308 (N_13308,N_13171,N_13142);
xor U13309 (N_13309,N_13170,N_13049);
nand U13310 (N_13310,N_13132,N_13133);
and U13311 (N_13311,N_13033,N_13139);
xor U13312 (N_13312,N_13002,N_13027);
and U13313 (N_13313,N_13150,N_13196);
or U13314 (N_13314,N_13168,N_13038);
nand U13315 (N_13315,N_13127,N_13033);
and U13316 (N_13316,N_13008,N_13125);
and U13317 (N_13317,N_13024,N_13194);
nor U13318 (N_13318,N_13093,N_13056);
nor U13319 (N_13319,N_13146,N_13066);
nor U13320 (N_13320,N_13154,N_13112);
nand U13321 (N_13321,N_13089,N_13185);
and U13322 (N_13322,N_13145,N_13093);
or U13323 (N_13323,N_13080,N_13131);
xnor U13324 (N_13324,N_13074,N_13143);
or U13325 (N_13325,N_13103,N_13143);
nor U13326 (N_13326,N_13100,N_13179);
nor U13327 (N_13327,N_13068,N_13070);
xor U13328 (N_13328,N_13102,N_13159);
and U13329 (N_13329,N_13040,N_13194);
xor U13330 (N_13330,N_13187,N_13144);
xnor U13331 (N_13331,N_13173,N_13086);
and U13332 (N_13332,N_13016,N_13122);
and U13333 (N_13333,N_13168,N_13075);
or U13334 (N_13334,N_13000,N_13088);
and U13335 (N_13335,N_13174,N_13150);
nand U13336 (N_13336,N_13012,N_13197);
nand U13337 (N_13337,N_13111,N_13173);
nor U13338 (N_13338,N_13195,N_13055);
or U13339 (N_13339,N_13183,N_13121);
and U13340 (N_13340,N_13079,N_13083);
nand U13341 (N_13341,N_13126,N_13144);
xnor U13342 (N_13342,N_13094,N_13018);
nor U13343 (N_13343,N_13144,N_13153);
xnor U13344 (N_13344,N_13049,N_13169);
nand U13345 (N_13345,N_13007,N_13156);
nand U13346 (N_13346,N_13183,N_13093);
nor U13347 (N_13347,N_13113,N_13163);
xor U13348 (N_13348,N_13026,N_13120);
and U13349 (N_13349,N_13033,N_13120);
and U13350 (N_13350,N_13161,N_13146);
nor U13351 (N_13351,N_13108,N_13145);
or U13352 (N_13352,N_13144,N_13074);
nor U13353 (N_13353,N_13082,N_13006);
nor U13354 (N_13354,N_13094,N_13106);
nor U13355 (N_13355,N_13102,N_13158);
nand U13356 (N_13356,N_13140,N_13021);
xor U13357 (N_13357,N_13146,N_13072);
nand U13358 (N_13358,N_13187,N_13129);
or U13359 (N_13359,N_13000,N_13077);
nand U13360 (N_13360,N_13165,N_13040);
nor U13361 (N_13361,N_13166,N_13144);
xor U13362 (N_13362,N_13081,N_13184);
or U13363 (N_13363,N_13158,N_13021);
or U13364 (N_13364,N_13078,N_13137);
or U13365 (N_13365,N_13131,N_13181);
or U13366 (N_13366,N_13164,N_13180);
and U13367 (N_13367,N_13136,N_13177);
nor U13368 (N_13368,N_13087,N_13018);
nor U13369 (N_13369,N_13081,N_13157);
nor U13370 (N_13370,N_13120,N_13132);
nor U13371 (N_13371,N_13093,N_13136);
nor U13372 (N_13372,N_13058,N_13160);
nand U13373 (N_13373,N_13049,N_13099);
nor U13374 (N_13374,N_13033,N_13135);
xor U13375 (N_13375,N_13046,N_13032);
or U13376 (N_13376,N_13129,N_13057);
nor U13377 (N_13377,N_13143,N_13193);
and U13378 (N_13378,N_13009,N_13131);
xor U13379 (N_13379,N_13075,N_13107);
nand U13380 (N_13380,N_13167,N_13011);
or U13381 (N_13381,N_13134,N_13152);
and U13382 (N_13382,N_13009,N_13003);
nand U13383 (N_13383,N_13007,N_13040);
xnor U13384 (N_13384,N_13022,N_13066);
and U13385 (N_13385,N_13167,N_13038);
nor U13386 (N_13386,N_13123,N_13031);
nand U13387 (N_13387,N_13157,N_13084);
or U13388 (N_13388,N_13104,N_13058);
nand U13389 (N_13389,N_13019,N_13156);
and U13390 (N_13390,N_13093,N_13137);
or U13391 (N_13391,N_13165,N_13161);
or U13392 (N_13392,N_13188,N_13111);
and U13393 (N_13393,N_13154,N_13099);
and U13394 (N_13394,N_13114,N_13196);
or U13395 (N_13395,N_13097,N_13189);
and U13396 (N_13396,N_13199,N_13170);
or U13397 (N_13397,N_13119,N_13072);
xor U13398 (N_13398,N_13118,N_13182);
and U13399 (N_13399,N_13034,N_13120);
nor U13400 (N_13400,N_13251,N_13224);
xnor U13401 (N_13401,N_13351,N_13205);
and U13402 (N_13402,N_13294,N_13382);
and U13403 (N_13403,N_13259,N_13365);
or U13404 (N_13404,N_13336,N_13341);
or U13405 (N_13405,N_13238,N_13300);
and U13406 (N_13406,N_13318,N_13323);
nand U13407 (N_13407,N_13279,N_13357);
nand U13408 (N_13408,N_13248,N_13376);
and U13409 (N_13409,N_13330,N_13317);
nand U13410 (N_13410,N_13230,N_13389);
xnor U13411 (N_13411,N_13367,N_13210);
or U13412 (N_13412,N_13354,N_13355);
and U13413 (N_13413,N_13260,N_13301);
or U13414 (N_13414,N_13325,N_13392);
nand U13415 (N_13415,N_13332,N_13227);
or U13416 (N_13416,N_13287,N_13253);
or U13417 (N_13417,N_13377,N_13207);
and U13418 (N_13418,N_13397,N_13274);
nand U13419 (N_13419,N_13211,N_13373);
nor U13420 (N_13420,N_13209,N_13304);
xor U13421 (N_13421,N_13270,N_13237);
nand U13422 (N_13422,N_13374,N_13347);
xnor U13423 (N_13423,N_13228,N_13222);
nand U13424 (N_13424,N_13288,N_13327);
and U13425 (N_13425,N_13329,N_13358);
or U13426 (N_13426,N_13362,N_13225);
nand U13427 (N_13427,N_13298,N_13240);
xnor U13428 (N_13428,N_13242,N_13349);
or U13429 (N_13429,N_13277,N_13396);
and U13430 (N_13430,N_13213,N_13223);
nand U13431 (N_13431,N_13345,N_13245);
and U13432 (N_13432,N_13276,N_13252);
or U13433 (N_13433,N_13200,N_13352);
nor U13434 (N_13434,N_13201,N_13388);
and U13435 (N_13435,N_13278,N_13387);
nor U13436 (N_13436,N_13319,N_13284);
or U13437 (N_13437,N_13293,N_13218);
xnor U13438 (N_13438,N_13206,N_13380);
and U13439 (N_13439,N_13333,N_13316);
nor U13440 (N_13440,N_13283,N_13232);
nand U13441 (N_13441,N_13220,N_13226);
xnor U13442 (N_13442,N_13309,N_13335);
and U13443 (N_13443,N_13272,N_13350);
and U13444 (N_13444,N_13202,N_13348);
nor U13445 (N_13445,N_13363,N_13398);
or U13446 (N_13446,N_13322,N_13372);
nor U13447 (N_13447,N_13315,N_13337);
and U13448 (N_13448,N_13244,N_13215);
and U13449 (N_13449,N_13399,N_13368);
and U13450 (N_13450,N_13250,N_13343);
nor U13451 (N_13451,N_13204,N_13370);
xor U13452 (N_13452,N_13271,N_13360);
and U13453 (N_13453,N_13263,N_13385);
nor U13454 (N_13454,N_13346,N_13353);
nand U13455 (N_13455,N_13262,N_13203);
nand U13456 (N_13456,N_13395,N_13269);
or U13457 (N_13457,N_13375,N_13312);
or U13458 (N_13458,N_13306,N_13378);
nor U13459 (N_13459,N_13321,N_13391);
nand U13460 (N_13460,N_13291,N_13273);
xnor U13461 (N_13461,N_13221,N_13390);
nor U13462 (N_13462,N_13310,N_13292);
and U13463 (N_13463,N_13265,N_13261);
and U13464 (N_13464,N_13383,N_13303);
or U13465 (N_13465,N_13246,N_13249);
xor U13466 (N_13466,N_13281,N_13256);
and U13467 (N_13467,N_13361,N_13216);
nor U13468 (N_13468,N_13324,N_13264);
nand U13469 (N_13469,N_13320,N_13296);
xor U13470 (N_13470,N_13254,N_13289);
or U13471 (N_13471,N_13231,N_13299);
nand U13472 (N_13472,N_13234,N_13229);
nand U13473 (N_13473,N_13290,N_13359);
nand U13474 (N_13474,N_13295,N_13338);
nor U13475 (N_13475,N_13371,N_13313);
xor U13476 (N_13476,N_13258,N_13255);
xor U13477 (N_13477,N_13302,N_13308);
nand U13478 (N_13478,N_13305,N_13340);
nor U13479 (N_13479,N_13339,N_13394);
nand U13480 (N_13480,N_13267,N_13369);
and U13481 (N_13481,N_13356,N_13241);
xor U13482 (N_13482,N_13236,N_13286);
and U13483 (N_13483,N_13280,N_13393);
xnor U13484 (N_13484,N_13235,N_13257);
nor U13485 (N_13485,N_13331,N_13282);
nor U13486 (N_13486,N_13334,N_13311);
xnor U13487 (N_13487,N_13268,N_13239);
xnor U13488 (N_13488,N_13344,N_13342);
xnor U13489 (N_13489,N_13364,N_13243);
and U13490 (N_13490,N_13285,N_13326);
and U13491 (N_13491,N_13307,N_13328);
nor U13492 (N_13492,N_13386,N_13219);
nand U13493 (N_13493,N_13214,N_13297);
and U13494 (N_13494,N_13379,N_13384);
nand U13495 (N_13495,N_13208,N_13212);
or U13496 (N_13496,N_13366,N_13217);
xor U13497 (N_13497,N_13233,N_13314);
nand U13498 (N_13498,N_13247,N_13381);
xor U13499 (N_13499,N_13266,N_13275);
xnor U13500 (N_13500,N_13391,N_13224);
and U13501 (N_13501,N_13273,N_13220);
nand U13502 (N_13502,N_13308,N_13211);
or U13503 (N_13503,N_13354,N_13344);
xor U13504 (N_13504,N_13343,N_13302);
and U13505 (N_13505,N_13290,N_13241);
and U13506 (N_13506,N_13207,N_13366);
nor U13507 (N_13507,N_13221,N_13212);
or U13508 (N_13508,N_13207,N_13356);
nor U13509 (N_13509,N_13346,N_13255);
or U13510 (N_13510,N_13275,N_13237);
nand U13511 (N_13511,N_13340,N_13375);
nor U13512 (N_13512,N_13302,N_13233);
or U13513 (N_13513,N_13213,N_13225);
nand U13514 (N_13514,N_13287,N_13275);
or U13515 (N_13515,N_13309,N_13378);
nand U13516 (N_13516,N_13287,N_13296);
xor U13517 (N_13517,N_13251,N_13352);
and U13518 (N_13518,N_13204,N_13305);
nor U13519 (N_13519,N_13260,N_13365);
nor U13520 (N_13520,N_13366,N_13345);
xor U13521 (N_13521,N_13207,N_13260);
or U13522 (N_13522,N_13397,N_13374);
xor U13523 (N_13523,N_13317,N_13320);
xnor U13524 (N_13524,N_13310,N_13330);
or U13525 (N_13525,N_13322,N_13387);
nand U13526 (N_13526,N_13253,N_13206);
and U13527 (N_13527,N_13274,N_13378);
nor U13528 (N_13528,N_13398,N_13346);
and U13529 (N_13529,N_13217,N_13256);
and U13530 (N_13530,N_13343,N_13294);
and U13531 (N_13531,N_13269,N_13226);
nor U13532 (N_13532,N_13266,N_13260);
and U13533 (N_13533,N_13349,N_13335);
or U13534 (N_13534,N_13258,N_13352);
xor U13535 (N_13535,N_13275,N_13353);
and U13536 (N_13536,N_13371,N_13242);
and U13537 (N_13537,N_13391,N_13392);
or U13538 (N_13538,N_13308,N_13224);
nand U13539 (N_13539,N_13219,N_13335);
and U13540 (N_13540,N_13356,N_13392);
xor U13541 (N_13541,N_13310,N_13248);
or U13542 (N_13542,N_13330,N_13236);
and U13543 (N_13543,N_13376,N_13356);
and U13544 (N_13544,N_13305,N_13346);
xnor U13545 (N_13545,N_13379,N_13378);
nand U13546 (N_13546,N_13266,N_13212);
xor U13547 (N_13547,N_13274,N_13233);
nor U13548 (N_13548,N_13285,N_13303);
or U13549 (N_13549,N_13307,N_13260);
and U13550 (N_13550,N_13297,N_13365);
xnor U13551 (N_13551,N_13238,N_13314);
and U13552 (N_13552,N_13279,N_13214);
or U13553 (N_13553,N_13392,N_13234);
nand U13554 (N_13554,N_13360,N_13266);
nor U13555 (N_13555,N_13318,N_13255);
or U13556 (N_13556,N_13349,N_13206);
or U13557 (N_13557,N_13323,N_13373);
nand U13558 (N_13558,N_13303,N_13238);
nand U13559 (N_13559,N_13342,N_13322);
and U13560 (N_13560,N_13275,N_13317);
nand U13561 (N_13561,N_13300,N_13289);
or U13562 (N_13562,N_13249,N_13224);
nor U13563 (N_13563,N_13211,N_13229);
and U13564 (N_13564,N_13216,N_13209);
xor U13565 (N_13565,N_13297,N_13295);
and U13566 (N_13566,N_13213,N_13202);
nor U13567 (N_13567,N_13323,N_13345);
and U13568 (N_13568,N_13225,N_13204);
nor U13569 (N_13569,N_13240,N_13375);
or U13570 (N_13570,N_13254,N_13298);
nand U13571 (N_13571,N_13247,N_13248);
nor U13572 (N_13572,N_13364,N_13379);
or U13573 (N_13573,N_13385,N_13376);
or U13574 (N_13574,N_13271,N_13263);
nor U13575 (N_13575,N_13397,N_13285);
and U13576 (N_13576,N_13211,N_13272);
nand U13577 (N_13577,N_13385,N_13350);
or U13578 (N_13578,N_13398,N_13214);
xnor U13579 (N_13579,N_13284,N_13276);
and U13580 (N_13580,N_13240,N_13307);
or U13581 (N_13581,N_13287,N_13245);
nand U13582 (N_13582,N_13357,N_13291);
xor U13583 (N_13583,N_13236,N_13276);
nand U13584 (N_13584,N_13346,N_13281);
nor U13585 (N_13585,N_13200,N_13289);
nand U13586 (N_13586,N_13305,N_13213);
or U13587 (N_13587,N_13308,N_13258);
and U13588 (N_13588,N_13223,N_13347);
and U13589 (N_13589,N_13305,N_13318);
nand U13590 (N_13590,N_13354,N_13254);
or U13591 (N_13591,N_13332,N_13235);
nand U13592 (N_13592,N_13284,N_13368);
xnor U13593 (N_13593,N_13328,N_13213);
or U13594 (N_13594,N_13333,N_13285);
nor U13595 (N_13595,N_13279,N_13325);
nand U13596 (N_13596,N_13237,N_13394);
xnor U13597 (N_13597,N_13218,N_13312);
nor U13598 (N_13598,N_13320,N_13319);
and U13599 (N_13599,N_13323,N_13325);
or U13600 (N_13600,N_13455,N_13525);
and U13601 (N_13601,N_13576,N_13423);
or U13602 (N_13602,N_13554,N_13591);
nand U13603 (N_13603,N_13549,N_13404);
or U13604 (N_13604,N_13542,N_13489);
nor U13605 (N_13605,N_13488,N_13460);
nor U13606 (N_13606,N_13413,N_13426);
or U13607 (N_13607,N_13563,N_13584);
xnor U13608 (N_13608,N_13573,N_13516);
xnor U13609 (N_13609,N_13529,N_13498);
and U13610 (N_13610,N_13578,N_13504);
nor U13611 (N_13611,N_13418,N_13595);
nor U13612 (N_13612,N_13402,N_13405);
or U13613 (N_13613,N_13515,N_13565);
and U13614 (N_13614,N_13523,N_13590);
and U13615 (N_13615,N_13519,N_13566);
or U13616 (N_13616,N_13527,N_13401);
or U13617 (N_13617,N_13530,N_13474);
xor U13618 (N_13618,N_13438,N_13459);
and U13619 (N_13619,N_13594,N_13431);
and U13620 (N_13620,N_13495,N_13425);
nand U13621 (N_13621,N_13482,N_13556);
nor U13622 (N_13622,N_13538,N_13453);
nand U13623 (N_13623,N_13572,N_13589);
nor U13624 (N_13624,N_13450,N_13437);
and U13625 (N_13625,N_13508,N_13592);
and U13626 (N_13626,N_13586,N_13585);
xor U13627 (N_13627,N_13408,N_13547);
and U13628 (N_13628,N_13507,N_13463);
nand U13629 (N_13629,N_13461,N_13492);
nand U13630 (N_13630,N_13448,N_13510);
nor U13631 (N_13631,N_13468,N_13419);
nand U13632 (N_13632,N_13567,N_13484);
nand U13633 (N_13633,N_13429,N_13475);
and U13634 (N_13634,N_13465,N_13535);
xnor U13635 (N_13635,N_13506,N_13551);
nor U13636 (N_13636,N_13575,N_13400);
xor U13637 (N_13637,N_13598,N_13456);
nor U13638 (N_13638,N_13564,N_13407);
nand U13639 (N_13639,N_13433,N_13502);
and U13640 (N_13640,N_13473,N_13597);
nand U13641 (N_13641,N_13593,N_13505);
and U13642 (N_13642,N_13517,N_13451);
nand U13643 (N_13643,N_13548,N_13533);
nor U13644 (N_13644,N_13560,N_13503);
or U13645 (N_13645,N_13553,N_13596);
xnor U13646 (N_13646,N_13480,N_13417);
nor U13647 (N_13647,N_13570,N_13546);
nor U13648 (N_13648,N_13490,N_13452);
nor U13649 (N_13649,N_13458,N_13531);
and U13650 (N_13650,N_13439,N_13557);
xnor U13651 (N_13651,N_13545,N_13583);
and U13652 (N_13652,N_13442,N_13559);
or U13653 (N_13653,N_13520,N_13562);
and U13654 (N_13654,N_13537,N_13409);
nand U13655 (N_13655,N_13462,N_13543);
and U13656 (N_13656,N_13513,N_13493);
nor U13657 (N_13657,N_13494,N_13412);
and U13658 (N_13658,N_13521,N_13470);
nor U13659 (N_13659,N_13441,N_13440);
nand U13660 (N_13660,N_13579,N_13541);
or U13661 (N_13661,N_13518,N_13436);
or U13662 (N_13662,N_13496,N_13485);
nor U13663 (N_13663,N_13561,N_13422);
or U13664 (N_13664,N_13581,N_13434);
or U13665 (N_13665,N_13569,N_13552);
xor U13666 (N_13666,N_13454,N_13501);
xor U13667 (N_13667,N_13432,N_13511);
nor U13668 (N_13668,N_13476,N_13544);
nand U13669 (N_13669,N_13500,N_13427);
and U13670 (N_13670,N_13558,N_13410);
and U13671 (N_13671,N_13528,N_13532);
nor U13672 (N_13672,N_13472,N_13477);
nor U13673 (N_13673,N_13464,N_13540);
xor U13674 (N_13674,N_13577,N_13514);
nand U13675 (N_13675,N_13449,N_13587);
nand U13676 (N_13676,N_13555,N_13479);
or U13677 (N_13677,N_13406,N_13446);
and U13678 (N_13678,N_13526,N_13512);
or U13679 (N_13679,N_13568,N_13411);
xnor U13680 (N_13680,N_13421,N_13478);
and U13681 (N_13681,N_13424,N_13580);
and U13682 (N_13682,N_13550,N_13457);
xnor U13683 (N_13683,N_13445,N_13467);
and U13684 (N_13684,N_13534,N_13486);
or U13685 (N_13685,N_13483,N_13481);
and U13686 (N_13686,N_13522,N_13509);
xor U13687 (N_13687,N_13491,N_13466);
and U13688 (N_13688,N_13536,N_13447);
nor U13689 (N_13689,N_13430,N_13499);
or U13690 (N_13690,N_13414,N_13435);
and U13691 (N_13691,N_13428,N_13571);
nor U13692 (N_13692,N_13444,N_13403);
or U13693 (N_13693,N_13497,N_13574);
or U13694 (N_13694,N_13524,N_13539);
or U13695 (N_13695,N_13487,N_13415);
nor U13696 (N_13696,N_13416,N_13588);
or U13697 (N_13697,N_13599,N_13420);
nor U13698 (N_13698,N_13469,N_13582);
and U13699 (N_13699,N_13443,N_13471);
or U13700 (N_13700,N_13467,N_13502);
and U13701 (N_13701,N_13405,N_13590);
and U13702 (N_13702,N_13570,N_13405);
nor U13703 (N_13703,N_13533,N_13526);
and U13704 (N_13704,N_13495,N_13465);
xnor U13705 (N_13705,N_13569,N_13486);
and U13706 (N_13706,N_13568,N_13524);
nand U13707 (N_13707,N_13579,N_13516);
nand U13708 (N_13708,N_13416,N_13559);
and U13709 (N_13709,N_13499,N_13496);
or U13710 (N_13710,N_13553,N_13406);
nand U13711 (N_13711,N_13458,N_13560);
nor U13712 (N_13712,N_13526,N_13473);
and U13713 (N_13713,N_13548,N_13416);
xnor U13714 (N_13714,N_13592,N_13467);
or U13715 (N_13715,N_13442,N_13568);
or U13716 (N_13716,N_13489,N_13451);
or U13717 (N_13717,N_13539,N_13407);
nand U13718 (N_13718,N_13496,N_13591);
nor U13719 (N_13719,N_13588,N_13515);
nor U13720 (N_13720,N_13532,N_13492);
nor U13721 (N_13721,N_13507,N_13501);
xor U13722 (N_13722,N_13462,N_13558);
nand U13723 (N_13723,N_13415,N_13474);
xor U13724 (N_13724,N_13517,N_13511);
nand U13725 (N_13725,N_13480,N_13553);
nor U13726 (N_13726,N_13416,N_13564);
nor U13727 (N_13727,N_13558,N_13494);
or U13728 (N_13728,N_13583,N_13521);
nand U13729 (N_13729,N_13595,N_13511);
or U13730 (N_13730,N_13565,N_13418);
xor U13731 (N_13731,N_13435,N_13563);
and U13732 (N_13732,N_13565,N_13557);
nor U13733 (N_13733,N_13542,N_13403);
nand U13734 (N_13734,N_13590,N_13434);
or U13735 (N_13735,N_13486,N_13578);
and U13736 (N_13736,N_13535,N_13501);
or U13737 (N_13737,N_13563,N_13531);
nand U13738 (N_13738,N_13430,N_13421);
nor U13739 (N_13739,N_13468,N_13480);
and U13740 (N_13740,N_13557,N_13431);
or U13741 (N_13741,N_13517,N_13510);
nor U13742 (N_13742,N_13577,N_13561);
xor U13743 (N_13743,N_13424,N_13525);
xnor U13744 (N_13744,N_13411,N_13450);
nor U13745 (N_13745,N_13433,N_13464);
or U13746 (N_13746,N_13512,N_13434);
or U13747 (N_13747,N_13475,N_13430);
and U13748 (N_13748,N_13533,N_13507);
xor U13749 (N_13749,N_13497,N_13528);
or U13750 (N_13750,N_13495,N_13515);
xnor U13751 (N_13751,N_13495,N_13445);
and U13752 (N_13752,N_13579,N_13504);
xor U13753 (N_13753,N_13482,N_13570);
and U13754 (N_13754,N_13458,N_13416);
nor U13755 (N_13755,N_13543,N_13572);
nand U13756 (N_13756,N_13536,N_13581);
and U13757 (N_13757,N_13548,N_13410);
nand U13758 (N_13758,N_13543,N_13459);
nor U13759 (N_13759,N_13586,N_13427);
nor U13760 (N_13760,N_13468,N_13566);
nor U13761 (N_13761,N_13545,N_13492);
xnor U13762 (N_13762,N_13417,N_13577);
nor U13763 (N_13763,N_13566,N_13420);
and U13764 (N_13764,N_13462,N_13541);
xor U13765 (N_13765,N_13418,N_13411);
nand U13766 (N_13766,N_13570,N_13492);
nand U13767 (N_13767,N_13597,N_13474);
nand U13768 (N_13768,N_13588,N_13424);
and U13769 (N_13769,N_13588,N_13459);
nor U13770 (N_13770,N_13502,N_13500);
and U13771 (N_13771,N_13455,N_13403);
or U13772 (N_13772,N_13409,N_13538);
xnor U13773 (N_13773,N_13549,N_13554);
and U13774 (N_13774,N_13532,N_13576);
and U13775 (N_13775,N_13591,N_13405);
xnor U13776 (N_13776,N_13517,N_13523);
or U13777 (N_13777,N_13429,N_13459);
and U13778 (N_13778,N_13416,N_13525);
nor U13779 (N_13779,N_13483,N_13581);
and U13780 (N_13780,N_13558,N_13434);
nand U13781 (N_13781,N_13481,N_13511);
xor U13782 (N_13782,N_13475,N_13413);
nand U13783 (N_13783,N_13492,N_13501);
or U13784 (N_13784,N_13428,N_13512);
xnor U13785 (N_13785,N_13436,N_13577);
nand U13786 (N_13786,N_13489,N_13417);
and U13787 (N_13787,N_13508,N_13409);
and U13788 (N_13788,N_13575,N_13550);
nor U13789 (N_13789,N_13417,N_13546);
xor U13790 (N_13790,N_13479,N_13599);
xnor U13791 (N_13791,N_13502,N_13534);
nor U13792 (N_13792,N_13446,N_13550);
and U13793 (N_13793,N_13544,N_13563);
xor U13794 (N_13794,N_13558,N_13457);
xor U13795 (N_13795,N_13451,N_13443);
or U13796 (N_13796,N_13478,N_13412);
nand U13797 (N_13797,N_13416,N_13501);
and U13798 (N_13798,N_13468,N_13479);
xnor U13799 (N_13799,N_13483,N_13405);
nor U13800 (N_13800,N_13756,N_13730);
xnor U13801 (N_13801,N_13773,N_13710);
nor U13802 (N_13802,N_13611,N_13604);
or U13803 (N_13803,N_13701,N_13724);
nor U13804 (N_13804,N_13765,N_13712);
or U13805 (N_13805,N_13763,N_13677);
xnor U13806 (N_13806,N_13680,N_13785);
nor U13807 (N_13807,N_13759,N_13670);
xor U13808 (N_13808,N_13729,N_13754);
or U13809 (N_13809,N_13771,N_13755);
nand U13810 (N_13810,N_13719,N_13702);
and U13811 (N_13811,N_13752,N_13634);
or U13812 (N_13812,N_13741,N_13711);
nand U13813 (N_13813,N_13660,N_13600);
nor U13814 (N_13814,N_13618,N_13659);
or U13815 (N_13815,N_13636,N_13744);
nand U13816 (N_13816,N_13794,N_13709);
and U13817 (N_13817,N_13775,N_13704);
and U13818 (N_13818,N_13691,N_13690);
and U13819 (N_13819,N_13657,N_13681);
or U13820 (N_13820,N_13747,N_13694);
nand U13821 (N_13821,N_13761,N_13776);
nor U13822 (N_13822,N_13654,N_13617);
and U13823 (N_13823,N_13679,N_13645);
nor U13824 (N_13824,N_13653,N_13602);
nand U13825 (N_13825,N_13609,N_13743);
nand U13826 (N_13826,N_13751,N_13778);
or U13827 (N_13827,N_13674,N_13766);
and U13828 (N_13828,N_13663,N_13772);
or U13829 (N_13829,N_13750,N_13760);
nor U13830 (N_13830,N_13769,N_13652);
nand U13831 (N_13831,N_13793,N_13638);
and U13832 (N_13832,N_13616,N_13783);
nand U13833 (N_13833,N_13629,N_13792);
and U13834 (N_13834,N_13768,N_13676);
and U13835 (N_13835,N_13736,N_13664);
xnor U13836 (N_13836,N_13738,N_13696);
nor U13837 (N_13837,N_13658,N_13728);
nand U13838 (N_13838,N_13671,N_13662);
nor U13839 (N_13839,N_13697,N_13699);
nand U13840 (N_13840,N_13779,N_13627);
xnor U13841 (N_13841,N_13610,N_13717);
xnor U13842 (N_13842,N_13705,N_13647);
or U13843 (N_13843,N_13720,N_13733);
nand U13844 (N_13844,N_13746,N_13685);
xnor U13845 (N_13845,N_13780,N_13740);
and U13846 (N_13846,N_13796,N_13624);
or U13847 (N_13847,N_13633,N_13787);
nor U13848 (N_13848,N_13642,N_13613);
nand U13849 (N_13849,N_13684,N_13742);
nor U13850 (N_13850,N_13621,N_13622);
nor U13851 (N_13851,N_13789,N_13607);
or U13852 (N_13852,N_13639,N_13673);
xnor U13853 (N_13853,N_13641,N_13737);
xor U13854 (N_13854,N_13716,N_13669);
nand U13855 (N_13855,N_13644,N_13732);
xor U13856 (N_13856,N_13631,N_13667);
nand U13857 (N_13857,N_13665,N_13608);
xnor U13858 (N_13858,N_13715,N_13781);
nand U13859 (N_13859,N_13795,N_13749);
xnor U13860 (N_13860,N_13626,N_13603);
or U13861 (N_13861,N_13767,N_13703);
or U13862 (N_13862,N_13630,N_13675);
nand U13863 (N_13863,N_13797,N_13695);
xor U13864 (N_13864,N_13687,N_13706);
or U13865 (N_13865,N_13799,N_13605);
xor U13866 (N_13866,N_13788,N_13718);
and U13867 (N_13867,N_13722,N_13693);
and U13868 (N_13868,N_13601,N_13655);
xnor U13869 (N_13869,N_13656,N_13734);
nor U13870 (N_13870,N_13615,N_13646);
or U13871 (N_13871,N_13757,N_13774);
or U13872 (N_13872,N_13790,N_13708);
nor U13873 (N_13873,N_13640,N_13688);
and U13874 (N_13874,N_13683,N_13707);
nor U13875 (N_13875,N_13682,N_13764);
nand U13876 (N_13876,N_13666,N_13758);
nor U13877 (N_13877,N_13762,N_13625);
and U13878 (N_13878,N_13723,N_13721);
and U13879 (N_13879,N_13727,N_13606);
or U13880 (N_13880,N_13753,N_13798);
and U13881 (N_13881,N_13619,N_13739);
or U13882 (N_13882,N_13649,N_13731);
nor U13883 (N_13883,N_13784,N_13686);
nor U13884 (N_13884,N_13692,N_13648);
or U13885 (N_13885,N_13620,N_13770);
xor U13886 (N_13886,N_13698,N_13672);
and U13887 (N_13887,N_13714,N_13786);
or U13888 (N_13888,N_13748,N_13635);
xor U13889 (N_13889,N_13725,N_13713);
nor U13890 (N_13890,N_13726,N_13623);
and U13891 (N_13891,N_13650,N_13614);
nor U13892 (N_13892,N_13678,N_13700);
nand U13893 (N_13893,N_13661,N_13668);
and U13894 (N_13894,N_13643,N_13777);
and U13895 (N_13895,N_13689,N_13791);
or U13896 (N_13896,N_13651,N_13637);
or U13897 (N_13897,N_13782,N_13612);
nand U13898 (N_13898,N_13632,N_13628);
and U13899 (N_13899,N_13745,N_13735);
or U13900 (N_13900,N_13690,N_13797);
or U13901 (N_13901,N_13685,N_13769);
or U13902 (N_13902,N_13721,N_13753);
nor U13903 (N_13903,N_13757,N_13635);
xnor U13904 (N_13904,N_13760,N_13736);
or U13905 (N_13905,N_13680,N_13732);
nor U13906 (N_13906,N_13700,N_13738);
nand U13907 (N_13907,N_13607,N_13778);
and U13908 (N_13908,N_13757,N_13736);
and U13909 (N_13909,N_13610,N_13794);
nor U13910 (N_13910,N_13626,N_13652);
or U13911 (N_13911,N_13680,N_13737);
nand U13912 (N_13912,N_13750,N_13765);
xnor U13913 (N_13913,N_13650,N_13696);
nor U13914 (N_13914,N_13767,N_13720);
xor U13915 (N_13915,N_13644,N_13673);
xor U13916 (N_13916,N_13617,N_13661);
or U13917 (N_13917,N_13742,N_13761);
or U13918 (N_13918,N_13724,N_13612);
and U13919 (N_13919,N_13615,N_13682);
and U13920 (N_13920,N_13601,N_13715);
and U13921 (N_13921,N_13688,N_13614);
nand U13922 (N_13922,N_13731,N_13640);
and U13923 (N_13923,N_13741,N_13714);
nor U13924 (N_13924,N_13643,N_13676);
nor U13925 (N_13925,N_13691,N_13633);
nand U13926 (N_13926,N_13727,N_13694);
nor U13927 (N_13927,N_13609,N_13771);
nor U13928 (N_13928,N_13625,N_13751);
nor U13929 (N_13929,N_13694,N_13676);
nand U13930 (N_13930,N_13665,N_13686);
nor U13931 (N_13931,N_13783,N_13716);
xnor U13932 (N_13932,N_13703,N_13680);
nand U13933 (N_13933,N_13687,N_13704);
nand U13934 (N_13934,N_13731,N_13683);
and U13935 (N_13935,N_13612,N_13748);
nand U13936 (N_13936,N_13684,N_13658);
or U13937 (N_13937,N_13732,N_13685);
xor U13938 (N_13938,N_13693,N_13623);
or U13939 (N_13939,N_13698,N_13782);
xnor U13940 (N_13940,N_13748,N_13663);
nor U13941 (N_13941,N_13662,N_13695);
nand U13942 (N_13942,N_13629,N_13689);
and U13943 (N_13943,N_13661,N_13680);
nor U13944 (N_13944,N_13793,N_13635);
nor U13945 (N_13945,N_13663,N_13712);
nand U13946 (N_13946,N_13615,N_13789);
nor U13947 (N_13947,N_13787,N_13600);
and U13948 (N_13948,N_13759,N_13710);
and U13949 (N_13949,N_13642,N_13716);
nor U13950 (N_13950,N_13732,N_13717);
nand U13951 (N_13951,N_13683,N_13770);
and U13952 (N_13952,N_13668,N_13691);
xor U13953 (N_13953,N_13758,N_13751);
nand U13954 (N_13954,N_13785,N_13687);
nor U13955 (N_13955,N_13693,N_13789);
or U13956 (N_13956,N_13725,N_13775);
nor U13957 (N_13957,N_13691,N_13644);
xor U13958 (N_13958,N_13610,N_13778);
xnor U13959 (N_13959,N_13723,N_13793);
nor U13960 (N_13960,N_13755,N_13648);
nand U13961 (N_13961,N_13621,N_13617);
nand U13962 (N_13962,N_13759,N_13623);
or U13963 (N_13963,N_13782,N_13723);
xor U13964 (N_13964,N_13696,N_13725);
nand U13965 (N_13965,N_13723,N_13744);
or U13966 (N_13966,N_13791,N_13767);
nor U13967 (N_13967,N_13620,N_13721);
or U13968 (N_13968,N_13662,N_13661);
xor U13969 (N_13969,N_13755,N_13700);
or U13970 (N_13970,N_13623,N_13728);
xor U13971 (N_13971,N_13618,N_13747);
xnor U13972 (N_13972,N_13772,N_13650);
nand U13973 (N_13973,N_13687,N_13655);
nand U13974 (N_13974,N_13736,N_13628);
and U13975 (N_13975,N_13622,N_13752);
nand U13976 (N_13976,N_13723,N_13618);
nor U13977 (N_13977,N_13609,N_13638);
and U13978 (N_13978,N_13671,N_13610);
and U13979 (N_13979,N_13745,N_13757);
xnor U13980 (N_13980,N_13695,N_13689);
xnor U13981 (N_13981,N_13661,N_13697);
and U13982 (N_13982,N_13602,N_13703);
and U13983 (N_13983,N_13638,N_13644);
and U13984 (N_13984,N_13787,N_13658);
or U13985 (N_13985,N_13650,N_13761);
nand U13986 (N_13986,N_13756,N_13760);
xnor U13987 (N_13987,N_13688,N_13797);
nand U13988 (N_13988,N_13690,N_13715);
xnor U13989 (N_13989,N_13741,N_13627);
nand U13990 (N_13990,N_13648,N_13797);
xnor U13991 (N_13991,N_13780,N_13668);
or U13992 (N_13992,N_13711,N_13627);
xnor U13993 (N_13993,N_13710,N_13646);
xnor U13994 (N_13994,N_13742,N_13648);
nor U13995 (N_13995,N_13671,N_13708);
xnor U13996 (N_13996,N_13640,N_13748);
nor U13997 (N_13997,N_13696,N_13712);
nand U13998 (N_13998,N_13753,N_13670);
nand U13999 (N_13999,N_13610,N_13692);
nor U14000 (N_14000,N_13816,N_13960);
xnor U14001 (N_14001,N_13906,N_13947);
xnor U14002 (N_14002,N_13895,N_13877);
nand U14003 (N_14003,N_13832,N_13875);
xor U14004 (N_14004,N_13928,N_13942);
or U14005 (N_14005,N_13818,N_13978);
xnor U14006 (N_14006,N_13855,N_13952);
nor U14007 (N_14007,N_13915,N_13900);
and U14008 (N_14008,N_13974,N_13968);
nand U14009 (N_14009,N_13812,N_13980);
nand U14010 (N_14010,N_13874,N_13940);
xor U14011 (N_14011,N_13831,N_13857);
nor U14012 (N_14012,N_13834,N_13901);
nand U14013 (N_14013,N_13944,N_13969);
xnor U14014 (N_14014,N_13884,N_13837);
and U14015 (N_14015,N_13820,N_13945);
and U14016 (N_14016,N_13970,N_13918);
xnor U14017 (N_14017,N_13989,N_13836);
nor U14018 (N_14018,N_13859,N_13894);
nor U14019 (N_14019,N_13885,N_13999);
and U14020 (N_14020,N_13956,N_13809);
xnor U14021 (N_14021,N_13811,N_13943);
and U14022 (N_14022,N_13876,N_13890);
xnor U14023 (N_14023,N_13807,N_13971);
nor U14024 (N_14024,N_13897,N_13997);
and U14025 (N_14025,N_13994,N_13983);
and U14026 (N_14026,N_13804,N_13886);
or U14027 (N_14027,N_13925,N_13988);
and U14028 (N_14028,N_13949,N_13920);
nand U14029 (N_14029,N_13854,N_13826);
and U14030 (N_14030,N_13976,N_13991);
nor U14031 (N_14031,N_13935,N_13995);
nand U14032 (N_14032,N_13810,N_13815);
nor U14033 (N_14033,N_13987,N_13898);
nor U14034 (N_14034,N_13904,N_13870);
nor U14035 (N_14035,N_13993,N_13938);
xor U14036 (N_14036,N_13902,N_13930);
xor U14037 (N_14037,N_13800,N_13998);
and U14038 (N_14038,N_13825,N_13977);
or U14039 (N_14039,N_13914,N_13973);
xnor U14040 (N_14040,N_13959,N_13931);
nand U14041 (N_14041,N_13964,N_13821);
nor U14042 (N_14042,N_13916,N_13802);
xnor U14043 (N_14043,N_13957,N_13850);
nand U14044 (N_14044,N_13882,N_13907);
and U14045 (N_14045,N_13941,N_13879);
nor U14046 (N_14046,N_13862,N_13853);
nand U14047 (N_14047,N_13801,N_13979);
or U14048 (N_14048,N_13806,N_13873);
and U14049 (N_14049,N_13847,N_13828);
nand U14050 (N_14050,N_13954,N_13933);
xnor U14051 (N_14051,N_13972,N_13965);
and U14052 (N_14052,N_13858,N_13844);
or U14053 (N_14053,N_13909,N_13922);
or U14054 (N_14054,N_13867,N_13975);
or U14055 (N_14055,N_13888,N_13990);
xnor U14056 (N_14056,N_13927,N_13866);
xor U14057 (N_14057,N_13937,N_13871);
nand U14058 (N_14058,N_13848,N_13814);
nand U14059 (N_14059,N_13936,N_13946);
or U14060 (N_14060,N_13986,N_13852);
nand U14061 (N_14061,N_13839,N_13824);
nor U14062 (N_14062,N_13803,N_13808);
xnor U14063 (N_14063,N_13929,N_13917);
xnor U14064 (N_14064,N_13840,N_13924);
nand U14065 (N_14065,N_13910,N_13865);
nor U14066 (N_14066,N_13966,N_13851);
or U14067 (N_14067,N_13827,N_13950);
nand U14068 (N_14068,N_13843,N_13984);
xor U14069 (N_14069,N_13992,N_13948);
nand U14070 (N_14070,N_13953,N_13863);
xnor U14071 (N_14071,N_13893,N_13962);
xor U14072 (N_14072,N_13958,N_13805);
or U14073 (N_14073,N_13919,N_13899);
or U14074 (N_14074,N_13905,N_13860);
nand U14075 (N_14075,N_13881,N_13817);
nand U14076 (N_14076,N_13981,N_13932);
nor U14077 (N_14077,N_13813,N_13856);
nand U14078 (N_14078,N_13985,N_13982);
nor U14079 (N_14079,N_13835,N_13845);
nor U14080 (N_14080,N_13967,N_13903);
and U14081 (N_14081,N_13819,N_13878);
nand U14082 (N_14082,N_13913,N_13939);
nor U14083 (N_14083,N_13955,N_13880);
nand U14084 (N_14084,N_13951,N_13846);
nand U14085 (N_14085,N_13833,N_13864);
nand U14086 (N_14086,N_13829,N_13861);
xor U14087 (N_14087,N_13823,N_13889);
or U14088 (N_14088,N_13822,N_13923);
nor U14089 (N_14089,N_13963,N_13926);
and U14090 (N_14090,N_13896,N_13934);
nand U14091 (N_14091,N_13887,N_13891);
xor U14092 (N_14092,N_13868,N_13842);
nor U14093 (N_14093,N_13911,N_13996);
xor U14094 (N_14094,N_13883,N_13830);
xor U14095 (N_14095,N_13961,N_13908);
xor U14096 (N_14096,N_13892,N_13872);
and U14097 (N_14097,N_13849,N_13921);
nor U14098 (N_14098,N_13841,N_13838);
nor U14099 (N_14099,N_13869,N_13912);
xor U14100 (N_14100,N_13994,N_13886);
xor U14101 (N_14101,N_13978,N_13840);
or U14102 (N_14102,N_13927,N_13920);
or U14103 (N_14103,N_13831,N_13984);
xnor U14104 (N_14104,N_13941,N_13819);
xnor U14105 (N_14105,N_13815,N_13855);
nand U14106 (N_14106,N_13980,N_13849);
nand U14107 (N_14107,N_13906,N_13880);
or U14108 (N_14108,N_13801,N_13984);
nor U14109 (N_14109,N_13815,N_13881);
and U14110 (N_14110,N_13963,N_13818);
nor U14111 (N_14111,N_13832,N_13936);
nor U14112 (N_14112,N_13974,N_13813);
xor U14113 (N_14113,N_13906,N_13930);
xnor U14114 (N_14114,N_13948,N_13945);
or U14115 (N_14115,N_13988,N_13935);
nand U14116 (N_14116,N_13838,N_13815);
nor U14117 (N_14117,N_13824,N_13811);
nor U14118 (N_14118,N_13991,N_13867);
and U14119 (N_14119,N_13836,N_13859);
or U14120 (N_14120,N_13974,N_13939);
nor U14121 (N_14121,N_13892,N_13906);
nor U14122 (N_14122,N_13922,N_13808);
nand U14123 (N_14123,N_13937,N_13908);
or U14124 (N_14124,N_13997,N_13982);
nand U14125 (N_14125,N_13835,N_13925);
or U14126 (N_14126,N_13934,N_13815);
xor U14127 (N_14127,N_13820,N_13826);
nand U14128 (N_14128,N_13973,N_13910);
xor U14129 (N_14129,N_13982,N_13915);
nand U14130 (N_14130,N_13839,N_13875);
and U14131 (N_14131,N_13860,N_13979);
or U14132 (N_14132,N_13926,N_13881);
nand U14133 (N_14133,N_13855,N_13841);
nand U14134 (N_14134,N_13965,N_13849);
xnor U14135 (N_14135,N_13998,N_13897);
or U14136 (N_14136,N_13881,N_13895);
nand U14137 (N_14137,N_13948,N_13849);
nand U14138 (N_14138,N_13985,N_13953);
and U14139 (N_14139,N_13925,N_13927);
nand U14140 (N_14140,N_13865,N_13922);
and U14141 (N_14141,N_13813,N_13841);
xor U14142 (N_14142,N_13976,N_13994);
and U14143 (N_14143,N_13868,N_13885);
xor U14144 (N_14144,N_13804,N_13965);
xor U14145 (N_14145,N_13839,N_13993);
nand U14146 (N_14146,N_13886,N_13853);
xor U14147 (N_14147,N_13980,N_13863);
nand U14148 (N_14148,N_13920,N_13950);
or U14149 (N_14149,N_13862,N_13945);
nor U14150 (N_14150,N_13895,N_13922);
xnor U14151 (N_14151,N_13911,N_13855);
or U14152 (N_14152,N_13920,N_13970);
and U14153 (N_14153,N_13903,N_13881);
or U14154 (N_14154,N_13948,N_13839);
or U14155 (N_14155,N_13808,N_13915);
nor U14156 (N_14156,N_13802,N_13981);
and U14157 (N_14157,N_13817,N_13846);
and U14158 (N_14158,N_13868,N_13858);
nor U14159 (N_14159,N_13842,N_13827);
nor U14160 (N_14160,N_13990,N_13998);
and U14161 (N_14161,N_13944,N_13962);
nand U14162 (N_14162,N_13899,N_13840);
nor U14163 (N_14163,N_13859,N_13963);
or U14164 (N_14164,N_13853,N_13996);
or U14165 (N_14165,N_13805,N_13929);
nand U14166 (N_14166,N_13886,N_13867);
nand U14167 (N_14167,N_13856,N_13906);
nor U14168 (N_14168,N_13963,N_13955);
xnor U14169 (N_14169,N_13920,N_13972);
nor U14170 (N_14170,N_13985,N_13875);
nand U14171 (N_14171,N_13911,N_13977);
and U14172 (N_14172,N_13856,N_13931);
or U14173 (N_14173,N_13980,N_13895);
xor U14174 (N_14174,N_13953,N_13813);
nor U14175 (N_14175,N_13824,N_13919);
nand U14176 (N_14176,N_13961,N_13953);
or U14177 (N_14177,N_13992,N_13873);
and U14178 (N_14178,N_13949,N_13900);
nor U14179 (N_14179,N_13847,N_13951);
or U14180 (N_14180,N_13816,N_13812);
and U14181 (N_14181,N_13861,N_13909);
nand U14182 (N_14182,N_13800,N_13953);
and U14183 (N_14183,N_13970,N_13809);
or U14184 (N_14184,N_13867,N_13914);
nand U14185 (N_14185,N_13899,N_13961);
nand U14186 (N_14186,N_13813,N_13883);
xnor U14187 (N_14187,N_13895,N_13869);
or U14188 (N_14188,N_13856,N_13957);
nand U14189 (N_14189,N_13961,N_13924);
or U14190 (N_14190,N_13958,N_13885);
nand U14191 (N_14191,N_13964,N_13804);
and U14192 (N_14192,N_13974,N_13872);
and U14193 (N_14193,N_13833,N_13916);
nor U14194 (N_14194,N_13910,N_13909);
xor U14195 (N_14195,N_13988,N_13970);
xnor U14196 (N_14196,N_13904,N_13935);
nand U14197 (N_14197,N_13987,N_13962);
nor U14198 (N_14198,N_13822,N_13879);
and U14199 (N_14199,N_13958,N_13985);
and U14200 (N_14200,N_14155,N_14147);
nor U14201 (N_14201,N_14064,N_14108);
or U14202 (N_14202,N_14140,N_14080);
or U14203 (N_14203,N_14011,N_14076);
xnor U14204 (N_14204,N_14189,N_14186);
nand U14205 (N_14205,N_14170,N_14010);
and U14206 (N_14206,N_14000,N_14124);
xnor U14207 (N_14207,N_14184,N_14031);
or U14208 (N_14208,N_14195,N_14020);
nor U14209 (N_14209,N_14171,N_14117);
and U14210 (N_14210,N_14086,N_14062);
nand U14211 (N_14211,N_14002,N_14103);
and U14212 (N_14212,N_14027,N_14192);
or U14213 (N_14213,N_14055,N_14053);
xor U14214 (N_14214,N_14178,N_14029);
nand U14215 (N_14215,N_14058,N_14167);
or U14216 (N_14216,N_14074,N_14169);
nand U14217 (N_14217,N_14004,N_14081);
xor U14218 (N_14218,N_14090,N_14061);
or U14219 (N_14219,N_14163,N_14135);
xnor U14220 (N_14220,N_14159,N_14119);
nor U14221 (N_14221,N_14110,N_14068);
or U14222 (N_14222,N_14154,N_14183);
or U14223 (N_14223,N_14123,N_14038);
nor U14224 (N_14224,N_14036,N_14032);
nor U14225 (N_14225,N_14072,N_14084);
xnor U14226 (N_14226,N_14132,N_14087);
nand U14227 (N_14227,N_14129,N_14179);
nor U14228 (N_14228,N_14125,N_14035);
or U14229 (N_14229,N_14174,N_14180);
nand U14230 (N_14230,N_14156,N_14014);
xnor U14231 (N_14231,N_14148,N_14191);
nand U14232 (N_14232,N_14199,N_14030);
nor U14233 (N_14233,N_14175,N_14005);
xor U14234 (N_14234,N_14099,N_14047);
and U14235 (N_14235,N_14146,N_14012);
or U14236 (N_14236,N_14059,N_14187);
nor U14237 (N_14237,N_14115,N_14024);
nor U14238 (N_14238,N_14121,N_14094);
and U14239 (N_14239,N_14193,N_14168);
xor U14240 (N_14240,N_14083,N_14131);
or U14241 (N_14241,N_14134,N_14105);
nand U14242 (N_14242,N_14116,N_14065);
and U14243 (N_14243,N_14037,N_14127);
or U14244 (N_14244,N_14197,N_14126);
or U14245 (N_14245,N_14046,N_14172);
nor U14246 (N_14246,N_14075,N_14130);
nor U14247 (N_14247,N_14088,N_14138);
or U14248 (N_14248,N_14142,N_14111);
nor U14249 (N_14249,N_14098,N_14161);
xor U14250 (N_14250,N_14128,N_14085);
nor U14251 (N_14251,N_14021,N_14151);
xor U14252 (N_14252,N_14145,N_14101);
and U14253 (N_14253,N_14091,N_14139);
xnor U14254 (N_14254,N_14157,N_14019);
nor U14255 (N_14255,N_14066,N_14079);
xnor U14256 (N_14256,N_14071,N_14039);
xor U14257 (N_14257,N_14096,N_14023);
nand U14258 (N_14258,N_14095,N_14164);
xnor U14259 (N_14259,N_14173,N_14026);
and U14260 (N_14260,N_14144,N_14149);
nand U14261 (N_14261,N_14120,N_14158);
nand U14262 (N_14262,N_14143,N_14141);
and U14263 (N_14263,N_14051,N_14078);
nor U14264 (N_14264,N_14133,N_14177);
nand U14265 (N_14265,N_14054,N_14048);
and U14266 (N_14266,N_14050,N_14100);
and U14267 (N_14267,N_14063,N_14057);
xor U14268 (N_14268,N_14093,N_14070);
or U14269 (N_14269,N_14016,N_14185);
or U14270 (N_14270,N_14007,N_14045);
nor U14271 (N_14271,N_14009,N_14082);
nand U14272 (N_14272,N_14028,N_14015);
nor U14273 (N_14273,N_14001,N_14162);
xnor U14274 (N_14274,N_14018,N_14041);
xor U14275 (N_14275,N_14089,N_14069);
xnor U14276 (N_14276,N_14097,N_14073);
or U14277 (N_14277,N_14160,N_14153);
xor U14278 (N_14278,N_14114,N_14017);
or U14279 (N_14279,N_14102,N_14104);
and U14280 (N_14280,N_14106,N_14113);
nor U14281 (N_14281,N_14112,N_14188);
and U14282 (N_14282,N_14166,N_14176);
xor U14283 (N_14283,N_14198,N_14067);
nor U14284 (N_14284,N_14022,N_14034);
and U14285 (N_14285,N_14136,N_14006);
nor U14286 (N_14286,N_14042,N_14049);
nand U14287 (N_14287,N_14118,N_14003);
and U14288 (N_14288,N_14060,N_14077);
nand U14289 (N_14289,N_14196,N_14008);
or U14290 (N_14290,N_14152,N_14040);
nor U14291 (N_14291,N_14150,N_14092);
and U14292 (N_14292,N_14107,N_14137);
nand U14293 (N_14293,N_14043,N_14165);
nand U14294 (N_14294,N_14025,N_14190);
nand U14295 (N_14295,N_14194,N_14122);
xor U14296 (N_14296,N_14052,N_14181);
nand U14297 (N_14297,N_14044,N_14182);
and U14298 (N_14298,N_14013,N_14109);
xnor U14299 (N_14299,N_14056,N_14033);
nand U14300 (N_14300,N_14174,N_14070);
nor U14301 (N_14301,N_14091,N_14193);
nor U14302 (N_14302,N_14169,N_14129);
and U14303 (N_14303,N_14033,N_14096);
nor U14304 (N_14304,N_14117,N_14158);
xnor U14305 (N_14305,N_14061,N_14025);
and U14306 (N_14306,N_14125,N_14171);
and U14307 (N_14307,N_14090,N_14176);
and U14308 (N_14308,N_14149,N_14165);
xnor U14309 (N_14309,N_14076,N_14100);
xor U14310 (N_14310,N_14062,N_14191);
xor U14311 (N_14311,N_14083,N_14008);
nor U14312 (N_14312,N_14032,N_14099);
or U14313 (N_14313,N_14113,N_14024);
nand U14314 (N_14314,N_14093,N_14046);
nand U14315 (N_14315,N_14123,N_14190);
and U14316 (N_14316,N_14005,N_14075);
xor U14317 (N_14317,N_14014,N_14148);
nand U14318 (N_14318,N_14040,N_14051);
xor U14319 (N_14319,N_14130,N_14174);
or U14320 (N_14320,N_14132,N_14097);
xnor U14321 (N_14321,N_14151,N_14112);
xnor U14322 (N_14322,N_14082,N_14104);
nand U14323 (N_14323,N_14073,N_14118);
and U14324 (N_14324,N_14012,N_14149);
xnor U14325 (N_14325,N_14080,N_14015);
nor U14326 (N_14326,N_14015,N_14167);
or U14327 (N_14327,N_14058,N_14066);
xnor U14328 (N_14328,N_14138,N_14075);
and U14329 (N_14329,N_14173,N_14130);
and U14330 (N_14330,N_14144,N_14062);
and U14331 (N_14331,N_14113,N_14093);
xnor U14332 (N_14332,N_14009,N_14100);
and U14333 (N_14333,N_14053,N_14196);
or U14334 (N_14334,N_14140,N_14101);
xnor U14335 (N_14335,N_14143,N_14160);
nand U14336 (N_14336,N_14001,N_14048);
or U14337 (N_14337,N_14096,N_14055);
nand U14338 (N_14338,N_14024,N_14040);
or U14339 (N_14339,N_14036,N_14088);
and U14340 (N_14340,N_14157,N_14040);
xnor U14341 (N_14341,N_14165,N_14064);
nand U14342 (N_14342,N_14177,N_14170);
and U14343 (N_14343,N_14167,N_14162);
or U14344 (N_14344,N_14044,N_14175);
nand U14345 (N_14345,N_14016,N_14156);
or U14346 (N_14346,N_14054,N_14068);
or U14347 (N_14347,N_14127,N_14049);
xor U14348 (N_14348,N_14074,N_14165);
xnor U14349 (N_14349,N_14115,N_14182);
nor U14350 (N_14350,N_14078,N_14190);
or U14351 (N_14351,N_14021,N_14130);
and U14352 (N_14352,N_14025,N_14184);
nand U14353 (N_14353,N_14142,N_14156);
and U14354 (N_14354,N_14131,N_14031);
or U14355 (N_14355,N_14048,N_14130);
and U14356 (N_14356,N_14004,N_14037);
and U14357 (N_14357,N_14020,N_14005);
nand U14358 (N_14358,N_14054,N_14094);
nand U14359 (N_14359,N_14047,N_14005);
nand U14360 (N_14360,N_14110,N_14121);
or U14361 (N_14361,N_14122,N_14158);
and U14362 (N_14362,N_14045,N_14047);
or U14363 (N_14363,N_14140,N_14111);
or U14364 (N_14364,N_14069,N_14008);
nor U14365 (N_14365,N_14001,N_14104);
nor U14366 (N_14366,N_14044,N_14180);
or U14367 (N_14367,N_14017,N_14190);
and U14368 (N_14368,N_14076,N_14041);
nor U14369 (N_14369,N_14010,N_14133);
nand U14370 (N_14370,N_14146,N_14124);
nand U14371 (N_14371,N_14166,N_14153);
and U14372 (N_14372,N_14071,N_14186);
nor U14373 (N_14373,N_14151,N_14064);
or U14374 (N_14374,N_14139,N_14050);
nand U14375 (N_14375,N_14002,N_14097);
and U14376 (N_14376,N_14181,N_14147);
and U14377 (N_14377,N_14100,N_14143);
nand U14378 (N_14378,N_14079,N_14119);
and U14379 (N_14379,N_14080,N_14135);
nor U14380 (N_14380,N_14143,N_14117);
nor U14381 (N_14381,N_14069,N_14117);
and U14382 (N_14382,N_14009,N_14043);
or U14383 (N_14383,N_14161,N_14077);
and U14384 (N_14384,N_14039,N_14022);
nand U14385 (N_14385,N_14198,N_14072);
nand U14386 (N_14386,N_14139,N_14036);
nand U14387 (N_14387,N_14083,N_14021);
xnor U14388 (N_14388,N_14138,N_14129);
xor U14389 (N_14389,N_14095,N_14044);
and U14390 (N_14390,N_14120,N_14122);
nor U14391 (N_14391,N_14163,N_14112);
nor U14392 (N_14392,N_14096,N_14115);
xnor U14393 (N_14393,N_14036,N_14064);
and U14394 (N_14394,N_14180,N_14017);
xnor U14395 (N_14395,N_14083,N_14175);
nor U14396 (N_14396,N_14155,N_14077);
nor U14397 (N_14397,N_14051,N_14036);
and U14398 (N_14398,N_14003,N_14031);
nor U14399 (N_14399,N_14142,N_14092);
or U14400 (N_14400,N_14246,N_14257);
xnor U14401 (N_14401,N_14335,N_14342);
xor U14402 (N_14402,N_14368,N_14319);
xnor U14403 (N_14403,N_14226,N_14317);
and U14404 (N_14404,N_14337,N_14315);
and U14405 (N_14405,N_14268,N_14297);
nand U14406 (N_14406,N_14225,N_14375);
nand U14407 (N_14407,N_14380,N_14304);
or U14408 (N_14408,N_14330,N_14347);
xor U14409 (N_14409,N_14252,N_14237);
nor U14410 (N_14410,N_14314,N_14366);
or U14411 (N_14411,N_14200,N_14322);
nand U14412 (N_14412,N_14270,N_14321);
xnor U14413 (N_14413,N_14288,N_14229);
or U14414 (N_14414,N_14370,N_14326);
nand U14415 (N_14415,N_14308,N_14381);
nand U14416 (N_14416,N_14272,N_14302);
nor U14417 (N_14417,N_14286,N_14269);
xor U14418 (N_14418,N_14359,N_14307);
xor U14419 (N_14419,N_14350,N_14376);
nand U14420 (N_14420,N_14334,N_14336);
xnor U14421 (N_14421,N_14377,N_14239);
and U14422 (N_14422,N_14224,N_14203);
or U14423 (N_14423,N_14367,N_14389);
nor U14424 (N_14424,N_14396,N_14274);
nand U14425 (N_14425,N_14294,N_14217);
nand U14426 (N_14426,N_14213,N_14369);
or U14427 (N_14427,N_14220,N_14289);
xnor U14428 (N_14428,N_14324,N_14249);
xor U14429 (N_14429,N_14360,N_14339);
and U14430 (N_14430,N_14348,N_14373);
nand U14431 (N_14431,N_14386,N_14344);
nor U14432 (N_14432,N_14327,N_14388);
nand U14433 (N_14433,N_14259,N_14205);
or U14434 (N_14434,N_14346,N_14357);
nor U14435 (N_14435,N_14341,N_14230);
nor U14436 (N_14436,N_14299,N_14320);
or U14437 (N_14437,N_14206,N_14210);
and U14438 (N_14438,N_14353,N_14323);
nor U14439 (N_14439,N_14345,N_14361);
xor U14440 (N_14440,N_14312,N_14214);
or U14441 (N_14441,N_14232,N_14236);
xnor U14442 (N_14442,N_14278,N_14248);
or U14443 (N_14443,N_14378,N_14394);
or U14444 (N_14444,N_14242,N_14265);
xor U14445 (N_14445,N_14309,N_14395);
nor U14446 (N_14446,N_14250,N_14301);
or U14447 (N_14447,N_14273,N_14384);
xnor U14448 (N_14448,N_14393,N_14260);
or U14449 (N_14449,N_14362,N_14247);
and U14450 (N_14450,N_14328,N_14219);
and U14451 (N_14451,N_14208,N_14218);
or U14452 (N_14452,N_14284,N_14343);
nor U14453 (N_14453,N_14329,N_14238);
nor U14454 (N_14454,N_14349,N_14383);
or U14455 (N_14455,N_14233,N_14262);
or U14456 (N_14456,N_14385,N_14223);
and U14457 (N_14457,N_14333,N_14338);
xnor U14458 (N_14458,N_14212,N_14331);
nor U14459 (N_14459,N_14311,N_14363);
or U14460 (N_14460,N_14228,N_14234);
nor U14461 (N_14461,N_14221,N_14399);
xor U14462 (N_14462,N_14251,N_14372);
or U14463 (N_14463,N_14261,N_14258);
or U14464 (N_14464,N_14227,N_14209);
xnor U14465 (N_14465,N_14244,N_14392);
nor U14466 (N_14466,N_14266,N_14241);
and U14467 (N_14467,N_14263,N_14243);
xnor U14468 (N_14468,N_14313,N_14293);
nand U14469 (N_14469,N_14310,N_14295);
and U14470 (N_14470,N_14277,N_14254);
nand U14471 (N_14471,N_14398,N_14365);
and U14472 (N_14472,N_14255,N_14291);
and U14473 (N_14473,N_14292,N_14207);
xor U14474 (N_14474,N_14235,N_14300);
or U14475 (N_14475,N_14390,N_14264);
nor U14476 (N_14476,N_14256,N_14325);
or U14477 (N_14477,N_14283,N_14318);
xor U14478 (N_14478,N_14201,N_14316);
nand U14479 (N_14479,N_14276,N_14280);
and U14480 (N_14480,N_14374,N_14231);
or U14481 (N_14481,N_14211,N_14379);
xor U14482 (N_14482,N_14290,N_14303);
and U14483 (N_14483,N_14271,N_14281);
nor U14484 (N_14484,N_14354,N_14306);
nand U14485 (N_14485,N_14298,N_14371);
or U14486 (N_14486,N_14364,N_14282);
xnor U14487 (N_14487,N_14387,N_14204);
nand U14488 (N_14488,N_14279,N_14305);
xnor U14489 (N_14489,N_14382,N_14351);
nor U14490 (N_14490,N_14340,N_14356);
or U14491 (N_14491,N_14222,N_14245);
or U14492 (N_14492,N_14287,N_14216);
or U14493 (N_14493,N_14358,N_14332);
xnor U14494 (N_14494,N_14352,N_14391);
and U14495 (N_14495,N_14285,N_14267);
nor U14496 (N_14496,N_14397,N_14240);
and U14497 (N_14497,N_14355,N_14275);
nor U14498 (N_14498,N_14253,N_14296);
nand U14499 (N_14499,N_14202,N_14215);
and U14500 (N_14500,N_14338,N_14230);
or U14501 (N_14501,N_14352,N_14282);
nor U14502 (N_14502,N_14386,N_14304);
nand U14503 (N_14503,N_14261,N_14297);
nor U14504 (N_14504,N_14353,N_14236);
nand U14505 (N_14505,N_14380,N_14343);
or U14506 (N_14506,N_14383,N_14278);
or U14507 (N_14507,N_14357,N_14219);
xor U14508 (N_14508,N_14385,N_14216);
and U14509 (N_14509,N_14278,N_14345);
or U14510 (N_14510,N_14228,N_14239);
or U14511 (N_14511,N_14299,N_14237);
nor U14512 (N_14512,N_14247,N_14355);
nand U14513 (N_14513,N_14210,N_14250);
or U14514 (N_14514,N_14302,N_14364);
or U14515 (N_14515,N_14250,N_14345);
nand U14516 (N_14516,N_14204,N_14256);
xor U14517 (N_14517,N_14325,N_14226);
xnor U14518 (N_14518,N_14318,N_14294);
and U14519 (N_14519,N_14314,N_14284);
xor U14520 (N_14520,N_14206,N_14393);
nand U14521 (N_14521,N_14293,N_14288);
and U14522 (N_14522,N_14393,N_14268);
nor U14523 (N_14523,N_14285,N_14313);
and U14524 (N_14524,N_14388,N_14350);
and U14525 (N_14525,N_14244,N_14237);
and U14526 (N_14526,N_14392,N_14245);
nor U14527 (N_14527,N_14243,N_14350);
or U14528 (N_14528,N_14297,N_14274);
nor U14529 (N_14529,N_14393,N_14203);
xor U14530 (N_14530,N_14219,N_14334);
or U14531 (N_14531,N_14215,N_14356);
nor U14532 (N_14532,N_14203,N_14243);
or U14533 (N_14533,N_14236,N_14249);
or U14534 (N_14534,N_14363,N_14325);
nand U14535 (N_14535,N_14231,N_14288);
or U14536 (N_14536,N_14385,N_14322);
xnor U14537 (N_14537,N_14338,N_14292);
or U14538 (N_14538,N_14381,N_14391);
nand U14539 (N_14539,N_14294,N_14239);
and U14540 (N_14540,N_14393,N_14311);
and U14541 (N_14541,N_14339,N_14312);
nor U14542 (N_14542,N_14270,N_14286);
nand U14543 (N_14543,N_14376,N_14203);
xnor U14544 (N_14544,N_14302,N_14357);
xor U14545 (N_14545,N_14339,N_14286);
nand U14546 (N_14546,N_14293,N_14399);
nor U14547 (N_14547,N_14276,N_14271);
and U14548 (N_14548,N_14210,N_14287);
nand U14549 (N_14549,N_14298,N_14365);
xnor U14550 (N_14550,N_14265,N_14384);
nor U14551 (N_14551,N_14285,N_14291);
and U14552 (N_14552,N_14210,N_14319);
or U14553 (N_14553,N_14339,N_14357);
nor U14554 (N_14554,N_14207,N_14310);
nor U14555 (N_14555,N_14238,N_14259);
xnor U14556 (N_14556,N_14297,N_14276);
and U14557 (N_14557,N_14287,N_14259);
and U14558 (N_14558,N_14208,N_14226);
xnor U14559 (N_14559,N_14326,N_14344);
and U14560 (N_14560,N_14238,N_14282);
nor U14561 (N_14561,N_14389,N_14289);
and U14562 (N_14562,N_14295,N_14313);
xor U14563 (N_14563,N_14223,N_14370);
xor U14564 (N_14564,N_14347,N_14246);
nor U14565 (N_14565,N_14276,N_14334);
nand U14566 (N_14566,N_14342,N_14300);
nor U14567 (N_14567,N_14323,N_14233);
and U14568 (N_14568,N_14234,N_14223);
xor U14569 (N_14569,N_14299,N_14235);
and U14570 (N_14570,N_14214,N_14222);
or U14571 (N_14571,N_14238,N_14219);
nor U14572 (N_14572,N_14301,N_14331);
nor U14573 (N_14573,N_14221,N_14307);
or U14574 (N_14574,N_14360,N_14312);
nor U14575 (N_14575,N_14259,N_14378);
xnor U14576 (N_14576,N_14216,N_14266);
nor U14577 (N_14577,N_14282,N_14307);
nand U14578 (N_14578,N_14317,N_14217);
or U14579 (N_14579,N_14259,N_14279);
xnor U14580 (N_14580,N_14350,N_14266);
nand U14581 (N_14581,N_14313,N_14209);
and U14582 (N_14582,N_14303,N_14316);
or U14583 (N_14583,N_14260,N_14225);
and U14584 (N_14584,N_14346,N_14354);
and U14585 (N_14585,N_14280,N_14264);
and U14586 (N_14586,N_14378,N_14385);
xor U14587 (N_14587,N_14210,N_14321);
and U14588 (N_14588,N_14292,N_14277);
and U14589 (N_14589,N_14258,N_14380);
nand U14590 (N_14590,N_14367,N_14349);
xnor U14591 (N_14591,N_14310,N_14274);
and U14592 (N_14592,N_14339,N_14226);
nor U14593 (N_14593,N_14247,N_14376);
nand U14594 (N_14594,N_14318,N_14228);
nor U14595 (N_14595,N_14333,N_14295);
nand U14596 (N_14596,N_14252,N_14248);
and U14597 (N_14597,N_14204,N_14232);
and U14598 (N_14598,N_14346,N_14272);
and U14599 (N_14599,N_14258,N_14256);
nor U14600 (N_14600,N_14417,N_14454);
or U14601 (N_14601,N_14523,N_14515);
nor U14602 (N_14602,N_14536,N_14555);
nor U14603 (N_14603,N_14548,N_14576);
and U14604 (N_14604,N_14457,N_14443);
nor U14605 (N_14605,N_14505,N_14442);
or U14606 (N_14606,N_14456,N_14403);
nor U14607 (N_14607,N_14549,N_14534);
and U14608 (N_14608,N_14563,N_14430);
nor U14609 (N_14609,N_14463,N_14537);
nor U14610 (N_14610,N_14528,N_14583);
or U14611 (N_14611,N_14424,N_14479);
nor U14612 (N_14612,N_14402,N_14520);
nor U14613 (N_14613,N_14480,N_14513);
nand U14614 (N_14614,N_14579,N_14511);
xor U14615 (N_14615,N_14438,N_14452);
nor U14616 (N_14616,N_14478,N_14444);
and U14617 (N_14617,N_14560,N_14406);
or U14618 (N_14618,N_14578,N_14539);
xor U14619 (N_14619,N_14545,N_14447);
nor U14620 (N_14620,N_14477,N_14464);
xnor U14621 (N_14621,N_14497,N_14459);
nand U14622 (N_14622,N_14556,N_14519);
nand U14623 (N_14623,N_14569,N_14493);
and U14624 (N_14624,N_14400,N_14449);
nand U14625 (N_14625,N_14518,N_14465);
nor U14626 (N_14626,N_14461,N_14469);
nor U14627 (N_14627,N_14504,N_14485);
nand U14628 (N_14628,N_14582,N_14496);
or U14629 (N_14629,N_14408,N_14494);
or U14630 (N_14630,N_14423,N_14506);
or U14631 (N_14631,N_14595,N_14597);
or U14632 (N_14632,N_14517,N_14557);
xnor U14633 (N_14633,N_14592,N_14572);
nor U14634 (N_14634,N_14413,N_14487);
nor U14635 (N_14635,N_14470,N_14587);
nor U14636 (N_14636,N_14552,N_14481);
nor U14637 (N_14637,N_14498,N_14410);
nand U14638 (N_14638,N_14492,N_14526);
or U14639 (N_14639,N_14577,N_14516);
nor U14640 (N_14640,N_14596,N_14524);
nand U14641 (N_14641,N_14483,N_14565);
nand U14642 (N_14642,N_14467,N_14441);
nand U14643 (N_14643,N_14472,N_14440);
nand U14644 (N_14644,N_14588,N_14418);
nand U14645 (N_14645,N_14414,N_14509);
nand U14646 (N_14646,N_14439,N_14409);
and U14647 (N_14647,N_14405,N_14566);
or U14648 (N_14648,N_14431,N_14543);
nor U14649 (N_14649,N_14574,N_14546);
nor U14650 (N_14650,N_14571,N_14599);
or U14651 (N_14651,N_14491,N_14471);
xor U14652 (N_14652,N_14458,N_14422);
nand U14653 (N_14653,N_14550,N_14529);
and U14654 (N_14654,N_14462,N_14475);
or U14655 (N_14655,N_14562,N_14530);
and U14656 (N_14656,N_14553,N_14538);
xnor U14657 (N_14657,N_14581,N_14584);
nor U14658 (N_14658,N_14434,N_14568);
nand U14659 (N_14659,N_14598,N_14547);
or U14660 (N_14660,N_14446,N_14567);
nor U14661 (N_14661,N_14535,N_14476);
nor U14662 (N_14662,N_14450,N_14484);
or U14663 (N_14663,N_14429,N_14580);
nor U14664 (N_14664,N_14575,N_14489);
or U14665 (N_14665,N_14416,N_14522);
or U14666 (N_14666,N_14542,N_14426);
xnor U14667 (N_14667,N_14503,N_14420);
and U14668 (N_14668,N_14512,N_14573);
nor U14669 (N_14669,N_14590,N_14499);
or U14670 (N_14670,N_14533,N_14421);
or U14671 (N_14671,N_14564,N_14482);
nand U14672 (N_14672,N_14593,N_14558);
nand U14673 (N_14673,N_14428,N_14521);
or U14674 (N_14674,N_14453,N_14540);
nand U14675 (N_14675,N_14466,N_14591);
nand U14676 (N_14676,N_14570,N_14433);
nor U14677 (N_14677,N_14488,N_14427);
or U14678 (N_14678,N_14527,N_14445);
nor U14679 (N_14679,N_14525,N_14532);
xnor U14680 (N_14680,N_14561,N_14554);
nand U14681 (N_14681,N_14436,N_14486);
xnor U14682 (N_14682,N_14551,N_14586);
nand U14683 (N_14683,N_14412,N_14455);
nor U14684 (N_14684,N_14502,N_14425);
and U14685 (N_14685,N_14507,N_14490);
nor U14686 (N_14686,N_14589,N_14585);
and U14687 (N_14687,N_14468,N_14435);
or U14688 (N_14688,N_14473,N_14411);
nor U14689 (N_14689,N_14401,N_14501);
xnor U14690 (N_14690,N_14415,N_14531);
nand U14691 (N_14691,N_14419,N_14508);
xnor U14692 (N_14692,N_14544,N_14500);
xor U14693 (N_14693,N_14432,N_14448);
nor U14694 (N_14694,N_14594,N_14404);
nor U14695 (N_14695,N_14474,N_14495);
or U14696 (N_14696,N_14541,N_14407);
xor U14697 (N_14697,N_14559,N_14510);
nor U14698 (N_14698,N_14460,N_14514);
nand U14699 (N_14699,N_14451,N_14437);
and U14700 (N_14700,N_14464,N_14469);
nand U14701 (N_14701,N_14509,N_14524);
nand U14702 (N_14702,N_14571,N_14417);
nor U14703 (N_14703,N_14518,N_14466);
xor U14704 (N_14704,N_14591,N_14595);
nand U14705 (N_14705,N_14497,N_14471);
nor U14706 (N_14706,N_14480,N_14581);
nand U14707 (N_14707,N_14487,N_14525);
or U14708 (N_14708,N_14498,N_14462);
or U14709 (N_14709,N_14431,N_14598);
xnor U14710 (N_14710,N_14486,N_14574);
and U14711 (N_14711,N_14590,N_14418);
and U14712 (N_14712,N_14596,N_14435);
or U14713 (N_14713,N_14552,N_14569);
and U14714 (N_14714,N_14571,N_14513);
xnor U14715 (N_14715,N_14432,N_14576);
or U14716 (N_14716,N_14497,N_14540);
xnor U14717 (N_14717,N_14497,N_14587);
and U14718 (N_14718,N_14480,N_14520);
xnor U14719 (N_14719,N_14585,N_14503);
and U14720 (N_14720,N_14563,N_14493);
nand U14721 (N_14721,N_14553,N_14440);
xnor U14722 (N_14722,N_14596,N_14463);
or U14723 (N_14723,N_14402,N_14504);
and U14724 (N_14724,N_14544,N_14485);
nand U14725 (N_14725,N_14489,N_14502);
nor U14726 (N_14726,N_14551,N_14573);
xor U14727 (N_14727,N_14488,N_14452);
and U14728 (N_14728,N_14464,N_14448);
nor U14729 (N_14729,N_14459,N_14480);
and U14730 (N_14730,N_14525,N_14478);
or U14731 (N_14731,N_14400,N_14548);
or U14732 (N_14732,N_14583,N_14525);
or U14733 (N_14733,N_14559,N_14419);
xnor U14734 (N_14734,N_14552,N_14532);
nand U14735 (N_14735,N_14554,N_14572);
or U14736 (N_14736,N_14462,N_14465);
and U14737 (N_14737,N_14549,N_14494);
xnor U14738 (N_14738,N_14533,N_14491);
or U14739 (N_14739,N_14418,N_14475);
xor U14740 (N_14740,N_14512,N_14417);
and U14741 (N_14741,N_14464,N_14400);
nor U14742 (N_14742,N_14437,N_14554);
or U14743 (N_14743,N_14497,N_14461);
or U14744 (N_14744,N_14440,N_14546);
and U14745 (N_14745,N_14584,N_14403);
xnor U14746 (N_14746,N_14430,N_14558);
and U14747 (N_14747,N_14505,N_14477);
nand U14748 (N_14748,N_14477,N_14409);
and U14749 (N_14749,N_14547,N_14562);
and U14750 (N_14750,N_14422,N_14441);
or U14751 (N_14751,N_14519,N_14467);
nand U14752 (N_14752,N_14419,N_14536);
nand U14753 (N_14753,N_14428,N_14534);
nand U14754 (N_14754,N_14535,N_14401);
nor U14755 (N_14755,N_14460,N_14498);
nor U14756 (N_14756,N_14418,N_14477);
xnor U14757 (N_14757,N_14512,N_14548);
and U14758 (N_14758,N_14501,N_14515);
xor U14759 (N_14759,N_14495,N_14528);
xor U14760 (N_14760,N_14559,N_14452);
xnor U14761 (N_14761,N_14559,N_14470);
nand U14762 (N_14762,N_14474,N_14575);
or U14763 (N_14763,N_14453,N_14459);
nand U14764 (N_14764,N_14580,N_14442);
nor U14765 (N_14765,N_14453,N_14429);
nor U14766 (N_14766,N_14534,N_14556);
and U14767 (N_14767,N_14474,N_14589);
xnor U14768 (N_14768,N_14457,N_14413);
and U14769 (N_14769,N_14598,N_14571);
nand U14770 (N_14770,N_14405,N_14471);
nand U14771 (N_14771,N_14517,N_14550);
or U14772 (N_14772,N_14435,N_14478);
nor U14773 (N_14773,N_14595,N_14546);
xnor U14774 (N_14774,N_14560,N_14516);
nand U14775 (N_14775,N_14582,N_14476);
xor U14776 (N_14776,N_14551,N_14470);
nor U14777 (N_14777,N_14455,N_14553);
or U14778 (N_14778,N_14474,N_14502);
xnor U14779 (N_14779,N_14555,N_14566);
xnor U14780 (N_14780,N_14584,N_14438);
nor U14781 (N_14781,N_14407,N_14445);
nor U14782 (N_14782,N_14480,N_14468);
xnor U14783 (N_14783,N_14460,N_14453);
and U14784 (N_14784,N_14554,N_14505);
or U14785 (N_14785,N_14427,N_14467);
or U14786 (N_14786,N_14544,N_14482);
nand U14787 (N_14787,N_14567,N_14419);
nor U14788 (N_14788,N_14509,N_14578);
xor U14789 (N_14789,N_14471,N_14579);
nor U14790 (N_14790,N_14472,N_14599);
xnor U14791 (N_14791,N_14549,N_14544);
xnor U14792 (N_14792,N_14451,N_14456);
or U14793 (N_14793,N_14478,N_14496);
xor U14794 (N_14794,N_14544,N_14574);
nand U14795 (N_14795,N_14472,N_14423);
and U14796 (N_14796,N_14587,N_14570);
or U14797 (N_14797,N_14580,N_14582);
nand U14798 (N_14798,N_14584,N_14598);
xor U14799 (N_14799,N_14550,N_14504);
or U14800 (N_14800,N_14706,N_14771);
nand U14801 (N_14801,N_14776,N_14740);
xnor U14802 (N_14802,N_14753,N_14622);
xnor U14803 (N_14803,N_14674,N_14619);
and U14804 (N_14804,N_14640,N_14729);
or U14805 (N_14805,N_14726,N_14767);
nor U14806 (N_14806,N_14617,N_14690);
xnor U14807 (N_14807,N_14708,N_14782);
nand U14808 (N_14808,N_14737,N_14724);
nand U14809 (N_14809,N_14607,N_14645);
and U14810 (N_14810,N_14697,N_14676);
or U14811 (N_14811,N_14758,N_14765);
or U14812 (N_14812,N_14675,N_14734);
or U14813 (N_14813,N_14716,N_14602);
or U14814 (N_14814,N_14732,N_14608);
nor U14815 (N_14815,N_14727,N_14793);
nand U14816 (N_14816,N_14777,N_14685);
nand U14817 (N_14817,N_14651,N_14684);
or U14818 (N_14818,N_14789,N_14760);
nand U14819 (N_14819,N_14612,N_14621);
and U14820 (N_14820,N_14717,N_14719);
and U14821 (N_14821,N_14795,N_14731);
and U14822 (N_14822,N_14628,N_14683);
and U14823 (N_14823,N_14616,N_14764);
nand U14824 (N_14824,N_14714,N_14720);
nand U14825 (N_14825,N_14643,N_14703);
or U14826 (N_14826,N_14604,N_14678);
nor U14827 (N_14827,N_14794,N_14680);
xor U14828 (N_14828,N_14610,N_14664);
and U14829 (N_14829,N_14766,N_14774);
or U14830 (N_14830,N_14712,N_14642);
and U14831 (N_14831,N_14759,N_14723);
nand U14832 (N_14832,N_14705,N_14701);
or U14833 (N_14833,N_14606,N_14728);
xor U14834 (N_14834,N_14632,N_14745);
nor U14835 (N_14835,N_14788,N_14662);
nor U14836 (N_14836,N_14634,N_14641);
nand U14837 (N_14837,N_14689,N_14784);
nor U14838 (N_14838,N_14688,N_14786);
and U14839 (N_14839,N_14624,N_14707);
xnor U14840 (N_14840,N_14635,N_14778);
nand U14841 (N_14841,N_14791,N_14768);
and U14842 (N_14842,N_14633,N_14679);
xor U14843 (N_14843,N_14785,N_14748);
and U14844 (N_14844,N_14646,N_14755);
or U14845 (N_14845,N_14751,N_14790);
xor U14846 (N_14846,N_14709,N_14681);
or U14847 (N_14847,N_14620,N_14653);
nor U14848 (N_14848,N_14658,N_14629);
xor U14849 (N_14849,N_14715,N_14711);
nor U14850 (N_14850,N_14757,N_14738);
nor U14851 (N_14851,N_14743,N_14770);
or U14852 (N_14852,N_14694,N_14747);
or U14853 (N_14853,N_14603,N_14721);
nand U14854 (N_14854,N_14781,N_14625);
nand U14855 (N_14855,N_14611,N_14601);
nand U14856 (N_14856,N_14605,N_14775);
and U14857 (N_14857,N_14704,N_14691);
or U14858 (N_14858,N_14735,N_14693);
or U14859 (N_14859,N_14773,N_14700);
nand U14860 (N_14860,N_14698,N_14673);
nand U14861 (N_14861,N_14600,N_14626);
xnor U14862 (N_14862,N_14722,N_14744);
nor U14863 (N_14863,N_14687,N_14739);
or U14864 (N_14864,N_14761,N_14670);
or U14865 (N_14865,N_14615,N_14686);
and U14866 (N_14866,N_14654,N_14779);
or U14867 (N_14867,N_14730,N_14652);
nand U14868 (N_14868,N_14677,N_14752);
nand U14869 (N_14869,N_14710,N_14613);
or U14870 (N_14870,N_14798,N_14783);
nand U14871 (N_14871,N_14671,N_14682);
xor U14872 (N_14872,N_14647,N_14754);
and U14873 (N_14873,N_14756,N_14648);
nor U14874 (N_14874,N_14742,N_14787);
xnor U14875 (N_14875,N_14702,N_14725);
nand U14876 (N_14876,N_14733,N_14746);
xnor U14877 (N_14877,N_14796,N_14660);
nor U14878 (N_14878,N_14762,N_14695);
nand U14879 (N_14879,N_14638,N_14659);
nor U14880 (N_14880,N_14699,N_14665);
nand U14881 (N_14881,N_14792,N_14780);
or U14882 (N_14882,N_14772,N_14799);
or U14883 (N_14883,N_14750,N_14672);
xor U14884 (N_14884,N_14741,N_14630);
xor U14885 (N_14885,N_14639,N_14644);
xnor U14886 (N_14886,N_14713,N_14657);
nor U14887 (N_14887,N_14627,N_14696);
nor U14888 (N_14888,N_14614,N_14769);
nor U14889 (N_14889,N_14669,N_14797);
nor U14890 (N_14890,N_14623,N_14668);
or U14891 (N_14891,N_14656,N_14667);
or U14892 (N_14892,N_14763,N_14649);
nor U14893 (N_14893,N_14655,N_14661);
nor U14894 (N_14894,N_14663,N_14692);
nor U14895 (N_14895,N_14666,N_14650);
nor U14896 (N_14896,N_14718,N_14736);
xnor U14897 (N_14897,N_14631,N_14749);
nand U14898 (N_14898,N_14637,N_14609);
or U14899 (N_14899,N_14618,N_14636);
or U14900 (N_14900,N_14722,N_14781);
nor U14901 (N_14901,N_14642,N_14696);
xor U14902 (N_14902,N_14642,N_14682);
or U14903 (N_14903,N_14603,N_14632);
and U14904 (N_14904,N_14705,N_14609);
xor U14905 (N_14905,N_14798,N_14732);
and U14906 (N_14906,N_14770,N_14722);
and U14907 (N_14907,N_14722,N_14608);
or U14908 (N_14908,N_14627,N_14640);
nand U14909 (N_14909,N_14755,N_14635);
or U14910 (N_14910,N_14679,N_14645);
nand U14911 (N_14911,N_14651,N_14647);
xnor U14912 (N_14912,N_14744,N_14794);
or U14913 (N_14913,N_14770,N_14677);
nand U14914 (N_14914,N_14768,N_14770);
and U14915 (N_14915,N_14699,N_14661);
or U14916 (N_14916,N_14685,N_14761);
xnor U14917 (N_14917,N_14659,N_14793);
nor U14918 (N_14918,N_14709,N_14707);
nor U14919 (N_14919,N_14629,N_14716);
or U14920 (N_14920,N_14674,N_14740);
nand U14921 (N_14921,N_14762,N_14655);
xnor U14922 (N_14922,N_14640,N_14775);
and U14923 (N_14923,N_14681,N_14767);
nor U14924 (N_14924,N_14745,N_14656);
and U14925 (N_14925,N_14675,N_14639);
and U14926 (N_14926,N_14758,N_14707);
nor U14927 (N_14927,N_14792,N_14679);
nand U14928 (N_14928,N_14691,N_14709);
nand U14929 (N_14929,N_14687,N_14778);
xnor U14930 (N_14930,N_14749,N_14694);
nor U14931 (N_14931,N_14678,N_14725);
or U14932 (N_14932,N_14781,N_14708);
and U14933 (N_14933,N_14775,N_14756);
nor U14934 (N_14934,N_14745,N_14648);
and U14935 (N_14935,N_14731,N_14791);
nor U14936 (N_14936,N_14641,N_14796);
and U14937 (N_14937,N_14716,N_14679);
or U14938 (N_14938,N_14617,N_14619);
xor U14939 (N_14939,N_14649,N_14772);
xor U14940 (N_14940,N_14664,N_14696);
nor U14941 (N_14941,N_14620,N_14708);
and U14942 (N_14942,N_14612,N_14783);
and U14943 (N_14943,N_14768,N_14625);
nor U14944 (N_14944,N_14767,N_14600);
nand U14945 (N_14945,N_14619,N_14676);
xnor U14946 (N_14946,N_14699,N_14771);
nor U14947 (N_14947,N_14727,N_14652);
or U14948 (N_14948,N_14772,N_14715);
xor U14949 (N_14949,N_14713,N_14641);
nand U14950 (N_14950,N_14705,N_14789);
and U14951 (N_14951,N_14683,N_14711);
xor U14952 (N_14952,N_14620,N_14717);
nor U14953 (N_14953,N_14750,N_14690);
and U14954 (N_14954,N_14796,N_14795);
nor U14955 (N_14955,N_14757,N_14771);
nand U14956 (N_14956,N_14666,N_14619);
or U14957 (N_14957,N_14757,N_14634);
xnor U14958 (N_14958,N_14696,N_14782);
xor U14959 (N_14959,N_14613,N_14614);
nor U14960 (N_14960,N_14764,N_14608);
and U14961 (N_14961,N_14778,N_14791);
or U14962 (N_14962,N_14693,N_14633);
nand U14963 (N_14963,N_14670,N_14750);
nor U14964 (N_14964,N_14711,N_14648);
and U14965 (N_14965,N_14650,N_14750);
or U14966 (N_14966,N_14666,N_14636);
or U14967 (N_14967,N_14625,N_14760);
nand U14968 (N_14968,N_14786,N_14737);
and U14969 (N_14969,N_14652,N_14742);
nor U14970 (N_14970,N_14775,N_14690);
nand U14971 (N_14971,N_14619,N_14682);
xor U14972 (N_14972,N_14653,N_14702);
xor U14973 (N_14973,N_14733,N_14615);
and U14974 (N_14974,N_14735,N_14668);
nand U14975 (N_14975,N_14628,N_14675);
nand U14976 (N_14976,N_14766,N_14670);
nand U14977 (N_14977,N_14736,N_14784);
nand U14978 (N_14978,N_14631,N_14752);
or U14979 (N_14979,N_14625,N_14670);
nor U14980 (N_14980,N_14634,N_14769);
xnor U14981 (N_14981,N_14771,N_14664);
and U14982 (N_14982,N_14623,N_14797);
and U14983 (N_14983,N_14674,N_14638);
xor U14984 (N_14984,N_14715,N_14641);
nand U14985 (N_14985,N_14747,N_14775);
nor U14986 (N_14986,N_14648,N_14762);
and U14987 (N_14987,N_14760,N_14657);
nor U14988 (N_14988,N_14635,N_14740);
or U14989 (N_14989,N_14643,N_14787);
and U14990 (N_14990,N_14641,N_14624);
nand U14991 (N_14991,N_14687,N_14645);
nand U14992 (N_14992,N_14659,N_14709);
xnor U14993 (N_14993,N_14639,N_14728);
nor U14994 (N_14994,N_14741,N_14715);
nor U14995 (N_14995,N_14639,N_14770);
nor U14996 (N_14996,N_14728,N_14772);
nor U14997 (N_14997,N_14686,N_14614);
or U14998 (N_14998,N_14690,N_14666);
or U14999 (N_14999,N_14707,N_14628);
or U15000 (N_15000,N_14813,N_14881);
nor U15001 (N_15001,N_14822,N_14895);
xnor U15002 (N_15002,N_14913,N_14814);
or U15003 (N_15003,N_14876,N_14852);
and U15004 (N_15004,N_14992,N_14968);
nand U15005 (N_15005,N_14937,N_14975);
nor U15006 (N_15006,N_14931,N_14907);
or U15007 (N_15007,N_14888,N_14811);
nor U15008 (N_15008,N_14862,N_14824);
xnor U15009 (N_15009,N_14879,N_14863);
nor U15010 (N_15010,N_14982,N_14926);
and U15011 (N_15011,N_14976,N_14987);
or U15012 (N_15012,N_14918,N_14851);
nand U15013 (N_15013,N_14939,N_14991);
nand U15014 (N_15014,N_14836,N_14981);
or U15015 (N_15015,N_14940,N_14845);
and U15016 (N_15016,N_14864,N_14807);
or U15017 (N_15017,N_14848,N_14821);
nand U15018 (N_15018,N_14949,N_14816);
and U15019 (N_15019,N_14901,N_14817);
nand U15020 (N_15020,N_14983,N_14887);
nand U15021 (N_15021,N_14819,N_14954);
nor U15022 (N_15022,N_14833,N_14906);
xor U15023 (N_15023,N_14815,N_14843);
nor U15024 (N_15024,N_14962,N_14915);
xnor U15025 (N_15025,N_14800,N_14917);
nand U15026 (N_15026,N_14969,N_14927);
nand U15027 (N_15027,N_14946,N_14856);
nor U15028 (N_15028,N_14990,N_14827);
nor U15029 (N_15029,N_14844,N_14942);
nand U15030 (N_15030,N_14932,N_14920);
and U15031 (N_15031,N_14874,N_14938);
nand U15032 (N_15032,N_14867,N_14994);
nand U15033 (N_15033,N_14870,N_14979);
or U15034 (N_15034,N_14802,N_14829);
and U15035 (N_15035,N_14971,N_14997);
or U15036 (N_15036,N_14914,N_14869);
or U15037 (N_15037,N_14880,N_14803);
nor U15038 (N_15038,N_14999,N_14903);
xor U15039 (N_15039,N_14908,N_14995);
and U15040 (N_15040,N_14890,N_14849);
nand U15041 (N_15041,N_14952,N_14871);
or U15042 (N_15042,N_14825,N_14974);
xor U15043 (N_15043,N_14893,N_14985);
nand U15044 (N_15044,N_14841,N_14905);
nand U15045 (N_15045,N_14978,N_14839);
xnor U15046 (N_15046,N_14892,N_14910);
nor U15047 (N_15047,N_14970,N_14959);
nor U15048 (N_15048,N_14935,N_14897);
nor U15049 (N_15049,N_14808,N_14947);
xor U15050 (N_15050,N_14891,N_14826);
xor U15051 (N_15051,N_14916,N_14872);
nand U15052 (N_15052,N_14837,N_14957);
nor U15053 (N_15053,N_14878,N_14933);
and U15054 (N_15054,N_14928,N_14885);
nand U15055 (N_15055,N_14919,N_14832);
nor U15056 (N_15056,N_14823,N_14854);
or U15057 (N_15057,N_14934,N_14865);
nor U15058 (N_15058,N_14973,N_14801);
or U15059 (N_15059,N_14896,N_14950);
or U15060 (N_15060,N_14830,N_14923);
xor U15061 (N_15061,N_14964,N_14853);
nand U15062 (N_15062,N_14929,N_14850);
nand U15063 (N_15063,N_14912,N_14840);
xnor U15064 (N_15064,N_14894,N_14804);
nand U15065 (N_15065,N_14967,N_14868);
xor U15066 (N_15066,N_14960,N_14948);
nor U15067 (N_15067,N_14805,N_14904);
or U15068 (N_15068,N_14831,N_14882);
nor U15069 (N_15069,N_14922,N_14941);
and U15070 (N_15070,N_14958,N_14810);
and U15071 (N_15071,N_14911,N_14921);
or U15072 (N_15072,N_14861,N_14834);
and U15073 (N_15073,N_14989,N_14838);
and U15074 (N_15074,N_14820,N_14944);
or U15075 (N_15075,N_14902,N_14961);
and U15076 (N_15076,N_14980,N_14998);
xnor U15077 (N_15077,N_14889,N_14835);
nand U15078 (N_15078,N_14809,N_14812);
or U15079 (N_15079,N_14873,N_14858);
nor U15080 (N_15080,N_14988,N_14936);
xnor U15081 (N_15081,N_14886,N_14866);
or U15082 (N_15082,N_14984,N_14898);
nand U15083 (N_15083,N_14828,N_14818);
nor U15084 (N_15084,N_14884,N_14966);
or U15085 (N_15085,N_14925,N_14875);
nand U15086 (N_15086,N_14924,N_14842);
nor U15087 (N_15087,N_14956,N_14846);
nor U15088 (N_15088,N_14972,N_14806);
nand U15089 (N_15089,N_14859,N_14977);
xnor U15090 (N_15090,N_14945,N_14996);
xor U15091 (N_15091,N_14951,N_14857);
or U15092 (N_15092,N_14955,N_14855);
nand U15093 (N_15093,N_14953,N_14963);
xor U15094 (N_15094,N_14883,N_14930);
nand U15095 (N_15095,N_14900,N_14877);
xnor U15096 (N_15096,N_14847,N_14909);
nand U15097 (N_15097,N_14899,N_14943);
nor U15098 (N_15098,N_14860,N_14986);
xor U15099 (N_15099,N_14965,N_14993);
nand U15100 (N_15100,N_14960,N_14812);
nor U15101 (N_15101,N_14807,N_14921);
nand U15102 (N_15102,N_14822,N_14851);
xor U15103 (N_15103,N_14847,N_14984);
nand U15104 (N_15104,N_14933,N_14842);
nand U15105 (N_15105,N_14981,N_14976);
nand U15106 (N_15106,N_14998,N_14883);
and U15107 (N_15107,N_14964,N_14899);
nor U15108 (N_15108,N_14812,N_14800);
nor U15109 (N_15109,N_14953,N_14986);
or U15110 (N_15110,N_14942,N_14990);
nor U15111 (N_15111,N_14882,N_14822);
nand U15112 (N_15112,N_14878,N_14829);
nand U15113 (N_15113,N_14850,N_14807);
or U15114 (N_15114,N_14888,N_14804);
xnor U15115 (N_15115,N_14811,N_14920);
nor U15116 (N_15116,N_14961,N_14863);
xor U15117 (N_15117,N_14947,N_14826);
xnor U15118 (N_15118,N_14954,N_14912);
nand U15119 (N_15119,N_14996,N_14863);
xor U15120 (N_15120,N_14915,N_14946);
xnor U15121 (N_15121,N_14953,N_14867);
nand U15122 (N_15122,N_14809,N_14895);
xnor U15123 (N_15123,N_14946,N_14880);
xnor U15124 (N_15124,N_14903,N_14957);
or U15125 (N_15125,N_14968,N_14976);
and U15126 (N_15126,N_14980,N_14971);
nor U15127 (N_15127,N_14828,N_14842);
or U15128 (N_15128,N_14804,N_14830);
nand U15129 (N_15129,N_14901,N_14863);
nor U15130 (N_15130,N_14989,N_14900);
or U15131 (N_15131,N_14915,N_14846);
or U15132 (N_15132,N_14852,N_14866);
nor U15133 (N_15133,N_14974,N_14870);
and U15134 (N_15134,N_14975,N_14953);
nand U15135 (N_15135,N_14911,N_14828);
nor U15136 (N_15136,N_14954,N_14888);
or U15137 (N_15137,N_14933,N_14911);
xnor U15138 (N_15138,N_14928,N_14956);
nand U15139 (N_15139,N_14830,N_14956);
or U15140 (N_15140,N_14930,N_14841);
xnor U15141 (N_15141,N_14826,N_14945);
nor U15142 (N_15142,N_14941,N_14934);
and U15143 (N_15143,N_14963,N_14895);
or U15144 (N_15144,N_14853,N_14888);
nor U15145 (N_15145,N_14813,N_14820);
nand U15146 (N_15146,N_14896,N_14918);
xnor U15147 (N_15147,N_14954,N_14898);
or U15148 (N_15148,N_14824,N_14983);
nor U15149 (N_15149,N_14992,N_14827);
nor U15150 (N_15150,N_14961,N_14901);
nor U15151 (N_15151,N_14960,N_14973);
nand U15152 (N_15152,N_14861,N_14987);
xnor U15153 (N_15153,N_14834,N_14805);
and U15154 (N_15154,N_14802,N_14862);
xnor U15155 (N_15155,N_14823,N_14948);
nor U15156 (N_15156,N_14854,N_14803);
and U15157 (N_15157,N_14841,N_14885);
xor U15158 (N_15158,N_14819,N_14843);
xor U15159 (N_15159,N_14910,N_14847);
nor U15160 (N_15160,N_14972,N_14905);
and U15161 (N_15161,N_14941,N_14801);
nand U15162 (N_15162,N_14841,N_14842);
or U15163 (N_15163,N_14902,N_14904);
and U15164 (N_15164,N_14989,N_14998);
xnor U15165 (N_15165,N_14887,N_14839);
nand U15166 (N_15166,N_14829,N_14819);
xnor U15167 (N_15167,N_14998,N_14840);
xor U15168 (N_15168,N_14953,N_14808);
nand U15169 (N_15169,N_14967,N_14845);
nor U15170 (N_15170,N_14839,N_14958);
and U15171 (N_15171,N_14932,N_14843);
nand U15172 (N_15172,N_14953,N_14928);
nor U15173 (N_15173,N_14904,N_14847);
nand U15174 (N_15174,N_14944,N_14889);
and U15175 (N_15175,N_14891,N_14881);
nand U15176 (N_15176,N_14934,N_14848);
nor U15177 (N_15177,N_14900,N_14815);
nand U15178 (N_15178,N_14819,N_14854);
or U15179 (N_15179,N_14898,N_14861);
nor U15180 (N_15180,N_14809,N_14948);
nor U15181 (N_15181,N_14953,N_14945);
nand U15182 (N_15182,N_14941,N_14903);
xnor U15183 (N_15183,N_14938,N_14822);
nor U15184 (N_15184,N_14881,N_14939);
xnor U15185 (N_15185,N_14893,N_14854);
or U15186 (N_15186,N_14818,N_14922);
nor U15187 (N_15187,N_14840,N_14922);
xnor U15188 (N_15188,N_14899,N_14824);
or U15189 (N_15189,N_14816,N_14839);
nand U15190 (N_15190,N_14952,N_14856);
nor U15191 (N_15191,N_14826,N_14930);
nand U15192 (N_15192,N_14903,N_14938);
or U15193 (N_15193,N_14988,N_14917);
nand U15194 (N_15194,N_14821,N_14938);
and U15195 (N_15195,N_14980,N_14871);
xnor U15196 (N_15196,N_14999,N_14824);
nand U15197 (N_15197,N_14813,N_14839);
or U15198 (N_15198,N_14822,N_14923);
nand U15199 (N_15199,N_14899,N_14981);
and U15200 (N_15200,N_15165,N_15111);
nor U15201 (N_15201,N_15002,N_15058);
and U15202 (N_15202,N_15145,N_15160);
or U15203 (N_15203,N_15095,N_15161);
xor U15204 (N_15204,N_15078,N_15043);
and U15205 (N_15205,N_15031,N_15101);
nor U15206 (N_15206,N_15060,N_15036);
or U15207 (N_15207,N_15026,N_15173);
xnor U15208 (N_15208,N_15088,N_15087);
or U15209 (N_15209,N_15077,N_15110);
or U15210 (N_15210,N_15039,N_15146);
nor U15211 (N_15211,N_15148,N_15038);
or U15212 (N_15212,N_15041,N_15167);
xor U15213 (N_15213,N_15090,N_15169);
or U15214 (N_15214,N_15108,N_15092);
nor U15215 (N_15215,N_15125,N_15079);
nand U15216 (N_15216,N_15183,N_15109);
xor U15217 (N_15217,N_15118,N_15071);
nor U15218 (N_15218,N_15047,N_15127);
xor U15219 (N_15219,N_15054,N_15184);
and U15220 (N_15220,N_15138,N_15164);
and U15221 (N_15221,N_15018,N_15170);
or U15222 (N_15222,N_15176,N_15191);
and U15223 (N_15223,N_15162,N_15102);
xor U15224 (N_15224,N_15012,N_15010);
or U15225 (N_15225,N_15113,N_15051);
and U15226 (N_15226,N_15032,N_15159);
and U15227 (N_15227,N_15030,N_15197);
or U15228 (N_15228,N_15153,N_15003);
nand U15229 (N_15229,N_15104,N_15186);
xor U15230 (N_15230,N_15130,N_15139);
nor U15231 (N_15231,N_15048,N_15099);
nor U15232 (N_15232,N_15196,N_15199);
or U15233 (N_15233,N_15067,N_15185);
nand U15234 (N_15234,N_15016,N_15068);
or U15235 (N_15235,N_15024,N_15076);
or U15236 (N_15236,N_15055,N_15154);
nor U15237 (N_15237,N_15120,N_15124);
xnor U15238 (N_15238,N_15001,N_15187);
xnor U15239 (N_15239,N_15112,N_15045);
nor U15240 (N_15240,N_15056,N_15128);
or U15241 (N_15241,N_15157,N_15117);
xnor U15242 (N_15242,N_15082,N_15115);
or U15243 (N_15243,N_15141,N_15171);
and U15244 (N_15244,N_15000,N_15155);
nor U15245 (N_15245,N_15168,N_15144);
xnor U15246 (N_15246,N_15089,N_15073);
nor U15247 (N_15247,N_15094,N_15091);
nand U15248 (N_15248,N_15037,N_15059);
nor U15249 (N_15249,N_15074,N_15093);
nor U15250 (N_15250,N_15033,N_15062);
and U15251 (N_15251,N_15006,N_15052);
and U15252 (N_15252,N_15023,N_15121);
or U15253 (N_15253,N_15150,N_15080);
nand U15254 (N_15254,N_15057,N_15119);
xnor U15255 (N_15255,N_15181,N_15123);
nor U15256 (N_15256,N_15179,N_15049);
xor U15257 (N_15257,N_15004,N_15042);
nand U15258 (N_15258,N_15175,N_15014);
xor U15259 (N_15259,N_15100,N_15005);
or U15260 (N_15260,N_15063,N_15028);
nor U15261 (N_15261,N_15069,N_15135);
and U15262 (N_15262,N_15065,N_15046);
nor U15263 (N_15263,N_15195,N_15019);
or U15264 (N_15264,N_15137,N_15190);
and U15265 (N_15265,N_15152,N_15131);
nor U15266 (N_15266,N_15075,N_15105);
nand U15267 (N_15267,N_15061,N_15103);
or U15268 (N_15268,N_15025,N_15116);
and U15269 (N_15269,N_15053,N_15050);
xor U15270 (N_15270,N_15177,N_15134);
and U15271 (N_15271,N_15158,N_15129);
or U15272 (N_15272,N_15029,N_15156);
or U15273 (N_15273,N_15017,N_15114);
and U15274 (N_15274,N_15149,N_15126);
xor U15275 (N_15275,N_15189,N_15163);
nor U15276 (N_15276,N_15085,N_15142);
nor U15277 (N_15277,N_15034,N_15133);
or U15278 (N_15278,N_15122,N_15107);
nor U15279 (N_15279,N_15009,N_15044);
nor U15280 (N_15280,N_15022,N_15178);
nor U15281 (N_15281,N_15072,N_15015);
and U15282 (N_15282,N_15027,N_15084);
xnor U15283 (N_15283,N_15011,N_15081);
or U15284 (N_15284,N_15020,N_15188);
xor U15285 (N_15285,N_15007,N_15098);
xor U15286 (N_15286,N_15066,N_15166);
xnor U15287 (N_15287,N_15140,N_15040);
nand U15288 (N_15288,N_15147,N_15106);
and U15289 (N_15289,N_15151,N_15035);
and U15290 (N_15290,N_15172,N_15174);
and U15291 (N_15291,N_15182,N_15194);
nand U15292 (N_15292,N_15193,N_15132);
nand U15293 (N_15293,N_15064,N_15008);
and U15294 (N_15294,N_15180,N_15096);
and U15295 (N_15295,N_15198,N_15083);
and U15296 (N_15296,N_15143,N_15097);
nand U15297 (N_15297,N_15086,N_15192);
or U15298 (N_15298,N_15136,N_15013);
and U15299 (N_15299,N_15021,N_15070);
and U15300 (N_15300,N_15017,N_15025);
xor U15301 (N_15301,N_15009,N_15085);
nor U15302 (N_15302,N_15040,N_15064);
or U15303 (N_15303,N_15034,N_15075);
and U15304 (N_15304,N_15071,N_15021);
nor U15305 (N_15305,N_15015,N_15146);
nand U15306 (N_15306,N_15034,N_15069);
or U15307 (N_15307,N_15184,N_15071);
xnor U15308 (N_15308,N_15165,N_15058);
nand U15309 (N_15309,N_15148,N_15149);
and U15310 (N_15310,N_15094,N_15084);
nor U15311 (N_15311,N_15165,N_15088);
nor U15312 (N_15312,N_15094,N_15191);
and U15313 (N_15313,N_15078,N_15123);
nand U15314 (N_15314,N_15022,N_15090);
or U15315 (N_15315,N_15057,N_15191);
nor U15316 (N_15316,N_15135,N_15037);
and U15317 (N_15317,N_15066,N_15054);
or U15318 (N_15318,N_15050,N_15180);
and U15319 (N_15319,N_15118,N_15112);
nor U15320 (N_15320,N_15189,N_15054);
or U15321 (N_15321,N_15116,N_15135);
xnor U15322 (N_15322,N_15047,N_15092);
nand U15323 (N_15323,N_15143,N_15122);
nor U15324 (N_15324,N_15129,N_15041);
nor U15325 (N_15325,N_15009,N_15002);
and U15326 (N_15326,N_15080,N_15106);
nor U15327 (N_15327,N_15161,N_15145);
xor U15328 (N_15328,N_15091,N_15164);
and U15329 (N_15329,N_15003,N_15016);
nor U15330 (N_15330,N_15146,N_15085);
nand U15331 (N_15331,N_15164,N_15118);
and U15332 (N_15332,N_15120,N_15078);
and U15333 (N_15333,N_15139,N_15125);
nor U15334 (N_15334,N_15154,N_15148);
and U15335 (N_15335,N_15026,N_15176);
nand U15336 (N_15336,N_15183,N_15148);
nand U15337 (N_15337,N_15121,N_15190);
or U15338 (N_15338,N_15038,N_15011);
nor U15339 (N_15339,N_15192,N_15012);
and U15340 (N_15340,N_15180,N_15132);
nor U15341 (N_15341,N_15150,N_15071);
nand U15342 (N_15342,N_15042,N_15184);
xnor U15343 (N_15343,N_15012,N_15011);
or U15344 (N_15344,N_15171,N_15043);
nor U15345 (N_15345,N_15147,N_15175);
nor U15346 (N_15346,N_15007,N_15148);
and U15347 (N_15347,N_15115,N_15147);
xor U15348 (N_15348,N_15091,N_15143);
nand U15349 (N_15349,N_15168,N_15024);
nand U15350 (N_15350,N_15195,N_15103);
or U15351 (N_15351,N_15194,N_15120);
nand U15352 (N_15352,N_15028,N_15035);
xnor U15353 (N_15353,N_15164,N_15185);
or U15354 (N_15354,N_15102,N_15001);
nor U15355 (N_15355,N_15122,N_15014);
xnor U15356 (N_15356,N_15080,N_15021);
and U15357 (N_15357,N_15079,N_15022);
and U15358 (N_15358,N_15174,N_15092);
and U15359 (N_15359,N_15036,N_15157);
and U15360 (N_15360,N_15145,N_15164);
nor U15361 (N_15361,N_15133,N_15054);
and U15362 (N_15362,N_15181,N_15047);
nor U15363 (N_15363,N_15052,N_15058);
or U15364 (N_15364,N_15130,N_15140);
nor U15365 (N_15365,N_15168,N_15012);
and U15366 (N_15366,N_15152,N_15190);
nor U15367 (N_15367,N_15035,N_15186);
xnor U15368 (N_15368,N_15191,N_15119);
nand U15369 (N_15369,N_15092,N_15171);
xnor U15370 (N_15370,N_15032,N_15139);
or U15371 (N_15371,N_15004,N_15191);
nand U15372 (N_15372,N_15163,N_15066);
xor U15373 (N_15373,N_15173,N_15160);
xnor U15374 (N_15374,N_15115,N_15016);
or U15375 (N_15375,N_15066,N_15093);
nor U15376 (N_15376,N_15072,N_15034);
and U15377 (N_15377,N_15000,N_15122);
xor U15378 (N_15378,N_15010,N_15089);
xnor U15379 (N_15379,N_15005,N_15093);
and U15380 (N_15380,N_15184,N_15175);
nand U15381 (N_15381,N_15039,N_15068);
nor U15382 (N_15382,N_15164,N_15070);
or U15383 (N_15383,N_15119,N_15043);
xor U15384 (N_15384,N_15164,N_15028);
nor U15385 (N_15385,N_15081,N_15093);
nor U15386 (N_15386,N_15066,N_15014);
nor U15387 (N_15387,N_15185,N_15131);
xnor U15388 (N_15388,N_15158,N_15088);
or U15389 (N_15389,N_15102,N_15082);
or U15390 (N_15390,N_15118,N_15088);
or U15391 (N_15391,N_15040,N_15051);
xor U15392 (N_15392,N_15015,N_15109);
nand U15393 (N_15393,N_15186,N_15136);
and U15394 (N_15394,N_15036,N_15114);
or U15395 (N_15395,N_15106,N_15176);
nor U15396 (N_15396,N_15097,N_15040);
nor U15397 (N_15397,N_15069,N_15012);
nor U15398 (N_15398,N_15191,N_15111);
xnor U15399 (N_15399,N_15195,N_15080);
xnor U15400 (N_15400,N_15354,N_15225);
and U15401 (N_15401,N_15337,N_15399);
and U15402 (N_15402,N_15222,N_15289);
nor U15403 (N_15403,N_15208,N_15232);
nand U15404 (N_15404,N_15278,N_15256);
and U15405 (N_15405,N_15341,N_15262);
nand U15406 (N_15406,N_15235,N_15257);
or U15407 (N_15407,N_15316,N_15327);
xnor U15408 (N_15408,N_15258,N_15296);
or U15409 (N_15409,N_15213,N_15231);
xor U15410 (N_15410,N_15260,N_15263);
xnor U15411 (N_15411,N_15383,N_15224);
xor U15412 (N_15412,N_15261,N_15339);
nand U15413 (N_15413,N_15398,N_15202);
xor U15414 (N_15414,N_15335,N_15298);
nand U15415 (N_15415,N_15265,N_15227);
xor U15416 (N_15416,N_15370,N_15228);
and U15417 (N_15417,N_15217,N_15294);
xnor U15418 (N_15418,N_15363,N_15272);
nand U15419 (N_15419,N_15285,N_15391);
nor U15420 (N_15420,N_15209,N_15317);
xor U15421 (N_15421,N_15393,N_15374);
or U15422 (N_15422,N_15279,N_15216);
and U15423 (N_15423,N_15361,N_15322);
and U15424 (N_15424,N_15266,N_15223);
nand U15425 (N_15425,N_15308,N_15379);
nand U15426 (N_15426,N_15366,N_15274);
xor U15427 (N_15427,N_15237,N_15333);
nand U15428 (N_15428,N_15245,N_15269);
xnor U15429 (N_15429,N_15203,N_15302);
nor U15430 (N_15430,N_15214,N_15369);
nand U15431 (N_15431,N_15375,N_15338);
nand U15432 (N_15432,N_15349,N_15259);
xor U15433 (N_15433,N_15382,N_15355);
or U15434 (N_15434,N_15277,N_15357);
xor U15435 (N_15435,N_15310,N_15377);
or U15436 (N_15436,N_15204,N_15252);
xor U15437 (N_15437,N_15211,N_15395);
nand U15438 (N_15438,N_15300,N_15323);
nor U15439 (N_15439,N_15314,N_15291);
nand U15440 (N_15440,N_15242,N_15387);
nor U15441 (N_15441,N_15320,N_15385);
xnor U15442 (N_15442,N_15336,N_15297);
or U15443 (N_15443,N_15388,N_15276);
nand U15444 (N_15444,N_15348,N_15358);
and U15445 (N_15445,N_15234,N_15301);
xor U15446 (N_15446,N_15283,N_15284);
nor U15447 (N_15447,N_15206,N_15249);
nor U15448 (N_15448,N_15319,N_15286);
and U15449 (N_15449,N_15306,N_15332);
nor U15450 (N_15450,N_15389,N_15334);
nand U15451 (N_15451,N_15288,N_15230);
nor U15452 (N_15452,N_15293,N_15326);
or U15453 (N_15453,N_15392,N_15324);
nand U15454 (N_15454,N_15303,N_15384);
nor U15455 (N_15455,N_15321,N_15253);
nand U15456 (N_15456,N_15376,N_15312);
or U15457 (N_15457,N_15215,N_15292);
nor U15458 (N_15458,N_15220,N_15290);
and U15459 (N_15459,N_15246,N_15251);
xor U15460 (N_15460,N_15305,N_15318);
xnor U15461 (N_15461,N_15347,N_15218);
and U15462 (N_15462,N_15299,N_15344);
xor U15463 (N_15463,N_15394,N_15250);
nor U15464 (N_15464,N_15313,N_15205);
nand U15465 (N_15465,N_15309,N_15201);
xor U15466 (N_15466,N_15340,N_15255);
and U15467 (N_15467,N_15397,N_15352);
nand U15468 (N_15468,N_15244,N_15273);
and U15469 (N_15469,N_15381,N_15325);
nand U15470 (N_15470,N_15373,N_15210);
nand U15471 (N_15471,N_15241,N_15287);
or U15472 (N_15472,N_15345,N_15219);
nor U15473 (N_15473,N_15390,N_15343);
or U15474 (N_15474,N_15270,N_15346);
xor U15475 (N_15475,N_15267,N_15329);
nand U15476 (N_15476,N_15243,N_15380);
and U15477 (N_15477,N_15365,N_15330);
nor U15478 (N_15478,N_15378,N_15364);
or U15479 (N_15479,N_15328,N_15304);
and U15480 (N_15480,N_15353,N_15271);
xnor U15481 (N_15481,N_15221,N_15372);
or U15482 (N_15482,N_15315,N_15386);
and U15483 (N_15483,N_15275,N_15371);
nor U15484 (N_15484,N_15238,N_15362);
xor U15485 (N_15485,N_15236,N_15233);
nor U15486 (N_15486,N_15248,N_15226);
and U15487 (N_15487,N_15281,N_15264);
or U15488 (N_15488,N_15356,N_15342);
nor U15489 (N_15489,N_15254,N_15396);
or U15490 (N_15490,N_15331,N_15311);
nand U15491 (N_15491,N_15307,N_15351);
xor U15492 (N_15492,N_15359,N_15212);
or U15493 (N_15493,N_15207,N_15240);
or U15494 (N_15494,N_15295,N_15268);
and U15495 (N_15495,N_15282,N_15280);
and U15496 (N_15496,N_15239,N_15360);
nor U15497 (N_15497,N_15350,N_15200);
nor U15498 (N_15498,N_15367,N_15229);
nand U15499 (N_15499,N_15247,N_15368);
and U15500 (N_15500,N_15370,N_15202);
nor U15501 (N_15501,N_15204,N_15370);
nand U15502 (N_15502,N_15399,N_15382);
xor U15503 (N_15503,N_15204,N_15324);
and U15504 (N_15504,N_15276,N_15222);
nor U15505 (N_15505,N_15274,N_15288);
nor U15506 (N_15506,N_15204,N_15337);
xor U15507 (N_15507,N_15314,N_15257);
nor U15508 (N_15508,N_15386,N_15263);
nand U15509 (N_15509,N_15317,N_15206);
and U15510 (N_15510,N_15207,N_15349);
xnor U15511 (N_15511,N_15206,N_15214);
nor U15512 (N_15512,N_15296,N_15359);
and U15513 (N_15513,N_15281,N_15311);
or U15514 (N_15514,N_15310,N_15246);
nand U15515 (N_15515,N_15238,N_15386);
nand U15516 (N_15516,N_15237,N_15266);
and U15517 (N_15517,N_15303,N_15309);
nor U15518 (N_15518,N_15389,N_15252);
nor U15519 (N_15519,N_15340,N_15264);
and U15520 (N_15520,N_15227,N_15361);
xnor U15521 (N_15521,N_15340,N_15280);
xor U15522 (N_15522,N_15218,N_15223);
and U15523 (N_15523,N_15292,N_15311);
or U15524 (N_15524,N_15302,N_15343);
xor U15525 (N_15525,N_15258,N_15222);
and U15526 (N_15526,N_15250,N_15285);
or U15527 (N_15527,N_15369,N_15333);
nand U15528 (N_15528,N_15245,N_15285);
nand U15529 (N_15529,N_15387,N_15340);
or U15530 (N_15530,N_15209,N_15303);
or U15531 (N_15531,N_15363,N_15281);
and U15532 (N_15532,N_15386,N_15352);
nor U15533 (N_15533,N_15222,N_15205);
xnor U15534 (N_15534,N_15313,N_15357);
and U15535 (N_15535,N_15325,N_15300);
nor U15536 (N_15536,N_15286,N_15380);
xnor U15537 (N_15537,N_15397,N_15291);
nand U15538 (N_15538,N_15353,N_15355);
xor U15539 (N_15539,N_15355,N_15251);
nor U15540 (N_15540,N_15312,N_15207);
nor U15541 (N_15541,N_15303,N_15332);
and U15542 (N_15542,N_15345,N_15348);
nand U15543 (N_15543,N_15236,N_15287);
nand U15544 (N_15544,N_15319,N_15391);
nand U15545 (N_15545,N_15364,N_15200);
xor U15546 (N_15546,N_15302,N_15283);
nor U15547 (N_15547,N_15271,N_15204);
nor U15548 (N_15548,N_15209,N_15356);
or U15549 (N_15549,N_15254,N_15369);
or U15550 (N_15550,N_15208,N_15345);
and U15551 (N_15551,N_15304,N_15336);
or U15552 (N_15552,N_15368,N_15358);
nand U15553 (N_15553,N_15235,N_15251);
nor U15554 (N_15554,N_15324,N_15285);
and U15555 (N_15555,N_15308,N_15287);
or U15556 (N_15556,N_15358,N_15385);
nand U15557 (N_15557,N_15225,N_15217);
xnor U15558 (N_15558,N_15344,N_15238);
nand U15559 (N_15559,N_15213,N_15276);
and U15560 (N_15560,N_15337,N_15294);
nand U15561 (N_15561,N_15225,N_15289);
xor U15562 (N_15562,N_15294,N_15239);
nand U15563 (N_15563,N_15361,N_15228);
or U15564 (N_15564,N_15303,N_15268);
nor U15565 (N_15565,N_15242,N_15375);
xor U15566 (N_15566,N_15241,N_15347);
nor U15567 (N_15567,N_15366,N_15352);
and U15568 (N_15568,N_15210,N_15317);
xnor U15569 (N_15569,N_15225,N_15348);
nor U15570 (N_15570,N_15264,N_15252);
nand U15571 (N_15571,N_15267,N_15331);
and U15572 (N_15572,N_15387,N_15399);
or U15573 (N_15573,N_15304,N_15235);
and U15574 (N_15574,N_15220,N_15238);
xnor U15575 (N_15575,N_15304,N_15396);
and U15576 (N_15576,N_15322,N_15206);
or U15577 (N_15577,N_15269,N_15243);
and U15578 (N_15578,N_15204,N_15202);
xnor U15579 (N_15579,N_15339,N_15375);
xnor U15580 (N_15580,N_15210,N_15338);
or U15581 (N_15581,N_15369,N_15314);
nand U15582 (N_15582,N_15396,N_15397);
or U15583 (N_15583,N_15355,N_15210);
xnor U15584 (N_15584,N_15335,N_15270);
nand U15585 (N_15585,N_15372,N_15299);
nor U15586 (N_15586,N_15268,N_15310);
nand U15587 (N_15587,N_15341,N_15399);
or U15588 (N_15588,N_15262,N_15231);
nor U15589 (N_15589,N_15268,N_15236);
nor U15590 (N_15590,N_15279,N_15303);
and U15591 (N_15591,N_15216,N_15298);
nand U15592 (N_15592,N_15276,N_15381);
nand U15593 (N_15593,N_15350,N_15207);
and U15594 (N_15594,N_15340,N_15215);
and U15595 (N_15595,N_15277,N_15222);
or U15596 (N_15596,N_15365,N_15235);
and U15597 (N_15597,N_15286,N_15293);
xor U15598 (N_15598,N_15306,N_15240);
xnor U15599 (N_15599,N_15344,N_15359);
xnor U15600 (N_15600,N_15462,N_15582);
nand U15601 (N_15601,N_15443,N_15400);
nor U15602 (N_15602,N_15589,N_15501);
or U15603 (N_15603,N_15482,N_15597);
or U15604 (N_15604,N_15453,N_15430);
xnor U15605 (N_15605,N_15468,N_15480);
or U15606 (N_15606,N_15523,N_15455);
or U15607 (N_15607,N_15515,N_15489);
and U15608 (N_15608,N_15529,N_15472);
nor U15609 (N_15609,N_15580,N_15421);
and U15610 (N_15610,N_15479,N_15512);
xor U15611 (N_15611,N_15484,N_15578);
xor U15612 (N_15612,N_15475,N_15596);
nand U15613 (N_15613,N_15517,N_15571);
xor U15614 (N_15614,N_15513,N_15545);
xnor U15615 (N_15615,N_15599,N_15527);
or U15616 (N_15616,N_15460,N_15549);
nor U15617 (N_15617,N_15587,N_15476);
xnor U15618 (N_15618,N_15494,N_15465);
nor U15619 (N_15619,N_15520,N_15579);
and U15620 (N_15620,N_15541,N_15450);
or U15621 (N_15621,N_15410,N_15429);
xnor U15622 (N_15622,N_15406,N_15525);
xnor U15623 (N_15623,N_15426,N_15486);
or U15624 (N_15624,N_15487,N_15546);
and U15625 (N_15625,N_15411,N_15509);
or U15626 (N_15626,N_15598,N_15540);
nor U15627 (N_15627,N_15403,N_15417);
xor U15628 (N_15628,N_15467,N_15446);
nand U15629 (N_15629,N_15466,N_15436);
nand U15630 (N_15630,N_15555,N_15594);
xor U15631 (N_15631,N_15550,N_15535);
nand U15632 (N_15632,N_15528,N_15469);
and U15633 (N_15633,N_15577,N_15510);
and U15634 (N_15634,N_15408,N_15564);
xnor U15635 (N_15635,N_15519,N_15507);
nor U15636 (N_15636,N_15551,N_15473);
xor U15637 (N_15637,N_15434,N_15454);
and U15638 (N_15638,N_15524,N_15413);
nand U15639 (N_15639,N_15435,N_15561);
and U15640 (N_15640,N_15463,N_15585);
or U15641 (N_15641,N_15447,N_15566);
or U15642 (N_15642,N_15415,N_15448);
or U15643 (N_15643,N_15478,N_15569);
nand U15644 (N_15644,N_15452,N_15474);
nand U15645 (N_15645,N_15425,N_15495);
and U15646 (N_15646,N_15537,N_15511);
and U15647 (N_15647,N_15573,N_15534);
nor U15648 (N_15648,N_15418,N_15522);
and U15649 (N_15649,N_15536,N_15428);
nor U15650 (N_15650,N_15481,N_15538);
nand U15651 (N_15651,N_15456,N_15457);
and U15652 (N_15652,N_15544,N_15412);
and U15653 (N_15653,N_15542,N_15552);
or U15654 (N_15654,N_15490,N_15458);
xnor U15655 (N_15655,N_15539,N_15592);
and U15656 (N_15656,N_15563,N_15565);
and U15657 (N_15657,N_15548,N_15464);
and U15658 (N_15658,N_15444,N_15562);
or U15659 (N_15659,N_15574,N_15407);
nor U15660 (N_15660,N_15414,N_15438);
nand U15661 (N_15661,N_15405,N_15493);
or U15662 (N_15662,N_15581,N_15575);
xor U15663 (N_15663,N_15595,N_15572);
xor U15664 (N_15664,N_15437,N_15431);
or U15665 (N_15665,N_15439,N_15409);
xor U15666 (N_15666,N_15583,N_15518);
and U15667 (N_15667,N_15459,N_15505);
nand U15668 (N_15668,N_15432,N_15588);
nand U15669 (N_15669,N_15554,N_15516);
xor U15670 (N_15670,N_15442,N_15401);
xnor U15671 (N_15671,N_15433,N_15461);
nand U15672 (N_15672,N_15553,N_15568);
nor U15673 (N_15673,N_15591,N_15557);
or U15674 (N_15674,N_15500,N_15559);
xor U15675 (N_15675,N_15499,N_15449);
or U15676 (N_15676,N_15593,N_15530);
nand U15677 (N_15677,N_15451,N_15532);
nand U15678 (N_15678,N_15504,N_15502);
or U15679 (N_15679,N_15427,N_15531);
or U15680 (N_15680,N_15497,N_15424);
nand U15681 (N_15681,N_15488,N_15496);
nand U15682 (N_15682,N_15570,N_15567);
and U15683 (N_15683,N_15560,N_15483);
and U15684 (N_15684,N_15508,N_15521);
and U15685 (N_15685,N_15471,N_15492);
nand U15686 (N_15686,N_15477,N_15543);
and U15687 (N_15687,N_15506,N_15558);
xor U15688 (N_15688,N_15590,N_15423);
and U15689 (N_15689,N_15440,N_15420);
xnor U15690 (N_15690,N_15441,N_15503);
xnor U15691 (N_15691,N_15514,N_15586);
nand U15692 (N_15692,N_15584,N_15576);
nor U15693 (N_15693,N_15556,N_15416);
nor U15694 (N_15694,N_15402,N_15470);
and U15695 (N_15695,N_15404,N_15498);
nand U15696 (N_15696,N_15422,N_15491);
and U15697 (N_15697,N_15526,N_15533);
or U15698 (N_15698,N_15445,N_15419);
and U15699 (N_15699,N_15485,N_15547);
and U15700 (N_15700,N_15484,N_15592);
xor U15701 (N_15701,N_15473,N_15472);
xnor U15702 (N_15702,N_15483,N_15544);
xor U15703 (N_15703,N_15419,N_15519);
nand U15704 (N_15704,N_15589,N_15569);
and U15705 (N_15705,N_15472,N_15498);
xnor U15706 (N_15706,N_15482,N_15506);
nor U15707 (N_15707,N_15519,N_15575);
or U15708 (N_15708,N_15561,N_15529);
or U15709 (N_15709,N_15447,N_15431);
nand U15710 (N_15710,N_15444,N_15440);
nand U15711 (N_15711,N_15513,N_15514);
nand U15712 (N_15712,N_15457,N_15592);
or U15713 (N_15713,N_15412,N_15530);
nand U15714 (N_15714,N_15508,N_15538);
nand U15715 (N_15715,N_15472,N_15563);
xnor U15716 (N_15716,N_15438,N_15539);
nor U15717 (N_15717,N_15518,N_15416);
nor U15718 (N_15718,N_15571,N_15581);
and U15719 (N_15719,N_15565,N_15437);
and U15720 (N_15720,N_15402,N_15584);
xor U15721 (N_15721,N_15581,N_15543);
or U15722 (N_15722,N_15414,N_15544);
xnor U15723 (N_15723,N_15449,N_15555);
xor U15724 (N_15724,N_15439,N_15472);
nand U15725 (N_15725,N_15583,N_15425);
and U15726 (N_15726,N_15432,N_15464);
xor U15727 (N_15727,N_15439,N_15457);
and U15728 (N_15728,N_15580,N_15422);
and U15729 (N_15729,N_15519,N_15523);
nor U15730 (N_15730,N_15423,N_15598);
and U15731 (N_15731,N_15511,N_15516);
or U15732 (N_15732,N_15555,N_15551);
nand U15733 (N_15733,N_15510,N_15479);
or U15734 (N_15734,N_15509,N_15516);
xor U15735 (N_15735,N_15567,N_15410);
and U15736 (N_15736,N_15409,N_15462);
or U15737 (N_15737,N_15479,N_15453);
nand U15738 (N_15738,N_15515,N_15551);
and U15739 (N_15739,N_15495,N_15455);
nand U15740 (N_15740,N_15427,N_15559);
or U15741 (N_15741,N_15427,N_15463);
nand U15742 (N_15742,N_15598,N_15445);
and U15743 (N_15743,N_15405,N_15518);
xnor U15744 (N_15744,N_15469,N_15499);
or U15745 (N_15745,N_15509,N_15487);
nor U15746 (N_15746,N_15571,N_15407);
nor U15747 (N_15747,N_15416,N_15496);
and U15748 (N_15748,N_15548,N_15570);
or U15749 (N_15749,N_15490,N_15489);
or U15750 (N_15750,N_15533,N_15402);
nor U15751 (N_15751,N_15480,N_15594);
nor U15752 (N_15752,N_15551,N_15569);
xor U15753 (N_15753,N_15407,N_15418);
nand U15754 (N_15754,N_15435,N_15461);
nand U15755 (N_15755,N_15510,N_15465);
nand U15756 (N_15756,N_15586,N_15486);
or U15757 (N_15757,N_15488,N_15458);
xor U15758 (N_15758,N_15463,N_15566);
nor U15759 (N_15759,N_15427,N_15504);
nand U15760 (N_15760,N_15400,N_15425);
xnor U15761 (N_15761,N_15553,N_15569);
nor U15762 (N_15762,N_15528,N_15446);
and U15763 (N_15763,N_15533,N_15479);
or U15764 (N_15764,N_15473,N_15433);
xor U15765 (N_15765,N_15530,N_15550);
nor U15766 (N_15766,N_15532,N_15475);
and U15767 (N_15767,N_15547,N_15509);
nand U15768 (N_15768,N_15456,N_15453);
nor U15769 (N_15769,N_15474,N_15538);
nand U15770 (N_15770,N_15482,N_15417);
xor U15771 (N_15771,N_15486,N_15461);
or U15772 (N_15772,N_15557,N_15478);
xnor U15773 (N_15773,N_15501,N_15449);
nor U15774 (N_15774,N_15522,N_15464);
or U15775 (N_15775,N_15402,N_15580);
xnor U15776 (N_15776,N_15566,N_15545);
nand U15777 (N_15777,N_15588,N_15498);
and U15778 (N_15778,N_15406,N_15561);
xor U15779 (N_15779,N_15591,N_15446);
and U15780 (N_15780,N_15541,N_15486);
xnor U15781 (N_15781,N_15474,N_15414);
nor U15782 (N_15782,N_15406,N_15495);
nor U15783 (N_15783,N_15590,N_15531);
or U15784 (N_15784,N_15573,N_15497);
nand U15785 (N_15785,N_15593,N_15451);
and U15786 (N_15786,N_15474,N_15472);
or U15787 (N_15787,N_15506,N_15574);
and U15788 (N_15788,N_15470,N_15403);
nand U15789 (N_15789,N_15534,N_15535);
xor U15790 (N_15790,N_15474,N_15557);
and U15791 (N_15791,N_15457,N_15519);
or U15792 (N_15792,N_15474,N_15486);
nor U15793 (N_15793,N_15594,N_15409);
nor U15794 (N_15794,N_15570,N_15526);
nand U15795 (N_15795,N_15522,N_15566);
or U15796 (N_15796,N_15473,N_15529);
xnor U15797 (N_15797,N_15432,N_15541);
nor U15798 (N_15798,N_15486,N_15524);
nor U15799 (N_15799,N_15531,N_15575);
nand U15800 (N_15800,N_15786,N_15713);
xor U15801 (N_15801,N_15688,N_15664);
nor U15802 (N_15802,N_15769,N_15729);
nand U15803 (N_15803,N_15620,N_15706);
nand U15804 (N_15804,N_15700,N_15617);
nand U15805 (N_15805,N_15641,N_15690);
and U15806 (N_15806,N_15672,N_15738);
nand U15807 (N_15807,N_15724,N_15683);
or U15808 (N_15808,N_15737,N_15774);
nor U15809 (N_15809,N_15630,N_15798);
and U15810 (N_15810,N_15741,N_15651);
xor U15811 (N_15811,N_15719,N_15623);
and U15812 (N_15812,N_15662,N_15707);
nand U15813 (N_15813,N_15681,N_15760);
nand U15814 (N_15814,N_15742,N_15708);
xnor U15815 (N_15815,N_15710,N_15601);
nand U15816 (N_15816,N_15747,N_15763);
nand U15817 (N_15817,N_15771,N_15604);
or U15818 (N_15818,N_15775,N_15733);
xnor U15819 (N_15819,N_15615,N_15725);
and U15820 (N_15820,N_15756,N_15715);
nor U15821 (N_15821,N_15634,N_15671);
or U15822 (N_15822,N_15793,N_15768);
or U15823 (N_15823,N_15697,N_15799);
xor U15824 (N_15824,N_15693,N_15609);
or U15825 (N_15825,N_15782,N_15665);
or U15826 (N_15826,N_15629,N_15640);
and U15827 (N_15827,N_15692,N_15663);
or U15828 (N_15828,N_15780,N_15703);
nor U15829 (N_15829,N_15701,N_15602);
nand U15830 (N_15830,N_15722,N_15759);
and U15831 (N_15831,N_15734,N_15625);
xor U15832 (N_15832,N_15748,N_15772);
xnor U15833 (N_15833,N_15614,N_15773);
or U15834 (N_15834,N_15643,N_15740);
nor U15835 (N_15835,N_15777,N_15755);
nor U15836 (N_15836,N_15789,N_15680);
nand U15837 (N_15837,N_15730,N_15785);
nor U15838 (N_15838,N_15660,N_15612);
or U15839 (N_15839,N_15749,N_15721);
nand U15840 (N_15840,N_15649,N_15744);
or U15841 (N_15841,N_15605,N_15762);
and U15842 (N_15842,N_15687,N_15675);
and U15843 (N_15843,N_15669,N_15647);
and U15844 (N_15844,N_15752,N_15642);
nor U15845 (N_15845,N_15637,N_15699);
xnor U15846 (N_15846,N_15757,N_15611);
nor U15847 (N_15847,N_15732,N_15776);
and U15848 (N_15848,N_15691,N_15606);
nor U15849 (N_15849,N_15767,N_15761);
xnor U15850 (N_15850,N_15731,N_15686);
xnor U15851 (N_15851,N_15636,N_15736);
nand U15852 (N_15852,N_15695,N_15779);
and U15853 (N_15853,N_15626,N_15783);
or U15854 (N_15854,N_15627,N_15682);
or U15855 (N_15855,N_15603,N_15610);
nand U15856 (N_15856,N_15766,N_15650);
and U15857 (N_15857,N_15600,N_15754);
nand U15858 (N_15858,N_15678,N_15778);
nor U15859 (N_15859,N_15619,N_15745);
nor U15860 (N_15860,N_15702,N_15633);
nand U15861 (N_15861,N_15726,N_15618);
nor U15862 (N_15862,N_15613,N_15656);
xor U15863 (N_15863,N_15670,N_15628);
and U15864 (N_15864,N_15677,N_15751);
xnor U15865 (N_15865,N_15790,N_15717);
or U15866 (N_15866,N_15781,N_15621);
nor U15867 (N_15867,N_15797,N_15709);
nor U15868 (N_15868,N_15654,N_15652);
and U15869 (N_15869,N_15739,N_15784);
nor U15870 (N_15870,N_15674,N_15788);
nand U15871 (N_15871,N_15705,N_15795);
and U15872 (N_15872,N_15765,N_15658);
nor U15873 (N_15873,N_15787,N_15750);
nand U15874 (N_15874,N_15796,N_15791);
and U15875 (N_15875,N_15711,N_15685);
nor U15876 (N_15876,N_15792,N_15668);
xor U15877 (N_15877,N_15694,N_15657);
nor U15878 (N_15878,N_15631,N_15632);
and U15879 (N_15879,N_15716,N_15667);
xor U15880 (N_15880,N_15644,N_15653);
or U15881 (N_15881,N_15794,N_15723);
xnor U15882 (N_15882,N_15666,N_15638);
nand U15883 (N_15883,N_15684,N_15735);
xnor U15884 (N_15884,N_15712,N_15608);
or U15885 (N_15885,N_15696,N_15743);
nor U15886 (N_15886,N_15655,N_15676);
and U15887 (N_15887,N_15645,N_15758);
or U15888 (N_15888,N_15728,N_15679);
and U15889 (N_15889,N_15720,N_15659);
xnor U15890 (N_15890,N_15714,N_15727);
and U15891 (N_15891,N_15753,N_15624);
or U15892 (N_15892,N_15689,N_15718);
xnor U15893 (N_15893,N_15635,N_15607);
xnor U15894 (N_15894,N_15746,N_15646);
nand U15895 (N_15895,N_15698,N_15639);
nor U15896 (N_15896,N_15648,N_15622);
xor U15897 (N_15897,N_15704,N_15673);
nand U15898 (N_15898,N_15770,N_15616);
xnor U15899 (N_15899,N_15661,N_15764);
nand U15900 (N_15900,N_15662,N_15618);
nor U15901 (N_15901,N_15691,N_15718);
and U15902 (N_15902,N_15616,N_15720);
xor U15903 (N_15903,N_15751,N_15794);
nor U15904 (N_15904,N_15658,N_15688);
nor U15905 (N_15905,N_15786,N_15728);
or U15906 (N_15906,N_15733,N_15781);
nor U15907 (N_15907,N_15646,N_15609);
or U15908 (N_15908,N_15708,N_15752);
nor U15909 (N_15909,N_15766,N_15623);
xor U15910 (N_15910,N_15658,N_15748);
nand U15911 (N_15911,N_15782,N_15652);
xor U15912 (N_15912,N_15691,N_15654);
xor U15913 (N_15913,N_15786,N_15636);
or U15914 (N_15914,N_15648,N_15783);
xnor U15915 (N_15915,N_15685,N_15726);
nor U15916 (N_15916,N_15637,N_15647);
nand U15917 (N_15917,N_15707,N_15653);
or U15918 (N_15918,N_15790,N_15766);
nand U15919 (N_15919,N_15773,N_15707);
or U15920 (N_15920,N_15697,N_15672);
nor U15921 (N_15921,N_15719,N_15665);
or U15922 (N_15922,N_15690,N_15720);
xnor U15923 (N_15923,N_15796,N_15685);
xor U15924 (N_15924,N_15639,N_15718);
xor U15925 (N_15925,N_15722,N_15745);
or U15926 (N_15926,N_15750,N_15673);
nand U15927 (N_15927,N_15774,N_15618);
nor U15928 (N_15928,N_15685,N_15640);
and U15929 (N_15929,N_15652,N_15732);
or U15930 (N_15930,N_15646,N_15674);
nand U15931 (N_15931,N_15744,N_15703);
and U15932 (N_15932,N_15622,N_15775);
and U15933 (N_15933,N_15609,N_15662);
xnor U15934 (N_15934,N_15648,N_15640);
nand U15935 (N_15935,N_15746,N_15606);
nand U15936 (N_15936,N_15604,N_15687);
nor U15937 (N_15937,N_15637,N_15733);
nor U15938 (N_15938,N_15692,N_15721);
and U15939 (N_15939,N_15729,N_15791);
or U15940 (N_15940,N_15767,N_15756);
and U15941 (N_15941,N_15616,N_15656);
nand U15942 (N_15942,N_15613,N_15787);
nor U15943 (N_15943,N_15735,N_15615);
or U15944 (N_15944,N_15720,N_15639);
and U15945 (N_15945,N_15717,N_15668);
nor U15946 (N_15946,N_15654,N_15719);
and U15947 (N_15947,N_15667,N_15751);
nor U15948 (N_15948,N_15635,N_15785);
and U15949 (N_15949,N_15611,N_15633);
xnor U15950 (N_15950,N_15637,N_15710);
nor U15951 (N_15951,N_15744,N_15605);
and U15952 (N_15952,N_15606,N_15653);
xor U15953 (N_15953,N_15671,N_15687);
nor U15954 (N_15954,N_15763,N_15706);
nand U15955 (N_15955,N_15651,N_15785);
or U15956 (N_15956,N_15656,N_15762);
or U15957 (N_15957,N_15789,N_15670);
nand U15958 (N_15958,N_15714,N_15622);
and U15959 (N_15959,N_15763,N_15741);
nor U15960 (N_15960,N_15668,N_15736);
and U15961 (N_15961,N_15734,N_15786);
nand U15962 (N_15962,N_15658,N_15758);
nor U15963 (N_15963,N_15769,N_15695);
xnor U15964 (N_15964,N_15771,N_15663);
and U15965 (N_15965,N_15608,N_15687);
and U15966 (N_15966,N_15612,N_15730);
and U15967 (N_15967,N_15719,N_15661);
or U15968 (N_15968,N_15775,N_15754);
nand U15969 (N_15969,N_15755,N_15729);
and U15970 (N_15970,N_15645,N_15672);
xnor U15971 (N_15971,N_15684,N_15755);
or U15972 (N_15972,N_15681,N_15618);
nor U15973 (N_15973,N_15779,N_15780);
xnor U15974 (N_15974,N_15623,N_15629);
or U15975 (N_15975,N_15609,N_15622);
and U15976 (N_15976,N_15745,N_15747);
xnor U15977 (N_15977,N_15776,N_15600);
or U15978 (N_15978,N_15697,N_15631);
and U15979 (N_15979,N_15617,N_15670);
nor U15980 (N_15980,N_15781,N_15640);
or U15981 (N_15981,N_15656,N_15610);
nand U15982 (N_15982,N_15666,N_15795);
and U15983 (N_15983,N_15749,N_15713);
xor U15984 (N_15984,N_15729,N_15711);
or U15985 (N_15985,N_15627,N_15636);
nor U15986 (N_15986,N_15661,N_15716);
xnor U15987 (N_15987,N_15746,N_15737);
xor U15988 (N_15988,N_15639,N_15702);
nor U15989 (N_15989,N_15707,N_15605);
xor U15990 (N_15990,N_15664,N_15624);
nand U15991 (N_15991,N_15739,N_15758);
nor U15992 (N_15992,N_15630,N_15746);
and U15993 (N_15993,N_15655,N_15650);
or U15994 (N_15994,N_15671,N_15716);
xnor U15995 (N_15995,N_15694,N_15606);
nor U15996 (N_15996,N_15624,N_15638);
nand U15997 (N_15997,N_15607,N_15700);
or U15998 (N_15998,N_15789,N_15630);
or U15999 (N_15999,N_15658,N_15620);
or U16000 (N_16000,N_15985,N_15926);
or U16001 (N_16001,N_15945,N_15847);
or U16002 (N_16002,N_15989,N_15922);
or U16003 (N_16003,N_15936,N_15881);
nor U16004 (N_16004,N_15800,N_15884);
nand U16005 (N_16005,N_15959,N_15972);
and U16006 (N_16006,N_15934,N_15999);
and U16007 (N_16007,N_15839,N_15904);
nor U16008 (N_16008,N_15919,N_15942);
or U16009 (N_16009,N_15844,N_15961);
and U16010 (N_16010,N_15949,N_15906);
or U16011 (N_16011,N_15981,N_15903);
nand U16012 (N_16012,N_15875,N_15946);
or U16013 (N_16013,N_15995,N_15829);
and U16014 (N_16014,N_15824,N_15914);
xnor U16015 (N_16015,N_15909,N_15809);
and U16016 (N_16016,N_15862,N_15965);
and U16017 (N_16017,N_15849,N_15840);
xor U16018 (N_16018,N_15939,N_15810);
xnor U16019 (N_16019,N_15852,N_15905);
nand U16020 (N_16020,N_15864,N_15951);
or U16021 (N_16021,N_15878,N_15900);
xnor U16022 (N_16022,N_15950,N_15843);
or U16023 (N_16023,N_15870,N_15837);
nand U16024 (N_16024,N_15929,N_15987);
and U16025 (N_16025,N_15963,N_15943);
nand U16026 (N_16026,N_15804,N_15937);
and U16027 (N_16027,N_15892,N_15865);
xor U16028 (N_16028,N_15826,N_15967);
and U16029 (N_16029,N_15899,N_15979);
nand U16030 (N_16030,N_15997,N_15984);
and U16031 (N_16031,N_15815,N_15910);
or U16032 (N_16032,N_15994,N_15883);
and U16033 (N_16033,N_15938,N_15832);
or U16034 (N_16034,N_15841,N_15858);
and U16035 (N_16035,N_15908,N_15986);
xnor U16036 (N_16036,N_15948,N_15834);
nand U16037 (N_16037,N_15998,N_15953);
nor U16038 (N_16038,N_15818,N_15867);
nor U16039 (N_16039,N_15857,N_15872);
or U16040 (N_16040,N_15918,N_15932);
or U16041 (N_16041,N_15813,N_15923);
or U16042 (N_16042,N_15893,N_15833);
xnor U16043 (N_16043,N_15928,N_15853);
and U16044 (N_16044,N_15868,N_15952);
xnor U16045 (N_16045,N_15819,N_15808);
nand U16046 (N_16046,N_15876,N_15966);
nand U16047 (N_16047,N_15947,N_15980);
nand U16048 (N_16048,N_15902,N_15917);
nor U16049 (N_16049,N_15887,N_15898);
xor U16050 (N_16050,N_15859,N_15933);
nand U16051 (N_16051,N_15891,N_15978);
nand U16052 (N_16052,N_15988,N_15856);
and U16053 (N_16053,N_15816,N_15885);
nand U16054 (N_16054,N_15968,N_15940);
nor U16055 (N_16055,N_15993,N_15901);
and U16056 (N_16056,N_15845,N_15823);
nand U16057 (N_16057,N_15861,N_15931);
nand U16058 (N_16058,N_15869,N_15846);
or U16059 (N_16059,N_15806,N_15830);
or U16060 (N_16060,N_15977,N_15921);
and U16061 (N_16061,N_15895,N_15956);
xor U16062 (N_16062,N_15836,N_15992);
xnor U16063 (N_16063,N_15880,N_15822);
xor U16064 (N_16064,N_15803,N_15969);
nand U16065 (N_16065,N_15842,N_15851);
and U16066 (N_16066,N_15976,N_15915);
and U16067 (N_16067,N_15801,N_15882);
and U16068 (N_16068,N_15955,N_15896);
xnor U16069 (N_16069,N_15888,N_15925);
and U16070 (N_16070,N_15802,N_15831);
nor U16071 (N_16071,N_15874,N_15886);
xnor U16072 (N_16072,N_15920,N_15873);
xor U16073 (N_16073,N_15897,N_15848);
and U16074 (N_16074,N_15958,N_15941);
nand U16075 (N_16075,N_15807,N_15973);
or U16076 (N_16076,N_15983,N_15954);
nor U16077 (N_16077,N_15821,N_15911);
and U16078 (N_16078,N_15991,N_15962);
xnor U16079 (N_16079,N_15974,N_15990);
and U16080 (N_16080,N_15970,N_15889);
xnor U16081 (N_16081,N_15811,N_15912);
nor U16082 (N_16082,N_15855,N_15850);
nand U16083 (N_16083,N_15924,N_15996);
and U16084 (N_16084,N_15854,N_15825);
nor U16085 (N_16085,N_15838,N_15964);
nand U16086 (N_16086,N_15812,N_15894);
or U16087 (N_16087,N_15820,N_15863);
or U16088 (N_16088,N_15805,N_15957);
and U16089 (N_16089,N_15835,N_15890);
or U16090 (N_16090,N_15982,N_15871);
xnor U16091 (N_16091,N_15960,N_15944);
or U16092 (N_16092,N_15930,N_15907);
and U16093 (N_16093,N_15814,N_15975);
nand U16094 (N_16094,N_15927,N_15866);
or U16095 (N_16095,N_15971,N_15913);
and U16096 (N_16096,N_15935,N_15817);
and U16097 (N_16097,N_15916,N_15879);
and U16098 (N_16098,N_15860,N_15827);
nand U16099 (N_16099,N_15828,N_15877);
nand U16100 (N_16100,N_15867,N_15893);
and U16101 (N_16101,N_15933,N_15987);
xnor U16102 (N_16102,N_15924,N_15849);
nand U16103 (N_16103,N_15986,N_15844);
nor U16104 (N_16104,N_15816,N_15979);
nand U16105 (N_16105,N_15804,N_15892);
and U16106 (N_16106,N_15926,N_15931);
or U16107 (N_16107,N_15815,N_15872);
xnor U16108 (N_16108,N_15900,N_15835);
or U16109 (N_16109,N_15850,N_15974);
or U16110 (N_16110,N_15889,N_15842);
nand U16111 (N_16111,N_15863,N_15823);
nor U16112 (N_16112,N_15926,N_15998);
and U16113 (N_16113,N_15816,N_15986);
or U16114 (N_16114,N_15986,N_15992);
or U16115 (N_16115,N_15861,N_15909);
and U16116 (N_16116,N_15813,N_15845);
nand U16117 (N_16117,N_15943,N_15900);
nand U16118 (N_16118,N_15833,N_15801);
and U16119 (N_16119,N_15873,N_15899);
or U16120 (N_16120,N_15925,N_15993);
xor U16121 (N_16121,N_15944,N_15800);
xnor U16122 (N_16122,N_15820,N_15851);
nor U16123 (N_16123,N_15953,N_15855);
xnor U16124 (N_16124,N_15881,N_15857);
nor U16125 (N_16125,N_15976,N_15840);
or U16126 (N_16126,N_15851,N_15945);
or U16127 (N_16127,N_15808,N_15966);
or U16128 (N_16128,N_15826,N_15931);
or U16129 (N_16129,N_15846,N_15945);
nand U16130 (N_16130,N_15875,N_15930);
and U16131 (N_16131,N_15990,N_15858);
nor U16132 (N_16132,N_15820,N_15980);
nor U16133 (N_16133,N_15874,N_15880);
nand U16134 (N_16134,N_15949,N_15809);
nand U16135 (N_16135,N_15837,N_15991);
nor U16136 (N_16136,N_15891,N_15869);
or U16137 (N_16137,N_15934,N_15953);
xnor U16138 (N_16138,N_15965,N_15870);
or U16139 (N_16139,N_15995,N_15943);
nand U16140 (N_16140,N_15956,N_15858);
or U16141 (N_16141,N_15832,N_15823);
xnor U16142 (N_16142,N_15868,N_15885);
xor U16143 (N_16143,N_15995,N_15920);
nand U16144 (N_16144,N_15958,N_15836);
or U16145 (N_16145,N_15843,N_15817);
nand U16146 (N_16146,N_15950,N_15890);
and U16147 (N_16147,N_15824,N_15862);
nand U16148 (N_16148,N_15865,N_15969);
nor U16149 (N_16149,N_15994,N_15897);
and U16150 (N_16150,N_15930,N_15831);
nor U16151 (N_16151,N_15879,N_15994);
nand U16152 (N_16152,N_15996,N_15913);
or U16153 (N_16153,N_15891,N_15921);
xor U16154 (N_16154,N_15890,N_15884);
xnor U16155 (N_16155,N_15977,N_15824);
nand U16156 (N_16156,N_15973,N_15867);
nor U16157 (N_16157,N_15859,N_15831);
xnor U16158 (N_16158,N_15839,N_15911);
nor U16159 (N_16159,N_15908,N_15928);
nand U16160 (N_16160,N_15858,N_15907);
or U16161 (N_16161,N_15832,N_15942);
nor U16162 (N_16162,N_15981,N_15964);
xor U16163 (N_16163,N_15802,N_15932);
xnor U16164 (N_16164,N_15966,N_15993);
or U16165 (N_16165,N_15977,N_15931);
xnor U16166 (N_16166,N_15979,N_15920);
xor U16167 (N_16167,N_15918,N_15833);
nor U16168 (N_16168,N_15871,N_15813);
nor U16169 (N_16169,N_15863,N_15933);
xnor U16170 (N_16170,N_15828,N_15845);
nand U16171 (N_16171,N_15867,N_15900);
and U16172 (N_16172,N_15815,N_15883);
and U16173 (N_16173,N_15826,N_15818);
or U16174 (N_16174,N_15967,N_15991);
nor U16175 (N_16175,N_15824,N_15814);
nor U16176 (N_16176,N_15929,N_15998);
or U16177 (N_16177,N_15891,N_15913);
or U16178 (N_16178,N_15812,N_15856);
nand U16179 (N_16179,N_15887,N_15826);
nor U16180 (N_16180,N_15914,N_15898);
and U16181 (N_16181,N_15887,N_15812);
or U16182 (N_16182,N_15873,N_15985);
nor U16183 (N_16183,N_15922,N_15808);
nor U16184 (N_16184,N_15906,N_15845);
xnor U16185 (N_16185,N_15932,N_15977);
and U16186 (N_16186,N_15936,N_15873);
nor U16187 (N_16187,N_15925,N_15923);
xnor U16188 (N_16188,N_15905,N_15942);
xor U16189 (N_16189,N_15980,N_15966);
nand U16190 (N_16190,N_15844,N_15946);
nand U16191 (N_16191,N_15862,N_15883);
xor U16192 (N_16192,N_15836,N_15922);
and U16193 (N_16193,N_15997,N_15900);
nand U16194 (N_16194,N_15819,N_15941);
nand U16195 (N_16195,N_15853,N_15978);
nor U16196 (N_16196,N_15853,N_15867);
xnor U16197 (N_16197,N_15849,N_15975);
nor U16198 (N_16198,N_15966,N_15953);
nor U16199 (N_16199,N_15967,N_15910);
nor U16200 (N_16200,N_16179,N_16165);
or U16201 (N_16201,N_16115,N_16177);
nor U16202 (N_16202,N_16016,N_16045);
nor U16203 (N_16203,N_16094,N_16060);
xor U16204 (N_16204,N_16131,N_16031);
nand U16205 (N_16205,N_16176,N_16089);
nor U16206 (N_16206,N_16019,N_16057);
or U16207 (N_16207,N_16024,N_16123);
nor U16208 (N_16208,N_16059,N_16146);
or U16209 (N_16209,N_16041,N_16196);
nor U16210 (N_16210,N_16053,N_16051);
nor U16211 (N_16211,N_16187,N_16022);
and U16212 (N_16212,N_16056,N_16084);
nor U16213 (N_16213,N_16033,N_16172);
nand U16214 (N_16214,N_16110,N_16171);
or U16215 (N_16215,N_16182,N_16015);
or U16216 (N_16216,N_16096,N_16004);
nor U16217 (N_16217,N_16132,N_16030);
nor U16218 (N_16218,N_16032,N_16023);
xor U16219 (N_16219,N_16077,N_16193);
xor U16220 (N_16220,N_16046,N_16087);
or U16221 (N_16221,N_16166,N_16168);
nor U16222 (N_16222,N_16078,N_16050);
nor U16223 (N_16223,N_16184,N_16109);
and U16224 (N_16224,N_16076,N_16066);
and U16225 (N_16225,N_16070,N_16155);
nor U16226 (N_16226,N_16007,N_16067);
nor U16227 (N_16227,N_16020,N_16080);
and U16228 (N_16228,N_16150,N_16192);
xnor U16229 (N_16229,N_16163,N_16140);
xor U16230 (N_16230,N_16125,N_16174);
xnor U16231 (N_16231,N_16114,N_16058);
xor U16232 (N_16232,N_16002,N_16017);
xor U16233 (N_16233,N_16064,N_16164);
xnor U16234 (N_16234,N_16069,N_16111);
and U16235 (N_16235,N_16180,N_16061);
nand U16236 (N_16236,N_16122,N_16037);
and U16237 (N_16237,N_16011,N_16021);
or U16238 (N_16238,N_16044,N_16175);
nor U16239 (N_16239,N_16082,N_16107);
and U16240 (N_16240,N_16097,N_16026);
and U16241 (N_16241,N_16065,N_16185);
or U16242 (N_16242,N_16008,N_16113);
and U16243 (N_16243,N_16199,N_16048);
or U16244 (N_16244,N_16142,N_16014);
and U16245 (N_16245,N_16034,N_16012);
nor U16246 (N_16246,N_16093,N_16152);
or U16247 (N_16247,N_16038,N_16160);
nor U16248 (N_16248,N_16091,N_16001);
and U16249 (N_16249,N_16103,N_16198);
and U16250 (N_16250,N_16181,N_16112);
and U16251 (N_16251,N_16191,N_16124);
xor U16252 (N_16252,N_16137,N_16063);
xor U16253 (N_16253,N_16157,N_16042);
xnor U16254 (N_16254,N_16079,N_16104);
and U16255 (N_16255,N_16013,N_16105);
nor U16256 (N_16256,N_16086,N_16158);
or U16257 (N_16257,N_16153,N_16095);
or U16258 (N_16258,N_16144,N_16108);
and U16259 (N_16259,N_16043,N_16183);
xor U16260 (N_16260,N_16161,N_16003);
and U16261 (N_16261,N_16100,N_16075);
nand U16262 (N_16262,N_16098,N_16128);
xnor U16263 (N_16263,N_16085,N_16047);
nor U16264 (N_16264,N_16025,N_16138);
xor U16265 (N_16265,N_16149,N_16039);
xor U16266 (N_16266,N_16029,N_16169);
and U16267 (N_16267,N_16072,N_16197);
nand U16268 (N_16268,N_16006,N_16190);
and U16269 (N_16269,N_16143,N_16073);
xnor U16270 (N_16270,N_16134,N_16186);
xor U16271 (N_16271,N_16055,N_16136);
nand U16272 (N_16272,N_16092,N_16126);
xnor U16273 (N_16273,N_16083,N_16167);
xor U16274 (N_16274,N_16178,N_16195);
nor U16275 (N_16275,N_16071,N_16018);
xnor U16276 (N_16276,N_16088,N_16005);
or U16277 (N_16277,N_16090,N_16156);
and U16278 (N_16278,N_16074,N_16099);
xnor U16279 (N_16279,N_16119,N_16117);
nor U16280 (N_16280,N_16102,N_16062);
and U16281 (N_16281,N_16148,N_16054);
nor U16282 (N_16282,N_16130,N_16154);
nand U16283 (N_16283,N_16120,N_16000);
or U16284 (N_16284,N_16027,N_16118);
xor U16285 (N_16285,N_16036,N_16101);
and U16286 (N_16286,N_16170,N_16081);
nand U16287 (N_16287,N_16121,N_16159);
or U16288 (N_16288,N_16068,N_16127);
nor U16289 (N_16289,N_16139,N_16010);
nand U16290 (N_16290,N_16129,N_16188);
or U16291 (N_16291,N_16133,N_16173);
and U16292 (N_16292,N_16049,N_16145);
nand U16293 (N_16293,N_16141,N_16106);
nor U16294 (N_16294,N_16135,N_16147);
nand U16295 (N_16295,N_16052,N_16035);
xor U16296 (N_16296,N_16151,N_16040);
and U16297 (N_16297,N_16028,N_16162);
and U16298 (N_16298,N_16116,N_16189);
nor U16299 (N_16299,N_16009,N_16194);
xor U16300 (N_16300,N_16134,N_16116);
nor U16301 (N_16301,N_16107,N_16068);
nor U16302 (N_16302,N_16047,N_16169);
nor U16303 (N_16303,N_16175,N_16132);
and U16304 (N_16304,N_16080,N_16034);
nand U16305 (N_16305,N_16023,N_16072);
xnor U16306 (N_16306,N_16006,N_16063);
or U16307 (N_16307,N_16155,N_16105);
xnor U16308 (N_16308,N_16057,N_16030);
nor U16309 (N_16309,N_16123,N_16006);
nand U16310 (N_16310,N_16117,N_16052);
nor U16311 (N_16311,N_16026,N_16017);
xor U16312 (N_16312,N_16017,N_16147);
and U16313 (N_16313,N_16017,N_16095);
or U16314 (N_16314,N_16075,N_16069);
or U16315 (N_16315,N_16119,N_16044);
nand U16316 (N_16316,N_16174,N_16154);
nor U16317 (N_16317,N_16118,N_16016);
and U16318 (N_16318,N_16051,N_16106);
and U16319 (N_16319,N_16170,N_16089);
and U16320 (N_16320,N_16053,N_16010);
nor U16321 (N_16321,N_16087,N_16196);
and U16322 (N_16322,N_16193,N_16162);
nand U16323 (N_16323,N_16116,N_16062);
nor U16324 (N_16324,N_16125,N_16138);
nor U16325 (N_16325,N_16069,N_16191);
and U16326 (N_16326,N_16053,N_16101);
nand U16327 (N_16327,N_16068,N_16027);
nand U16328 (N_16328,N_16043,N_16078);
xnor U16329 (N_16329,N_16017,N_16033);
nor U16330 (N_16330,N_16040,N_16094);
xor U16331 (N_16331,N_16154,N_16014);
and U16332 (N_16332,N_16192,N_16066);
xor U16333 (N_16333,N_16049,N_16188);
nand U16334 (N_16334,N_16077,N_16143);
and U16335 (N_16335,N_16004,N_16127);
or U16336 (N_16336,N_16048,N_16131);
or U16337 (N_16337,N_16058,N_16043);
and U16338 (N_16338,N_16147,N_16016);
nand U16339 (N_16339,N_16151,N_16097);
or U16340 (N_16340,N_16057,N_16091);
and U16341 (N_16341,N_16045,N_16023);
or U16342 (N_16342,N_16193,N_16168);
or U16343 (N_16343,N_16169,N_16100);
nor U16344 (N_16344,N_16071,N_16169);
xnor U16345 (N_16345,N_16174,N_16009);
nand U16346 (N_16346,N_16069,N_16154);
nor U16347 (N_16347,N_16087,N_16193);
xor U16348 (N_16348,N_16042,N_16081);
nor U16349 (N_16349,N_16075,N_16073);
nand U16350 (N_16350,N_16150,N_16149);
nor U16351 (N_16351,N_16120,N_16181);
nand U16352 (N_16352,N_16143,N_16119);
or U16353 (N_16353,N_16063,N_16044);
xnor U16354 (N_16354,N_16149,N_16109);
xnor U16355 (N_16355,N_16025,N_16185);
nand U16356 (N_16356,N_16140,N_16173);
or U16357 (N_16357,N_16086,N_16064);
and U16358 (N_16358,N_16017,N_16157);
and U16359 (N_16359,N_16049,N_16110);
or U16360 (N_16360,N_16005,N_16098);
and U16361 (N_16361,N_16153,N_16131);
and U16362 (N_16362,N_16007,N_16025);
nand U16363 (N_16363,N_16130,N_16075);
nor U16364 (N_16364,N_16135,N_16096);
and U16365 (N_16365,N_16185,N_16180);
nor U16366 (N_16366,N_16194,N_16176);
and U16367 (N_16367,N_16077,N_16170);
nand U16368 (N_16368,N_16060,N_16185);
nor U16369 (N_16369,N_16049,N_16138);
xor U16370 (N_16370,N_16076,N_16037);
xnor U16371 (N_16371,N_16028,N_16137);
nor U16372 (N_16372,N_16013,N_16010);
or U16373 (N_16373,N_16091,N_16018);
or U16374 (N_16374,N_16058,N_16153);
nor U16375 (N_16375,N_16123,N_16105);
or U16376 (N_16376,N_16022,N_16147);
xnor U16377 (N_16377,N_16001,N_16104);
xnor U16378 (N_16378,N_16178,N_16042);
and U16379 (N_16379,N_16190,N_16046);
nand U16380 (N_16380,N_16098,N_16159);
nand U16381 (N_16381,N_16068,N_16185);
nand U16382 (N_16382,N_16059,N_16034);
nand U16383 (N_16383,N_16192,N_16162);
nor U16384 (N_16384,N_16100,N_16006);
nand U16385 (N_16385,N_16174,N_16072);
or U16386 (N_16386,N_16133,N_16018);
or U16387 (N_16387,N_16008,N_16058);
nor U16388 (N_16388,N_16170,N_16164);
or U16389 (N_16389,N_16081,N_16161);
and U16390 (N_16390,N_16076,N_16009);
nand U16391 (N_16391,N_16002,N_16154);
nor U16392 (N_16392,N_16185,N_16123);
nand U16393 (N_16393,N_16193,N_16030);
or U16394 (N_16394,N_16018,N_16006);
nor U16395 (N_16395,N_16108,N_16156);
nor U16396 (N_16396,N_16121,N_16111);
and U16397 (N_16397,N_16117,N_16183);
and U16398 (N_16398,N_16096,N_16009);
nand U16399 (N_16399,N_16142,N_16103);
xnor U16400 (N_16400,N_16265,N_16258);
and U16401 (N_16401,N_16313,N_16317);
or U16402 (N_16402,N_16341,N_16217);
or U16403 (N_16403,N_16200,N_16314);
and U16404 (N_16404,N_16228,N_16243);
nor U16405 (N_16405,N_16209,N_16336);
nor U16406 (N_16406,N_16304,N_16367);
nand U16407 (N_16407,N_16281,N_16215);
or U16408 (N_16408,N_16349,N_16241);
nor U16409 (N_16409,N_16284,N_16350);
or U16410 (N_16410,N_16214,N_16262);
and U16411 (N_16411,N_16259,N_16379);
xor U16412 (N_16412,N_16376,N_16357);
or U16413 (N_16413,N_16371,N_16225);
nor U16414 (N_16414,N_16295,N_16245);
and U16415 (N_16415,N_16252,N_16325);
and U16416 (N_16416,N_16239,N_16279);
and U16417 (N_16417,N_16315,N_16308);
and U16418 (N_16418,N_16227,N_16303);
nand U16419 (N_16419,N_16251,N_16360);
xnor U16420 (N_16420,N_16226,N_16391);
and U16421 (N_16421,N_16397,N_16362);
and U16422 (N_16422,N_16318,N_16211);
xnor U16423 (N_16423,N_16203,N_16261);
nor U16424 (N_16424,N_16329,N_16378);
and U16425 (N_16425,N_16338,N_16264);
nand U16426 (N_16426,N_16267,N_16277);
xor U16427 (N_16427,N_16319,N_16322);
or U16428 (N_16428,N_16298,N_16216);
or U16429 (N_16429,N_16290,N_16202);
xor U16430 (N_16430,N_16353,N_16271);
and U16431 (N_16431,N_16233,N_16399);
nor U16432 (N_16432,N_16289,N_16328);
nand U16433 (N_16433,N_16345,N_16201);
nor U16434 (N_16434,N_16230,N_16242);
xor U16435 (N_16435,N_16356,N_16244);
and U16436 (N_16436,N_16301,N_16263);
and U16437 (N_16437,N_16392,N_16310);
nor U16438 (N_16438,N_16358,N_16393);
nand U16439 (N_16439,N_16237,N_16282);
nor U16440 (N_16440,N_16285,N_16381);
nand U16441 (N_16441,N_16223,N_16294);
xor U16442 (N_16442,N_16316,N_16394);
xor U16443 (N_16443,N_16292,N_16246);
or U16444 (N_16444,N_16388,N_16369);
or U16445 (N_16445,N_16339,N_16343);
or U16446 (N_16446,N_16275,N_16361);
or U16447 (N_16447,N_16248,N_16299);
nor U16448 (N_16448,N_16221,N_16309);
nor U16449 (N_16449,N_16398,N_16347);
or U16450 (N_16450,N_16354,N_16320);
nand U16451 (N_16451,N_16365,N_16324);
or U16452 (N_16452,N_16218,N_16331);
nand U16453 (N_16453,N_16302,N_16213);
nor U16454 (N_16454,N_16236,N_16384);
nand U16455 (N_16455,N_16288,N_16344);
or U16456 (N_16456,N_16368,N_16250);
nor U16457 (N_16457,N_16300,N_16395);
nand U16458 (N_16458,N_16208,N_16386);
nand U16459 (N_16459,N_16312,N_16274);
nand U16460 (N_16460,N_16297,N_16293);
and U16461 (N_16461,N_16366,N_16206);
nor U16462 (N_16462,N_16340,N_16351);
and U16463 (N_16463,N_16387,N_16273);
nor U16464 (N_16464,N_16210,N_16337);
or U16465 (N_16465,N_16305,N_16330);
or U16466 (N_16466,N_16270,N_16253);
xnor U16467 (N_16467,N_16334,N_16272);
nand U16468 (N_16468,N_16377,N_16222);
xor U16469 (N_16469,N_16238,N_16260);
and U16470 (N_16470,N_16342,N_16254);
or U16471 (N_16471,N_16326,N_16355);
or U16472 (N_16472,N_16364,N_16219);
nor U16473 (N_16473,N_16224,N_16257);
nor U16474 (N_16474,N_16352,N_16380);
nor U16475 (N_16475,N_16291,N_16268);
and U16476 (N_16476,N_16348,N_16255);
or U16477 (N_16477,N_16389,N_16327);
nand U16478 (N_16478,N_16383,N_16247);
xor U16479 (N_16479,N_16269,N_16373);
nor U16480 (N_16480,N_16212,N_16359);
nand U16481 (N_16481,N_16286,N_16363);
nor U16482 (N_16482,N_16278,N_16375);
and U16483 (N_16483,N_16280,N_16266);
or U16484 (N_16484,N_16390,N_16333);
nand U16485 (N_16485,N_16220,N_16287);
and U16486 (N_16486,N_16306,N_16307);
xor U16487 (N_16487,N_16204,N_16249);
and U16488 (N_16488,N_16396,N_16374);
xor U16489 (N_16489,N_16332,N_16296);
and U16490 (N_16490,N_16372,N_16240);
nand U16491 (N_16491,N_16335,N_16205);
nor U16492 (N_16492,N_16229,N_16231);
or U16493 (N_16493,N_16323,N_16370);
nand U16494 (N_16494,N_16321,N_16232);
xnor U16495 (N_16495,N_16311,N_16276);
nand U16496 (N_16496,N_16234,N_16346);
or U16497 (N_16497,N_16283,N_16235);
nor U16498 (N_16498,N_16385,N_16207);
nand U16499 (N_16499,N_16382,N_16256);
nand U16500 (N_16500,N_16224,N_16339);
or U16501 (N_16501,N_16210,N_16347);
xnor U16502 (N_16502,N_16244,N_16387);
or U16503 (N_16503,N_16272,N_16280);
or U16504 (N_16504,N_16248,N_16298);
and U16505 (N_16505,N_16354,N_16355);
nor U16506 (N_16506,N_16338,N_16381);
nand U16507 (N_16507,N_16337,N_16357);
nand U16508 (N_16508,N_16227,N_16322);
xnor U16509 (N_16509,N_16341,N_16316);
nor U16510 (N_16510,N_16208,N_16244);
xor U16511 (N_16511,N_16201,N_16322);
xnor U16512 (N_16512,N_16296,N_16338);
or U16513 (N_16513,N_16225,N_16237);
xnor U16514 (N_16514,N_16332,N_16308);
and U16515 (N_16515,N_16390,N_16241);
xnor U16516 (N_16516,N_16205,N_16279);
xor U16517 (N_16517,N_16313,N_16341);
nand U16518 (N_16518,N_16342,N_16308);
xnor U16519 (N_16519,N_16290,N_16342);
xnor U16520 (N_16520,N_16282,N_16269);
and U16521 (N_16521,N_16267,N_16384);
nor U16522 (N_16522,N_16399,N_16360);
nor U16523 (N_16523,N_16321,N_16248);
and U16524 (N_16524,N_16398,N_16326);
nor U16525 (N_16525,N_16329,N_16353);
and U16526 (N_16526,N_16219,N_16282);
and U16527 (N_16527,N_16229,N_16257);
or U16528 (N_16528,N_16338,N_16258);
nand U16529 (N_16529,N_16311,N_16384);
xnor U16530 (N_16530,N_16287,N_16384);
xnor U16531 (N_16531,N_16205,N_16299);
nor U16532 (N_16532,N_16370,N_16394);
nor U16533 (N_16533,N_16366,N_16232);
xor U16534 (N_16534,N_16234,N_16291);
nand U16535 (N_16535,N_16325,N_16381);
or U16536 (N_16536,N_16307,N_16234);
nand U16537 (N_16537,N_16347,N_16394);
and U16538 (N_16538,N_16200,N_16387);
nor U16539 (N_16539,N_16236,N_16337);
xnor U16540 (N_16540,N_16315,N_16374);
xnor U16541 (N_16541,N_16273,N_16240);
and U16542 (N_16542,N_16329,N_16262);
and U16543 (N_16543,N_16376,N_16244);
nand U16544 (N_16544,N_16247,N_16273);
or U16545 (N_16545,N_16309,N_16338);
nor U16546 (N_16546,N_16210,N_16300);
or U16547 (N_16547,N_16380,N_16339);
or U16548 (N_16548,N_16263,N_16234);
and U16549 (N_16549,N_16362,N_16237);
xor U16550 (N_16550,N_16313,N_16242);
and U16551 (N_16551,N_16252,N_16307);
and U16552 (N_16552,N_16278,N_16267);
nor U16553 (N_16553,N_16300,N_16272);
and U16554 (N_16554,N_16288,N_16393);
or U16555 (N_16555,N_16395,N_16271);
nand U16556 (N_16556,N_16211,N_16309);
nand U16557 (N_16557,N_16271,N_16291);
nor U16558 (N_16558,N_16369,N_16206);
xnor U16559 (N_16559,N_16379,N_16254);
xnor U16560 (N_16560,N_16236,N_16230);
nand U16561 (N_16561,N_16316,N_16274);
or U16562 (N_16562,N_16370,N_16236);
nor U16563 (N_16563,N_16267,N_16223);
and U16564 (N_16564,N_16395,N_16371);
nand U16565 (N_16565,N_16241,N_16311);
xnor U16566 (N_16566,N_16312,N_16264);
or U16567 (N_16567,N_16263,N_16295);
nor U16568 (N_16568,N_16280,N_16257);
and U16569 (N_16569,N_16291,N_16317);
nand U16570 (N_16570,N_16262,N_16316);
and U16571 (N_16571,N_16255,N_16332);
nor U16572 (N_16572,N_16332,N_16289);
xnor U16573 (N_16573,N_16284,N_16220);
nand U16574 (N_16574,N_16375,N_16248);
nor U16575 (N_16575,N_16234,N_16288);
nand U16576 (N_16576,N_16206,N_16385);
nor U16577 (N_16577,N_16284,N_16330);
xnor U16578 (N_16578,N_16389,N_16291);
nand U16579 (N_16579,N_16327,N_16267);
xor U16580 (N_16580,N_16321,N_16281);
xnor U16581 (N_16581,N_16276,N_16290);
nand U16582 (N_16582,N_16378,N_16355);
nor U16583 (N_16583,N_16285,N_16294);
or U16584 (N_16584,N_16312,N_16325);
nand U16585 (N_16585,N_16282,N_16223);
or U16586 (N_16586,N_16374,N_16357);
nor U16587 (N_16587,N_16329,N_16283);
and U16588 (N_16588,N_16273,N_16282);
or U16589 (N_16589,N_16351,N_16308);
nor U16590 (N_16590,N_16335,N_16248);
or U16591 (N_16591,N_16278,N_16342);
nor U16592 (N_16592,N_16308,N_16386);
and U16593 (N_16593,N_16230,N_16388);
nor U16594 (N_16594,N_16299,N_16382);
or U16595 (N_16595,N_16324,N_16240);
xor U16596 (N_16596,N_16315,N_16369);
nand U16597 (N_16597,N_16288,N_16241);
or U16598 (N_16598,N_16307,N_16394);
nand U16599 (N_16599,N_16318,N_16381);
nor U16600 (N_16600,N_16424,N_16414);
or U16601 (N_16601,N_16530,N_16503);
and U16602 (N_16602,N_16411,N_16553);
nor U16603 (N_16603,N_16513,N_16481);
xor U16604 (N_16604,N_16408,N_16573);
xnor U16605 (N_16605,N_16592,N_16574);
nand U16606 (N_16606,N_16404,N_16580);
nor U16607 (N_16607,N_16551,N_16474);
nor U16608 (N_16608,N_16599,N_16577);
or U16609 (N_16609,N_16486,N_16462);
or U16610 (N_16610,N_16479,N_16536);
nand U16611 (N_16611,N_16526,N_16512);
xnor U16612 (N_16612,N_16522,N_16423);
xnor U16613 (N_16613,N_16409,N_16500);
xnor U16614 (N_16614,N_16528,N_16436);
nand U16615 (N_16615,N_16435,N_16588);
nor U16616 (N_16616,N_16446,N_16562);
nor U16617 (N_16617,N_16456,N_16568);
nor U16618 (N_16618,N_16549,N_16590);
and U16619 (N_16619,N_16506,N_16478);
xor U16620 (N_16620,N_16485,N_16405);
nand U16621 (N_16621,N_16468,N_16412);
or U16622 (N_16622,N_16450,N_16529);
or U16623 (N_16623,N_16463,N_16586);
xnor U16624 (N_16624,N_16587,N_16507);
and U16625 (N_16625,N_16417,N_16516);
and U16626 (N_16626,N_16487,N_16499);
or U16627 (N_16627,N_16439,N_16473);
and U16628 (N_16628,N_16504,N_16482);
nor U16629 (N_16629,N_16469,N_16401);
and U16630 (N_16630,N_16451,N_16440);
xnor U16631 (N_16631,N_16567,N_16497);
and U16632 (N_16632,N_16565,N_16581);
and U16633 (N_16633,N_16496,N_16596);
nand U16634 (N_16634,N_16544,N_16537);
and U16635 (N_16635,N_16552,N_16557);
xnor U16636 (N_16636,N_16492,N_16445);
and U16637 (N_16637,N_16548,N_16584);
nor U16638 (N_16638,N_16515,N_16476);
xor U16639 (N_16639,N_16470,N_16595);
or U16640 (N_16640,N_16457,N_16461);
nor U16641 (N_16641,N_16583,N_16525);
or U16642 (N_16642,N_16533,N_16410);
or U16643 (N_16643,N_16523,N_16582);
nand U16644 (N_16644,N_16421,N_16542);
or U16645 (N_16645,N_16501,N_16598);
nand U16646 (N_16646,N_16594,N_16493);
or U16647 (N_16647,N_16495,N_16402);
or U16648 (N_16648,N_16466,N_16420);
and U16649 (N_16649,N_16431,N_16475);
xnor U16650 (N_16650,N_16422,N_16494);
nor U16651 (N_16651,N_16521,N_16453);
nand U16652 (N_16652,N_16407,N_16449);
and U16653 (N_16653,N_16563,N_16419);
or U16654 (N_16654,N_16576,N_16467);
nand U16655 (N_16655,N_16550,N_16403);
nand U16656 (N_16656,N_16535,N_16491);
nand U16657 (N_16657,N_16532,N_16559);
nand U16658 (N_16658,N_16441,N_16418);
xor U16659 (N_16659,N_16593,N_16508);
or U16660 (N_16660,N_16538,N_16442);
nor U16661 (N_16661,N_16460,N_16502);
nor U16662 (N_16662,N_16444,N_16558);
nor U16663 (N_16663,N_16406,N_16517);
xor U16664 (N_16664,N_16540,N_16527);
xor U16665 (N_16665,N_16471,N_16572);
xnor U16666 (N_16666,N_16570,N_16531);
or U16667 (N_16667,N_16545,N_16430);
nor U16668 (N_16668,N_16556,N_16585);
and U16669 (N_16669,N_16589,N_16452);
or U16670 (N_16670,N_16413,N_16429);
or U16671 (N_16671,N_16541,N_16564);
xor U16672 (N_16672,N_16561,N_16575);
xor U16673 (N_16673,N_16597,N_16591);
nand U16674 (N_16674,N_16448,N_16509);
xnor U16675 (N_16675,N_16438,N_16543);
nand U16676 (N_16676,N_16510,N_16578);
and U16677 (N_16677,N_16459,N_16511);
and U16678 (N_16678,N_16498,N_16505);
nor U16679 (N_16679,N_16400,N_16554);
nor U16680 (N_16680,N_16428,N_16569);
xnor U16681 (N_16681,N_16484,N_16579);
or U16682 (N_16682,N_16518,N_16514);
nor U16683 (N_16683,N_16483,N_16454);
or U16684 (N_16684,N_16534,N_16519);
nor U16685 (N_16685,N_16480,N_16546);
nand U16686 (N_16686,N_16425,N_16472);
nand U16687 (N_16687,N_16571,N_16433);
or U16688 (N_16688,N_16520,N_16539);
nand U16689 (N_16689,N_16434,N_16489);
xor U16690 (N_16690,N_16547,N_16427);
nand U16691 (N_16691,N_16415,N_16458);
xor U16692 (N_16692,N_16555,N_16465);
or U16693 (N_16693,N_16432,N_16437);
nor U16694 (N_16694,N_16488,N_16443);
xnor U16695 (N_16695,N_16416,N_16464);
nor U16696 (N_16696,N_16566,N_16426);
xnor U16697 (N_16697,N_16560,N_16524);
and U16698 (N_16698,N_16490,N_16447);
nand U16699 (N_16699,N_16477,N_16455);
or U16700 (N_16700,N_16438,N_16584);
or U16701 (N_16701,N_16507,N_16549);
xor U16702 (N_16702,N_16475,N_16505);
or U16703 (N_16703,N_16465,N_16475);
xor U16704 (N_16704,N_16435,N_16595);
and U16705 (N_16705,N_16484,N_16585);
nor U16706 (N_16706,N_16477,N_16528);
and U16707 (N_16707,N_16559,N_16428);
and U16708 (N_16708,N_16507,N_16404);
or U16709 (N_16709,N_16516,N_16546);
nor U16710 (N_16710,N_16482,N_16525);
and U16711 (N_16711,N_16546,N_16515);
nand U16712 (N_16712,N_16535,N_16457);
nor U16713 (N_16713,N_16503,N_16490);
and U16714 (N_16714,N_16438,N_16408);
nand U16715 (N_16715,N_16501,N_16506);
or U16716 (N_16716,N_16558,N_16462);
nor U16717 (N_16717,N_16502,N_16416);
nor U16718 (N_16718,N_16461,N_16545);
nand U16719 (N_16719,N_16497,N_16458);
or U16720 (N_16720,N_16416,N_16535);
and U16721 (N_16721,N_16464,N_16461);
or U16722 (N_16722,N_16567,N_16539);
or U16723 (N_16723,N_16503,N_16580);
nand U16724 (N_16724,N_16462,N_16530);
and U16725 (N_16725,N_16427,N_16403);
and U16726 (N_16726,N_16422,N_16581);
and U16727 (N_16727,N_16494,N_16530);
or U16728 (N_16728,N_16548,N_16586);
nor U16729 (N_16729,N_16559,N_16571);
nand U16730 (N_16730,N_16532,N_16536);
nor U16731 (N_16731,N_16403,N_16460);
or U16732 (N_16732,N_16599,N_16498);
nor U16733 (N_16733,N_16406,N_16495);
nand U16734 (N_16734,N_16524,N_16579);
nor U16735 (N_16735,N_16556,N_16404);
xor U16736 (N_16736,N_16463,N_16493);
nand U16737 (N_16737,N_16412,N_16495);
nor U16738 (N_16738,N_16577,N_16440);
nand U16739 (N_16739,N_16496,N_16564);
nor U16740 (N_16740,N_16528,N_16598);
nor U16741 (N_16741,N_16493,N_16488);
nand U16742 (N_16742,N_16586,N_16487);
xnor U16743 (N_16743,N_16424,N_16546);
xor U16744 (N_16744,N_16532,N_16491);
or U16745 (N_16745,N_16552,N_16427);
and U16746 (N_16746,N_16494,N_16548);
nand U16747 (N_16747,N_16477,N_16493);
nor U16748 (N_16748,N_16597,N_16446);
or U16749 (N_16749,N_16506,N_16596);
nor U16750 (N_16750,N_16423,N_16437);
or U16751 (N_16751,N_16490,N_16487);
or U16752 (N_16752,N_16433,N_16543);
xnor U16753 (N_16753,N_16544,N_16469);
nor U16754 (N_16754,N_16545,N_16423);
nor U16755 (N_16755,N_16468,N_16591);
nand U16756 (N_16756,N_16486,N_16593);
nand U16757 (N_16757,N_16573,N_16421);
or U16758 (N_16758,N_16424,N_16490);
and U16759 (N_16759,N_16513,N_16461);
and U16760 (N_16760,N_16430,N_16587);
nand U16761 (N_16761,N_16502,N_16569);
and U16762 (N_16762,N_16555,N_16452);
and U16763 (N_16763,N_16501,N_16522);
xor U16764 (N_16764,N_16444,N_16598);
and U16765 (N_16765,N_16442,N_16434);
or U16766 (N_16766,N_16446,N_16504);
nor U16767 (N_16767,N_16443,N_16564);
nand U16768 (N_16768,N_16474,N_16552);
nand U16769 (N_16769,N_16406,N_16492);
xor U16770 (N_16770,N_16582,N_16599);
nand U16771 (N_16771,N_16582,N_16487);
or U16772 (N_16772,N_16485,N_16578);
nor U16773 (N_16773,N_16596,N_16429);
nand U16774 (N_16774,N_16456,N_16416);
xnor U16775 (N_16775,N_16513,N_16512);
nor U16776 (N_16776,N_16503,N_16441);
nand U16777 (N_16777,N_16436,N_16495);
and U16778 (N_16778,N_16504,N_16530);
or U16779 (N_16779,N_16503,N_16495);
nand U16780 (N_16780,N_16529,N_16564);
or U16781 (N_16781,N_16422,N_16476);
and U16782 (N_16782,N_16546,N_16437);
nor U16783 (N_16783,N_16550,N_16448);
and U16784 (N_16784,N_16594,N_16581);
xor U16785 (N_16785,N_16461,N_16427);
nand U16786 (N_16786,N_16432,N_16459);
or U16787 (N_16787,N_16408,N_16550);
or U16788 (N_16788,N_16565,N_16505);
and U16789 (N_16789,N_16533,N_16581);
and U16790 (N_16790,N_16573,N_16419);
nor U16791 (N_16791,N_16400,N_16409);
nor U16792 (N_16792,N_16472,N_16561);
nor U16793 (N_16793,N_16533,N_16573);
nand U16794 (N_16794,N_16530,N_16529);
or U16795 (N_16795,N_16513,N_16551);
and U16796 (N_16796,N_16429,N_16425);
nor U16797 (N_16797,N_16465,N_16526);
nor U16798 (N_16798,N_16511,N_16439);
or U16799 (N_16799,N_16472,N_16533);
xor U16800 (N_16800,N_16646,N_16704);
nor U16801 (N_16801,N_16670,N_16642);
and U16802 (N_16802,N_16621,N_16743);
nor U16803 (N_16803,N_16639,N_16707);
or U16804 (N_16804,N_16647,N_16784);
nand U16805 (N_16805,N_16659,N_16702);
and U16806 (N_16806,N_16628,N_16788);
nand U16807 (N_16807,N_16715,N_16780);
nor U16808 (N_16808,N_16769,N_16636);
and U16809 (N_16809,N_16705,N_16732);
or U16810 (N_16810,N_16783,N_16701);
nand U16811 (N_16811,N_16664,N_16717);
or U16812 (N_16812,N_16722,N_16785);
nand U16813 (N_16813,N_16624,N_16608);
xor U16814 (N_16814,N_16792,N_16626);
xor U16815 (N_16815,N_16612,N_16610);
and U16816 (N_16816,N_16652,N_16791);
nand U16817 (N_16817,N_16625,N_16775);
nand U16818 (N_16818,N_16727,N_16607);
and U16819 (N_16819,N_16677,N_16728);
or U16820 (N_16820,N_16657,N_16737);
or U16821 (N_16821,N_16772,N_16739);
nor U16822 (N_16822,N_16620,N_16731);
nor U16823 (N_16823,N_16766,N_16640);
nand U16824 (N_16824,N_16662,N_16763);
nor U16825 (N_16825,N_16755,N_16684);
xor U16826 (N_16826,N_16767,N_16648);
nor U16827 (N_16827,N_16712,N_16794);
or U16828 (N_16828,N_16760,N_16713);
nor U16829 (N_16829,N_16771,N_16759);
and U16830 (N_16830,N_16683,N_16645);
xnor U16831 (N_16831,N_16603,N_16706);
or U16832 (N_16832,N_16623,N_16663);
or U16833 (N_16833,N_16693,N_16700);
nor U16834 (N_16834,N_16616,N_16619);
or U16835 (N_16835,N_16776,N_16793);
and U16836 (N_16836,N_16615,N_16708);
or U16837 (N_16837,N_16740,N_16653);
xor U16838 (N_16838,N_16751,N_16724);
nand U16839 (N_16839,N_16644,N_16643);
xnor U16840 (N_16840,N_16609,N_16752);
nor U16841 (N_16841,N_16696,N_16742);
nand U16842 (N_16842,N_16757,N_16638);
or U16843 (N_16843,N_16611,N_16736);
and U16844 (N_16844,N_16668,N_16667);
nor U16845 (N_16845,N_16754,N_16725);
and U16846 (N_16846,N_16673,N_16654);
and U16847 (N_16847,N_16779,N_16730);
or U16848 (N_16848,N_16600,N_16681);
xnor U16849 (N_16849,N_16789,N_16690);
and U16850 (N_16850,N_16686,N_16768);
xnor U16851 (N_16851,N_16680,N_16658);
and U16852 (N_16852,N_16738,N_16689);
and U16853 (N_16853,N_16735,N_16637);
nor U16854 (N_16854,N_16634,N_16633);
nor U16855 (N_16855,N_16666,N_16632);
xor U16856 (N_16856,N_16758,N_16782);
and U16857 (N_16857,N_16765,N_16714);
and U16858 (N_16858,N_16606,N_16698);
and U16859 (N_16859,N_16674,N_16691);
and U16860 (N_16860,N_16795,N_16719);
nand U16861 (N_16861,N_16744,N_16641);
nor U16862 (N_16862,N_16720,N_16650);
and U16863 (N_16863,N_16747,N_16786);
and U16864 (N_16864,N_16799,N_16622);
or U16865 (N_16865,N_16679,N_16703);
nand U16866 (N_16866,N_16687,N_16798);
xor U16867 (N_16867,N_16797,N_16790);
nor U16868 (N_16868,N_16692,N_16614);
nor U16869 (N_16869,N_16726,N_16605);
nand U16870 (N_16870,N_16694,N_16675);
nand U16871 (N_16871,N_16729,N_16734);
nor U16872 (N_16872,N_16672,N_16709);
or U16873 (N_16873,N_16749,N_16750);
nor U16874 (N_16874,N_16723,N_16601);
nor U16875 (N_16875,N_16651,N_16629);
xnor U16876 (N_16876,N_16796,N_16617);
xor U16877 (N_16877,N_16656,N_16669);
xor U16878 (N_16878,N_16746,N_16613);
and U16879 (N_16879,N_16774,N_16745);
and U16880 (N_16880,N_16718,N_16604);
or U16881 (N_16881,N_16685,N_16741);
xor U16882 (N_16882,N_16762,N_16753);
and U16883 (N_16883,N_16661,N_16655);
nor U16884 (N_16884,N_16787,N_16770);
xnor U16885 (N_16885,N_16781,N_16716);
nand U16886 (N_16886,N_16682,N_16773);
and U16887 (N_16887,N_16602,N_16695);
nor U16888 (N_16888,N_16630,N_16721);
xor U16889 (N_16889,N_16777,N_16618);
and U16890 (N_16890,N_16748,N_16711);
and U16891 (N_16891,N_16676,N_16627);
nor U16892 (N_16892,N_16660,N_16710);
xor U16893 (N_16893,N_16697,N_16756);
or U16894 (N_16894,N_16733,N_16635);
and U16895 (N_16895,N_16678,N_16699);
or U16896 (N_16896,N_16778,N_16764);
and U16897 (N_16897,N_16688,N_16631);
nand U16898 (N_16898,N_16649,N_16665);
nand U16899 (N_16899,N_16671,N_16761);
nand U16900 (N_16900,N_16614,N_16766);
and U16901 (N_16901,N_16648,N_16665);
nand U16902 (N_16902,N_16709,N_16736);
nand U16903 (N_16903,N_16732,N_16763);
xnor U16904 (N_16904,N_16747,N_16642);
and U16905 (N_16905,N_16777,N_16747);
xnor U16906 (N_16906,N_16622,N_16627);
xnor U16907 (N_16907,N_16728,N_16672);
nor U16908 (N_16908,N_16744,N_16741);
or U16909 (N_16909,N_16730,N_16757);
xor U16910 (N_16910,N_16615,N_16608);
or U16911 (N_16911,N_16760,N_16745);
xor U16912 (N_16912,N_16757,N_16678);
and U16913 (N_16913,N_16791,N_16748);
and U16914 (N_16914,N_16626,N_16634);
nand U16915 (N_16915,N_16717,N_16611);
nand U16916 (N_16916,N_16697,N_16685);
nand U16917 (N_16917,N_16615,N_16638);
nand U16918 (N_16918,N_16703,N_16604);
nor U16919 (N_16919,N_16676,N_16730);
nand U16920 (N_16920,N_16784,N_16738);
or U16921 (N_16921,N_16775,N_16724);
and U16922 (N_16922,N_16648,N_16620);
xnor U16923 (N_16923,N_16714,N_16672);
or U16924 (N_16924,N_16653,N_16729);
and U16925 (N_16925,N_16604,N_16686);
and U16926 (N_16926,N_16642,N_16787);
nor U16927 (N_16927,N_16663,N_16622);
nor U16928 (N_16928,N_16796,N_16795);
or U16929 (N_16929,N_16688,N_16685);
nor U16930 (N_16930,N_16762,N_16735);
nand U16931 (N_16931,N_16742,N_16688);
and U16932 (N_16932,N_16749,N_16624);
nor U16933 (N_16933,N_16773,N_16736);
nand U16934 (N_16934,N_16622,N_16600);
xor U16935 (N_16935,N_16633,N_16659);
xnor U16936 (N_16936,N_16604,N_16622);
or U16937 (N_16937,N_16775,N_16742);
xor U16938 (N_16938,N_16640,N_16611);
nand U16939 (N_16939,N_16770,N_16671);
or U16940 (N_16940,N_16629,N_16635);
xnor U16941 (N_16941,N_16693,N_16694);
or U16942 (N_16942,N_16647,N_16623);
or U16943 (N_16943,N_16665,N_16675);
or U16944 (N_16944,N_16665,N_16667);
or U16945 (N_16945,N_16640,N_16616);
or U16946 (N_16946,N_16713,N_16734);
xor U16947 (N_16947,N_16687,N_16650);
nand U16948 (N_16948,N_16721,N_16775);
nand U16949 (N_16949,N_16671,N_16798);
and U16950 (N_16950,N_16795,N_16613);
and U16951 (N_16951,N_16670,N_16664);
xor U16952 (N_16952,N_16605,N_16736);
and U16953 (N_16953,N_16787,N_16650);
and U16954 (N_16954,N_16604,N_16644);
or U16955 (N_16955,N_16682,N_16668);
xnor U16956 (N_16956,N_16723,N_16776);
nor U16957 (N_16957,N_16682,N_16748);
nand U16958 (N_16958,N_16739,N_16691);
nand U16959 (N_16959,N_16736,N_16761);
xor U16960 (N_16960,N_16634,N_16692);
nor U16961 (N_16961,N_16782,N_16776);
nand U16962 (N_16962,N_16660,N_16770);
xor U16963 (N_16963,N_16625,N_16794);
xnor U16964 (N_16964,N_16683,N_16796);
xor U16965 (N_16965,N_16623,N_16766);
nand U16966 (N_16966,N_16657,N_16782);
and U16967 (N_16967,N_16619,N_16653);
nor U16968 (N_16968,N_16784,N_16638);
xnor U16969 (N_16969,N_16705,N_16613);
nand U16970 (N_16970,N_16761,N_16630);
and U16971 (N_16971,N_16611,N_16663);
and U16972 (N_16972,N_16756,N_16787);
nand U16973 (N_16973,N_16675,N_16769);
or U16974 (N_16974,N_16795,N_16746);
nand U16975 (N_16975,N_16605,N_16644);
or U16976 (N_16976,N_16664,N_16725);
or U16977 (N_16977,N_16706,N_16683);
nand U16978 (N_16978,N_16775,N_16681);
and U16979 (N_16979,N_16633,N_16636);
nor U16980 (N_16980,N_16629,N_16763);
nand U16981 (N_16981,N_16623,N_16705);
and U16982 (N_16982,N_16752,N_16695);
or U16983 (N_16983,N_16780,N_16649);
and U16984 (N_16984,N_16653,N_16610);
nor U16985 (N_16985,N_16789,N_16721);
nor U16986 (N_16986,N_16621,N_16734);
nor U16987 (N_16987,N_16703,N_16738);
xnor U16988 (N_16988,N_16665,N_16637);
or U16989 (N_16989,N_16635,N_16615);
xnor U16990 (N_16990,N_16619,N_16636);
nor U16991 (N_16991,N_16699,N_16670);
and U16992 (N_16992,N_16720,N_16768);
nor U16993 (N_16993,N_16737,N_16650);
xnor U16994 (N_16994,N_16799,N_16760);
and U16995 (N_16995,N_16617,N_16673);
and U16996 (N_16996,N_16690,N_16641);
or U16997 (N_16997,N_16772,N_16746);
nor U16998 (N_16998,N_16613,N_16676);
and U16999 (N_16999,N_16755,N_16661);
nor U17000 (N_17000,N_16928,N_16870);
xor U17001 (N_17001,N_16819,N_16834);
nor U17002 (N_17002,N_16926,N_16839);
or U17003 (N_17003,N_16816,N_16802);
nand U17004 (N_17004,N_16916,N_16821);
nand U17005 (N_17005,N_16950,N_16830);
and U17006 (N_17006,N_16866,N_16893);
nand U17007 (N_17007,N_16887,N_16898);
and U17008 (N_17008,N_16854,N_16925);
xor U17009 (N_17009,N_16997,N_16946);
nor U17010 (N_17010,N_16813,N_16879);
nand U17011 (N_17011,N_16954,N_16959);
nand U17012 (N_17012,N_16920,N_16840);
nand U17013 (N_17013,N_16858,N_16972);
and U17014 (N_17014,N_16951,N_16957);
and U17015 (N_17015,N_16810,N_16909);
or U17016 (N_17016,N_16968,N_16889);
or U17017 (N_17017,N_16941,N_16838);
or U17018 (N_17018,N_16938,N_16882);
and U17019 (N_17019,N_16930,N_16892);
and U17020 (N_17020,N_16970,N_16935);
or U17021 (N_17021,N_16912,N_16988);
or U17022 (N_17022,N_16921,N_16817);
and U17023 (N_17023,N_16986,N_16853);
xnor U17024 (N_17024,N_16875,N_16998);
or U17025 (N_17025,N_16848,N_16936);
nor U17026 (N_17026,N_16971,N_16828);
and U17027 (N_17027,N_16977,N_16901);
or U17028 (N_17028,N_16974,N_16845);
xnor U17029 (N_17029,N_16976,N_16984);
and U17030 (N_17030,N_16900,N_16857);
or U17031 (N_17031,N_16815,N_16823);
nor U17032 (N_17032,N_16805,N_16965);
xor U17033 (N_17033,N_16982,N_16963);
nor U17034 (N_17034,N_16964,N_16842);
xnor U17035 (N_17035,N_16924,N_16871);
xnor U17036 (N_17036,N_16876,N_16826);
and U17037 (N_17037,N_16904,N_16944);
or U17038 (N_17038,N_16983,N_16877);
xnor U17039 (N_17039,N_16843,N_16993);
nand U17040 (N_17040,N_16956,N_16814);
nor U17041 (N_17041,N_16915,N_16897);
xnor U17042 (N_17042,N_16937,N_16812);
xnor U17043 (N_17043,N_16911,N_16981);
xor U17044 (N_17044,N_16880,N_16960);
xnor U17045 (N_17045,N_16999,N_16829);
and U17046 (N_17046,N_16859,N_16894);
and U17047 (N_17047,N_16837,N_16991);
and U17048 (N_17048,N_16851,N_16811);
xor U17049 (N_17049,N_16989,N_16808);
nor U17050 (N_17050,N_16918,N_16992);
xnor U17051 (N_17051,N_16869,N_16940);
or U17052 (N_17052,N_16907,N_16932);
or U17053 (N_17053,N_16891,N_16995);
or U17054 (N_17054,N_16807,N_16899);
or U17055 (N_17055,N_16903,N_16927);
or U17056 (N_17056,N_16943,N_16919);
nand U17057 (N_17057,N_16990,N_16873);
or U17058 (N_17058,N_16906,N_16910);
and U17059 (N_17059,N_16867,N_16969);
or U17060 (N_17060,N_16905,N_16832);
xnor U17061 (N_17061,N_16888,N_16945);
xor U17062 (N_17062,N_16929,N_16953);
nand U17063 (N_17063,N_16881,N_16825);
and U17064 (N_17064,N_16962,N_16896);
and U17065 (N_17065,N_16978,N_16934);
and U17066 (N_17066,N_16985,N_16818);
nand U17067 (N_17067,N_16847,N_16958);
or U17068 (N_17068,N_16979,N_16966);
nor U17069 (N_17069,N_16856,N_16806);
xnor U17070 (N_17070,N_16931,N_16955);
and U17071 (N_17071,N_16886,N_16884);
and U17072 (N_17072,N_16947,N_16874);
xor U17073 (N_17073,N_16827,N_16987);
nor U17074 (N_17074,N_16824,N_16849);
xor U17075 (N_17075,N_16850,N_16895);
nand U17076 (N_17076,N_16861,N_16868);
nor U17077 (N_17077,N_16980,N_16800);
and U17078 (N_17078,N_16942,N_16801);
xnor U17079 (N_17079,N_16860,N_16878);
nor U17080 (N_17080,N_16933,N_16831);
and U17081 (N_17081,N_16809,N_16820);
nand U17082 (N_17082,N_16833,N_16865);
nand U17083 (N_17083,N_16914,N_16917);
nor U17084 (N_17084,N_16952,N_16862);
nand U17085 (N_17085,N_16846,N_16949);
and U17086 (N_17086,N_16835,N_16913);
and U17087 (N_17087,N_16923,N_16902);
or U17088 (N_17088,N_16961,N_16822);
xnor U17089 (N_17089,N_16863,N_16803);
or U17090 (N_17090,N_16967,N_16883);
or U17091 (N_17091,N_16855,N_16864);
and U17092 (N_17092,N_16948,N_16890);
xnor U17093 (N_17093,N_16804,N_16836);
and U17094 (N_17094,N_16939,N_16996);
nand U17095 (N_17095,N_16852,N_16872);
and U17096 (N_17096,N_16841,N_16908);
nor U17097 (N_17097,N_16973,N_16994);
and U17098 (N_17098,N_16975,N_16922);
or U17099 (N_17099,N_16885,N_16844);
or U17100 (N_17100,N_16853,N_16975);
nand U17101 (N_17101,N_16833,N_16850);
and U17102 (N_17102,N_16906,N_16845);
nand U17103 (N_17103,N_16963,N_16984);
or U17104 (N_17104,N_16801,N_16889);
nor U17105 (N_17105,N_16884,N_16936);
nand U17106 (N_17106,N_16837,N_16939);
nand U17107 (N_17107,N_16801,N_16880);
or U17108 (N_17108,N_16904,N_16855);
xnor U17109 (N_17109,N_16801,N_16987);
and U17110 (N_17110,N_16874,N_16910);
nand U17111 (N_17111,N_16817,N_16821);
nand U17112 (N_17112,N_16858,N_16981);
nand U17113 (N_17113,N_16899,N_16944);
xor U17114 (N_17114,N_16831,N_16871);
or U17115 (N_17115,N_16819,N_16971);
xor U17116 (N_17116,N_16829,N_16987);
or U17117 (N_17117,N_16864,N_16860);
and U17118 (N_17118,N_16824,N_16877);
or U17119 (N_17119,N_16895,N_16851);
and U17120 (N_17120,N_16919,N_16829);
nand U17121 (N_17121,N_16852,N_16853);
or U17122 (N_17122,N_16920,N_16846);
or U17123 (N_17123,N_16906,N_16900);
and U17124 (N_17124,N_16923,N_16913);
and U17125 (N_17125,N_16837,N_16993);
and U17126 (N_17126,N_16871,N_16884);
xnor U17127 (N_17127,N_16841,N_16946);
or U17128 (N_17128,N_16828,N_16915);
or U17129 (N_17129,N_16997,N_16851);
or U17130 (N_17130,N_16812,N_16988);
or U17131 (N_17131,N_16923,N_16839);
xnor U17132 (N_17132,N_16833,N_16945);
xnor U17133 (N_17133,N_16865,N_16849);
xnor U17134 (N_17134,N_16849,N_16885);
xor U17135 (N_17135,N_16998,N_16922);
nand U17136 (N_17136,N_16800,N_16970);
xor U17137 (N_17137,N_16893,N_16940);
nor U17138 (N_17138,N_16812,N_16983);
and U17139 (N_17139,N_16979,N_16909);
xor U17140 (N_17140,N_16992,N_16825);
nand U17141 (N_17141,N_16831,N_16893);
nor U17142 (N_17142,N_16994,N_16828);
xor U17143 (N_17143,N_16801,N_16888);
and U17144 (N_17144,N_16946,N_16964);
nor U17145 (N_17145,N_16983,N_16824);
nor U17146 (N_17146,N_16938,N_16819);
nor U17147 (N_17147,N_16838,N_16875);
nor U17148 (N_17148,N_16943,N_16886);
xnor U17149 (N_17149,N_16946,N_16982);
nor U17150 (N_17150,N_16918,N_16871);
xnor U17151 (N_17151,N_16935,N_16827);
nor U17152 (N_17152,N_16868,N_16871);
or U17153 (N_17153,N_16994,N_16811);
and U17154 (N_17154,N_16943,N_16838);
and U17155 (N_17155,N_16828,N_16945);
or U17156 (N_17156,N_16862,N_16899);
nand U17157 (N_17157,N_16995,N_16897);
nand U17158 (N_17158,N_16855,N_16947);
nor U17159 (N_17159,N_16842,N_16807);
or U17160 (N_17160,N_16899,N_16907);
xor U17161 (N_17161,N_16858,N_16837);
and U17162 (N_17162,N_16870,N_16909);
and U17163 (N_17163,N_16902,N_16871);
xor U17164 (N_17164,N_16926,N_16821);
or U17165 (N_17165,N_16868,N_16985);
xnor U17166 (N_17166,N_16917,N_16830);
xnor U17167 (N_17167,N_16820,N_16875);
and U17168 (N_17168,N_16839,N_16883);
and U17169 (N_17169,N_16886,N_16833);
nand U17170 (N_17170,N_16966,N_16821);
nor U17171 (N_17171,N_16931,N_16842);
nand U17172 (N_17172,N_16821,N_16801);
and U17173 (N_17173,N_16899,N_16804);
xnor U17174 (N_17174,N_16874,N_16951);
nor U17175 (N_17175,N_16823,N_16961);
xnor U17176 (N_17176,N_16861,N_16962);
xnor U17177 (N_17177,N_16959,N_16967);
or U17178 (N_17178,N_16980,N_16847);
xor U17179 (N_17179,N_16882,N_16887);
nand U17180 (N_17180,N_16820,N_16889);
xor U17181 (N_17181,N_16862,N_16800);
nor U17182 (N_17182,N_16829,N_16883);
nor U17183 (N_17183,N_16918,N_16829);
and U17184 (N_17184,N_16898,N_16913);
nand U17185 (N_17185,N_16819,N_16916);
nor U17186 (N_17186,N_16912,N_16976);
nor U17187 (N_17187,N_16836,N_16814);
and U17188 (N_17188,N_16808,N_16893);
nand U17189 (N_17189,N_16848,N_16987);
and U17190 (N_17190,N_16813,N_16944);
nor U17191 (N_17191,N_16938,N_16979);
xor U17192 (N_17192,N_16991,N_16908);
or U17193 (N_17193,N_16811,N_16856);
nand U17194 (N_17194,N_16861,N_16990);
nor U17195 (N_17195,N_16835,N_16858);
and U17196 (N_17196,N_16847,N_16825);
and U17197 (N_17197,N_16873,N_16804);
xor U17198 (N_17198,N_16931,N_16856);
nand U17199 (N_17199,N_16966,N_16910);
nor U17200 (N_17200,N_17027,N_17093);
xor U17201 (N_17201,N_17006,N_17089);
or U17202 (N_17202,N_17132,N_17026);
nor U17203 (N_17203,N_17141,N_17036);
and U17204 (N_17204,N_17104,N_17011);
nand U17205 (N_17205,N_17168,N_17082);
and U17206 (N_17206,N_17126,N_17029);
nand U17207 (N_17207,N_17086,N_17019);
and U17208 (N_17208,N_17178,N_17025);
and U17209 (N_17209,N_17032,N_17102);
nor U17210 (N_17210,N_17066,N_17098);
nor U17211 (N_17211,N_17081,N_17007);
nand U17212 (N_17212,N_17047,N_17095);
nor U17213 (N_17213,N_17094,N_17055);
and U17214 (N_17214,N_17164,N_17101);
nand U17215 (N_17215,N_17062,N_17050);
and U17216 (N_17216,N_17107,N_17152);
and U17217 (N_17217,N_17021,N_17049);
nor U17218 (N_17218,N_17009,N_17175);
and U17219 (N_17219,N_17024,N_17059);
and U17220 (N_17220,N_17196,N_17124);
nor U17221 (N_17221,N_17070,N_17010);
xnor U17222 (N_17222,N_17184,N_17119);
nor U17223 (N_17223,N_17087,N_17060);
nand U17224 (N_17224,N_17197,N_17115);
or U17225 (N_17225,N_17003,N_17136);
and U17226 (N_17226,N_17022,N_17191);
nor U17227 (N_17227,N_17116,N_17143);
nand U17228 (N_17228,N_17150,N_17039);
xnor U17229 (N_17229,N_17088,N_17183);
and U17230 (N_17230,N_17016,N_17058);
and U17231 (N_17231,N_17048,N_17091);
xor U17232 (N_17232,N_17198,N_17075);
nor U17233 (N_17233,N_17065,N_17015);
nor U17234 (N_17234,N_17037,N_17077);
nor U17235 (N_17235,N_17166,N_17031);
nor U17236 (N_17236,N_17052,N_17071);
and U17237 (N_17237,N_17146,N_17138);
xnor U17238 (N_17238,N_17142,N_17108);
xor U17239 (N_17239,N_17100,N_17076);
and U17240 (N_17240,N_17174,N_17155);
or U17241 (N_17241,N_17160,N_17193);
nand U17242 (N_17242,N_17057,N_17148);
xor U17243 (N_17243,N_17000,N_17034);
nand U17244 (N_17244,N_17085,N_17192);
nand U17245 (N_17245,N_17035,N_17118);
xor U17246 (N_17246,N_17182,N_17061);
and U17247 (N_17247,N_17002,N_17188);
nor U17248 (N_17248,N_17144,N_17056);
or U17249 (N_17249,N_17195,N_17012);
nand U17250 (N_17250,N_17038,N_17109);
nor U17251 (N_17251,N_17171,N_17110);
and U17252 (N_17252,N_17131,N_17117);
or U17253 (N_17253,N_17004,N_17106);
nor U17254 (N_17254,N_17162,N_17063);
or U17255 (N_17255,N_17111,N_17170);
nor U17256 (N_17256,N_17185,N_17127);
and U17257 (N_17257,N_17134,N_17069);
or U17258 (N_17258,N_17033,N_17130);
or U17259 (N_17259,N_17123,N_17074);
nor U17260 (N_17260,N_17046,N_17092);
xor U17261 (N_17261,N_17054,N_17008);
and U17262 (N_17262,N_17041,N_17169);
xnor U17263 (N_17263,N_17137,N_17045);
xnor U17264 (N_17264,N_17157,N_17190);
nor U17265 (N_17265,N_17113,N_17112);
nand U17266 (N_17266,N_17140,N_17028);
xor U17267 (N_17267,N_17147,N_17149);
and U17268 (N_17268,N_17139,N_17001);
or U17269 (N_17269,N_17099,N_17125);
and U17270 (N_17270,N_17158,N_17153);
nor U17271 (N_17271,N_17189,N_17097);
nor U17272 (N_17272,N_17161,N_17173);
nor U17273 (N_17273,N_17163,N_17154);
and U17274 (N_17274,N_17179,N_17128);
nand U17275 (N_17275,N_17067,N_17051);
xnor U17276 (N_17276,N_17199,N_17105);
xnor U17277 (N_17277,N_17018,N_17151);
xnor U17278 (N_17278,N_17165,N_17096);
nor U17279 (N_17279,N_17042,N_17167);
xnor U17280 (N_17280,N_17156,N_17122);
nand U17281 (N_17281,N_17180,N_17176);
xor U17282 (N_17282,N_17043,N_17121);
and U17283 (N_17283,N_17133,N_17072);
nor U17284 (N_17284,N_17120,N_17053);
nand U17285 (N_17285,N_17083,N_17084);
xnor U17286 (N_17286,N_17040,N_17103);
nand U17287 (N_17287,N_17177,N_17090);
or U17288 (N_17288,N_17023,N_17020);
and U17289 (N_17289,N_17079,N_17044);
nor U17290 (N_17290,N_17145,N_17114);
and U17291 (N_17291,N_17080,N_17187);
xnor U17292 (N_17292,N_17017,N_17064);
xnor U17293 (N_17293,N_17030,N_17005);
or U17294 (N_17294,N_17014,N_17172);
and U17295 (N_17295,N_17194,N_17181);
nand U17296 (N_17296,N_17073,N_17186);
nand U17297 (N_17297,N_17159,N_17013);
nand U17298 (N_17298,N_17129,N_17078);
or U17299 (N_17299,N_17135,N_17068);
xnor U17300 (N_17300,N_17170,N_17086);
xnor U17301 (N_17301,N_17079,N_17166);
xnor U17302 (N_17302,N_17038,N_17037);
nand U17303 (N_17303,N_17104,N_17058);
nand U17304 (N_17304,N_17005,N_17154);
nor U17305 (N_17305,N_17138,N_17118);
nor U17306 (N_17306,N_17118,N_17088);
or U17307 (N_17307,N_17122,N_17100);
nand U17308 (N_17308,N_17116,N_17159);
and U17309 (N_17309,N_17045,N_17103);
xnor U17310 (N_17310,N_17100,N_17109);
nand U17311 (N_17311,N_17064,N_17058);
nand U17312 (N_17312,N_17079,N_17043);
nand U17313 (N_17313,N_17019,N_17080);
xor U17314 (N_17314,N_17135,N_17006);
nand U17315 (N_17315,N_17009,N_17123);
nor U17316 (N_17316,N_17073,N_17184);
nand U17317 (N_17317,N_17015,N_17188);
and U17318 (N_17318,N_17184,N_17037);
nand U17319 (N_17319,N_17116,N_17190);
nand U17320 (N_17320,N_17034,N_17105);
or U17321 (N_17321,N_17066,N_17156);
or U17322 (N_17322,N_17160,N_17050);
or U17323 (N_17323,N_17128,N_17091);
xor U17324 (N_17324,N_17070,N_17050);
xor U17325 (N_17325,N_17185,N_17054);
nor U17326 (N_17326,N_17033,N_17144);
and U17327 (N_17327,N_17110,N_17114);
or U17328 (N_17328,N_17045,N_17081);
or U17329 (N_17329,N_17072,N_17050);
nor U17330 (N_17330,N_17110,N_17038);
xnor U17331 (N_17331,N_17127,N_17081);
nand U17332 (N_17332,N_17068,N_17156);
xor U17333 (N_17333,N_17126,N_17132);
nor U17334 (N_17334,N_17186,N_17124);
or U17335 (N_17335,N_17154,N_17046);
nor U17336 (N_17336,N_17181,N_17000);
and U17337 (N_17337,N_17170,N_17177);
nand U17338 (N_17338,N_17184,N_17170);
xor U17339 (N_17339,N_17074,N_17141);
or U17340 (N_17340,N_17007,N_17172);
and U17341 (N_17341,N_17036,N_17035);
or U17342 (N_17342,N_17163,N_17085);
nand U17343 (N_17343,N_17132,N_17142);
or U17344 (N_17344,N_17072,N_17083);
nor U17345 (N_17345,N_17071,N_17177);
or U17346 (N_17346,N_17006,N_17194);
xnor U17347 (N_17347,N_17061,N_17080);
nand U17348 (N_17348,N_17126,N_17005);
nor U17349 (N_17349,N_17068,N_17095);
or U17350 (N_17350,N_17058,N_17131);
nor U17351 (N_17351,N_17105,N_17078);
nand U17352 (N_17352,N_17164,N_17087);
or U17353 (N_17353,N_17186,N_17034);
xnor U17354 (N_17354,N_17197,N_17112);
and U17355 (N_17355,N_17039,N_17189);
or U17356 (N_17356,N_17135,N_17196);
or U17357 (N_17357,N_17193,N_17188);
nand U17358 (N_17358,N_17141,N_17137);
and U17359 (N_17359,N_17155,N_17124);
nand U17360 (N_17360,N_17169,N_17121);
xnor U17361 (N_17361,N_17005,N_17182);
and U17362 (N_17362,N_17032,N_17178);
nor U17363 (N_17363,N_17097,N_17150);
nand U17364 (N_17364,N_17016,N_17149);
and U17365 (N_17365,N_17075,N_17080);
xnor U17366 (N_17366,N_17146,N_17190);
xnor U17367 (N_17367,N_17119,N_17139);
or U17368 (N_17368,N_17115,N_17134);
nor U17369 (N_17369,N_17064,N_17111);
xnor U17370 (N_17370,N_17013,N_17039);
nand U17371 (N_17371,N_17090,N_17074);
or U17372 (N_17372,N_17042,N_17017);
and U17373 (N_17373,N_17028,N_17148);
nor U17374 (N_17374,N_17037,N_17030);
nand U17375 (N_17375,N_17050,N_17059);
xor U17376 (N_17376,N_17123,N_17134);
nand U17377 (N_17377,N_17074,N_17146);
xnor U17378 (N_17378,N_17156,N_17144);
and U17379 (N_17379,N_17076,N_17008);
xnor U17380 (N_17380,N_17114,N_17057);
or U17381 (N_17381,N_17088,N_17110);
and U17382 (N_17382,N_17053,N_17127);
xnor U17383 (N_17383,N_17146,N_17010);
nor U17384 (N_17384,N_17074,N_17075);
xnor U17385 (N_17385,N_17008,N_17066);
and U17386 (N_17386,N_17062,N_17134);
nor U17387 (N_17387,N_17129,N_17146);
xor U17388 (N_17388,N_17080,N_17186);
nand U17389 (N_17389,N_17045,N_17113);
xnor U17390 (N_17390,N_17153,N_17093);
nor U17391 (N_17391,N_17092,N_17089);
nor U17392 (N_17392,N_17135,N_17162);
nand U17393 (N_17393,N_17105,N_17043);
nor U17394 (N_17394,N_17025,N_17090);
nand U17395 (N_17395,N_17193,N_17088);
xor U17396 (N_17396,N_17053,N_17006);
nor U17397 (N_17397,N_17087,N_17190);
xnor U17398 (N_17398,N_17072,N_17065);
nand U17399 (N_17399,N_17014,N_17190);
or U17400 (N_17400,N_17305,N_17282);
nand U17401 (N_17401,N_17243,N_17269);
xor U17402 (N_17402,N_17369,N_17289);
or U17403 (N_17403,N_17375,N_17261);
and U17404 (N_17404,N_17215,N_17275);
xor U17405 (N_17405,N_17217,N_17283);
or U17406 (N_17406,N_17249,N_17201);
nor U17407 (N_17407,N_17290,N_17300);
nor U17408 (N_17408,N_17214,N_17341);
xnor U17409 (N_17409,N_17237,N_17245);
nand U17410 (N_17410,N_17250,N_17228);
and U17411 (N_17411,N_17265,N_17385);
and U17412 (N_17412,N_17251,N_17203);
nand U17413 (N_17413,N_17239,N_17291);
nor U17414 (N_17414,N_17313,N_17252);
nand U17415 (N_17415,N_17364,N_17386);
and U17416 (N_17416,N_17200,N_17306);
nor U17417 (N_17417,N_17336,N_17370);
and U17418 (N_17418,N_17349,N_17363);
xnor U17419 (N_17419,N_17294,N_17389);
nor U17420 (N_17420,N_17351,N_17244);
xnor U17421 (N_17421,N_17267,N_17222);
nand U17422 (N_17422,N_17253,N_17212);
or U17423 (N_17423,N_17382,N_17246);
xnor U17424 (N_17424,N_17224,N_17235);
or U17425 (N_17425,N_17219,N_17395);
nand U17426 (N_17426,N_17333,N_17285);
xnor U17427 (N_17427,N_17338,N_17208);
or U17428 (N_17428,N_17205,N_17391);
nor U17429 (N_17429,N_17286,N_17209);
and U17430 (N_17430,N_17397,N_17334);
nand U17431 (N_17431,N_17392,N_17218);
nor U17432 (N_17432,N_17278,N_17276);
nor U17433 (N_17433,N_17358,N_17259);
and U17434 (N_17434,N_17279,N_17207);
xor U17435 (N_17435,N_17374,N_17347);
nand U17436 (N_17436,N_17309,N_17229);
nor U17437 (N_17437,N_17272,N_17284);
nor U17438 (N_17438,N_17398,N_17303);
xnor U17439 (N_17439,N_17264,N_17225);
nor U17440 (N_17440,N_17321,N_17383);
nor U17441 (N_17441,N_17213,N_17233);
xnor U17442 (N_17442,N_17371,N_17307);
nor U17443 (N_17443,N_17257,N_17262);
nor U17444 (N_17444,N_17339,N_17357);
nor U17445 (N_17445,N_17346,N_17316);
and U17446 (N_17446,N_17240,N_17377);
xor U17447 (N_17447,N_17221,N_17393);
nor U17448 (N_17448,N_17335,N_17308);
or U17449 (N_17449,N_17216,N_17356);
xor U17450 (N_17450,N_17337,N_17320);
and U17451 (N_17451,N_17361,N_17223);
or U17452 (N_17452,N_17211,N_17355);
xnor U17453 (N_17453,N_17248,N_17234);
and U17454 (N_17454,N_17328,N_17317);
nand U17455 (N_17455,N_17365,N_17232);
nor U17456 (N_17456,N_17372,N_17381);
or U17457 (N_17457,N_17315,N_17292);
and U17458 (N_17458,N_17254,N_17311);
nor U17459 (N_17459,N_17297,N_17255);
nand U17460 (N_17460,N_17323,N_17241);
nor U17461 (N_17461,N_17202,N_17345);
and U17462 (N_17462,N_17376,N_17399);
and U17463 (N_17463,N_17368,N_17280);
xor U17464 (N_17464,N_17390,N_17273);
nand U17465 (N_17465,N_17312,N_17206);
xnor U17466 (N_17466,N_17295,N_17324);
nor U17467 (N_17467,N_17299,N_17343);
and U17468 (N_17468,N_17367,N_17301);
and U17469 (N_17469,N_17352,N_17263);
nand U17470 (N_17470,N_17210,N_17379);
nand U17471 (N_17471,N_17258,N_17387);
nand U17472 (N_17472,N_17342,N_17304);
nor U17473 (N_17473,N_17236,N_17359);
xor U17474 (N_17474,N_17227,N_17353);
and U17475 (N_17475,N_17274,N_17326);
nand U17476 (N_17476,N_17281,N_17318);
nor U17477 (N_17477,N_17226,N_17230);
xor U17478 (N_17478,N_17287,N_17220);
xor U17479 (N_17479,N_17268,N_17350);
and U17480 (N_17480,N_17247,N_17322);
and U17481 (N_17481,N_17266,N_17354);
or U17482 (N_17482,N_17296,N_17298);
and U17483 (N_17483,N_17314,N_17231);
or U17484 (N_17484,N_17331,N_17348);
xor U17485 (N_17485,N_17242,N_17340);
or U17486 (N_17486,N_17293,N_17388);
nor U17487 (N_17487,N_17277,N_17360);
xor U17488 (N_17488,N_17256,N_17325);
and U17489 (N_17489,N_17302,N_17362);
xor U17490 (N_17490,N_17378,N_17384);
or U17491 (N_17491,N_17380,N_17330);
xnor U17492 (N_17492,N_17327,N_17204);
nor U17493 (N_17493,N_17332,N_17394);
or U17494 (N_17494,N_17271,N_17329);
nor U17495 (N_17495,N_17260,N_17310);
nor U17496 (N_17496,N_17344,N_17238);
and U17497 (N_17497,N_17396,N_17319);
xnor U17498 (N_17498,N_17270,N_17366);
or U17499 (N_17499,N_17288,N_17373);
and U17500 (N_17500,N_17278,N_17347);
xnor U17501 (N_17501,N_17235,N_17352);
or U17502 (N_17502,N_17247,N_17270);
nand U17503 (N_17503,N_17277,N_17256);
or U17504 (N_17504,N_17258,N_17266);
nor U17505 (N_17505,N_17259,N_17293);
and U17506 (N_17506,N_17285,N_17207);
xor U17507 (N_17507,N_17261,N_17241);
and U17508 (N_17508,N_17311,N_17226);
nand U17509 (N_17509,N_17253,N_17376);
or U17510 (N_17510,N_17234,N_17303);
or U17511 (N_17511,N_17306,N_17238);
nand U17512 (N_17512,N_17317,N_17216);
or U17513 (N_17513,N_17276,N_17257);
nor U17514 (N_17514,N_17218,N_17306);
nor U17515 (N_17515,N_17272,N_17362);
and U17516 (N_17516,N_17387,N_17281);
and U17517 (N_17517,N_17286,N_17324);
xor U17518 (N_17518,N_17337,N_17269);
nand U17519 (N_17519,N_17291,N_17283);
nand U17520 (N_17520,N_17249,N_17379);
and U17521 (N_17521,N_17397,N_17308);
nor U17522 (N_17522,N_17288,N_17338);
or U17523 (N_17523,N_17349,N_17229);
and U17524 (N_17524,N_17311,N_17333);
xor U17525 (N_17525,N_17296,N_17284);
or U17526 (N_17526,N_17235,N_17268);
or U17527 (N_17527,N_17320,N_17264);
xnor U17528 (N_17528,N_17214,N_17324);
xnor U17529 (N_17529,N_17331,N_17323);
or U17530 (N_17530,N_17285,N_17221);
and U17531 (N_17531,N_17386,N_17365);
xnor U17532 (N_17532,N_17275,N_17281);
nor U17533 (N_17533,N_17363,N_17269);
nand U17534 (N_17534,N_17220,N_17370);
and U17535 (N_17535,N_17301,N_17297);
nor U17536 (N_17536,N_17242,N_17253);
nand U17537 (N_17537,N_17284,N_17236);
xor U17538 (N_17538,N_17275,N_17345);
nand U17539 (N_17539,N_17308,N_17328);
or U17540 (N_17540,N_17342,N_17220);
nand U17541 (N_17541,N_17359,N_17345);
nand U17542 (N_17542,N_17363,N_17362);
nand U17543 (N_17543,N_17278,N_17358);
nor U17544 (N_17544,N_17248,N_17313);
and U17545 (N_17545,N_17240,N_17202);
and U17546 (N_17546,N_17210,N_17204);
nor U17547 (N_17547,N_17345,N_17233);
and U17548 (N_17548,N_17399,N_17395);
or U17549 (N_17549,N_17215,N_17367);
nand U17550 (N_17550,N_17312,N_17226);
or U17551 (N_17551,N_17221,N_17379);
and U17552 (N_17552,N_17262,N_17242);
xor U17553 (N_17553,N_17325,N_17218);
nand U17554 (N_17554,N_17206,N_17345);
and U17555 (N_17555,N_17263,N_17383);
xnor U17556 (N_17556,N_17259,N_17256);
or U17557 (N_17557,N_17219,N_17308);
and U17558 (N_17558,N_17349,N_17306);
and U17559 (N_17559,N_17257,N_17355);
nand U17560 (N_17560,N_17263,N_17353);
or U17561 (N_17561,N_17385,N_17368);
xor U17562 (N_17562,N_17383,N_17252);
or U17563 (N_17563,N_17374,N_17269);
and U17564 (N_17564,N_17337,N_17278);
xnor U17565 (N_17565,N_17271,N_17392);
nand U17566 (N_17566,N_17203,N_17219);
nor U17567 (N_17567,N_17330,N_17335);
xnor U17568 (N_17568,N_17354,N_17262);
nor U17569 (N_17569,N_17366,N_17375);
nand U17570 (N_17570,N_17308,N_17242);
or U17571 (N_17571,N_17348,N_17318);
and U17572 (N_17572,N_17316,N_17273);
and U17573 (N_17573,N_17213,N_17384);
nand U17574 (N_17574,N_17207,N_17257);
nor U17575 (N_17575,N_17330,N_17373);
xor U17576 (N_17576,N_17260,N_17371);
xor U17577 (N_17577,N_17382,N_17332);
nand U17578 (N_17578,N_17264,N_17393);
nor U17579 (N_17579,N_17260,N_17298);
xor U17580 (N_17580,N_17262,N_17259);
nor U17581 (N_17581,N_17299,N_17234);
nand U17582 (N_17582,N_17329,N_17236);
or U17583 (N_17583,N_17355,N_17206);
nor U17584 (N_17584,N_17341,N_17275);
xor U17585 (N_17585,N_17348,N_17363);
or U17586 (N_17586,N_17321,N_17282);
nor U17587 (N_17587,N_17243,N_17294);
xor U17588 (N_17588,N_17375,N_17341);
xor U17589 (N_17589,N_17251,N_17361);
nor U17590 (N_17590,N_17218,N_17286);
nand U17591 (N_17591,N_17312,N_17262);
xnor U17592 (N_17592,N_17286,N_17201);
and U17593 (N_17593,N_17256,N_17324);
or U17594 (N_17594,N_17208,N_17367);
xor U17595 (N_17595,N_17368,N_17348);
and U17596 (N_17596,N_17346,N_17264);
or U17597 (N_17597,N_17375,N_17328);
or U17598 (N_17598,N_17272,N_17255);
or U17599 (N_17599,N_17300,N_17306);
nand U17600 (N_17600,N_17504,N_17443);
and U17601 (N_17601,N_17440,N_17505);
or U17602 (N_17602,N_17531,N_17575);
nand U17603 (N_17603,N_17498,N_17435);
and U17604 (N_17604,N_17454,N_17516);
xor U17605 (N_17605,N_17553,N_17404);
and U17606 (N_17606,N_17476,N_17548);
and U17607 (N_17607,N_17500,N_17533);
or U17608 (N_17608,N_17570,N_17431);
xnor U17609 (N_17609,N_17563,N_17420);
or U17610 (N_17610,N_17410,N_17423);
nand U17611 (N_17611,N_17587,N_17477);
xnor U17612 (N_17612,N_17486,N_17450);
and U17613 (N_17613,N_17492,N_17406);
nor U17614 (N_17614,N_17532,N_17428);
or U17615 (N_17615,N_17453,N_17513);
nand U17616 (N_17616,N_17408,N_17503);
nor U17617 (N_17617,N_17529,N_17552);
xor U17618 (N_17618,N_17469,N_17528);
nand U17619 (N_17619,N_17530,N_17596);
nand U17620 (N_17620,N_17400,N_17535);
and U17621 (N_17621,N_17482,N_17433);
and U17622 (N_17622,N_17401,N_17554);
nor U17623 (N_17623,N_17422,N_17430);
or U17624 (N_17624,N_17475,N_17510);
nand U17625 (N_17625,N_17455,N_17542);
nor U17626 (N_17626,N_17460,N_17582);
and U17627 (N_17627,N_17429,N_17446);
and U17628 (N_17628,N_17470,N_17544);
nand U17629 (N_17629,N_17484,N_17508);
and U17630 (N_17630,N_17425,N_17466);
or U17631 (N_17631,N_17567,N_17525);
and U17632 (N_17632,N_17556,N_17471);
nor U17633 (N_17633,N_17547,N_17468);
or U17634 (N_17634,N_17562,N_17487);
or U17635 (N_17635,N_17561,N_17481);
nor U17636 (N_17636,N_17576,N_17541);
nor U17637 (N_17637,N_17434,N_17559);
or U17638 (N_17638,N_17478,N_17507);
and U17639 (N_17639,N_17540,N_17557);
or U17640 (N_17640,N_17413,N_17402);
nor U17641 (N_17641,N_17518,N_17591);
xor U17642 (N_17642,N_17412,N_17577);
xnor U17643 (N_17643,N_17493,N_17524);
and U17644 (N_17644,N_17467,N_17545);
or U17645 (N_17645,N_17491,N_17517);
nor U17646 (N_17646,N_17588,N_17439);
or U17647 (N_17647,N_17457,N_17480);
xor U17648 (N_17648,N_17580,N_17501);
nand U17649 (N_17649,N_17573,N_17586);
nor U17650 (N_17650,N_17441,N_17403);
nor U17651 (N_17651,N_17485,N_17526);
xor U17652 (N_17652,N_17496,N_17549);
or U17653 (N_17653,N_17437,N_17512);
or U17654 (N_17654,N_17527,N_17521);
or U17655 (N_17655,N_17495,N_17418);
and U17656 (N_17656,N_17565,N_17594);
xor U17657 (N_17657,N_17488,N_17432);
or U17658 (N_17658,N_17424,N_17449);
nor U17659 (N_17659,N_17519,N_17497);
nor U17660 (N_17660,N_17590,N_17574);
nand U17661 (N_17661,N_17566,N_17479);
nand U17662 (N_17662,N_17502,N_17593);
nand U17663 (N_17663,N_17555,N_17419);
or U17664 (N_17664,N_17564,N_17458);
and U17665 (N_17665,N_17595,N_17489);
nand U17666 (N_17666,N_17522,N_17427);
xor U17667 (N_17667,N_17536,N_17589);
nor U17668 (N_17668,N_17483,N_17599);
and U17669 (N_17669,N_17583,N_17474);
or U17670 (N_17670,N_17472,N_17451);
xnor U17671 (N_17671,N_17417,N_17514);
xnor U17672 (N_17672,N_17490,N_17523);
or U17673 (N_17673,N_17578,N_17592);
nand U17674 (N_17674,N_17585,N_17569);
nand U17675 (N_17675,N_17473,N_17494);
nor U17676 (N_17676,N_17598,N_17551);
and U17677 (N_17677,N_17456,N_17465);
or U17678 (N_17678,N_17405,N_17550);
nand U17679 (N_17679,N_17444,N_17442);
and U17680 (N_17680,N_17572,N_17414);
or U17681 (N_17681,N_17560,N_17436);
and U17682 (N_17682,N_17571,N_17459);
nand U17683 (N_17683,N_17515,N_17409);
nor U17684 (N_17684,N_17407,N_17506);
and U17685 (N_17685,N_17511,N_17537);
xnor U17686 (N_17686,N_17448,N_17539);
xor U17687 (N_17687,N_17426,N_17534);
xor U17688 (N_17688,N_17520,N_17581);
xnor U17689 (N_17689,N_17568,N_17461);
or U17690 (N_17690,N_17464,N_17463);
or U17691 (N_17691,N_17597,N_17415);
xnor U17692 (N_17692,N_17438,N_17462);
nor U17693 (N_17693,N_17416,N_17447);
nand U17694 (N_17694,N_17579,N_17499);
or U17695 (N_17695,N_17445,N_17538);
nand U17696 (N_17696,N_17546,N_17411);
nor U17697 (N_17697,N_17558,N_17543);
nand U17698 (N_17698,N_17421,N_17509);
and U17699 (N_17699,N_17452,N_17584);
and U17700 (N_17700,N_17443,N_17480);
nand U17701 (N_17701,N_17565,N_17578);
or U17702 (N_17702,N_17459,N_17559);
nand U17703 (N_17703,N_17598,N_17528);
or U17704 (N_17704,N_17503,N_17483);
nand U17705 (N_17705,N_17503,N_17405);
and U17706 (N_17706,N_17530,N_17511);
nand U17707 (N_17707,N_17471,N_17508);
and U17708 (N_17708,N_17536,N_17566);
nor U17709 (N_17709,N_17496,N_17461);
or U17710 (N_17710,N_17571,N_17512);
and U17711 (N_17711,N_17489,N_17497);
nand U17712 (N_17712,N_17506,N_17439);
xor U17713 (N_17713,N_17444,N_17443);
and U17714 (N_17714,N_17575,N_17511);
nand U17715 (N_17715,N_17480,N_17461);
and U17716 (N_17716,N_17562,N_17594);
or U17717 (N_17717,N_17529,N_17406);
xor U17718 (N_17718,N_17485,N_17563);
xor U17719 (N_17719,N_17477,N_17451);
xnor U17720 (N_17720,N_17481,N_17591);
or U17721 (N_17721,N_17436,N_17549);
nand U17722 (N_17722,N_17473,N_17532);
nand U17723 (N_17723,N_17439,N_17545);
nand U17724 (N_17724,N_17456,N_17542);
nor U17725 (N_17725,N_17566,N_17504);
xnor U17726 (N_17726,N_17579,N_17556);
xor U17727 (N_17727,N_17410,N_17499);
or U17728 (N_17728,N_17559,N_17413);
or U17729 (N_17729,N_17574,N_17579);
nor U17730 (N_17730,N_17476,N_17592);
and U17731 (N_17731,N_17488,N_17447);
nand U17732 (N_17732,N_17472,N_17440);
nand U17733 (N_17733,N_17428,N_17478);
and U17734 (N_17734,N_17439,N_17594);
and U17735 (N_17735,N_17416,N_17454);
xor U17736 (N_17736,N_17427,N_17433);
nand U17737 (N_17737,N_17528,N_17535);
nand U17738 (N_17738,N_17525,N_17592);
and U17739 (N_17739,N_17430,N_17562);
nor U17740 (N_17740,N_17444,N_17478);
and U17741 (N_17741,N_17573,N_17579);
nor U17742 (N_17742,N_17437,N_17522);
or U17743 (N_17743,N_17525,N_17442);
xnor U17744 (N_17744,N_17549,N_17597);
and U17745 (N_17745,N_17531,N_17597);
nand U17746 (N_17746,N_17576,N_17581);
nand U17747 (N_17747,N_17502,N_17511);
nand U17748 (N_17748,N_17574,N_17477);
xnor U17749 (N_17749,N_17541,N_17563);
nand U17750 (N_17750,N_17597,N_17412);
or U17751 (N_17751,N_17417,N_17460);
xor U17752 (N_17752,N_17594,N_17559);
nand U17753 (N_17753,N_17543,N_17410);
nand U17754 (N_17754,N_17550,N_17515);
or U17755 (N_17755,N_17552,N_17421);
or U17756 (N_17756,N_17501,N_17506);
or U17757 (N_17757,N_17596,N_17413);
xnor U17758 (N_17758,N_17588,N_17538);
or U17759 (N_17759,N_17419,N_17528);
and U17760 (N_17760,N_17534,N_17403);
xor U17761 (N_17761,N_17417,N_17539);
or U17762 (N_17762,N_17598,N_17440);
xor U17763 (N_17763,N_17432,N_17551);
nand U17764 (N_17764,N_17585,N_17469);
xor U17765 (N_17765,N_17519,N_17424);
and U17766 (N_17766,N_17494,N_17503);
and U17767 (N_17767,N_17460,N_17526);
or U17768 (N_17768,N_17444,N_17440);
nand U17769 (N_17769,N_17506,N_17563);
or U17770 (N_17770,N_17407,N_17481);
or U17771 (N_17771,N_17467,N_17481);
and U17772 (N_17772,N_17430,N_17594);
xnor U17773 (N_17773,N_17437,N_17480);
nand U17774 (N_17774,N_17449,N_17537);
nand U17775 (N_17775,N_17491,N_17530);
xor U17776 (N_17776,N_17595,N_17449);
nor U17777 (N_17777,N_17584,N_17448);
and U17778 (N_17778,N_17510,N_17569);
xnor U17779 (N_17779,N_17499,N_17434);
xor U17780 (N_17780,N_17433,N_17535);
nor U17781 (N_17781,N_17505,N_17584);
nand U17782 (N_17782,N_17565,N_17552);
nor U17783 (N_17783,N_17575,N_17425);
or U17784 (N_17784,N_17585,N_17526);
xor U17785 (N_17785,N_17411,N_17480);
and U17786 (N_17786,N_17591,N_17521);
or U17787 (N_17787,N_17437,N_17413);
and U17788 (N_17788,N_17402,N_17442);
or U17789 (N_17789,N_17419,N_17472);
xor U17790 (N_17790,N_17533,N_17454);
xnor U17791 (N_17791,N_17555,N_17563);
and U17792 (N_17792,N_17428,N_17514);
or U17793 (N_17793,N_17437,N_17521);
nor U17794 (N_17794,N_17500,N_17476);
xnor U17795 (N_17795,N_17534,N_17473);
and U17796 (N_17796,N_17434,N_17466);
or U17797 (N_17797,N_17437,N_17403);
nor U17798 (N_17798,N_17521,N_17552);
nand U17799 (N_17799,N_17522,N_17584);
or U17800 (N_17800,N_17601,N_17673);
or U17801 (N_17801,N_17710,N_17709);
and U17802 (N_17802,N_17787,N_17674);
nand U17803 (N_17803,N_17666,N_17613);
and U17804 (N_17804,N_17735,N_17694);
and U17805 (N_17805,N_17671,N_17720);
or U17806 (N_17806,N_17799,N_17762);
and U17807 (N_17807,N_17772,N_17707);
or U17808 (N_17808,N_17751,N_17771);
or U17809 (N_17809,N_17794,N_17629);
xnor U17810 (N_17810,N_17606,N_17616);
xnor U17811 (N_17811,N_17702,N_17656);
or U17812 (N_17812,N_17767,N_17756);
nor U17813 (N_17813,N_17734,N_17643);
nor U17814 (N_17814,N_17792,N_17786);
nor U17815 (N_17815,N_17649,N_17663);
nor U17816 (N_17816,N_17680,N_17660);
xor U17817 (N_17817,N_17714,N_17733);
or U17818 (N_17818,N_17638,N_17703);
xnor U17819 (N_17819,N_17778,N_17639);
nand U17820 (N_17820,N_17679,N_17727);
xor U17821 (N_17821,N_17798,N_17789);
nor U17822 (N_17822,N_17620,N_17698);
xor U17823 (N_17823,N_17741,N_17724);
nand U17824 (N_17824,N_17610,N_17737);
xnor U17825 (N_17825,N_17775,N_17717);
or U17826 (N_17826,N_17791,N_17659);
and U17827 (N_17827,N_17711,N_17745);
nor U17828 (N_17828,N_17614,N_17706);
and U17829 (N_17829,N_17774,N_17652);
or U17830 (N_17830,N_17642,N_17681);
nand U17831 (N_17831,N_17740,N_17777);
xor U17832 (N_17832,N_17640,N_17788);
and U17833 (N_17833,N_17701,N_17631);
or U17834 (N_17834,N_17688,N_17672);
xnor U17835 (N_17835,N_17764,N_17625);
or U17836 (N_17836,N_17618,N_17721);
nand U17837 (N_17837,N_17732,N_17723);
or U17838 (N_17838,N_17684,N_17634);
nand U17839 (N_17839,N_17646,N_17615);
nor U17840 (N_17840,N_17766,N_17667);
nor U17841 (N_17841,N_17622,N_17783);
nor U17842 (N_17842,N_17776,N_17604);
nand U17843 (N_17843,N_17655,N_17669);
nand U17844 (N_17844,N_17738,N_17651);
nand U17845 (N_17845,N_17728,N_17782);
and U17846 (N_17846,N_17708,N_17670);
and U17847 (N_17847,N_17687,N_17780);
xnor U17848 (N_17848,N_17695,N_17785);
and U17849 (N_17849,N_17657,N_17699);
or U17850 (N_17850,N_17790,N_17661);
and U17851 (N_17851,N_17715,N_17612);
xor U17852 (N_17852,N_17665,N_17630);
or U17853 (N_17853,N_17683,N_17760);
and U17854 (N_17854,N_17696,N_17609);
xnor U17855 (N_17855,N_17624,N_17752);
nand U17856 (N_17856,N_17689,N_17619);
nor U17857 (N_17857,N_17633,N_17758);
and U17858 (N_17858,N_17705,N_17763);
nor U17859 (N_17859,N_17682,N_17725);
nor U17860 (N_17860,N_17765,N_17685);
and U17861 (N_17861,N_17627,N_17749);
nand U17862 (N_17862,N_17731,N_17692);
or U17863 (N_17863,N_17668,N_17796);
nand U17864 (N_17864,N_17704,N_17754);
nor U17865 (N_17865,N_17693,N_17600);
nor U17866 (N_17866,N_17716,N_17626);
nand U17867 (N_17867,N_17755,N_17753);
and U17868 (N_17868,N_17781,N_17605);
nand U17869 (N_17869,N_17628,N_17722);
nand U17870 (N_17870,N_17748,N_17691);
xnor U17871 (N_17871,N_17797,N_17719);
nor U17872 (N_17872,N_17759,N_17784);
and U17873 (N_17873,N_17632,N_17743);
xor U17874 (N_17874,N_17718,N_17637);
and U17875 (N_17875,N_17726,N_17636);
nor U17876 (N_17876,N_17739,N_17761);
or U17877 (N_17877,N_17678,N_17769);
nand U17878 (N_17878,N_17650,N_17779);
and U17879 (N_17879,N_17700,N_17676);
nand U17880 (N_17880,N_17653,N_17675);
nor U17881 (N_17881,N_17742,N_17768);
nor U17882 (N_17882,N_17607,N_17602);
or U17883 (N_17883,N_17736,N_17603);
or U17884 (N_17884,N_17697,N_17729);
xnor U17885 (N_17885,N_17623,N_17647);
and U17886 (N_17886,N_17658,N_17744);
or U17887 (N_17887,N_17662,N_17712);
or U17888 (N_17888,N_17793,N_17730);
or U17889 (N_17889,N_17757,N_17621);
nand U17890 (N_17890,N_17690,N_17635);
nor U17891 (N_17891,N_17654,N_17713);
xnor U17892 (N_17892,N_17795,N_17747);
nand U17893 (N_17893,N_17750,N_17770);
and U17894 (N_17894,N_17645,N_17608);
and U17895 (N_17895,N_17641,N_17611);
nand U17896 (N_17896,N_17686,N_17648);
nor U17897 (N_17897,N_17746,N_17664);
nor U17898 (N_17898,N_17773,N_17644);
nor U17899 (N_17899,N_17617,N_17677);
or U17900 (N_17900,N_17707,N_17657);
or U17901 (N_17901,N_17762,N_17684);
and U17902 (N_17902,N_17666,N_17685);
nor U17903 (N_17903,N_17691,N_17736);
nor U17904 (N_17904,N_17605,N_17646);
and U17905 (N_17905,N_17609,N_17629);
and U17906 (N_17906,N_17678,N_17799);
xnor U17907 (N_17907,N_17682,N_17666);
or U17908 (N_17908,N_17646,N_17782);
or U17909 (N_17909,N_17626,N_17631);
and U17910 (N_17910,N_17609,N_17719);
xor U17911 (N_17911,N_17642,N_17631);
and U17912 (N_17912,N_17734,N_17784);
and U17913 (N_17913,N_17645,N_17609);
and U17914 (N_17914,N_17788,N_17711);
nand U17915 (N_17915,N_17643,N_17693);
nand U17916 (N_17916,N_17705,N_17647);
nor U17917 (N_17917,N_17642,N_17702);
and U17918 (N_17918,N_17744,N_17717);
or U17919 (N_17919,N_17760,N_17622);
or U17920 (N_17920,N_17785,N_17774);
and U17921 (N_17921,N_17632,N_17718);
and U17922 (N_17922,N_17755,N_17610);
nand U17923 (N_17923,N_17605,N_17743);
or U17924 (N_17924,N_17758,N_17683);
xnor U17925 (N_17925,N_17752,N_17758);
xor U17926 (N_17926,N_17786,N_17788);
nor U17927 (N_17927,N_17695,N_17628);
and U17928 (N_17928,N_17693,N_17777);
or U17929 (N_17929,N_17725,N_17754);
or U17930 (N_17930,N_17663,N_17725);
nand U17931 (N_17931,N_17659,N_17700);
and U17932 (N_17932,N_17685,N_17744);
and U17933 (N_17933,N_17794,N_17652);
nand U17934 (N_17934,N_17699,N_17780);
nor U17935 (N_17935,N_17655,N_17767);
or U17936 (N_17936,N_17621,N_17771);
nand U17937 (N_17937,N_17706,N_17719);
nor U17938 (N_17938,N_17692,N_17666);
and U17939 (N_17939,N_17769,N_17700);
nor U17940 (N_17940,N_17602,N_17780);
or U17941 (N_17941,N_17794,N_17724);
nor U17942 (N_17942,N_17784,N_17606);
and U17943 (N_17943,N_17644,N_17743);
and U17944 (N_17944,N_17736,N_17687);
nand U17945 (N_17945,N_17714,N_17741);
xnor U17946 (N_17946,N_17730,N_17608);
nor U17947 (N_17947,N_17793,N_17696);
and U17948 (N_17948,N_17624,N_17728);
xor U17949 (N_17949,N_17727,N_17709);
nor U17950 (N_17950,N_17651,N_17671);
nand U17951 (N_17951,N_17778,N_17793);
and U17952 (N_17952,N_17611,N_17723);
or U17953 (N_17953,N_17720,N_17618);
and U17954 (N_17954,N_17642,N_17727);
and U17955 (N_17955,N_17746,N_17769);
nand U17956 (N_17956,N_17701,N_17694);
xor U17957 (N_17957,N_17617,N_17661);
nand U17958 (N_17958,N_17608,N_17694);
xor U17959 (N_17959,N_17735,N_17684);
or U17960 (N_17960,N_17609,N_17637);
nand U17961 (N_17961,N_17686,N_17629);
nor U17962 (N_17962,N_17743,N_17694);
xnor U17963 (N_17963,N_17720,N_17707);
xor U17964 (N_17964,N_17787,N_17615);
xor U17965 (N_17965,N_17645,N_17721);
and U17966 (N_17966,N_17633,N_17745);
nor U17967 (N_17967,N_17637,N_17701);
xnor U17968 (N_17968,N_17759,N_17772);
xnor U17969 (N_17969,N_17664,N_17699);
or U17970 (N_17970,N_17754,N_17732);
nand U17971 (N_17971,N_17674,N_17642);
nor U17972 (N_17972,N_17698,N_17622);
nor U17973 (N_17973,N_17756,N_17723);
nor U17974 (N_17974,N_17780,N_17760);
nor U17975 (N_17975,N_17695,N_17625);
xnor U17976 (N_17976,N_17600,N_17797);
and U17977 (N_17977,N_17750,N_17626);
nor U17978 (N_17978,N_17711,N_17609);
and U17979 (N_17979,N_17602,N_17683);
nand U17980 (N_17980,N_17703,N_17721);
or U17981 (N_17981,N_17772,N_17740);
or U17982 (N_17982,N_17757,N_17636);
nor U17983 (N_17983,N_17618,N_17751);
nand U17984 (N_17984,N_17643,N_17611);
nor U17985 (N_17985,N_17606,N_17653);
nor U17986 (N_17986,N_17745,N_17701);
nor U17987 (N_17987,N_17691,N_17646);
nor U17988 (N_17988,N_17665,N_17614);
nand U17989 (N_17989,N_17709,N_17638);
xnor U17990 (N_17990,N_17697,N_17773);
xnor U17991 (N_17991,N_17704,N_17616);
xnor U17992 (N_17992,N_17712,N_17698);
or U17993 (N_17993,N_17698,N_17785);
or U17994 (N_17994,N_17778,N_17643);
nor U17995 (N_17995,N_17723,N_17629);
xnor U17996 (N_17996,N_17600,N_17646);
and U17997 (N_17997,N_17736,N_17651);
nor U17998 (N_17998,N_17684,N_17772);
nand U17999 (N_17999,N_17601,N_17738);
xor U18000 (N_18000,N_17888,N_17842);
and U18001 (N_18001,N_17977,N_17804);
or U18002 (N_18002,N_17844,N_17961);
and U18003 (N_18003,N_17958,N_17914);
xor U18004 (N_18004,N_17889,N_17987);
or U18005 (N_18005,N_17860,N_17922);
or U18006 (N_18006,N_17873,N_17821);
or U18007 (N_18007,N_17859,N_17965);
nand U18008 (N_18008,N_17926,N_17916);
nand U18009 (N_18009,N_17837,N_17923);
nor U18010 (N_18010,N_17852,N_17827);
nor U18011 (N_18011,N_17876,N_17855);
nand U18012 (N_18012,N_17910,N_17813);
nor U18013 (N_18013,N_17887,N_17880);
nand U18014 (N_18014,N_17935,N_17810);
xnor U18015 (N_18015,N_17823,N_17997);
xnor U18016 (N_18016,N_17815,N_17982);
xor U18017 (N_18017,N_17862,N_17963);
or U18018 (N_18018,N_17964,N_17816);
and U18019 (N_18019,N_17854,N_17847);
or U18020 (N_18020,N_17994,N_17996);
nand U18021 (N_18021,N_17901,N_17867);
and U18022 (N_18022,N_17956,N_17865);
and U18023 (N_18023,N_17918,N_17925);
and U18024 (N_18024,N_17834,N_17853);
nand U18025 (N_18025,N_17906,N_17843);
nor U18026 (N_18026,N_17917,N_17942);
xnor U18027 (N_18027,N_17838,N_17975);
and U18028 (N_18028,N_17990,N_17970);
and U18029 (N_18029,N_17902,N_17904);
and U18030 (N_18030,N_17828,N_17911);
nor U18031 (N_18031,N_17930,N_17851);
nand U18032 (N_18032,N_17920,N_17937);
and U18033 (N_18033,N_17919,N_17995);
or U18034 (N_18034,N_17875,N_17802);
nand U18035 (N_18035,N_17985,N_17869);
nand U18036 (N_18036,N_17900,N_17874);
nand U18037 (N_18037,N_17966,N_17915);
and U18038 (N_18038,N_17870,N_17962);
xor U18039 (N_18039,N_17836,N_17898);
xnor U18040 (N_18040,N_17814,N_17803);
nor U18041 (N_18041,N_17941,N_17992);
nand U18042 (N_18042,N_17973,N_17895);
or U18043 (N_18043,N_17864,N_17893);
nor U18044 (N_18044,N_17896,N_17885);
and U18045 (N_18045,N_17899,N_17955);
xnor U18046 (N_18046,N_17974,N_17801);
nor U18047 (N_18047,N_17981,N_17929);
and U18048 (N_18048,N_17856,N_17872);
or U18049 (N_18049,N_17831,N_17938);
or U18050 (N_18050,N_17909,N_17943);
nand U18051 (N_18051,N_17877,N_17811);
or U18052 (N_18052,N_17879,N_17806);
nand U18053 (N_18053,N_17863,N_17967);
nand U18054 (N_18054,N_17984,N_17945);
nor U18055 (N_18055,N_17905,N_17928);
nor U18056 (N_18056,N_17959,N_17969);
xor U18057 (N_18057,N_17934,N_17829);
xor U18058 (N_18058,N_17886,N_17932);
or U18059 (N_18059,N_17993,N_17971);
or U18060 (N_18060,N_17998,N_17857);
or U18061 (N_18061,N_17868,N_17809);
nor U18062 (N_18062,N_17991,N_17954);
and U18063 (N_18063,N_17936,N_17826);
or U18064 (N_18064,N_17949,N_17940);
nor U18065 (N_18065,N_17931,N_17912);
or U18066 (N_18066,N_17848,N_17908);
nor U18067 (N_18067,N_17927,N_17849);
xor U18068 (N_18068,N_17978,N_17946);
nand U18069 (N_18069,N_17881,N_17878);
xnor U18070 (N_18070,N_17824,N_17960);
xnor U18071 (N_18071,N_17825,N_17924);
nor U18072 (N_18072,N_17988,N_17953);
and U18073 (N_18073,N_17897,N_17957);
and U18074 (N_18074,N_17850,N_17832);
nand U18075 (N_18075,N_17819,N_17950);
nand U18076 (N_18076,N_17861,N_17818);
and U18077 (N_18077,N_17947,N_17808);
xor U18078 (N_18078,N_17907,N_17820);
nor U18079 (N_18079,N_17866,N_17817);
nand U18080 (N_18080,N_17979,N_17989);
nor U18081 (N_18081,N_17835,N_17841);
and U18082 (N_18082,N_17986,N_17840);
nor U18083 (N_18083,N_17976,N_17858);
or U18084 (N_18084,N_17805,N_17845);
xor U18085 (N_18085,N_17903,N_17921);
nand U18086 (N_18086,N_17972,N_17807);
nor U18087 (N_18087,N_17800,N_17871);
nand U18088 (N_18088,N_17822,N_17980);
nand U18089 (N_18089,N_17939,N_17882);
xor U18090 (N_18090,N_17952,N_17839);
nand U18091 (N_18091,N_17846,N_17951);
xnor U18092 (N_18092,N_17913,N_17891);
or U18093 (N_18093,N_17948,N_17944);
xor U18094 (N_18094,N_17890,N_17830);
xor U18095 (N_18095,N_17883,N_17999);
or U18096 (N_18096,N_17884,N_17968);
nand U18097 (N_18097,N_17894,N_17983);
nor U18098 (N_18098,N_17833,N_17933);
xor U18099 (N_18099,N_17812,N_17892);
or U18100 (N_18100,N_17848,N_17887);
nand U18101 (N_18101,N_17805,N_17967);
and U18102 (N_18102,N_17900,N_17977);
nor U18103 (N_18103,N_17927,N_17820);
or U18104 (N_18104,N_17893,N_17914);
xor U18105 (N_18105,N_17915,N_17815);
or U18106 (N_18106,N_17993,N_17912);
nor U18107 (N_18107,N_17896,N_17823);
xor U18108 (N_18108,N_17894,N_17866);
nand U18109 (N_18109,N_17905,N_17911);
or U18110 (N_18110,N_17831,N_17955);
nand U18111 (N_18111,N_17836,N_17811);
nor U18112 (N_18112,N_17969,N_17930);
and U18113 (N_18113,N_17928,N_17971);
nor U18114 (N_18114,N_17872,N_17982);
and U18115 (N_18115,N_17871,N_17997);
and U18116 (N_18116,N_17809,N_17941);
or U18117 (N_18117,N_17956,N_17875);
or U18118 (N_18118,N_17999,N_17853);
nand U18119 (N_18119,N_17856,N_17930);
or U18120 (N_18120,N_17984,N_17868);
xor U18121 (N_18121,N_17975,N_17817);
nand U18122 (N_18122,N_17913,N_17890);
and U18123 (N_18123,N_17914,N_17934);
nand U18124 (N_18124,N_17941,N_17813);
nand U18125 (N_18125,N_17832,N_17890);
or U18126 (N_18126,N_17996,N_17999);
xnor U18127 (N_18127,N_17903,N_17832);
xnor U18128 (N_18128,N_17829,N_17830);
and U18129 (N_18129,N_17975,N_17937);
or U18130 (N_18130,N_17888,N_17972);
nor U18131 (N_18131,N_17920,N_17860);
and U18132 (N_18132,N_17988,N_17836);
or U18133 (N_18133,N_17933,N_17992);
and U18134 (N_18134,N_17949,N_17848);
xor U18135 (N_18135,N_17899,N_17992);
nand U18136 (N_18136,N_17971,N_17819);
nor U18137 (N_18137,N_17807,N_17873);
or U18138 (N_18138,N_17935,N_17901);
nand U18139 (N_18139,N_17885,N_17996);
nor U18140 (N_18140,N_17958,N_17839);
nor U18141 (N_18141,N_17982,N_17892);
xnor U18142 (N_18142,N_17862,N_17933);
and U18143 (N_18143,N_17846,N_17991);
or U18144 (N_18144,N_17900,N_17983);
and U18145 (N_18145,N_17996,N_17923);
nor U18146 (N_18146,N_17910,N_17896);
xor U18147 (N_18147,N_17973,N_17832);
and U18148 (N_18148,N_17860,N_17818);
nor U18149 (N_18149,N_17887,N_17934);
xnor U18150 (N_18150,N_17908,N_17932);
nand U18151 (N_18151,N_17802,N_17821);
nand U18152 (N_18152,N_17901,N_17953);
or U18153 (N_18153,N_17969,N_17837);
xnor U18154 (N_18154,N_17926,N_17807);
or U18155 (N_18155,N_17914,N_17991);
nand U18156 (N_18156,N_17822,N_17962);
nor U18157 (N_18157,N_17983,N_17992);
nor U18158 (N_18158,N_17903,N_17886);
xor U18159 (N_18159,N_17905,N_17993);
and U18160 (N_18160,N_17839,N_17830);
xor U18161 (N_18161,N_17938,N_17950);
nand U18162 (N_18162,N_17957,N_17974);
nor U18163 (N_18163,N_17905,N_17830);
and U18164 (N_18164,N_17830,N_17901);
nor U18165 (N_18165,N_17801,N_17948);
and U18166 (N_18166,N_17982,N_17908);
or U18167 (N_18167,N_17912,N_17949);
or U18168 (N_18168,N_17848,N_17809);
xnor U18169 (N_18169,N_17934,N_17809);
and U18170 (N_18170,N_17819,N_17938);
and U18171 (N_18171,N_17982,N_17867);
and U18172 (N_18172,N_17923,N_17942);
and U18173 (N_18173,N_17953,N_17970);
nand U18174 (N_18174,N_17898,N_17975);
and U18175 (N_18175,N_17956,N_17992);
nor U18176 (N_18176,N_17869,N_17913);
nand U18177 (N_18177,N_17815,N_17970);
nand U18178 (N_18178,N_17902,N_17924);
or U18179 (N_18179,N_17983,N_17809);
nand U18180 (N_18180,N_17927,N_17901);
and U18181 (N_18181,N_17879,N_17813);
xor U18182 (N_18182,N_17989,N_17899);
nand U18183 (N_18183,N_17853,N_17862);
nand U18184 (N_18184,N_17901,N_17899);
xnor U18185 (N_18185,N_17946,N_17896);
nor U18186 (N_18186,N_17987,N_17849);
nand U18187 (N_18187,N_17978,N_17911);
and U18188 (N_18188,N_17825,N_17904);
or U18189 (N_18189,N_17850,N_17862);
nor U18190 (N_18190,N_17852,N_17960);
or U18191 (N_18191,N_17941,N_17868);
nor U18192 (N_18192,N_17890,N_17854);
nand U18193 (N_18193,N_17869,N_17975);
or U18194 (N_18194,N_17895,N_17893);
nand U18195 (N_18195,N_17803,N_17914);
nor U18196 (N_18196,N_17965,N_17805);
and U18197 (N_18197,N_17972,N_17929);
xor U18198 (N_18198,N_17994,N_17951);
xnor U18199 (N_18199,N_17911,N_17800);
xnor U18200 (N_18200,N_18034,N_18006);
or U18201 (N_18201,N_18184,N_18106);
or U18202 (N_18202,N_18031,N_18121);
or U18203 (N_18203,N_18064,N_18118);
nand U18204 (N_18204,N_18063,N_18197);
or U18205 (N_18205,N_18138,N_18093);
nand U18206 (N_18206,N_18182,N_18120);
or U18207 (N_18207,N_18147,N_18167);
xor U18208 (N_18208,N_18192,N_18042);
xnor U18209 (N_18209,N_18081,N_18011);
and U18210 (N_18210,N_18024,N_18040);
xor U18211 (N_18211,N_18170,N_18149);
xor U18212 (N_18212,N_18038,N_18073);
and U18213 (N_18213,N_18190,N_18001);
nand U18214 (N_18214,N_18126,N_18023);
nand U18215 (N_18215,N_18079,N_18015);
nand U18216 (N_18216,N_18030,N_18088);
nand U18217 (N_18217,N_18189,N_18092);
nand U18218 (N_18218,N_18020,N_18036);
nand U18219 (N_18219,N_18055,N_18198);
xnor U18220 (N_18220,N_18084,N_18179);
nor U18221 (N_18221,N_18112,N_18083);
and U18222 (N_18222,N_18123,N_18154);
xnor U18223 (N_18223,N_18012,N_18095);
xor U18224 (N_18224,N_18159,N_18098);
xnor U18225 (N_18225,N_18199,N_18109);
xnor U18226 (N_18226,N_18094,N_18003);
nor U18227 (N_18227,N_18186,N_18115);
nand U18228 (N_18228,N_18162,N_18168);
or U18229 (N_18229,N_18145,N_18061);
nand U18230 (N_18230,N_18177,N_18188);
or U18231 (N_18231,N_18049,N_18032);
or U18232 (N_18232,N_18193,N_18046);
nand U18233 (N_18233,N_18056,N_18181);
or U18234 (N_18234,N_18009,N_18130);
or U18235 (N_18235,N_18078,N_18157);
nor U18236 (N_18236,N_18074,N_18069);
nand U18237 (N_18237,N_18097,N_18103);
and U18238 (N_18238,N_18039,N_18060);
nor U18239 (N_18239,N_18171,N_18027);
and U18240 (N_18240,N_18143,N_18185);
or U18241 (N_18241,N_18110,N_18000);
and U18242 (N_18242,N_18122,N_18173);
xnor U18243 (N_18243,N_18137,N_18107);
nor U18244 (N_18244,N_18002,N_18178);
or U18245 (N_18245,N_18072,N_18071);
nand U18246 (N_18246,N_18175,N_18111);
nand U18247 (N_18247,N_18041,N_18017);
nand U18248 (N_18248,N_18057,N_18033);
or U18249 (N_18249,N_18028,N_18104);
or U18250 (N_18250,N_18007,N_18108);
nand U18251 (N_18251,N_18050,N_18187);
and U18252 (N_18252,N_18005,N_18144);
nand U18253 (N_18253,N_18051,N_18163);
and U18254 (N_18254,N_18116,N_18174);
xor U18255 (N_18255,N_18085,N_18180);
nand U18256 (N_18256,N_18066,N_18010);
nor U18257 (N_18257,N_18075,N_18004);
nor U18258 (N_18258,N_18129,N_18102);
nor U18259 (N_18259,N_18135,N_18166);
nor U18260 (N_18260,N_18052,N_18141);
or U18261 (N_18261,N_18195,N_18099);
nor U18262 (N_18262,N_18029,N_18068);
nor U18263 (N_18263,N_18043,N_18080);
nand U18264 (N_18264,N_18091,N_18044);
nand U18265 (N_18265,N_18113,N_18018);
nand U18266 (N_18266,N_18035,N_18059);
nand U18267 (N_18267,N_18152,N_18155);
nor U18268 (N_18268,N_18089,N_18128);
nand U18269 (N_18269,N_18082,N_18070);
and U18270 (N_18270,N_18158,N_18025);
or U18271 (N_18271,N_18100,N_18161);
or U18272 (N_18272,N_18191,N_18169);
and U18273 (N_18273,N_18148,N_18054);
xor U18274 (N_18274,N_18132,N_18134);
and U18275 (N_18275,N_18048,N_18140);
nor U18276 (N_18276,N_18150,N_18136);
nor U18277 (N_18277,N_18019,N_18176);
nor U18278 (N_18278,N_18172,N_18153);
nand U18279 (N_18279,N_18142,N_18067);
nand U18280 (N_18280,N_18062,N_18160);
or U18281 (N_18281,N_18183,N_18139);
or U18282 (N_18282,N_18096,N_18086);
nor U18283 (N_18283,N_18124,N_18058);
xor U18284 (N_18284,N_18013,N_18156);
or U18285 (N_18285,N_18008,N_18194);
and U18286 (N_18286,N_18133,N_18016);
nand U18287 (N_18287,N_18151,N_18114);
nand U18288 (N_18288,N_18196,N_18101);
or U18289 (N_18289,N_18077,N_18076);
nand U18290 (N_18290,N_18119,N_18021);
xor U18291 (N_18291,N_18065,N_18127);
xnor U18292 (N_18292,N_18146,N_18087);
xnor U18293 (N_18293,N_18131,N_18026);
or U18294 (N_18294,N_18053,N_18125);
and U18295 (N_18295,N_18014,N_18045);
xor U18296 (N_18296,N_18117,N_18164);
nand U18297 (N_18297,N_18037,N_18165);
nor U18298 (N_18298,N_18090,N_18022);
and U18299 (N_18299,N_18105,N_18047);
xor U18300 (N_18300,N_18139,N_18160);
or U18301 (N_18301,N_18063,N_18176);
nor U18302 (N_18302,N_18033,N_18124);
and U18303 (N_18303,N_18070,N_18116);
nor U18304 (N_18304,N_18191,N_18180);
nor U18305 (N_18305,N_18097,N_18161);
and U18306 (N_18306,N_18066,N_18053);
nor U18307 (N_18307,N_18160,N_18157);
nand U18308 (N_18308,N_18045,N_18142);
nand U18309 (N_18309,N_18089,N_18142);
and U18310 (N_18310,N_18093,N_18047);
xnor U18311 (N_18311,N_18077,N_18036);
xnor U18312 (N_18312,N_18059,N_18003);
and U18313 (N_18313,N_18019,N_18144);
and U18314 (N_18314,N_18065,N_18160);
xnor U18315 (N_18315,N_18113,N_18066);
xor U18316 (N_18316,N_18006,N_18004);
and U18317 (N_18317,N_18010,N_18181);
xnor U18318 (N_18318,N_18072,N_18125);
nand U18319 (N_18319,N_18129,N_18183);
and U18320 (N_18320,N_18050,N_18044);
nor U18321 (N_18321,N_18057,N_18024);
nand U18322 (N_18322,N_18198,N_18045);
xnor U18323 (N_18323,N_18161,N_18018);
and U18324 (N_18324,N_18158,N_18065);
and U18325 (N_18325,N_18112,N_18018);
or U18326 (N_18326,N_18088,N_18148);
nand U18327 (N_18327,N_18156,N_18047);
and U18328 (N_18328,N_18153,N_18116);
xor U18329 (N_18329,N_18068,N_18050);
and U18330 (N_18330,N_18048,N_18079);
nor U18331 (N_18331,N_18021,N_18185);
nand U18332 (N_18332,N_18102,N_18112);
nor U18333 (N_18333,N_18126,N_18028);
nor U18334 (N_18334,N_18061,N_18196);
xor U18335 (N_18335,N_18065,N_18121);
nand U18336 (N_18336,N_18138,N_18011);
xor U18337 (N_18337,N_18142,N_18131);
nor U18338 (N_18338,N_18141,N_18145);
nor U18339 (N_18339,N_18100,N_18084);
nor U18340 (N_18340,N_18031,N_18054);
nor U18341 (N_18341,N_18081,N_18046);
nor U18342 (N_18342,N_18030,N_18049);
nand U18343 (N_18343,N_18033,N_18178);
and U18344 (N_18344,N_18147,N_18068);
and U18345 (N_18345,N_18054,N_18176);
xnor U18346 (N_18346,N_18139,N_18185);
or U18347 (N_18347,N_18025,N_18193);
and U18348 (N_18348,N_18067,N_18166);
xor U18349 (N_18349,N_18151,N_18100);
nor U18350 (N_18350,N_18017,N_18172);
and U18351 (N_18351,N_18182,N_18165);
nor U18352 (N_18352,N_18143,N_18191);
and U18353 (N_18353,N_18165,N_18061);
and U18354 (N_18354,N_18192,N_18090);
xor U18355 (N_18355,N_18068,N_18055);
nor U18356 (N_18356,N_18087,N_18065);
xor U18357 (N_18357,N_18119,N_18129);
or U18358 (N_18358,N_18179,N_18061);
or U18359 (N_18359,N_18019,N_18179);
nand U18360 (N_18360,N_18160,N_18154);
xor U18361 (N_18361,N_18120,N_18070);
nand U18362 (N_18362,N_18196,N_18165);
and U18363 (N_18363,N_18086,N_18058);
xnor U18364 (N_18364,N_18123,N_18090);
nor U18365 (N_18365,N_18120,N_18160);
nor U18366 (N_18366,N_18128,N_18113);
nand U18367 (N_18367,N_18100,N_18042);
nor U18368 (N_18368,N_18061,N_18091);
nor U18369 (N_18369,N_18170,N_18162);
nor U18370 (N_18370,N_18178,N_18147);
nor U18371 (N_18371,N_18128,N_18119);
nand U18372 (N_18372,N_18079,N_18076);
or U18373 (N_18373,N_18182,N_18112);
or U18374 (N_18374,N_18186,N_18150);
and U18375 (N_18375,N_18131,N_18185);
nand U18376 (N_18376,N_18169,N_18074);
xnor U18377 (N_18377,N_18062,N_18197);
nor U18378 (N_18378,N_18036,N_18149);
xnor U18379 (N_18379,N_18157,N_18000);
nor U18380 (N_18380,N_18052,N_18177);
nand U18381 (N_18381,N_18106,N_18095);
xor U18382 (N_18382,N_18192,N_18107);
and U18383 (N_18383,N_18109,N_18118);
nand U18384 (N_18384,N_18079,N_18081);
nor U18385 (N_18385,N_18144,N_18197);
or U18386 (N_18386,N_18001,N_18156);
xnor U18387 (N_18387,N_18156,N_18183);
nand U18388 (N_18388,N_18022,N_18084);
nand U18389 (N_18389,N_18080,N_18085);
xnor U18390 (N_18390,N_18010,N_18041);
and U18391 (N_18391,N_18011,N_18194);
nor U18392 (N_18392,N_18051,N_18115);
nor U18393 (N_18393,N_18001,N_18021);
or U18394 (N_18394,N_18059,N_18160);
nor U18395 (N_18395,N_18039,N_18131);
and U18396 (N_18396,N_18155,N_18015);
nor U18397 (N_18397,N_18121,N_18150);
nor U18398 (N_18398,N_18176,N_18060);
and U18399 (N_18399,N_18141,N_18147);
nand U18400 (N_18400,N_18224,N_18337);
or U18401 (N_18401,N_18218,N_18212);
nand U18402 (N_18402,N_18361,N_18234);
nand U18403 (N_18403,N_18399,N_18334);
and U18404 (N_18404,N_18211,N_18228);
nor U18405 (N_18405,N_18217,N_18338);
nand U18406 (N_18406,N_18229,N_18281);
nand U18407 (N_18407,N_18305,N_18355);
or U18408 (N_18408,N_18372,N_18389);
or U18409 (N_18409,N_18230,N_18297);
nor U18410 (N_18410,N_18356,N_18306);
or U18411 (N_18411,N_18261,N_18317);
nand U18412 (N_18412,N_18286,N_18383);
xnor U18413 (N_18413,N_18360,N_18394);
nand U18414 (N_18414,N_18248,N_18381);
xor U18415 (N_18415,N_18263,N_18295);
nor U18416 (N_18416,N_18287,N_18298);
and U18417 (N_18417,N_18221,N_18235);
xor U18418 (N_18418,N_18324,N_18209);
xnor U18419 (N_18419,N_18260,N_18215);
xor U18420 (N_18420,N_18366,N_18315);
and U18421 (N_18421,N_18213,N_18344);
nand U18422 (N_18422,N_18284,N_18398);
nand U18423 (N_18423,N_18343,N_18253);
nor U18424 (N_18424,N_18240,N_18220);
xnor U18425 (N_18425,N_18377,N_18252);
or U18426 (N_18426,N_18369,N_18251);
nor U18427 (N_18427,N_18307,N_18247);
and U18428 (N_18428,N_18274,N_18237);
nand U18429 (N_18429,N_18242,N_18336);
nor U18430 (N_18430,N_18325,N_18200);
xor U18431 (N_18431,N_18280,N_18386);
nor U18432 (N_18432,N_18288,N_18373);
nand U18433 (N_18433,N_18300,N_18226);
and U18434 (N_18434,N_18339,N_18244);
and U18435 (N_18435,N_18367,N_18269);
nor U18436 (N_18436,N_18208,N_18362);
nor U18437 (N_18437,N_18340,N_18272);
and U18438 (N_18438,N_18351,N_18341);
xnor U18439 (N_18439,N_18259,N_18349);
nand U18440 (N_18440,N_18204,N_18246);
or U18441 (N_18441,N_18222,N_18318);
nor U18442 (N_18442,N_18276,N_18282);
nand U18443 (N_18443,N_18268,N_18301);
or U18444 (N_18444,N_18292,N_18258);
or U18445 (N_18445,N_18379,N_18283);
or U18446 (N_18446,N_18236,N_18231);
nor U18447 (N_18447,N_18267,N_18391);
xnor U18448 (N_18448,N_18254,N_18302);
and U18449 (N_18449,N_18358,N_18322);
xnor U18450 (N_18450,N_18327,N_18291);
or U18451 (N_18451,N_18352,N_18357);
nor U18452 (N_18452,N_18397,N_18368);
or U18453 (N_18453,N_18271,N_18347);
or U18454 (N_18454,N_18304,N_18365);
and U18455 (N_18455,N_18359,N_18203);
or U18456 (N_18456,N_18332,N_18314);
nand U18457 (N_18457,N_18225,N_18294);
nor U18458 (N_18458,N_18239,N_18308);
xor U18459 (N_18459,N_18323,N_18371);
and U18460 (N_18460,N_18321,N_18333);
or U18461 (N_18461,N_18227,N_18255);
nand U18462 (N_18462,N_18296,N_18364);
and U18463 (N_18463,N_18375,N_18266);
nor U18464 (N_18464,N_18264,N_18316);
nor U18465 (N_18465,N_18326,N_18243);
or U18466 (N_18466,N_18265,N_18390);
xnor U18467 (N_18467,N_18320,N_18313);
and U18468 (N_18468,N_18393,N_18384);
and U18469 (N_18469,N_18223,N_18273);
nor U18470 (N_18470,N_18380,N_18310);
nor U18471 (N_18471,N_18387,N_18328);
nor U18472 (N_18472,N_18278,N_18311);
or U18473 (N_18473,N_18202,N_18279);
or U18474 (N_18474,N_18275,N_18330);
or U18475 (N_18475,N_18385,N_18331);
nor U18476 (N_18476,N_18219,N_18256);
xnor U18477 (N_18477,N_18376,N_18289);
and U18478 (N_18478,N_18249,N_18363);
or U18479 (N_18479,N_18233,N_18395);
or U18480 (N_18480,N_18214,N_18335);
and U18481 (N_18481,N_18348,N_18319);
xor U18482 (N_18482,N_18290,N_18257);
nand U18483 (N_18483,N_18245,N_18396);
and U18484 (N_18484,N_18312,N_18378);
and U18485 (N_18485,N_18270,N_18382);
or U18486 (N_18486,N_18210,N_18354);
nand U18487 (N_18487,N_18353,N_18388);
xor U18488 (N_18488,N_18201,N_18342);
or U18489 (N_18489,N_18232,N_18303);
xnor U18490 (N_18490,N_18350,N_18285);
or U18491 (N_18491,N_18238,N_18241);
xor U18492 (N_18492,N_18293,N_18205);
nor U18493 (N_18493,N_18392,N_18374);
or U18494 (N_18494,N_18345,N_18250);
nor U18495 (N_18495,N_18309,N_18207);
nor U18496 (N_18496,N_18277,N_18370);
xor U18497 (N_18497,N_18216,N_18299);
xnor U18498 (N_18498,N_18346,N_18262);
and U18499 (N_18499,N_18206,N_18329);
nand U18500 (N_18500,N_18312,N_18371);
or U18501 (N_18501,N_18244,N_18288);
nand U18502 (N_18502,N_18235,N_18311);
xnor U18503 (N_18503,N_18268,N_18359);
nor U18504 (N_18504,N_18373,N_18374);
and U18505 (N_18505,N_18212,N_18309);
xnor U18506 (N_18506,N_18342,N_18355);
nor U18507 (N_18507,N_18349,N_18215);
nand U18508 (N_18508,N_18358,N_18338);
and U18509 (N_18509,N_18272,N_18244);
nand U18510 (N_18510,N_18235,N_18340);
or U18511 (N_18511,N_18228,N_18216);
nor U18512 (N_18512,N_18352,N_18334);
or U18513 (N_18513,N_18206,N_18341);
and U18514 (N_18514,N_18292,N_18373);
and U18515 (N_18515,N_18330,N_18373);
and U18516 (N_18516,N_18339,N_18302);
and U18517 (N_18517,N_18241,N_18240);
xnor U18518 (N_18518,N_18335,N_18262);
or U18519 (N_18519,N_18231,N_18302);
nor U18520 (N_18520,N_18234,N_18268);
nor U18521 (N_18521,N_18334,N_18268);
nor U18522 (N_18522,N_18324,N_18309);
and U18523 (N_18523,N_18372,N_18309);
or U18524 (N_18524,N_18391,N_18228);
nor U18525 (N_18525,N_18259,N_18292);
and U18526 (N_18526,N_18369,N_18224);
nand U18527 (N_18527,N_18366,N_18378);
or U18528 (N_18528,N_18327,N_18275);
or U18529 (N_18529,N_18346,N_18214);
xor U18530 (N_18530,N_18272,N_18265);
nor U18531 (N_18531,N_18255,N_18203);
nor U18532 (N_18532,N_18273,N_18316);
nand U18533 (N_18533,N_18218,N_18308);
or U18534 (N_18534,N_18305,N_18283);
or U18535 (N_18535,N_18301,N_18304);
or U18536 (N_18536,N_18358,N_18233);
nor U18537 (N_18537,N_18200,N_18365);
nor U18538 (N_18538,N_18300,N_18322);
nand U18539 (N_18539,N_18362,N_18339);
or U18540 (N_18540,N_18358,N_18364);
nor U18541 (N_18541,N_18351,N_18333);
nor U18542 (N_18542,N_18300,N_18302);
xor U18543 (N_18543,N_18313,N_18270);
nor U18544 (N_18544,N_18341,N_18273);
and U18545 (N_18545,N_18257,N_18233);
or U18546 (N_18546,N_18381,N_18391);
and U18547 (N_18547,N_18380,N_18224);
and U18548 (N_18548,N_18367,N_18310);
or U18549 (N_18549,N_18261,N_18324);
or U18550 (N_18550,N_18246,N_18366);
and U18551 (N_18551,N_18347,N_18285);
xnor U18552 (N_18552,N_18226,N_18282);
xnor U18553 (N_18553,N_18273,N_18219);
and U18554 (N_18554,N_18372,N_18294);
or U18555 (N_18555,N_18368,N_18398);
nand U18556 (N_18556,N_18249,N_18216);
and U18557 (N_18557,N_18337,N_18318);
nor U18558 (N_18558,N_18304,N_18354);
or U18559 (N_18559,N_18240,N_18274);
nand U18560 (N_18560,N_18327,N_18365);
nor U18561 (N_18561,N_18329,N_18280);
or U18562 (N_18562,N_18399,N_18245);
or U18563 (N_18563,N_18356,N_18393);
and U18564 (N_18564,N_18237,N_18259);
or U18565 (N_18565,N_18273,N_18321);
and U18566 (N_18566,N_18302,N_18217);
xnor U18567 (N_18567,N_18239,N_18232);
or U18568 (N_18568,N_18287,N_18328);
or U18569 (N_18569,N_18287,N_18300);
and U18570 (N_18570,N_18305,N_18252);
nor U18571 (N_18571,N_18351,N_18353);
and U18572 (N_18572,N_18319,N_18270);
nor U18573 (N_18573,N_18376,N_18320);
nor U18574 (N_18574,N_18208,N_18282);
and U18575 (N_18575,N_18311,N_18227);
and U18576 (N_18576,N_18321,N_18304);
xor U18577 (N_18577,N_18234,N_18226);
or U18578 (N_18578,N_18367,N_18240);
and U18579 (N_18579,N_18286,N_18396);
nand U18580 (N_18580,N_18218,N_18244);
or U18581 (N_18581,N_18338,N_18365);
nand U18582 (N_18582,N_18310,N_18307);
nand U18583 (N_18583,N_18355,N_18375);
nor U18584 (N_18584,N_18225,N_18333);
and U18585 (N_18585,N_18287,N_18299);
nor U18586 (N_18586,N_18269,N_18328);
nand U18587 (N_18587,N_18225,N_18275);
xnor U18588 (N_18588,N_18361,N_18280);
or U18589 (N_18589,N_18342,N_18281);
nor U18590 (N_18590,N_18318,N_18246);
or U18591 (N_18591,N_18353,N_18352);
nor U18592 (N_18592,N_18376,N_18335);
xnor U18593 (N_18593,N_18355,N_18311);
nand U18594 (N_18594,N_18299,N_18390);
or U18595 (N_18595,N_18369,N_18378);
nand U18596 (N_18596,N_18365,N_18283);
xor U18597 (N_18597,N_18284,N_18358);
xnor U18598 (N_18598,N_18262,N_18275);
or U18599 (N_18599,N_18354,N_18369);
and U18600 (N_18600,N_18515,N_18511);
and U18601 (N_18601,N_18541,N_18514);
nor U18602 (N_18602,N_18440,N_18404);
or U18603 (N_18603,N_18465,N_18599);
nor U18604 (N_18604,N_18510,N_18466);
nor U18605 (N_18605,N_18509,N_18459);
or U18606 (N_18606,N_18431,N_18411);
or U18607 (N_18607,N_18566,N_18526);
nor U18608 (N_18608,N_18598,N_18549);
and U18609 (N_18609,N_18450,N_18527);
nor U18610 (N_18610,N_18528,N_18568);
xnor U18611 (N_18611,N_18533,N_18556);
xnor U18612 (N_18612,N_18506,N_18453);
and U18613 (N_18613,N_18493,N_18488);
nor U18614 (N_18614,N_18524,N_18570);
or U18615 (N_18615,N_18460,N_18552);
nand U18616 (N_18616,N_18408,N_18430);
or U18617 (N_18617,N_18495,N_18490);
or U18618 (N_18618,N_18512,N_18428);
and U18619 (N_18619,N_18584,N_18562);
and U18620 (N_18620,N_18530,N_18559);
nand U18621 (N_18621,N_18560,N_18580);
or U18622 (N_18622,N_18574,N_18547);
or U18623 (N_18623,N_18548,N_18554);
xor U18624 (N_18624,N_18498,N_18497);
xnor U18625 (N_18625,N_18487,N_18481);
nor U18626 (N_18626,N_18436,N_18478);
nand U18627 (N_18627,N_18457,N_18414);
nor U18628 (N_18628,N_18448,N_18523);
or U18629 (N_18629,N_18519,N_18444);
and U18630 (N_18630,N_18421,N_18434);
nor U18631 (N_18631,N_18593,N_18545);
xor U18632 (N_18632,N_18518,N_18420);
nor U18633 (N_18633,N_18484,N_18485);
nor U18634 (N_18634,N_18412,N_18447);
and U18635 (N_18635,N_18443,N_18502);
nor U18636 (N_18636,N_18463,N_18532);
nor U18637 (N_18637,N_18476,N_18551);
nor U18638 (N_18638,N_18494,N_18482);
xnor U18639 (N_18639,N_18480,N_18516);
nor U18640 (N_18640,N_18501,N_18521);
xnor U18641 (N_18641,N_18537,N_18536);
nand U18642 (N_18642,N_18413,N_18429);
nor U18643 (N_18643,N_18462,N_18486);
and U18644 (N_18644,N_18433,N_18555);
nor U18645 (N_18645,N_18472,N_18455);
xnor U18646 (N_18646,N_18407,N_18458);
nor U18647 (N_18647,N_18517,N_18569);
or U18648 (N_18648,N_18410,N_18577);
and U18649 (N_18649,N_18461,N_18417);
nor U18650 (N_18650,N_18492,N_18597);
xor U18651 (N_18651,N_18534,N_18578);
nor U18652 (N_18652,N_18550,N_18452);
nand U18653 (N_18653,N_18469,N_18572);
nor U18654 (N_18654,N_18573,N_18543);
or U18655 (N_18655,N_18542,N_18539);
nand U18656 (N_18656,N_18418,N_18576);
nor U18657 (N_18657,N_18507,N_18451);
and U18658 (N_18658,N_18595,N_18424);
and U18659 (N_18659,N_18504,N_18535);
and U18660 (N_18660,N_18435,N_18403);
nand U18661 (N_18661,N_18508,N_18406);
or U18662 (N_18662,N_18416,N_18553);
and U18663 (N_18663,N_18477,N_18432);
or U18664 (N_18664,N_18499,N_18473);
and U18665 (N_18665,N_18425,N_18505);
or U18666 (N_18666,N_18474,N_18590);
and U18667 (N_18667,N_18591,N_18563);
and U18668 (N_18668,N_18564,N_18585);
nand U18669 (N_18669,N_18500,N_18520);
and U18670 (N_18670,N_18583,N_18571);
or U18671 (N_18671,N_18575,N_18422);
nor U18672 (N_18672,N_18437,N_18423);
nand U18673 (N_18673,N_18561,N_18445);
and U18674 (N_18674,N_18454,N_18582);
and U18675 (N_18675,N_18449,N_18479);
or U18676 (N_18676,N_18439,N_18471);
xor U18677 (N_18677,N_18557,N_18525);
nand U18678 (N_18678,N_18513,N_18538);
nor U18679 (N_18679,N_18446,N_18579);
and U18680 (N_18680,N_18415,N_18401);
nand U18681 (N_18681,N_18419,N_18409);
nor U18682 (N_18682,N_18558,N_18470);
nand U18683 (N_18683,N_18565,N_18491);
nor U18684 (N_18684,N_18456,N_18442);
nor U18685 (N_18685,N_18405,N_18475);
or U18686 (N_18686,N_18586,N_18483);
xnor U18687 (N_18687,N_18468,N_18438);
or U18688 (N_18688,N_18529,N_18503);
or U18689 (N_18689,N_18426,N_18587);
xnor U18690 (N_18690,N_18427,N_18592);
and U18691 (N_18691,N_18544,N_18588);
xnor U18692 (N_18692,N_18540,N_18589);
nand U18693 (N_18693,N_18496,N_18400);
and U18694 (N_18694,N_18489,N_18567);
nand U18695 (N_18695,N_18546,N_18581);
nand U18696 (N_18696,N_18531,N_18402);
and U18697 (N_18697,N_18594,N_18467);
xor U18698 (N_18698,N_18522,N_18441);
xor U18699 (N_18699,N_18464,N_18596);
or U18700 (N_18700,N_18543,N_18481);
or U18701 (N_18701,N_18534,N_18509);
and U18702 (N_18702,N_18457,N_18504);
nor U18703 (N_18703,N_18574,N_18465);
xor U18704 (N_18704,N_18584,N_18404);
and U18705 (N_18705,N_18441,N_18549);
and U18706 (N_18706,N_18472,N_18562);
nor U18707 (N_18707,N_18460,N_18448);
or U18708 (N_18708,N_18415,N_18419);
or U18709 (N_18709,N_18507,N_18567);
and U18710 (N_18710,N_18463,N_18550);
xnor U18711 (N_18711,N_18471,N_18416);
nand U18712 (N_18712,N_18431,N_18468);
and U18713 (N_18713,N_18442,N_18567);
and U18714 (N_18714,N_18598,N_18410);
and U18715 (N_18715,N_18590,N_18411);
or U18716 (N_18716,N_18400,N_18436);
and U18717 (N_18717,N_18478,N_18567);
nor U18718 (N_18718,N_18405,N_18573);
or U18719 (N_18719,N_18519,N_18515);
and U18720 (N_18720,N_18469,N_18495);
and U18721 (N_18721,N_18538,N_18595);
or U18722 (N_18722,N_18586,N_18414);
nor U18723 (N_18723,N_18559,N_18554);
and U18724 (N_18724,N_18434,N_18517);
nand U18725 (N_18725,N_18435,N_18486);
nor U18726 (N_18726,N_18590,N_18559);
and U18727 (N_18727,N_18510,N_18527);
and U18728 (N_18728,N_18549,N_18400);
and U18729 (N_18729,N_18506,N_18478);
nand U18730 (N_18730,N_18402,N_18572);
or U18731 (N_18731,N_18400,N_18562);
nand U18732 (N_18732,N_18419,N_18440);
nor U18733 (N_18733,N_18543,N_18476);
xnor U18734 (N_18734,N_18401,N_18535);
nand U18735 (N_18735,N_18404,N_18543);
xnor U18736 (N_18736,N_18575,N_18459);
or U18737 (N_18737,N_18514,N_18443);
xor U18738 (N_18738,N_18544,N_18566);
xor U18739 (N_18739,N_18453,N_18484);
nor U18740 (N_18740,N_18500,N_18472);
xor U18741 (N_18741,N_18515,N_18434);
and U18742 (N_18742,N_18474,N_18527);
and U18743 (N_18743,N_18401,N_18562);
nor U18744 (N_18744,N_18475,N_18538);
and U18745 (N_18745,N_18544,N_18496);
nor U18746 (N_18746,N_18407,N_18437);
and U18747 (N_18747,N_18547,N_18549);
and U18748 (N_18748,N_18498,N_18521);
and U18749 (N_18749,N_18422,N_18546);
and U18750 (N_18750,N_18474,N_18457);
or U18751 (N_18751,N_18466,N_18448);
or U18752 (N_18752,N_18430,N_18517);
and U18753 (N_18753,N_18526,N_18579);
nand U18754 (N_18754,N_18476,N_18550);
and U18755 (N_18755,N_18597,N_18477);
and U18756 (N_18756,N_18419,N_18479);
nor U18757 (N_18757,N_18496,N_18541);
xnor U18758 (N_18758,N_18534,N_18596);
nand U18759 (N_18759,N_18561,N_18471);
and U18760 (N_18760,N_18590,N_18444);
and U18761 (N_18761,N_18584,N_18588);
nand U18762 (N_18762,N_18462,N_18526);
nor U18763 (N_18763,N_18506,N_18415);
and U18764 (N_18764,N_18402,N_18466);
xor U18765 (N_18765,N_18584,N_18435);
xnor U18766 (N_18766,N_18424,N_18549);
and U18767 (N_18767,N_18437,N_18516);
or U18768 (N_18768,N_18579,N_18405);
nand U18769 (N_18769,N_18591,N_18557);
and U18770 (N_18770,N_18431,N_18562);
xnor U18771 (N_18771,N_18404,N_18476);
nand U18772 (N_18772,N_18503,N_18452);
and U18773 (N_18773,N_18585,N_18595);
xnor U18774 (N_18774,N_18434,N_18563);
xor U18775 (N_18775,N_18552,N_18473);
xnor U18776 (N_18776,N_18480,N_18409);
nor U18777 (N_18777,N_18420,N_18504);
nand U18778 (N_18778,N_18400,N_18401);
and U18779 (N_18779,N_18599,N_18448);
nor U18780 (N_18780,N_18580,N_18565);
and U18781 (N_18781,N_18473,N_18435);
or U18782 (N_18782,N_18480,N_18523);
or U18783 (N_18783,N_18511,N_18545);
and U18784 (N_18784,N_18546,N_18447);
and U18785 (N_18785,N_18488,N_18526);
nor U18786 (N_18786,N_18541,N_18580);
nor U18787 (N_18787,N_18590,N_18573);
nor U18788 (N_18788,N_18551,N_18576);
nand U18789 (N_18789,N_18571,N_18435);
nand U18790 (N_18790,N_18504,N_18407);
and U18791 (N_18791,N_18401,N_18567);
nand U18792 (N_18792,N_18473,N_18509);
or U18793 (N_18793,N_18543,N_18451);
nor U18794 (N_18794,N_18552,N_18541);
nor U18795 (N_18795,N_18584,N_18420);
or U18796 (N_18796,N_18581,N_18427);
xnor U18797 (N_18797,N_18565,N_18534);
or U18798 (N_18798,N_18581,N_18405);
or U18799 (N_18799,N_18517,N_18548);
or U18800 (N_18800,N_18626,N_18660);
nor U18801 (N_18801,N_18786,N_18606);
nor U18802 (N_18802,N_18664,N_18738);
nor U18803 (N_18803,N_18777,N_18735);
xor U18804 (N_18804,N_18655,N_18602);
and U18805 (N_18805,N_18618,N_18717);
nand U18806 (N_18806,N_18760,N_18677);
xnor U18807 (N_18807,N_18728,N_18720);
nand U18808 (N_18808,N_18670,N_18752);
or U18809 (N_18809,N_18736,N_18770);
and U18810 (N_18810,N_18653,N_18632);
nand U18811 (N_18811,N_18780,N_18721);
nand U18812 (N_18812,N_18713,N_18689);
nor U18813 (N_18813,N_18666,N_18766);
nor U18814 (N_18814,N_18610,N_18649);
xor U18815 (N_18815,N_18672,N_18723);
nor U18816 (N_18816,N_18758,N_18709);
or U18817 (N_18817,N_18669,N_18749);
nor U18818 (N_18818,N_18698,N_18731);
nor U18819 (N_18819,N_18774,N_18707);
and U18820 (N_18820,N_18771,N_18600);
nor U18821 (N_18821,N_18718,N_18768);
nor U18822 (N_18822,N_18747,N_18782);
or U18823 (N_18823,N_18743,N_18612);
xor U18824 (N_18824,N_18609,N_18787);
nand U18825 (N_18825,N_18737,N_18688);
and U18826 (N_18826,N_18622,N_18734);
xnor U18827 (N_18827,N_18702,N_18754);
or U18828 (N_18828,N_18776,N_18783);
nand U18829 (N_18829,N_18781,N_18654);
xor U18830 (N_18830,N_18633,N_18712);
or U18831 (N_18831,N_18668,N_18701);
nor U18832 (N_18832,N_18762,N_18607);
or U18833 (N_18833,N_18695,N_18682);
nand U18834 (N_18834,N_18708,N_18643);
nor U18835 (N_18835,N_18663,N_18603);
or U18836 (N_18836,N_18732,N_18710);
nand U18837 (N_18837,N_18646,N_18725);
nand U18838 (N_18838,N_18763,N_18733);
or U18839 (N_18839,N_18785,N_18638);
xor U18840 (N_18840,N_18745,N_18631);
nand U18841 (N_18841,N_18630,N_18648);
or U18842 (N_18842,N_18635,N_18623);
nor U18843 (N_18843,N_18687,N_18639);
and U18844 (N_18844,N_18793,N_18773);
nor U18845 (N_18845,N_18661,N_18613);
and U18846 (N_18846,N_18790,N_18704);
xor U18847 (N_18847,N_18797,N_18759);
nand U18848 (N_18848,N_18751,N_18756);
nor U18849 (N_18849,N_18685,N_18617);
and U18850 (N_18850,N_18719,N_18727);
or U18851 (N_18851,N_18699,N_18694);
nand U18852 (N_18852,N_18680,N_18791);
nand U18853 (N_18853,N_18659,N_18729);
nand U18854 (N_18854,N_18605,N_18650);
or U18855 (N_18855,N_18764,N_18616);
nand U18856 (N_18856,N_18799,N_18641);
and U18857 (N_18857,N_18604,N_18679);
nand U18858 (N_18858,N_18674,N_18693);
and U18859 (N_18859,N_18724,N_18611);
nor U18860 (N_18860,N_18757,N_18665);
and U18861 (N_18861,N_18697,N_18722);
nor U18862 (N_18862,N_18620,N_18628);
nor U18863 (N_18863,N_18765,N_18656);
and U18864 (N_18864,N_18714,N_18608);
and U18865 (N_18865,N_18742,N_18741);
xnor U18866 (N_18866,N_18715,N_18746);
nand U18867 (N_18867,N_18644,N_18750);
xor U18868 (N_18868,N_18696,N_18676);
xor U18869 (N_18869,N_18711,N_18645);
xor U18870 (N_18870,N_18657,N_18636);
nor U18871 (N_18871,N_18658,N_18634);
nor U18872 (N_18872,N_18784,N_18703);
nor U18873 (N_18873,N_18788,N_18671);
nand U18874 (N_18874,N_18625,N_18642);
and U18875 (N_18875,N_18629,N_18601);
nor U18876 (N_18876,N_18614,N_18651);
nand U18877 (N_18877,N_18647,N_18681);
and U18878 (N_18878,N_18767,N_18673);
or U18879 (N_18879,N_18686,N_18615);
nand U18880 (N_18880,N_18789,N_18692);
or U18881 (N_18881,N_18706,N_18678);
and U18882 (N_18882,N_18772,N_18691);
xnor U18883 (N_18883,N_18621,N_18624);
or U18884 (N_18884,N_18675,N_18740);
nand U18885 (N_18885,N_18796,N_18619);
xnor U18886 (N_18886,N_18690,N_18778);
and U18887 (N_18887,N_18652,N_18716);
nand U18888 (N_18888,N_18627,N_18640);
and U18889 (N_18889,N_18700,N_18744);
nand U18890 (N_18890,N_18753,N_18667);
and U18891 (N_18891,N_18662,N_18795);
nand U18892 (N_18892,N_18769,N_18792);
and U18893 (N_18893,N_18637,N_18755);
or U18894 (N_18894,N_18779,N_18775);
nand U18895 (N_18895,N_18683,N_18730);
nor U18896 (N_18896,N_18684,N_18739);
or U18897 (N_18897,N_18726,N_18798);
nand U18898 (N_18898,N_18705,N_18748);
nand U18899 (N_18899,N_18794,N_18761);
nand U18900 (N_18900,N_18631,N_18665);
nand U18901 (N_18901,N_18609,N_18613);
nand U18902 (N_18902,N_18710,N_18761);
and U18903 (N_18903,N_18694,N_18771);
and U18904 (N_18904,N_18605,N_18732);
nand U18905 (N_18905,N_18603,N_18630);
nor U18906 (N_18906,N_18639,N_18669);
nor U18907 (N_18907,N_18767,N_18741);
and U18908 (N_18908,N_18791,N_18635);
and U18909 (N_18909,N_18758,N_18694);
nor U18910 (N_18910,N_18698,N_18723);
nand U18911 (N_18911,N_18604,N_18683);
or U18912 (N_18912,N_18760,N_18695);
or U18913 (N_18913,N_18749,N_18647);
xor U18914 (N_18914,N_18711,N_18693);
nand U18915 (N_18915,N_18751,N_18626);
or U18916 (N_18916,N_18673,N_18675);
nand U18917 (N_18917,N_18647,N_18662);
and U18918 (N_18918,N_18680,N_18693);
xnor U18919 (N_18919,N_18689,N_18601);
or U18920 (N_18920,N_18765,N_18761);
and U18921 (N_18921,N_18790,N_18753);
and U18922 (N_18922,N_18696,N_18791);
xnor U18923 (N_18923,N_18705,N_18607);
nand U18924 (N_18924,N_18631,N_18741);
xnor U18925 (N_18925,N_18790,N_18777);
nor U18926 (N_18926,N_18774,N_18600);
xnor U18927 (N_18927,N_18631,N_18688);
or U18928 (N_18928,N_18628,N_18765);
or U18929 (N_18929,N_18790,N_18682);
or U18930 (N_18930,N_18736,N_18625);
nand U18931 (N_18931,N_18742,N_18722);
and U18932 (N_18932,N_18695,N_18601);
nor U18933 (N_18933,N_18633,N_18648);
and U18934 (N_18934,N_18694,N_18736);
or U18935 (N_18935,N_18725,N_18716);
nand U18936 (N_18936,N_18731,N_18794);
nand U18937 (N_18937,N_18765,N_18699);
nand U18938 (N_18938,N_18622,N_18778);
and U18939 (N_18939,N_18630,N_18650);
nor U18940 (N_18940,N_18696,N_18686);
or U18941 (N_18941,N_18752,N_18711);
nand U18942 (N_18942,N_18739,N_18776);
nor U18943 (N_18943,N_18759,N_18727);
and U18944 (N_18944,N_18763,N_18652);
and U18945 (N_18945,N_18798,N_18661);
and U18946 (N_18946,N_18733,N_18663);
xor U18947 (N_18947,N_18765,N_18727);
or U18948 (N_18948,N_18687,N_18740);
xnor U18949 (N_18949,N_18750,N_18702);
nand U18950 (N_18950,N_18656,N_18648);
xor U18951 (N_18951,N_18681,N_18744);
nor U18952 (N_18952,N_18798,N_18717);
and U18953 (N_18953,N_18673,N_18700);
nand U18954 (N_18954,N_18605,N_18615);
or U18955 (N_18955,N_18797,N_18722);
xor U18956 (N_18956,N_18669,N_18707);
nand U18957 (N_18957,N_18734,N_18763);
nor U18958 (N_18958,N_18778,N_18693);
nor U18959 (N_18959,N_18786,N_18735);
xor U18960 (N_18960,N_18741,N_18797);
and U18961 (N_18961,N_18722,N_18620);
xor U18962 (N_18962,N_18619,N_18780);
xor U18963 (N_18963,N_18702,N_18757);
nor U18964 (N_18964,N_18621,N_18780);
or U18965 (N_18965,N_18704,N_18751);
nor U18966 (N_18966,N_18680,N_18758);
nand U18967 (N_18967,N_18603,N_18696);
or U18968 (N_18968,N_18799,N_18694);
nand U18969 (N_18969,N_18612,N_18709);
or U18970 (N_18970,N_18758,N_18684);
nor U18971 (N_18971,N_18622,N_18762);
nor U18972 (N_18972,N_18745,N_18701);
or U18973 (N_18973,N_18770,N_18769);
nor U18974 (N_18974,N_18641,N_18676);
and U18975 (N_18975,N_18735,N_18673);
or U18976 (N_18976,N_18739,N_18644);
nor U18977 (N_18977,N_18739,N_18790);
nor U18978 (N_18978,N_18776,N_18622);
xor U18979 (N_18979,N_18701,N_18607);
nand U18980 (N_18980,N_18714,N_18670);
and U18981 (N_18981,N_18632,N_18668);
or U18982 (N_18982,N_18630,N_18608);
nor U18983 (N_18983,N_18771,N_18728);
nand U18984 (N_18984,N_18792,N_18699);
or U18985 (N_18985,N_18720,N_18661);
xor U18986 (N_18986,N_18725,N_18740);
or U18987 (N_18987,N_18614,N_18640);
nor U18988 (N_18988,N_18731,N_18678);
nand U18989 (N_18989,N_18670,N_18772);
or U18990 (N_18990,N_18710,N_18603);
or U18991 (N_18991,N_18613,N_18704);
nand U18992 (N_18992,N_18714,N_18678);
or U18993 (N_18993,N_18709,N_18745);
nand U18994 (N_18994,N_18676,N_18679);
xor U18995 (N_18995,N_18795,N_18645);
nand U18996 (N_18996,N_18721,N_18720);
or U18997 (N_18997,N_18758,N_18706);
or U18998 (N_18998,N_18682,N_18637);
nand U18999 (N_18999,N_18779,N_18752);
xnor U19000 (N_19000,N_18897,N_18952);
nand U19001 (N_19001,N_18929,N_18915);
or U19002 (N_19002,N_18866,N_18891);
nor U19003 (N_19003,N_18961,N_18923);
and U19004 (N_19004,N_18874,N_18872);
nor U19005 (N_19005,N_18855,N_18917);
and U19006 (N_19006,N_18948,N_18999);
or U19007 (N_19007,N_18856,N_18958);
nand U19008 (N_19008,N_18946,N_18975);
and U19009 (N_19009,N_18899,N_18937);
xor U19010 (N_19010,N_18962,N_18911);
and U19011 (N_19011,N_18936,N_18880);
and U19012 (N_19012,N_18841,N_18802);
nor U19013 (N_19013,N_18951,N_18983);
or U19014 (N_19014,N_18844,N_18851);
or U19015 (N_19015,N_18875,N_18808);
or U19016 (N_19016,N_18956,N_18819);
or U19017 (N_19017,N_18868,N_18995);
xor U19018 (N_19018,N_18974,N_18896);
nor U19019 (N_19019,N_18998,N_18867);
or U19020 (N_19020,N_18893,N_18969);
nand U19021 (N_19021,N_18817,N_18992);
nand U19022 (N_19022,N_18950,N_18980);
or U19023 (N_19023,N_18850,N_18846);
or U19024 (N_19024,N_18895,N_18824);
xnor U19025 (N_19025,N_18925,N_18943);
or U19026 (N_19026,N_18907,N_18979);
or U19027 (N_19027,N_18905,N_18906);
and U19028 (N_19028,N_18885,N_18833);
nand U19029 (N_19029,N_18942,N_18914);
nor U19030 (N_19030,N_18908,N_18892);
or U19031 (N_19031,N_18830,N_18881);
and U19032 (N_19032,N_18834,N_18949);
nor U19033 (N_19033,N_18888,N_18967);
xnor U19034 (N_19034,N_18918,N_18933);
and U19035 (N_19035,N_18800,N_18924);
nand U19036 (N_19036,N_18941,N_18903);
xnor U19037 (N_19037,N_18988,N_18993);
nor U19038 (N_19038,N_18807,N_18864);
xnor U19039 (N_19039,N_18938,N_18816);
xnor U19040 (N_19040,N_18978,N_18871);
xor U19041 (N_19041,N_18876,N_18947);
and U19042 (N_19042,N_18968,N_18883);
nand U19043 (N_19043,N_18828,N_18832);
xor U19044 (N_19044,N_18994,N_18822);
xnor U19045 (N_19045,N_18966,N_18965);
and U19046 (N_19046,N_18814,N_18970);
or U19047 (N_19047,N_18863,N_18858);
nor U19048 (N_19048,N_18835,N_18873);
nor U19049 (N_19049,N_18825,N_18870);
xnor U19050 (N_19050,N_18957,N_18955);
and U19051 (N_19051,N_18944,N_18811);
nor U19052 (N_19052,N_18919,N_18991);
or U19053 (N_19053,N_18857,N_18954);
nand U19054 (N_19054,N_18960,N_18823);
and U19055 (N_19055,N_18976,N_18826);
and U19056 (N_19056,N_18934,N_18890);
and U19057 (N_19057,N_18803,N_18909);
nor U19058 (N_19058,N_18886,N_18813);
nand U19059 (N_19059,N_18981,N_18989);
nor U19060 (N_19060,N_18940,N_18939);
and U19061 (N_19061,N_18820,N_18831);
and U19062 (N_19062,N_18913,N_18901);
nor U19063 (N_19063,N_18898,N_18838);
xnor U19064 (N_19064,N_18845,N_18852);
or U19065 (N_19065,N_18930,N_18862);
nor U19066 (N_19066,N_18806,N_18985);
nor U19067 (N_19067,N_18935,N_18926);
xnor U19068 (N_19068,N_18847,N_18910);
xnor U19069 (N_19069,N_18921,N_18996);
and U19070 (N_19070,N_18963,N_18837);
xnor U19071 (N_19071,N_18843,N_18805);
and U19072 (N_19072,N_18879,N_18882);
or U19073 (N_19073,N_18972,N_18931);
nor U19074 (N_19074,N_18912,N_18916);
nand U19075 (N_19075,N_18854,N_18928);
or U19076 (N_19076,N_18986,N_18927);
nor U19077 (N_19077,N_18877,N_18977);
nor U19078 (N_19078,N_18869,N_18971);
nor U19079 (N_19079,N_18964,N_18887);
or U19080 (N_19080,N_18904,N_18804);
or U19081 (N_19081,N_18953,N_18878);
nand U19082 (N_19082,N_18840,N_18829);
and U19083 (N_19083,N_18859,N_18990);
or U19084 (N_19084,N_18810,N_18815);
nand U19085 (N_19085,N_18884,N_18973);
or U19086 (N_19086,N_18959,N_18987);
xnor U19087 (N_19087,N_18801,N_18853);
xnor U19088 (N_19088,N_18902,N_18984);
nor U19089 (N_19089,N_18818,N_18922);
or U19090 (N_19090,N_18812,N_18821);
nor U19091 (N_19091,N_18920,N_18842);
nand U19092 (N_19092,N_18860,N_18932);
nand U19093 (N_19093,N_18836,N_18865);
nor U19094 (N_19094,N_18997,N_18839);
xor U19095 (N_19095,N_18982,N_18861);
xnor U19096 (N_19096,N_18848,N_18827);
nand U19097 (N_19097,N_18889,N_18894);
and U19098 (N_19098,N_18809,N_18900);
and U19099 (N_19099,N_18849,N_18945);
nor U19100 (N_19100,N_18823,N_18853);
and U19101 (N_19101,N_18913,N_18837);
or U19102 (N_19102,N_18946,N_18823);
and U19103 (N_19103,N_18869,N_18839);
or U19104 (N_19104,N_18920,N_18913);
or U19105 (N_19105,N_18878,N_18869);
nor U19106 (N_19106,N_18827,N_18821);
nand U19107 (N_19107,N_18942,N_18987);
and U19108 (N_19108,N_18945,N_18820);
and U19109 (N_19109,N_18971,N_18929);
and U19110 (N_19110,N_18986,N_18849);
nor U19111 (N_19111,N_18998,N_18816);
or U19112 (N_19112,N_18913,N_18845);
and U19113 (N_19113,N_18964,N_18990);
nand U19114 (N_19114,N_18978,N_18983);
xnor U19115 (N_19115,N_18922,N_18880);
and U19116 (N_19116,N_18831,N_18830);
or U19117 (N_19117,N_18802,N_18923);
nand U19118 (N_19118,N_18862,N_18803);
xnor U19119 (N_19119,N_18827,N_18979);
nand U19120 (N_19120,N_18913,N_18891);
or U19121 (N_19121,N_18987,N_18906);
nor U19122 (N_19122,N_18876,N_18945);
nor U19123 (N_19123,N_18923,N_18868);
nand U19124 (N_19124,N_18965,N_18808);
or U19125 (N_19125,N_18922,N_18928);
or U19126 (N_19126,N_18891,N_18955);
xnor U19127 (N_19127,N_18906,N_18982);
nor U19128 (N_19128,N_18841,N_18898);
nor U19129 (N_19129,N_18964,N_18832);
and U19130 (N_19130,N_18963,N_18961);
nor U19131 (N_19131,N_18831,N_18886);
nor U19132 (N_19132,N_18877,N_18924);
nor U19133 (N_19133,N_18934,N_18858);
or U19134 (N_19134,N_18832,N_18903);
and U19135 (N_19135,N_18992,N_18922);
and U19136 (N_19136,N_18851,N_18860);
xnor U19137 (N_19137,N_18889,N_18984);
nor U19138 (N_19138,N_18945,N_18934);
nand U19139 (N_19139,N_18945,N_18932);
and U19140 (N_19140,N_18890,N_18810);
nand U19141 (N_19141,N_18816,N_18942);
and U19142 (N_19142,N_18847,N_18960);
and U19143 (N_19143,N_18916,N_18904);
xor U19144 (N_19144,N_18861,N_18936);
and U19145 (N_19145,N_18853,N_18942);
nand U19146 (N_19146,N_18803,N_18934);
xnor U19147 (N_19147,N_18947,N_18828);
nand U19148 (N_19148,N_18839,N_18967);
and U19149 (N_19149,N_18923,N_18910);
and U19150 (N_19150,N_18894,N_18982);
and U19151 (N_19151,N_18850,N_18844);
or U19152 (N_19152,N_18823,N_18993);
nor U19153 (N_19153,N_18926,N_18996);
nor U19154 (N_19154,N_18835,N_18993);
and U19155 (N_19155,N_18814,N_18938);
nand U19156 (N_19156,N_18816,N_18827);
and U19157 (N_19157,N_18948,N_18841);
xor U19158 (N_19158,N_18953,N_18966);
and U19159 (N_19159,N_18860,N_18945);
or U19160 (N_19160,N_18963,N_18921);
and U19161 (N_19161,N_18989,N_18936);
or U19162 (N_19162,N_18828,N_18991);
and U19163 (N_19163,N_18979,N_18923);
xnor U19164 (N_19164,N_18970,N_18802);
nor U19165 (N_19165,N_18841,N_18812);
and U19166 (N_19166,N_18882,N_18967);
xnor U19167 (N_19167,N_18814,N_18939);
xor U19168 (N_19168,N_18985,N_18960);
nor U19169 (N_19169,N_18969,N_18866);
xor U19170 (N_19170,N_18858,N_18826);
or U19171 (N_19171,N_18894,N_18896);
or U19172 (N_19172,N_18900,N_18976);
or U19173 (N_19173,N_18817,N_18851);
xnor U19174 (N_19174,N_18863,N_18839);
nand U19175 (N_19175,N_18904,N_18855);
xnor U19176 (N_19176,N_18904,N_18865);
xnor U19177 (N_19177,N_18941,N_18884);
nor U19178 (N_19178,N_18935,N_18892);
and U19179 (N_19179,N_18841,N_18820);
nand U19180 (N_19180,N_18913,N_18826);
or U19181 (N_19181,N_18959,N_18932);
nor U19182 (N_19182,N_18823,N_18910);
or U19183 (N_19183,N_18853,N_18932);
or U19184 (N_19184,N_18922,N_18926);
nor U19185 (N_19185,N_18838,N_18964);
or U19186 (N_19186,N_18965,N_18941);
or U19187 (N_19187,N_18931,N_18806);
nand U19188 (N_19188,N_18868,N_18898);
or U19189 (N_19189,N_18880,N_18821);
xnor U19190 (N_19190,N_18824,N_18836);
nand U19191 (N_19191,N_18995,N_18959);
xnor U19192 (N_19192,N_18979,N_18848);
and U19193 (N_19193,N_18944,N_18815);
and U19194 (N_19194,N_18984,N_18849);
nand U19195 (N_19195,N_18839,N_18809);
nand U19196 (N_19196,N_18984,N_18872);
nor U19197 (N_19197,N_18914,N_18991);
xor U19198 (N_19198,N_18805,N_18981);
xor U19199 (N_19199,N_18833,N_18964);
xnor U19200 (N_19200,N_19149,N_19138);
xor U19201 (N_19201,N_19111,N_19093);
and U19202 (N_19202,N_19192,N_19044);
nand U19203 (N_19203,N_19074,N_19167);
or U19204 (N_19204,N_19026,N_19053);
nand U19205 (N_19205,N_19136,N_19190);
or U19206 (N_19206,N_19112,N_19091);
xnor U19207 (N_19207,N_19067,N_19052);
and U19208 (N_19208,N_19147,N_19145);
xnor U19209 (N_19209,N_19049,N_19008);
nand U19210 (N_19210,N_19163,N_19082);
nand U19211 (N_19211,N_19064,N_19195);
or U19212 (N_19212,N_19103,N_19141);
nand U19213 (N_19213,N_19126,N_19086);
and U19214 (N_19214,N_19010,N_19023);
xnor U19215 (N_19215,N_19135,N_19000);
nand U19216 (N_19216,N_19160,N_19140);
xnor U19217 (N_19217,N_19031,N_19179);
and U19218 (N_19218,N_19172,N_19133);
or U19219 (N_19219,N_19063,N_19131);
and U19220 (N_19220,N_19094,N_19099);
and U19221 (N_19221,N_19118,N_19065);
and U19222 (N_19222,N_19050,N_19100);
nor U19223 (N_19223,N_19150,N_19077);
and U19224 (N_19224,N_19005,N_19117);
or U19225 (N_19225,N_19041,N_19196);
nand U19226 (N_19226,N_19075,N_19011);
or U19227 (N_19227,N_19051,N_19114);
or U19228 (N_19228,N_19018,N_19030);
nand U19229 (N_19229,N_19182,N_19102);
nor U19230 (N_19230,N_19106,N_19088);
nor U19231 (N_19231,N_19061,N_19153);
nor U19232 (N_19232,N_19076,N_19174);
nand U19233 (N_19233,N_19056,N_19062);
xnor U19234 (N_19234,N_19137,N_19134);
xnor U19235 (N_19235,N_19024,N_19171);
nand U19236 (N_19236,N_19142,N_19119);
or U19237 (N_19237,N_19027,N_19020);
xnor U19238 (N_19238,N_19156,N_19016);
nand U19239 (N_19239,N_19007,N_19198);
and U19240 (N_19240,N_19072,N_19068);
or U19241 (N_19241,N_19097,N_19038);
nor U19242 (N_19242,N_19183,N_19101);
or U19243 (N_19243,N_19170,N_19006);
nand U19244 (N_19244,N_19154,N_19022);
nand U19245 (N_19245,N_19021,N_19177);
or U19246 (N_19246,N_19098,N_19158);
nor U19247 (N_19247,N_19148,N_19151);
xnor U19248 (N_19248,N_19019,N_19178);
or U19249 (N_19249,N_19002,N_19092);
xnor U19250 (N_19250,N_19081,N_19071);
and U19251 (N_19251,N_19087,N_19042);
and U19252 (N_19252,N_19104,N_19194);
and U19253 (N_19253,N_19073,N_19189);
nand U19254 (N_19254,N_19169,N_19125);
or U19255 (N_19255,N_19034,N_19084);
nor U19256 (N_19256,N_19162,N_19128);
nor U19257 (N_19257,N_19124,N_19109);
nand U19258 (N_19258,N_19017,N_19180);
or U19259 (N_19259,N_19043,N_19079);
nand U19260 (N_19260,N_19040,N_19029);
or U19261 (N_19261,N_19009,N_19089);
xnor U19262 (N_19262,N_19161,N_19059);
or U19263 (N_19263,N_19120,N_19047);
xor U19264 (N_19264,N_19176,N_19152);
or U19265 (N_19265,N_19045,N_19181);
nand U19266 (N_19266,N_19013,N_19123);
xnor U19267 (N_19267,N_19083,N_19085);
nor U19268 (N_19268,N_19036,N_19070);
or U19269 (N_19269,N_19054,N_19115);
xnor U19270 (N_19270,N_19035,N_19129);
and U19271 (N_19271,N_19080,N_19069);
nor U19272 (N_19272,N_19055,N_19095);
xnor U19273 (N_19273,N_19004,N_19165);
or U19274 (N_19274,N_19107,N_19188);
nand U19275 (N_19275,N_19025,N_19146);
or U19276 (N_19276,N_19173,N_19057);
or U19277 (N_19277,N_19139,N_19130);
xor U19278 (N_19278,N_19168,N_19159);
xnor U19279 (N_19279,N_19186,N_19132);
xnor U19280 (N_19280,N_19037,N_19060);
nor U19281 (N_19281,N_19012,N_19033);
and U19282 (N_19282,N_19127,N_19184);
and U19283 (N_19283,N_19185,N_19121);
and U19284 (N_19284,N_19032,N_19122);
nor U19285 (N_19285,N_19155,N_19014);
xor U19286 (N_19286,N_19046,N_19113);
nand U19287 (N_19287,N_19096,N_19157);
or U19288 (N_19288,N_19175,N_19193);
nand U19289 (N_19289,N_19144,N_19058);
or U19290 (N_19290,N_19048,N_19143);
and U19291 (N_19291,N_19110,N_19066);
nor U19292 (N_19292,N_19003,N_19108);
or U19293 (N_19293,N_19039,N_19001);
nand U19294 (N_19294,N_19105,N_19199);
and U19295 (N_19295,N_19028,N_19187);
nand U19296 (N_19296,N_19197,N_19015);
nand U19297 (N_19297,N_19191,N_19164);
nand U19298 (N_19298,N_19090,N_19078);
xnor U19299 (N_19299,N_19166,N_19116);
xor U19300 (N_19300,N_19199,N_19075);
and U19301 (N_19301,N_19158,N_19060);
nand U19302 (N_19302,N_19128,N_19158);
nor U19303 (N_19303,N_19148,N_19025);
nand U19304 (N_19304,N_19028,N_19124);
xnor U19305 (N_19305,N_19189,N_19009);
xor U19306 (N_19306,N_19024,N_19157);
or U19307 (N_19307,N_19163,N_19119);
xor U19308 (N_19308,N_19100,N_19068);
nand U19309 (N_19309,N_19067,N_19012);
nor U19310 (N_19310,N_19027,N_19025);
or U19311 (N_19311,N_19195,N_19140);
or U19312 (N_19312,N_19167,N_19191);
nand U19313 (N_19313,N_19156,N_19180);
or U19314 (N_19314,N_19099,N_19181);
nand U19315 (N_19315,N_19099,N_19132);
nand U19316 (N_19316,N_19047,N_19138);
nand U19317 (N_19317,N_19118,N_19052);
nand U19318 (N_19318,N_19027,N_19112);
and U19319 (N_19319,N_19045,N_19113);
and U19320 (N_19320,N_19182,N_19173);
xnor U19321 (N_19321,N_19122,N_19104);
xnor U19322 (N_19322,N_19035,N_19065);
xnor U19323 (N_19323,N_19029,N_19060);
and U19324 (N_19324,N_19199,N_19018);
nor U19325 (N_19325,N_19042,N_19117);
and U19326 (N_19326,N_19153,N_19137);
and U19327 (N_19327,N_19162,N_19028);
nor U19328 (N_19328,N_19150,N_19055);
or U19329 (N_19329,N_19073,N_19078);
xnor U19330 (N_19330,N_19162,N_19030);
nand U19331 (N_19331,N_19195,N_19198);
xor U19332 (N_19332,N_19015,N_19107);
xor U19333 (N_19333,N_19053,N_19180);
nor U19334 (N_19334,N_19045,N_19130);
and U19335 (N_19335,N_19183,N_19142);
nor U19336 (N_19336,N_19045,N_19193);
and U19337 (N_19337,N_19133,N_19007);
or U19338 (N_19338,N_19141,N_19172);
or U19339 (N_19339,N_19175,N_19147);
and U19340 (N_19340,N_19163,N_19045);
or U19341 (N_19341,N_19172,N_19012);
nand U19342 (N_19342,N_19165,N_19023);
xnor U19343 (N_19343,N_19134,N_19126);
or U19344 (N_19344,N_19193,N_19127);
nand U19345 (N_19345,N_19008,N_19016);
nor U19346 (N_19346,N_19037,N_19042);
or U19347 (N_19347,N_19001,N_19174);
xnor U19348 (N_19348,N_19101,N_19025);
and U19349 (N_19349,N_19037,N_19077);
nand U19350 (N_19350,N_19043,N_19078);
and U19351 (N_19351,N_19072,N_19165);
nand U19352 (N_19352,N_19130,N_19055);
or U19353 (N_19353,N_19160,N_19017);
and U19354 (N_19354,N_19031,N_19191);
nor U19355 (N_19355,N_19111,N_19008);
or U19356 (N_19356,N_19150,N_19070);
nor U19357 (N_19357,N_19175,N_19011);
nand U19358 (N_19358,N_19022,N_19158);
or U19359 (N_19359,N_19026,N_19093);
nand U19360 (N_19360,N_19113,N_19020);
nand U19361 (N_19361,N_19157,N_19090);
and U19362 (N_19362,N_19070,N_19161);
nor U19363 (N_19363,N_19048,N_19070);
nor U19364 (N_19364,N_19095,N_19065);
and U19365 (N_19365,N_19037,N_19041);
nand U19366 (N_19366,N_19069,N_19099);
nor U19367 (N_19367,N_19075,N_19137);
xnor U19368 (N_19368,N_19014,N_19183);
and U19369 (N_19369,N_19179,N_19078);
or U19370 (N_19370,N_19056,N_19161);
xnor U19371 (N_19371,N_19119,N_19184);
and U19372 (N_19372,N_19001,N_19051);
nand U19373 (N_19373,N_19166,N_19157);
nor U19374 (N_19374,N_19012,N_19095);
nand U19375 (N_19375,N_19099,N_19139);
nor U19376 (N_19376,N_19006,N_19103);
and U19377 (N_19377,N_19159,N_19187);
and U19378 (N_19378,N_19158,N_19091);
and U19379 (N_19379,N_19133,N_19019);
nand U19380 (N_19380,N_19138,N_19069);
nand U19381 (N_19381,N_19107,N_19140);
xor U19382 (N_19382,N_19019,N_19010);
or U19383 (N_19383,N_19106,N_19109);
or U19384 (N_19384,N_19090,N_19102);
nor U19385 (N_19385,N_19112,N_19164);
and U19386 (N_19386,N_19168,N_19121);
or U19387 (N_19387,N_19123,N_19093);
and U19388 (N_19388,N_19120,N_19173);
or U19389 (N_19389,N_19150,N_19021);
xnor U19390 (N_19390,N_19163,N_19102);
nor U19391 (N_19391,N_19022,N_19052);
and U19392 (N_19392,N_19058,N_19044);
xor U19393 (N_19393,N_19118,N_19143);
and U19394 (N_19394,N_19063,N_19167);
xor U19395 (N_19395,N_19070,N_19197);
or U19396 (N_19396,N_19020,N_19036);
or U19397 (N_19397,N_19025,N_19123);
nor U19398 (N_19398,N_19031,N_19002);
and U19399 (N_19399,N_19110,N_19014);
nand U19400 (N_19400,N_19208,N_19325);
nand U19401 (N_19401,N_19344,N_19333);
xor U19402 (N_19402,N_19279,N_19374);
or U19403 (N_19403,N_19352,N_19353);
nor U19404 (N_19404,N_19350,N_19362);
and U19405 (N_19405,N_19226,N_19312);
nand U19406 (N_19406,N_19246,N_19258);
nor U19407 (N_19407,N_19268,N_19377);
nor U19408 (N_19408,N_19283,N_19367);
xor U19409 (N_19409,N_19340,N_19231);
or U19410 (N_19410,N_19274,N_19320);
nor U19411 (N_19411,N_19277,N_19330);
or U19412 (N_19412,N_19219,N_19372);
and U19413 (N_19413,N_19217,N_19381);
and U19414 (N_19414,N_19328,N_19270);
and U19415 (N_19415,N_19302,N_19289);
or U19416 (N_19416,N_19349,N_19318);
nor U19417 (N_19417,N_19201,N_19371);
xnor U19418 (N_19418,N_19384,N_19299);
xor U19419 (N_19419,N_19296,N_19308);
xor U19420 (N_19420,N_19248,N_19238);
and U19421 (N_19421,N_19388,N_19273);
xor U19422 (N_19422,N_19360,N_19310);
nand U19423 (N_19423,N_19244,N_19361);
and U19424 (N_19424,N_19233,N_19394);
and U19425 (N_19425,N_19383,N_19324);
and U19426 (N_19426,N_19234,N_19269);
nand U19427 (N_19427,N_19319,N_19306);
and U19428 (N_19428,N_19210,N_19316);
and U19429 (N_19429,N_19207,N_19313);
xor U19430 (N_19430,N_19245,N_19282);
nand U19431 (N_19431,N_19332,N_19376);
nand U19432 (N_19432,N_19253,N_19396);
nor U19433 (N_19433,N_19285,N_19323);
nand U19434 (N_19434,N_19251,N_19204);
or U19435 (N_19435,N_19221,N_19365);
and U19436 (N_19436,N_19202,N_19220);
nand U19437 (N_19437,N_19382,N_19255);
and U19438 (N_19438,N_19256,N_19264);
nand U19439 (N_19439,N_19375,N_19286);
or U19440 (N_19440,N_19366,N_19370);
or U19441 (N_19441,N_19398,N_19250);
or U19442 (N_19442,N_19363,N_19243);
or U19443 (N_19443,N_19291,N_19228);
nor U19444 (N_19444,N_19338,N_19364);
nor U19445 (N_19445,N_19281,N_19314);
nor U19446 (N_19446,N_19267,N_19395);
nor U19447 (N_19447,N_19378,N_19331);
or U19448 (N_19448,N_19290,N_19393);
xnor U19449 (N_19449,N_19347,N_19288);
xor U19450 (N_19450,N_19224,N_19303);
or U19451 (N_19451,N_19392,N_19214);
nor U19452 (N_19452,N_19239,N_19271);
xor U19453 (N_19453,N_19209,N_19240);
nor U19454 (N_19454,N_19227,N_19272);
or U19455 (N_19455,N_19345,N_19300);
or U19456 (N_19456,N_19295,N_19354);
xor U19457 (N_19457,N_19337,N_19351);
nand U19458 (N_19458,N_19358,N_19212);
xor U19459 (N_19459,N_19343,N_19322);
and U19460 (N_19460,N_19346,N_19397);
xor U19461 (N_19461,N_19311,N_19336);
nand U19462 (N_19462,N_19309,N_19293);
xnor U19463 (N_19463,N_19389,N_19297);
and U19464 (N_19464,N_19301,N_19284);
xnor U19465 (N_19465,N_19305,N_19379);
xnor U19466 (N_19466,N_19387,N_19278);
and U19467 (N_19467,N_19307,N_19298);
nor U19468 (N_19468,N_19380,N_19223);
xor U19469 (N_19469,N_19236,N_19335);
nor U19470 (N_19470,N_19242,N_19235);
nor U19471 (N_19471,N_19315,N_19215);
nand U19472 (N_19472,N_19211,N_19232);
nor U19473 (N_19473,N_19369,N_19222);
nand U19474 (N_19474,N_19200,N_19257);
or U19475 (N_19475,N_19342,N_19237);
nand U19476 (N_19476,N_19356,N_19359);
xnor U19477 (N_19477,N_19275,N_19292);
or U19478 (N_19478,N_19334,N_19326);
or U19479 (N_19479,N_19225,N_19249);
or U19480 (N_19480,N_19391,N_19386);
xnor U19481 (N_19481,N_19229,N_19357);
xor U19482 (N_19482,N_19304,N_19203);
nand U19483 (N_19483,N_19355,N_19260);
xnor U19484 (N_19484,N_19261,N_19294);
nand U19485 (N_19485,N_19321,N_19341);
or U19486 (N_19486,N_19213,N_19317);
or U19487 (N_19487,N_19373,N_19280);
xor U19488 (N_19488,N_19230,N_19266);
or U19489 (N_19489,N_19276,N_19329);
nand U19490 (N_19490,N_19390,N_19287);
xnor U19491 (N_19491,N_19241,N_19339);
nand U19492 (N_19492,N_19247,N_19348);
or U19493 (N_19493,N_19265,N_19216);
or U19494 (N_19494,N_19262,N_19218);
and U19495 (N_19495,N_19327,N_19263);
xor U19496 (N_19496,N_19259,N_19205);
nand U19497 (N_19497,N_19254,N_19368);
xnor U19498 (N_19498,N_19252,N_19385);
nand U19499 (N_19499,N_19206,N_19399);
and U19500 (N_19500,N_19249,N_19246);
or U19501 (N_19501,N_19350,N_19300);
xnor U19502 (N_19502,N_19379,N_19332);
nor U19503 (N_19503,N_19296,N_19350);
xor U19504 (N_19504,N_19236,N_19223);
xnor U19505 (N_19505,N_19399,N_19371);
xnor U19506 (N_19506,N_19374,N_19341);
nor U19507 (N_19507,N_19204,N_19280);
and U19508 (N_19508,N_19303,N_19228);
xor U19509 (N_19509,N_19329,N_19261);
nor U19510 (N_19510,N_19370,N_19299);
or U19511 (N_19511,N_19351,N_19363);
and U19512 (N_19512,N_19223,N_19384);
nand U19513 (N_19513,N_19208,N_19276);
nor U19514 (N_19514,N_19210,N_19349);
nor U19515 (N_19515,N_19384,N_19348);
and U19516 (N_19516,N_19339,N_19364);
xor U19517 (N_19517,N_19219,N_19291);
and U19518 (N_19518,N_19326,N_19206);
nor U19519 (N_19519,N_19301,N_19254);
nor U19520 (N_19520,N_19389,N_19377);
xor U19521 (N_19521,N_19276,N_19362);
xnor U19522 (N_19522,N_19352,N_19262);
and U19523 (N_19523,N_19374,N_19283);
or U19524 (N_19524,N_19286,N_19207);
or U19525 (N_19525,N_19283,N_19246);
or U19526 (N_19526,N_19332,N_19377);
nand U19527 (N_19527,N_19207,N_19213);
nor U19528 (N_19528,N_19263,N_19277);
or U19529 (N_19529,N_19227,N_19335);
nor U19530 (N_19530,N_19216,N_19307);
nor U19531 (N_19531,N_19324,N_19285);
or U19532 (N_19532,N_19210,N_19315);
nor U19533 (N_19533,N_19265,N_19203);
and U19534 (N_19534,N_19314,N_19232);
and U19535 (N_19535,N_19274,N_19391);
xnor U19536 (N_19536,N_19375,N_19261);
or U19537 (N_19537,N_19333,N_19294);
nor U19538 (N_19538,N_19379,N_19294);
and U19539 (N_19539,N_19219,N_19220);
xnor U19540 (N_19540,N_19239,N_19223);
nand U19541 (N_19541,N_19250,N_19383);
xnor U19542 (N_19542,N_19204,N_19255);
or U19543 (N_19543,N_19377,N_19204);
nor U19544 (N_19544,N_19396,N_19302);
and U19545 (N_19545,N_19291,N_19238);
or U19546 (N_19546,N_19354,N_19363);
or U19547 (N_19547,N_19235,N_19327);
and U19548 (N_19548,N_19273,N_19308);
xnor U19549 (N_19549,N_19396,N_19382);
or U19550 (N_19550,N_19221,N_19346);
nand U19551 (N_19551,N_19316,N_19264);
nand U19552 (N_19552,N_19359,N_19374);
xnor U19553 (N_19553,N_19360,N_19269);
and U19554 (N_19554,N_19301,N_19383);
nor U19555 (N_19555,N_19344,N_19307);
and U19556 (N_19556,N_19268,N_19340);
xnor U19557 (N_19557,N_19290,N_19213);
and U19558 (N_19558,N_19341,N_19221);
or U19559 (N_19559,N_19238,N_19214);
nand U19560 (N_19560,N_19232,N_19320);
and U19561 (N_19561,N_19368,N_19331);
xnor U19562 (N_19562,N_19213,N_19345);
and U19563 (N_19563,N_19355,N_19301);
or U19564 (N_19564,N_19254,N_19292);
xnor U19565 (N_19565,N_19262,N_19210);
nand U19566 (N_19566,N_19241,N_19205);
nand U19567 (N_19567,N_19350,N_19262);
nor U19568 (N_19568,N_19375,N_19270);
or U19569 (N_19569,N_19282,N_19391);
or U19570 (N_19570,N_19308,N_19374);
or U19571 (N_19571,N_19219,N_19376);
xor U19572 (N_19572,N_19398,N_19312);
or U19573 (N_19573,N_19288,N_19228);
nor U19574 (N_19574,N_19224,N_19235);
xnor U19575 (N_19575,N_19239,N_19380);
and U19576 (N_19576,N_19368,N_19248);
nand U19577 (N_19577,N_19200,N_19303);
nand U19578 (N_19578,N_19343,N_19388);
xor U19579 (N_19579,N_19289,N_19246);
xnor U19580 (N_19580,N_19250,N_19311);
or U19581 (N_19581,N_19343,N_19345);
and U19582 (N_19582,N_19282,N_19294);
and U19583 (N_19583,N_19266,N_19241);
and U19584 (N_19584,N_19288,N_19280);
nor U19585 (N_19585,N_19317,N_19329);
and U19586 (N_19586,N_19375,N_19314);
xor U19587 (N_19587,N_19294,N_19228);
or U19588 (N_19588,N_19381,N_19366);
and U19589 (N_19589,N_19291,N_19388);
or U19590 (N_19590,N_19240,N_19343);
nor U19591 (N_19591,N_19238,N_19343);
xor U19592 (N_19592,N_19394,N_19332);
xor U19593 (N_19593,N_19320,N_19234);
or U19594 (N_19594,N_19250,N_19202);
nor U19595 (N_19595,N_19372,N_19266);
xor U19596 (N_19596,N_19304,N_19383);
nor U19597 (N_19597,N_19213,N_19222);
xor U19598 (N_19598,N_19364,N_19348);
nor U19599 (N_19599,N_19326,N_19377);
or U19600 (N_19600,N_19402,N_19593);
nand U19601 (N_19601,N_19450,N_19509);
nor U19602 (N_19602,N_19455,N_19495);
and U19603 (N_19603,N_19416,N_19410);
xor U19604 (N_19604,N_19542,N_19513);
and U19605 (N_19605,N_19598,N_19506);
nor U19606 (N_19606,N_19556,N_19444);
nor U19607 (N_19607,N_19480,N_19445);
nand U19608 (N_19608,N_19572,N_19533);
nand U19609 (N_19609,N_19423,N_19515);
nand U19610 (N_19610,N_19493,N_19404);
nand U19611 (N_19611,N_19427,N_19528);
nor U19612 (N_19612,N_19578,N_19585);
and U19613 (N_19613,N_19459,N_19567);
xnor U19614 (N_19614,N_19541,N_19523);
and U19615 (N_19615,N_19453,N_19510);
or U19616 (N_19616,N_19486,N_19560);
or U19617 (N_19617,N_19597,N_19518);
and U19618 (N_19618,N_19573,N_19488);
xor U19619 (N_19619,N_19526,N_19463);
and U19620 (N_19620,N_19507,N_19530);
nand U19621 (N_19621,N_19456,N_19532);
xor U19622 (N_19622,N_19469,N_19487);
and U19623 (N_19623,N_19421,N_19483);
nand U19624 (N_19624,N_19589,N_19412);
nor U19625 (N_19625,N_19475,N_19409);
nand U19626 (N_19626,N_19545,N_19579);
and U19627 (N_19627,N_19477,N_19544);
xnor U19628 (N_19628,N_19595,N_19519);
nand U19629 (N_19629,N_19422,N_19552);
xnor U19630 (N_19630,N_19586,N_19537);
or U19631 (N_19631,N_19599,N_19529);
or U19632 (N_19632,N_19516,N_19464);
xnor U19633 (N_19633,N_19407,N_19505);
nand U19634 (N_19634,N_19558,N_19442);
and U19635 (N_19635,N_19562,N_19555);
and U19636 (N_19636,N_19446,N_19574);
xnor U19637 (N_19637,N_19548,N_19539);
nor U19638 (N_19638,N_19575,N_19522);
and U19639 (N_19639,N_19466,N_19411);
or U19640 (N_19640,N_19582,N_19594);
and U19641 (N_19641,N_19448,N_19429);
nor U19642 (N_19642,N_19403,N_19592);
and U19643 (N_19643,N_19476,N_19461);
nor U19644 (N_19644,N_19501,N_19497);
nand U19645 (N_19645,N_19540,N_19465);
nor U19646 (N_19646,N_19491,N_19568);
or U19647 (N_19647,N_19474,N_19470);
xor U19648 (N_19648,N_19449,N_19451);
nor U19649 (N_19649,N_19436,N_19581);
xnor U19650 (N_19650,N_19571,N_19524);
nand U19651 (N_19651,N_19473,N_19511);
nand U19652 (N_19652,N_19489,N_19547);
nor U19653 (N_19653,N_19479,N_19441);
nand U19654 (N_19654,N_19460,N_19462);
nand U19655 (N_19655,N_19431,N_19408);
xnor U19656 (N_19656,N_19433,N_19498);
nor U19657 (N_19657,N_19417,N_19428);
or U19658 (N_19658,N_19467,N_19484);
and U19659 (N_19659,N_19527,N_19517);
and U19660 (N_19660,N_19546,N_19485);
nand U19661 (N_19661,N_19536,N_19551);
xor U19662 (N_19662,N_19426,N_19419);
or U19663 (N_19663,N_19588,N_19434);
and U19664 (N_19664,N_19520,N_19554);
and U19665 (N_19665,N_19535,N_19468);
or U19666 (N_19666,N_19502,N_19439);
nand U19667 (N_19667,N_19525,N_19564);
and U19668 (N_19668,N_19482,N_19432);
nand U19669 (N_19669,N_19500,N_19563);
or U19670 (N_19670,N_19424,N_19472);
nand U19671 (N_19671,N_19457,N_19587);
nor U19672 (N_19672,N_19443,N_19580);
or U19673 (N_19673,N_19437,N_19406);
xnor U19674 (N_19674,N_19521,N_19591);
xor U19675 (N_19675,N_19413,N_19557);
and U19676 (N_19676,N_19452,N_19534);
nor U19677 (N_19677,N_19503,N_19584);
or U19678 (N_19678,N_19492,N_19415);
or U19679 (N_19679,N_19569,N_19550);
or U19680 (N_19680,N_19496,N_19420);
and U19681 (N_19681,N_19590,N_19401);
or U19682 (N_19682,N_19531,N_19565);
xnor U19683 (N_19683,N_19543,N_19440);
or U19684 (N_19684,N_19508,N_19447);
and U19685 (N_19685,N_19577,N_19576);
nor U19686 (N_19686,N_19596,N_19454);
and U19687 (N_19687,N_19400,N_19570);
nor U19688 (N_19688,N_19504,N_19490);
nor U19689 (N_19689,N_19481,N_19494);
xor U19690 (N_19690,N_19538,N_19583);
nand U19691 (N_19691,N_19499,N_19405);
or U19692 (N_19692,N_19418,N_19559);
or U19693 (N_19693,N_19430,N_19514);
and U19694 (N_19694,N_19425,N_19471);
and U19695 (N_19695,N_19458,N_19566);
and U19696 (N_19696,N_19414,N_19512);
xnor U19697 (N_19697,N_19438,N_19549);
nand U19698 (N_19698,N_19435,N_19561);
or U19699 (N_19699,N_19478,N_19553);
nand U19700 (N_19700,N_19491,N_19456);
or U19701 (N_19701,N_19542,N_19445);
nand U19702 (N_19702,N_19542,N_19437);
xnor U19703 (N_19703,N_19427,N_19407);
xnor U19704 (N_19704,N_19491,N_19554);
and U19705 (N_19705,N_19405,N_19446);
nor U19706 (N_19706,N_19456,N_19541);
xor U19707 (N_19707,N_19487,N_19516);
nor U19708 (N_19708,N_19525,N_19520);
xor U19709 (N_19709,N_19448,N_19520);
or U19710 (N_19710,N_19428,N_19414);
or U19711 (N_19711,N_19568,N_19479);
and U19712 (N_19712,N_19479,N_19503);
nor U19713 (N_19713,N_19531,N_19511);
nand U19714 (N_19714,N_19576,N_19457);
nor U19715 (N_19715,N_19474,N_19458);
nand U19716 (N_19716,N_19570,N_19547);
and U19717 (N_19717,N_19513,N_19576);
or U19718 (N_19718,N_19480,N_19467);
nand U19719 (N_19719,N_19552,N_19503);
xnor U19720 (N_19720,N_19571,N_19442);
nor U19721 (N_19721,N_19574,N_19404);
or U19722 (N_19722,N_19455,N_19409);
nor U19723 (N_19723,N_19571,N_19503);
and U19724 (N_19724,N_19427,N_19505);
nand U19725 (N_19725,N_19450,N_19522);
and U19726 (N_19726,N_19529,N_19591);
or U19727 (N_19727,N_19541,N_19589);
nand U19728 (N_19728,N_19554,N_19496);
xor U19729 (N_19729,N_19490,N_19445);
nand U19730 (N_19730,N_19535,N_19453);
xnor U19731 (N_19731,N_19470,N_19521);
or U19732 (N_19732,N_19511,N_19437);
xor U19733 (N_19733,N_19559,N_19558);
xor U19734 (N_19734,N_19573,N_19552);
and U19735 (N_19735,N_19471,N_19434);
nand U19736 (N_19736,N_19476,N_19432);
xnor U19737 (N_19737,N_19409,N_19589);
and U19738 (N_19738,N_19487,N_19533);
or U19739 (N_19739,N_19455,N_19552);
xor U19740 (N_19740,N_19472,N_19422);
xor U19741 (N_19741,N_19553,N_19502);
xnor U19742 (N_19742,N_19511,N_19472);
and U19743 (N_19743,N_19583,N_19474);
and U19744 (N_19744,N_19555,N_19456);
nor U19745 (N_19745,N_19456,N_19583);
xor U19746 (N_19746,N_19579,N_19445);
or U19747 (N_19747,N_19509,N_19433);
and U19748 (N_19748,N_19432,N_19523);
nor U19749 (N_19749,N_19440,N_19409);
nand U19750 (N_19750,N_19492,N_19586);
xor U19751 (N_19751,N_19561,N_19416);
or U19752 (N_19752,N_19515,N_19466);
or U19753 (N_19753,N_19589,N_19484);
xor U19754 (N_19754,N_19497,N_19576);
xor U19755 (N_19755,N_19589,N_19594);
xnor U19756 (N_19756,N_19558,N_19577);
and U19757 (N_19757,N_19594,N_19429);
nor U19758 (N_19758,N_19495,N_19535);
nand U19759 (N_19759,N_19573,N_19418);
nor U19760 (N_19760,N_19401,N_19456);
nand U19761 (N_19761,N_19428,N_19425);
xor U19762 (N_19762,N_19539,N_19453);
and U19763 (N_19763,N_19449,N_19477);
xor U19764 (N_19764,N_19536,N_19584);
and U19765 (N_19765,N_19486,N_19509);
xnor U19766 (N_19766,N_19428,N_19575);
or U19767 (N_19767,N_19460,N_19444);
and U19768 (N_19768,N_19474,N_19547);
nand U19769 (N_19769,N_19563,N_19531);
nand U19770 (N_19770,N_19420,N_19506);
nand U19771 (N_19771,N_19526,N_19445);
nand U19772 (N_19772,N_19498,N_19451);
or U19773 (N_19773,N_19493,N_19590);
nor U19774 (N_19774,N_19515,N_19500);
and U19775 (N_19775,N_19511,N_19466);
or U19776 (N_19776,N_19418,N_19531);
nand U19777 (N_19777,N_19503,N_19525);
xnor U19778 (N_19778,N_19588,N_19486);
nand U19779 (N_19779,N_19482,N_19445);
and U19780 (N_19780,N_19438,N_19587);
nand U19781 (N_19781,N_19544,N_19453);
and U19782 (N_19782,N_19471,N_19519);
nand U19783 (N_19783,N_19561,N_19420);
and U19784 (N_19784,N_19414,N_19545);
or U19785 (N_19785,N_19484,N_19452);
nand U19786 (N_19786,N_19513,N_19464);
or U19787 (N_19787,N_19553,N_19574);
nor U19788 (N_19788,N_19552,N_19505);
or U19789 (N_19789,N_19514,N_19502);
nor U19790 (N_19790,N_19542,N_19416);
nor U19791 (N_19791,N_19585,N_19513);
nand U19792 (N_19792,N_19587,N_19444);
nand U19793 (N_19793,N_19478,N_19534);
or U19794 (N_19794,N_19466,N_19497);
and U19795 (N_19795,N_19471,N_19526);
nand U19796 (N_19796,N_19444,N_19486);
xor U19797 (N_19797,N_19569,N_19520);
nand U19798 (N_19798,N_19466,N_19503);
or U19799 (N_19799,N_19470,N_19503);
nor U19800 (N_19800,N_19785,N_19666);
and U19801 (N_19801,N_19699,N_19679);
nand U19802 (N_19802,N_19766,N_19767);
nand U19803 (N_19803,N_19751,N_19788);
nand U19804 (N_19804,N_19704,N_19737);
or U19805 (N_19805,N_19692,N_19650);
nand U19806 (N_19806,N_19633,N_19774);
and U19807 (N_19807,N_19635,N_19670);
and U19808 (N_19808,N_19615,N_19778);
nor U19809 (N_19809,N_19651,N_19676);
and U19810 (N_19810,N_19682,N_19631);
or U19811 (N_19811,N_19758,N_19713);
and U19812 (N_19812,N_19753,N_19625);
or U19813 (N_19813,N_19773,N_19782);
xnor U19814 (N_19814,N_19762,N_19678);
nor U19815 (N_19815,N_19728,N_19603);
xor U19816 (N_19816,N_19746,N_19671);
nor U19817 (N_19817,N_19771,N_19664);
nor U19818 (N_19818,N_19777,N_19744);
xor U19819 (N_19819,N_19765,N_19747);
and U19820 (N_19820,N_19675,N_19695);
or U19821 (N_19821,N_19661,N_19677);
xor U19822 (N_19822,N_19764,N_19646);
xor U19823 (N_19823,N_19748,N_19623);
and U19824 (N_19824,N_19653,N_19601);
and U19825 (N_19825,N_19790,N_19725);
xor U19826 (N_19826,N_19688,N_19637);
or U19827 (N_19827,N_19609,N_19719);
nand U19828 (N_19828,N_19618,N_19647);
or U19829 (N_19829,N_19617,N_19648);
nand U19830 (N_19830,N_19693,N_19757);
or U19831 (N_19831,N_19644,N_19681);
nor U19832 (N_19832,N_19740,N_19684);
and U19833 (N_19833,N_19752,N_19750);
or U19834 (N_19834,N_19658,N_19720);
nor U19835 (N_19835,N_19768,N_19760);
and U19836 (N_19836,N_19745,N_19718);
or U19837 (N_19837,N_19660,N_19749);
and U19838 (N_19838,N_19795,N_19687);
or U19839 (N_19839,N_19792,N_19616);
and U19840 (N_19840,N_19781,N_19636);
xor U19841 (N_19841,N_19629,N_19686);
and U19842 (N_19842,N_19708,N_19736);
and U19843 (N_19843,N_19639,N_19717);
and U19844 (N_19844,N_19673,N_19657);
or U19845 (N_19845,N_19709,N_19667);
xor U19846 (N_19846,N_19793,N_19784);
nand U19847 (N_19847,N_19607,N_19685);
nor U19848 (N_19848,N_19712,N_19627);
or U19849 (N_19849,N_19789,N_19654);
or U19850 (N_19850,N_19630,N_19726);
nand U19851 (N_19851,N_19696,N_19761);
or U19852 (N_19852,N_19614,N_19705);
nand U19853 (N_19853,N_19714,N_19727);
and U19854 (N_19854,N_19626,N_19632);
nor U19855 (N_19855,N_19663,N_19783);
nor U19856 (N_19856,N_19770,N_19741);
and U19857 (N_19857,N_19703,N_19662);
and U19858 (N_19858,N_19743,N_19797);
and U19859 (N_19859,N_19642,N_19799);
nand U19860 (N_19860,N_19721,N_19796);
or U19861 (N_19861,N_19619,N_19780);
xnor U19862 (N_19862,N_19710,N_19612);
nor U19863 (N_19863,N_19772,N_19649);
nand U19864 (N_19864,N_19702,N_19742);
nand U19865 (N_19865,N_19643,N_19707);
and U19866 (N_19866,N_19739,N_19689);
and U19867 (N_19867,N_19624,N_19735);
or U19868 (N_19868,N_19754,N_19672);
nor U19869 (N_19869,N_19604,N_19638);
and U19870 (N_19870,N_19668,N_19763);
nand U19871 (N_19871,N_19716,N_19621);
or U19872 (N_19872,N_19690,N_19640);
nor U19873 (N_19873,N_19680,N_19794);
nand U19874 (N_19874,N_19715,N_19610);
xnor U19875 (N_19875,N_19620,N_19786);
and U19876 (N_19876,N_19641,N_19645);
nand U19877 (N_19877,N_19730,N_19652);
xor U19878 (N_19878,N_19613,N_19734);
nand U19879 (N_19879,N_19698,N_19759);
xor U19880 (N_19880,N_19634,N_19756);
or U19881 (N_19881,N_19606,N_19665);
or U19882 (N_19882,N_19722,N_19697);
xnor U19883 (N_19883,N_19724,N_19611);
nand U19884 (N_19884,N_19729,N_19655);
nand U19885 (N_19885,N_19700,N_19779);
xnor U19886 (N_19886,N_19691,N_19711);
xor U19887 (N_19887,N_19791,N_19600);
xor U19888 (N_19888,N_19608,N_19602);
or U19889 (N_19889,N_19694,N_19656);
or U19890 (N_19890,N_19723,N_19674);
or U19891 (N_19891,N_19628,N_19605);
or U19892 (N_19892,N_19659,N_19775);
xor U19893 (N_19893,N_19769,N_19776);
xor U19894 (N_19894,N_19798,N_19732);
or U19895 (N_19895,N_19701,N_19755);
nand U19896 (N_19896,N_19683,N_19731);
and U19897 (N_19897,N_19787,N_19669);
or U19898 (N_19898,N_19733,N_19622);
xnor U19899 (N_19899,N_19738,N_19706);
xnor U19900 (N_19900,N_19735,N_19762);
nor U19901 (N_19901,N_19612,N_19762);
xor U19902 (N_19902,N_19723,N_19616);
and U19903 (N_19903,N_19649,N_19620);
xor U19904 (N_19904,N_19714,N_19696);
nor U19905 (N_19905,N_19738,N_19628);
or U19906 (N_19906,N_19786,N_19666);
and U19907 (N_19907,N_19779,N_19678);
and U19908 (N_19908,N_19714,N_19692);
nor U19909 (N_19909,N_19789,N_19723);
nor U19910 (N_19910,N_19777,N_19689);
nor U19911 (N_19911,N_19701,N_19790);
nand U19912 (N_19912,N_19796,N_19694);
and U19913 (N_19913,N_19600,N_19696);
xor U19914 (N_19914,N_19724,N_19732);
and U19915 (N_19915,N_19618,N_19664);
xnor U19916 (N_19916,N_19628,N_19649);
or U19917 (N_19917,N_19761,N_19762);
or U19918 (N_19918,N_19645,N_19717);
or U19919 (N_19919,N_19741,N_19706);
and U19920 (N_19920,N_19696,N_19704);
nand U19921 (N_19921,N_19713,N_19730);
xnor U19922 (N_19922,N_19748,N_19618);
or U19923 (N_19923,N_19639,N_19745);
or U19924 (N_19924,N_19644,N_19719);
nor U19925 (N_19925,N_19702,N_19621);
nand U19926 (N_19926,N_19667,N_19660);
nor U19927 (N_19927,N_19602,N_19715);
or U19928 (N_19928,N_19693,N_19775);
or U19929 (N_19929,N_19623,N_19603);
xnor U19930 (N_19930,N_19629,N_19720);
nand U19931 (N_19931,N_19784,N_19725);
or U19932 (N_19932,N_19678,N_19765);
or U19933 (N_19933,N_19777,N_19713);
xnor U19934 (N_19934,N_19756,N_19701);
or U19935 (N_19935,N_19773,N_19753);
nor U19936 (N_19936,N_19614,N_19723);
xnor U19937 (N_19937,N_19617,N_19728);
nor U19938 (N_19938,N_19691,N_19654);
nor U19939 (N_19939,N_19631,N_19728);
and U19940 (N_19940,N_19658,N_19790);
or U19941 (N_19941,N_19720,N_19617);
xor U19942 (N_19942,N_19622,N_19649);
or U19943 (N_19943,N_19605,N_19690);
nand U19944 (N_19944,N_19749,N_19689);
nand U19945 (N_19945,N_19699,N_19775);
or U19946 (N_19946,N_19675,N_19721);
nor U19947 (N_19947,N_19627,N_19689);
nand U19948 (N_19948,N_19680,N_19688);
nor U19949 (N_19949,N_19708,N_19699);
or U19950 (N_19950,N_19602,N_19691);
nand U19951 (N_19951,N_19712,N_19634);
nor U19952 (N_19952,N_19654,N_19613);
xnor U19953 (N_19953,N_19743,N_19644);
xor U19954 (N_19954,N_19659,N_19799);
and U19955 (N_19955,N_19617,N_19650);
and U19956 (N_19956,N_19606,N_19708);
nor U19957 (N_19957,N_19633,N_19654);
or U19958 (N_19958,N_19771,N_19742);
or U19959 (N_19959,N_19703,N_19737);
nor U19960 (N_19960,N_19753,N_19759);
nand U19961 (N_19961,N_19719,N_19774);
and U19962 (N_19962,N_19722,N_19610);
nor U19963 (N_19963,N_19614,N_19626);
nor U19964 (N_19964,N_19733,N_19727);
nand U19965 (N_19965,N_19708,N_19754);
or U19966 (N_19966,N_19678,N_19749);
nor U19967 (N_19967,N_19629,N_19795);
or U19968 (N_19968,N_19760,N_19664);
and U19969 (N_19969,N_19711,N_19634);
or U19970 (N_19970,N_19631,N_19646);
nand U19971 (N_19971,N_19613,N_19653);
nor U19972 (N_19972,N_19746,N_19661);
or U19973 (N_19973,N_19733,N_19659);
nor U19974 (N_19974,N_19678,N_19771);
xnor U19975 (N_19975,N_19772,N_19754);
nor U19976 (N_19976,N_19646,N_19702);
xnor U19977 (N_19977,N_19759,N_19658);
xnor U19978 (N_19978,N_19753,N_19730);
and U19979 (N_19979,N_19659,N_19640);
nand U19980 (N_19980,N_19667,N_19665);
nand U19981 (N_19981,N_19637,N_19698);
and U19982 (N_19982,N_19689,N_19683);
xnor U19983 (N_19983,N_19773,N_19645);
nor U19984 (N_19984,N_19749,N_19692);
xor U19985 (N_19985,N_19640,N_19707);
nor U19986 (N_19986,N_19612,N_19674);
xor U19987 (N_19987,N_19719,N_19681);
nor U19988 (N_19988,N_19652,N_19610);
and U19989 (N_19989,N_19608,N_19772);
xor U19990 (N_19990,N_19611,N_19638);
nor U19991 (N_19991,N_19688,N_19678);
and U19992 (N_19992,N_19684,N_19630);
nand U19993 (N_19993,N_19646,N_19750);
xnor U19994 (N_19994,N_19737,N_19742);
and U19995 (N_19995,N_19716,N_19617);
or U19996 (N_19996,N_19752,N_19669);
and U19997 (N_19997,N_19622,N_19708);
nand U19998 (N_19998,N_19629,N_19768);
nor U19999 (N_19999,N_19663,N_19667);
and U20000 (N_20000,N_19987,N_19928);
nand U20001 (N_20001,N_19981,N_19903);
nand U20002 (N_20002,N_19976,N_19961);
nor U20003 (N_20003,N_19809,N_19955);
nand U20004 (N_20004,N_19868,N_19880);
xnor U20005 (N_20005,N_19890,N_19852);
xnor U20006 (N_20006,N_19877,N_19846);
nand U20007 (N_20007,N_19949,N_19966);
nor U20008 (N_20008,N_19950,N_19869);
nor U20009 (N_20009,N_19937,N_19896);
and U20010 (N_20010,N_19865,N_19849);
xor U20011 (N_20011,N_19963,N_19951);
nand U20012 (N_20012,N_19986,N_19901);
and U20013 (N_20013,N_19980,N_19945);
xnor U20014 (N_20014,N_19812,N_19837);
nand U20015 (N_20015,N_19983,N_19922);
xor U20016 (N_20016,N_19831,N_19806);
nor U20017 (N_20017,N_19910,N_19838);
or U20018 (N_20018,N_19925,N_19946);
nand U20019 (N_20019,N_19829,N_19904);
xnor U20020 (N_20020,N_19824,N_19940);
nor U20021 (N_20021,N_19832,N_19834);
or U20022 (N_20022,N_19825,N_19856);
or U20023 (N_20023,N_19914,N_19997);
nand U20024 (N_20024,N_19857,N_19858);
and U20025 (N_20025,N_19891,N_19969);
or U20026 (N_20026,N_19828,N_19855);
nand U20027 (N_20027,N_19820,N_19967);
nor U20028 (N_20028,N_19893,N_19885);
or U20029 (N_20029,N_19836,N_19962);
or U20030 (N_20030,N_19802,N_19916);
nand U20031 (N_20031,N_19985,N_19822);
or U20032 (N_20032,N_19841,N_19912);
or U20033 (N_20033,N_19804,N_19939);
nand U20034 (N_20034,N_19844,N_19948);
nand U20035 (N_20035,N_19860,N_19982);
and U20036 (N_20036,N_19821,N_19805);
nand U20037 (N_20037,N_19847,N_19861);
xor U20038 (N_20038,N_19813,N_19902);
nand U20039 (N_20039,N_19835,N_19935);
xor U20040 (N_20040,N_19971,N_19905);
or U20041 (N_20041,N_19895,N_19881);
nand U20042 (N_20042,N_19814,N_19898);
and U20043 (N_20043,N_19818,N_19990);
nor U20044 (N_20044,N_19899,N_19906);
and U20045 (N_20045,N_19974,N_19989);
nand U20046 (N_20046,N_19862,N_19871);
nand U20047 (N_20047,N_19840,N_19859);
or U20048 (N_20048,N_19992,N_19968);
or U20049 (N_20049,N_19897,N_19908);
nor U20050 (N_20050,N_19960,N_19873);
and U20051 (N_20051,N_19984,N_19882);
nor U20052 (N_20052,N_19938,N_19921);
or U20053 (N_20053,N_19920,N_19826);
or U20054 (N_20054,N_19915,N_19965);
or U20055 (N_20055,N_19995,N_19853);
or U20056 (N_20056,N_19907,N_19801);
nand U20057 (N_20057,N_19952,N_19917);
xnor U20058 (N_20058,N_19839,N_19878);
nor U20059 (N_20059,N_19867,N_19959);
nor U20060 (N_20060,N_19947,N_19927);
xor U20061 (N_20061,N_19964,N_19854);
nand U20062 (N_20062,N_19979,N_19886);
nand U20063 (N_20063,N_19972,N_19884);
xnor U20064 (N_20064,N_19936,N_19931);
nand U20065 (N_20065,N_19978,N_19944);
and U20066 (N_20066,N_19817,N_19816);
and U20067 (N_20067,N_19954,N_19930);
nor U20068 (N_20068,N_19845,N_19866);
nor U20069 (N_20069,N_19994,N_19870);
nand U20070 (N_20070,N_19888,N_19803);
and U20071 (N_20071,N_19843,N_19988);
xor U20072 (N_20072,N_19993,N_19811);
or U20073 (N_20073,N_19926,N_19833);
nand U20074 (N_20074,N_19887,N_19958);
nand U20075 (N_20075,N_19929,N_19932);
nor U20076 (N_20076,N_19991,N_19808);
nand U20077 (N_20077,N_19919,N_19924);
nor U20078 (N_20078,N_19874,N_19815);
or U20079 (N_20079,N_19943,N_19800);
or U20080 (N_20080,N_19883,N_19850);
xnor U20081 (N_20081,N_19911,N_19827);
nand U20082 (N_20082,N_19810,N_19819);
and U20083 (N_20083,N_19872,N_19996);
xnor U20084 (N_20084,N_19977,N_19913);
nor U20085 (N_20085,N_19953,N_19975);
nor U20086 (N_20086,N_19851,N_19892);
and U20087 (N_20087,N_19848,N_19942);
xor U20088 (N_20088,N_19889,N_19842);
nand U20089 (N_20089,N_19875,N_19918);
nor U20090 (N_20090,N_19957,N_19879);
nor U20091 (N_20091,N_19973,N_19933);
xor U20092 (N_20092,N_19999,N_19941);
nand U20093 (N_20093,N_19956,N_19970);
nor U20094 (N_20094,N_19823,N_19909);
nand U20095 (N_20095,N_19876,N_19807);
xnor U20096 (N_20096,N_19830,N_19998);
or U20097 (N_20097,N_19863,N_19864);
and U20098 (N_20098,N_19900,N_19894);
nor U20099 (N_20099,N_19923,N_19934);
and U20100 (N_20100,N_19949,N_19870);
xor U20101 (N_20101,N_19800,N_19925);
or U20102 (N_20102,N_19813,N_19969);
or U20103 (N_20103,N_19970,N_19878);
or U20104 (N_20104,N_19859,N_19831);
and U20105 (N_20105,N_19961,N_19809);
and U20106 (N_20106,N_19860,N_19888);
nand U20107 (N_20107,N_19899,N_19810);
or U20108 (N_20108,N_19827,N_19899);
or U20109 (N_20109,N_19809,N_19922);
xnor U20110 (N_20110,N_19974,N_19802);
xnor U20111 (N_20111,N_19818,N_19860);
nand U20112 (N_20112,N_19817,N_19825);
or U20113 (N_20113,N_19986,N_19884);
or U20114 (N_20114,N_19806,N_19920);
and U20115 (N_20115,N_19838,N_19908);
xnor U20116 (N_20116,N_19897,N_19823);
or U20117 (N_20117,N_19823,N_19896);
and U20118 (N_20118,N_19830,N_19922);
xnor U20119 (N_20119,N_19885,N_19824);
xor U20120 (N_20120,N_19867,N_19974);
nand U20121 (N_20121,N_19858,N_19892);
or U20122 (N_20122,N_19956,N_19816);
nand U20123 (N_20123,N_19957,N_19869);
nor U20124 (N_20124,N_19862,N_19849);
nor U20125 (N_20125,N_19855,N_19956);
or U20126 (N_20126,N_19911,N_19899);
nor U20127 (N_20127,N_19803,N_19899);
nand U20128 (N_20128,N_19805,N_19991);
xor U20129 (N_20129,N_19835,N_19989);
or U20130 (N_20130,N_19874,N_19842);
or U20131 (N_20131,N_19806,N_19939);
nor U20132 (N_20132,N_19808,N_19977);
or U20133 (N_20133,N_19937,N_19820);
xnor U20134 (N_20134,N_19900,N_19915);
nand U20135 (N_20135,N_19962,N_19950);
nand U20136 (N_20136,N_19989,N_19911);
xor U20137 (N_20137,N_19842,N_19963);
nand U20138 (N_20138,N_19887,N_19899);
nor U20139 (N_20139,N_19966,N_19910);
or U20140 (N_20140,N_19991,N_19814);
and U20141 (N_20141,N_19964,N_19884);
nand U20142 (N_20142,N_19828,N_19971);
nor U20143 (N_20143,N_19953,N_19943);
nand U20144 (N_20144,N_19974,N_19899);
xor U20145 (N_20145,N_19898,N_19992);
or U20146 (N_20146,N_19801,N_19875);
xor U20147 (N_20147,N_19990,N_19863);
xnor U20148 (N_20148,N_19935,N_19953);
nand U20149 (N_20149,N_19881,N_19993);
nand U20150 (N_20150,N_19834,N_19940);
xnor U20151 (N_20151,N_19981,N_19818);
or U20152 (N_20152,N_19972,N_19943);
and U20153 (N_20153,N_19973,N_19872);
or U20154 (N_20154,N_19803,N_19846);
nand U20155 (N_20155,N_19990,N_19893);
or U20156 (N_20156,N_19938,N_19908);
and U20157 (N_20157,N_19873,N_19993);
nor U20158 (N_20158,N_19965,N_19936);
nand U20159 (N_20159,N_19871,N_19912);
nand U20160 (N_20160,N_19950,N_19912);
or U20161 (N_20161,N_19844,N_19924);
xor U20162 (N_20162,N_19912,N_19882);
and U20163 (N_20163,N_19825,N_19901);
xor U20164 (N_20164,N_19948,N_19939);
and U20165 (N_20165,N_19919,N_19914);
nor U20166 (N_20166,N_19856,N_19884);
and U20167 (N_20167,N_19884,N_19808);
and U20168 (N_20168,N_19874,N_19966);
nor U20169 (N_20169,N_19971,N_19862);
nor U20170 (N_20170,N_19922,N_19992);
and U20171 (N_20171,N_19914,N_19968);
xor U20172 (N_20172,N_19905,N_19878);
and U20173 (N_20173,N_19965,N_19864);
and U20174 (N_20174,N_19845,N_19890);
xor U20175 (N_20175,N_19888,N_19880);
nand U20176 (N_20176,N_19979,N_19801);
and U20177 (N_20177,N_19805,N_19939);
nor U20178 (N_20178,N_19977,N_19931);
nand U20179 (N_20179,N_19869,N_19932);
xnor U20180 (N_20180,N_19857,N_19898);
and U20181 (N_20181,N_19969,N_19869);
xor U20182 (N_20182,N_19993,N_19897);
xnor U20183 (N_20183,N_19892,N_19957);
nand U20184 (N_20184,N_19852,N_19806);
or U20185 (N_20185,N_19991,N_19985);
nor U20186 (N_20186,N_19943,N_19870);
nor U20187 (N_20187,N_19954,N_19890);
xnor U20188 (N_20188,N_19997,N_19922);
or U20189 (N_20189,N_19932,N_19954);
or U20190 (N_20190,N_19937,N_19949);
or U20191 (N_20191,N_19814,N_19964);
or U20192 (N_20192,N_19974,N_19856);
nand U20193 (N_20193,N_19882,N_19917);
nand U20194 (N_20194,N_19920,N_19941);
nor U20195 (N_20195,N_19840,N_19846);
and U20196 (N_20196,N_19936,N_19967);
or U20197 (N_20197,N_19856,N_19848);
nand U20198 (N_20198,N_19919,N_19858);
nand U20199 (N_20199,N_19862,N_19914);
or U20200 (N_20200,N_20115,N_20022);
or U20201 (N_20201,N_20190,N_20169);
nor U20202 (N_20202,N_20107,N_20199);
nand U20203 (N_20203,N_20149,N_20043);
nor U20204 (N_20204,N_20028,N_20056);
xnor U20205 (N_20205,N_20013,N_20012);
and U20206 (N_20206,N_20057,N_20133);
and U20207 (N_20207,N_20126,N_20069);
nor U20208 (N_20208,N_20104,N_20196);
and U20209 (N_20209,N_20048,N_20054);
or U20210 (N_20210,N_20095,N_20111);
and U20211 (N_20211,N_20157,N_20154);
xnor U20212 (N_20212,N_20142,N_20038);
or U20213 (N_20213,N_20088,N_20040);
xor U20214 (N_20214,N_20101,N_20117);
or U20215 (N_20215,N_20106,N_20170);
or U20216 (N_20216,N_20179,N_20178);
nor U20217 (N_20217,N_20083,N_20034);
and U20218 (N_20218,N_20121,N_20118);
xnor U20219 (N_20219,N_20008,N_20172);
and U20220 (N_20220,N_20156,N_20145);
and U20221 (N_20221,N_20116,N_20073);
and U20222 (N_20222,N_20015,N_20182);
nor U20223 (N_20223,N_20122,N_20051);
and U20224 (N_20224,N_20176,N_20023);
and U20225 (N_20225,N_20194,N_20079);
nand U20226 (N_20226,N_20119,N_20123);
nor U20227 (N_20227,N_20080,N_20058);
nor U20228 (N_20228,N_20060,N_20053);
xnor U20229 (N_20229,N_20100,N_20006);
nand U20230 (N_20230,N_20067,N_20105);
nand U20231 (N_20231,N_20141,N_20184);
or U20232 (N_20232,N_20193,N_20129);
nand U20233 (N_20233,N_20084,N_20068);
nor U20234 (N_20234,N_20191,N_20150);
or U20235 (N_20235,N_20072,N_20020);
and U20236 (N_20236,N_20186,N_20163);
nand U20237 (N_20237,N_20081,N_20046);
xor U20238 (N_20238,N_20096,N_20114);
or U20239 (N_20239,N_20188,N_20174);
or U20240 (N_20240,N_20042,N_20134);
nand U20241 (N_20241,N_20098,N_20185);
nor U20242 (N_20242,N_20109,N_20148);
nand U20243 (N_20243,N_20161,N_20014);
and U20244 (N_20244,N_20047,N_20030);
or U20245 (N_20245,N_20103,N_20004);
or U20246 (N_20246,N_20125,N_20074);
nor U20247 (N_20247,N_20092,N_20025);
xor U20248 (N_20248,N_20160,N_20075);
or U20249 (N_20249,N_20187,N_20009);
nor U20250 (N_20250,N_20112,N_20087);
nand U20251 (N_20251,N_20183,N_20147);
nand U20252 (N_20252,N_20078,N_20102);
or U20253 (N_20253,N_20017,N_20144);
xnor U20254 (N_20254,N_20164,N_20130);
nor U20255 (N_20255,N_20167,N_20192);
and U20256 (N_20256,N_20029,N_20021);
or U20257 (N_20257,N_20173,N_20143);
xnor U20258 (N_20258,N_20035,N_20089);
or U20259 (N_20259,N_20099,N_20061);
nor U20260 (N_20260,N_20132,N_20151);
and U20261 (N_20261,N_20082,N_20000);
and U20262 (N_20262,N_20097,N_20165);
xor U20263 (N_20263,N_20110,N_20168);
xor U20264 (N_20264,N_20076,N_20064);
xnor U20265 (N_20265,N_20189,N_20065);
xnor U20266 (N_20266,N_20050,N_20032);
xnor U20267 (N_20267,N_20140,N_20019);
nor U20268 (N_20268,N_20007,N_20093);
and U20269 (N_20269,N_20001,N_20041);
and U20270 (N_20270,N_20036,N_20011);
or U20271 (N_20271,N_20085,N_20005);
and U20272 (N_20272,N_20152,N_20177);
and U20273 (N_20273,N_20044,N_20120);
nor U20274 (N_20274,N_20027,N_20090);
xor U20275 (N_20275,N_20108,N_20153);
xor U20276 (N_20276,N_20039,N_20002);
nor U20277 (N_20277,N_20059,N_20033);
or U20278 (N_20278,N_20198,N_20136);
nand U20279 (N_20279,N_20171,N_20113);
nor U20280 (N_20280,N_20086,N_20071);
nor U20281 (N_20281,N_20049,N_20045);
nor U20282 (N_20282,N_20155,N_20195);
and U20283 (N_20283,N_20062,N_20026);
or U20284 (N_20284,N_20138,N_20037);
nor U20285 (N_20285,N_20197,N_20162);
or U20286 (N_20286,N_20146,N_20175);
and U20287 (N_20287,N_20091,N_20128);
xnor U20288 (N_20288,N_20124,N_20159);
nor U20289 (N_20289,N_20180,N_20127);
and U20290 (N_20290,N_20070,N_20024);
and U20291 (N_20291,N_20055,N_20066);
or U20292 (N_20292,N_20063,N_20131);
or U20293 (N_20293,N_20003,N_20137);
xnor U20294 (N_20294,N_20094,N_20010);
xor U20295 (N_20295,N_20181,N_20018);
nand U20296 (N_20296,N_20077,N_20158);
xnor U20297 (N_20297,N_20016,N_20139);
or U20298 (N_20298,N_20166,N_20052);
or U20299 (N_20299,N_20031,N_20135);
and U20300 (N_20300,N_20053,N_20030);
or U20301 (N_20301,N_20159,N_20087);
or U20302 (N_20302,N_20176,N_20114);
and U20303 (N_20303,N_20141,N_20007);
xor U20304 (N_20304,N_20180,N_20075);
and U20305 (N_20305,N_20095,N_20129);
and U20306 (N_20306,N_20114,N_20115);
and U20307 (N_20307,N_20066,N_20097);
and U20308 (N_20308,N_20156,N_20109);
xnor U20309 (N_20309,N_20194,N_20020);
and U20310 (N_20310,N_20115,N_20017);
or U20311 (N_20311,N_20093,N_20175);
or U20312 (N_20312,N_20029,N_20077);
nor U20313 (N_20313,N_20186,N_20120);
and U20314 (N_20314,N_20007,N_20169);
nand U20315 (N_20315,N_20111,N_20073);
or U20316 (N_20316,N_20149,N_20048);
or U20317 (N_20317,N_20016,N_20070);
nor U20318 (N_20318,N_20063,N_20104);
and U20319 (N_20319,N_20037,N_20154);
xor U20320 (N_20320,N_20066,N_20013);
nand U20321 (N_20321,N_20140,N_20152);
nor U20322 (N_20322,N_20086,N_20074);
or U20323 (N_20323,N_20139,N_20076);
xor U20324 (N_20324,N_20024,N_20090);
nor U20325 (N_20325,N_20143,N_20010);
nor U20326 (N_20326,N_20059,N_20063);
nor U20327 (N_20327,N_20060,N_20052);
nor U20328 (N_20328,N_20184,N_20186);
nor U20329 (N_20329,N_20158,N_20197);
or U20330 (N_20330,N_20028,N_20129);
and U20331 (N_20331,N_20075,N_20027);
nand U20332 (N_20332,N_20154,N_20086);
or U20333 (N_20333,N_20133,N_20190);
nand U20334 (N_20334,N_20191,N_20076);
xnor U20335 (N_20335,N_20162,N_20192);
and U20336 (N_20336,N_20022,N_20172);
or U20337 (N_20337,N_20121,N_20015);
and U20338 (N_20338,N_20036,N_20048);
nand U20339 (N_20339,N_20055,N_20189);
and U20340 (N_20340,N_20079,N_20039);
nor U20341 (N_20341,N_20057,N_20115);
xnor U20342 (N_20342,N_20152,N_20123);
or U20343 (N_20343,N_20059,N_20055);
and U20344 (N_20344,N_20154,N_20114);
xor U20345 (N_20345,N_20023,N_20189);
nand U20346 (N_20346,N_20087,N_20149);
or U20347 (N_20347,N_20067,N_20172);
xnor U20348 (N_20348,N_20036,N_20044);
nor U20349 (N_20349,N_20133,N_20118);
or U20350 (N_20350,N_20114,N_20081);
nor U20351 (N_20351,N_20130,N_20156);
and U20352 (N_20352,N_20111,N_20083);
or U20353 (N_20353,N_20116,N_20099);
or U20354 (N_20354,N_20131,N_20170);
and U20355 (N_20355,N_20031,N_20024);
or U20356 (N_20356,N_20065,N_20049);
nand U20357 (N_20357,N_20081,N_20171);
or U20358 (N_20358,N_20116,N_20189);
and U20359 (N_20359,N_20095,N_20159);
xor U20360 (N_20360,N_20139,N_20021);
xor U20361 (N_20361,N_20120,N_20179);
nor U20362 (N_20362,N_20019,N_20029);
nand U20363 (N_20363,N_20176,N_20071);
xor U20364 (N_20364,N_20079,N_20154);
nor U20365 (N_20365,N_20024,N_20089);
nor U20366 (N_20366,N_20075,N_20035);
xnor U20367 (N_20367,N_20013,N_20192);
nor U20368 (N_20368,N_20149,N_20097);
nor U20369 (N_20369,N_20063,N_20000);
and U20370 (N_20370,N_20180,N_20024);
and U20371 (N_20371,N_20025,N_20157);
and U20372 (N_20372,N_20166,N_20049);
or U20373 (N_20373,N_20103,N_20136);
or U20374 (N_20374,N_20146,N_20123);
or U20375 (N_20375,N_20178,N_20100);
and U20376 (N_20376,N_20142,N_20184);
xor U20377 (N_20377,N_20112,N_20153);
or U20378 (N_20378,N_20086,N_20077);
or U20379 (N_20379,N_20106,N_20169);
nor U20380 (N_20380,N_20002,N_20028);
and U20381 (N_20381,N_20013,N_20130);
nand U20382 (N_20382,N_20061,N_20057);
and U20383 (N_20383,N_20008,N_20133);
and U20384 (N_20384,N_20161,N_20174);
nor U20385 (N_20385,N_20021,N_20127);
xor U20386 (N_20386,N_20068,N_20061);
xor U20387 (N_20387,N_20149,N_20074);
nor U20388 (N_20388,N_20133,N_20168);
nor U20389 (N_20389,N_20011,N_20069);
nand U20390 (N_20390,N_20165,N_20154);
and U20391 (N_20391,N_20084,N_20120);
xnor U20392 (N_20392,N_20153,N_20020);
xnor U20393 (N_20393,N_20128,N_20166);
or U20394 (N_20394,N_20195,N_20050);
and U20395 (N_20395,N_20019,N_20091);
and U20396 (N_20396,N_20084,N_20042);
xor U20397 (N_20397,N_20064,N_20020);
nand U20398 (N_20398,N_20186,N_20054);
and U20399 (N_20399,N_20179,N_20059);
nand U20400 (N_20400,N_20339,N_20278);
nor U20401 (N_20401,N_20237,N_20342);
xor U20402 (N_20402,N_20272,N_20382);
nand U20403 (N_20403,N_20200,N_20268);
xor U20404 (N_20404,N_20269,N_20258);
xor U20405 (N_20405,N_20201,N_20327);
nor U20406 (N_20406,N_20374,N_20241);
xor U20407 (N_20407,N_20338,N_20210);
and U20408 (N_20408,N_20256,N_20255);
nor U20409 (N_20409,N_20330,N_20251);
xnor U20410 (N_20410,N_20310,N_20261);
xor U20411 (N_20411,N_20383,N_20322);
nand U20412 (N_20412,N_20244,N_20329);
xnor U20413 (N_20413,N_20324,N_20264);
nand U20414 (N_20414,N_20325,N_20347);
or U20415 (N_20415,N_20368,N_20303);
or U20416 (N_20416,N_20289,N_20358);
or U20417 (N_20417,N_20316,N_20217);
nand U20418 (N_20418,N_20290,N_20300);
xnor U20419 (N_20419,N_20213,N_20384);
and U20420 (N_20420,N_20206,N_20355);
nor U20421 (N_20421,N_20248,N_20295);
nand U20422 (N_20422,N_20326,N_20247);
nand U20423 (N_20423,N_20218,N_20238);
and U20424 (N_20424,N_20340,N_20292);
xor U20425 (N_20425,N_20328,N_20380);
or U20426 (N_20426,N_20359,N_20392);
or U20427 (N_20427,N_20275,N_20281);
or U20428 (N_20428,N_20386,N_20335);
or U20429 (N_20429,N_20346,N_20288);
nand U20430 (N_20430,N_20345,N_20271);
xnor U20431 (N_20431,N_20293,N_20318);
xnor U20432 (N_20432,N_20224,N_20398);
or U20433 (N_20433,N_20221,N_20216);
nor U20434 (N_20434,N_20351,N_20262);
or U20435 (N_20435,N_20252,N_20321);
and U20436 (N_20436,N_20387,N_20378);
nand U20437 (N_20437,N_20309,N_20245);
and U20438 (N_20438,N_20302,N_20280);
or U20439 (N_20439,N_20211,N_20394);
and U20440 (N_20440,N_20337,N_20307);
nand U20441 (N_20441,N_20375,N_20323);
and U20442 (N_20442,N_20353,N_20365);
xor U20443 (N_20443,N_20209,N_20389);
and U20444 (N_20444,N_20220,N_20314);
nor U20445 (N_20445,N_20279,N_20265);
and U20446 (N_20446,N_20299,N_20348);
nand U20447 (N_20447,N_20242,N_20230);
nor U20448 (N_20448,N_20363,N_20249);
nand U20449 (N_20449,N_20390,N_20306);
or U20450 (N_20450,N_20219,N_20367);
nor U20451 (N_20451,N_20260,N_20395);
nor U20452 (N_20452,N_20222,N_20225);
and U20453 (N_20453,N_20298,N_20204);
nor U20454 (N_20454,N_20364,N_20385);
or U20455 (N_20455,N_20332,N_20287);
nand U20456 (N_20456,N_20253,N_20239);
or U20457 (N_20457,N_20285,N_20373);
nand U20458 (N_20458,N_20371,N_20313);
or U20459 (N_20459,N_20311,N_20250);
and U20460 (N_20460,N_20208,N_20229);
and U20461 (N_20461,N_20257,N_20254);
nand U20462 (N_20462,N_20240,N_20263);
or U20463 (N_20463,N_20361,N_20274);
or U20464 (N_20464,N_20344,N_20336);
xnor U20465 (N_20465,N_20372,N_20232);
nand U20466 (N_20466,N_20350,N_20354);
xnor U20467 (N_20467,N_20243,N_20388);
xnor U20468 (N_20468,N_20277,N_20282);
xnor U20469 (N_20469,N_20343,N_20369);
nand U20470 (N_20470,N_20319,N_20320);
and U20471 (N_20471,N_20397,N_20223);
nor U20472 (N_20472,N_20334,N_20266);
or U20473 (N_20473,N_20308,N_20270);
and U20474 (N_20474,N_20357,N_20341);
nand U20475 (N_20475,N_20377,N_20370);
and U20476 (N_20476,N_20205,N_20317);
nor U20477 (N_20477,N_20202,N_20284);
nand U20478 (N_20478,N_20333,N_20366);
nor U20479 (N_20479,N_20379,N_20297);
nor U20480 (N_20480,N_20393,N_20376);
or U20481 (N_20481,N_20286,N_20381);
or U20482 (N_20482,N_20267,N_20291);
nand U20483 (N_20483,N_20259,N_20235);
or U20484 (N_20484,N_20349,N_20305);
and U20485 (N_20485,N_20273,N_20315);
nor U20486 (N_20486,N_20231,N_20331);
nand U20487 (N_20487,N_20301,N_20304);
nor U20488 (N_20488,N_20356,N_20294);
or U20489 (N_20489,N_20312,N_20215);
nor U20490 (N_20490,N_20228,N_20276);
or U20491 (N_20491,N_20360,N_20296);
xor U20492 (N_20492,N_20227,N_20362);
or U20493 (N_20493,N_20236,N_20283);
or U20494 (N_20494,N_20246,N_20214);
nor U20495 (N_20495,N_20399,N_20352);
or U20496 (N_20496,N_20233,N_20203);
xnor U20497 (N_20497,N_20226,N_20207);
nor U20498 (N_20498,N_20234,N_20391);
and U20499 (N_20499,N_20396,N_20212);
nor U20500 (N_20500,N_20360,N_20369);
nor U20501 (N_20501,N_20378,N_20336);
nor U20502 (N_20502,N_20341,N_20249);
or U20503 (N_20503,N_20370,N_20313);
xor U20504 (N_20504,N_20360,N_20242);
or U20505 (N_20505,N_20376,N_20294);
xnor U20506 (N_20506,N_20336,N_20316);
and U20507 (N_20507,N_20393,N_20225);
or U20508 (N_20508,N_20322,N_20373);
xnor U20509 (N_20509,N_20239,N_20367);
xor U20510 (N_20510,N_20381,N_20230);
xor U20511 (N_20511,N_20237,N_20263);
nand U20512 (N_20512,N_20348,N_20372);
and U20513 (N_20513,N_20383,N_20305);
or U20514 (N_20514,N_20373,N_20293);
nand U20515 (N_20515,N_20216,N_20372);
and U20516 (N_20516,N_20370,N_20259);
xnor U20517 (N_20517,N_20378,N_20274);
and U20518 (N_20518,N_20219,N_20332);
nand U20519 (N_20519,N_20361,N_20305);
xor U20520 (N_20520,N_20215,N_20375);
and U20521 (N_20521,N_20231,N_20285);
nor U20522 (N_20522,N_20274,N_20349);
or U20523 (N_20523,N_20275,N_20285);
nor U20524 (N_20524,N_20222,N_20296);
or U20525 (N_20525,N_20309,N_20387);
xor U20526 (N_20526,N_20310,N_20223);
nor U20527 (N_20527,N_20217,N_20287);
nand U20528 (N_20528,N_20380,N_20218);
nor U20529 (N_20529,N_20318,N_20253);
and U20530 (N_20530,N_20393,N_20337);
and U20531 (N_20531,N_20309,N_20273);
or U20532 (N_20532,N_20288,N_20318);
or U20533 (N_20533,N_20398,N_20301);
nand U20534 (N_20534,N_20238,N_20253);
nand U20535 (N_20535,N_20202,N_20207);
nand U20536 (N_20536,N_20314,N_20348);
nand U20537 (N_20537,N_20357,N_20259);
xor U20538 (N_20538,N_20345,N_20355);
nand U20539 (N_20539,N_20267,N_20311);
and U20540 (N_20540,N_20294,N_20222);
xor U20541 (N_20541,N_20352,N_20318);
xnor U20542 (N_20542,N_20390,N_20249);
nand U20543 (N_20543,N_20297,N_20247);
or U20544 (N_20544,N_20232,N_20386);
or U20545 (N_20545,N_20260,N_20266);
nand U20546 (N_20546,N_20266,N_20215);
xor U20547 (N_20547,N_20278,N_20241);
nor U20548 (N_20548,N_20282,N_20208);
or U20549 (N_20549,N_20375,N_20227);
nor U20550 (N_20550,N_20359,N_20247);
nand U20551 (N_20551,N_20353,N_20304);
and U20552 (N_20552,N_20342,N_20278);
xor U20553 (N_20553,N_20368,N_20356);
nor U20554 (N_20554,N_20228,N_20239);
nand U20555 (N_20555,N_20383,N_20232);
nand U20556 (N_20556,N_20365,N_20274);
and U20557 (N_20557,N_20283,N_20268);
nor U20558 (N_20558,N_20367,N_20293);
and U20559 (N_20559,N_20293,N_20311);
nand U20560 (N_20560,N_20328,N_20394);
or U20561 (N_20561,N_20238,N_20321);
nor U20562 (N_20562,N_20371,N_20340);
xor U20563 (N_20563,N_20234,N_20332);
nor U20564 (N_20564,N_20397,N_20263);
or U20565 (N_20565,N_20299,N_20217);
or U20566 (N_20566,N_20297,N_20345);
nand U20567 (N_20567,N_20341,N_20244);
or U20568 (N_20568,N_20314,N_20223);
or U20569 (N_20569,N_20221,N_20325);
or U20570 (N_20570,N_20278,N_20273);
nand U20571 (N_20571,N_20358,N_20237);
xor U20572 (N_20572,N_20264,N_20289);
or U20573 (N_20573,N_20287,N_20336);
nand U20574 (N_20574,N_20383,N_20287);
nand U20575 (N_20575,N_20398,N_20239);
and U20576 (N_20576,N_20320,N_20299);
or U20577 (N_20577,N_20360,N_20293);
xor U20578 (N_20578,N_20297,N_20322);
and U20579 (N_20579,N_20245,N_20312);
and U20580 (N_20580,N_20217,N_20236);
xnor U20581 (N_20581,N_20313,N_20257);
xnor U20582 (N_20582,N_20357,N_20249);
nor U20583 (N_20583,N_20292,N_20396);
nor U20584 (N_20584,N_20293,N_20386);
or U20585 (N_20585,N_20360,N_20289);
xor U20586 (N_20586,N_20396,N_20266);
nand U20587 (N_20587,N_20387,N_20238);
or U20588 (N_20588,N_20219,N_20344);
xnor U20589 (N_20589,N_20237,N_20203);
or U20590 (N_20590,N_20302,N_20369);
or U20591 (N_20591,N_20344,N_20246);
nor U20592 (N_20592,N_20239,N_20352);
xnor U20593 (N_20593,N_20358,N_20232);
nand U20594 (N_20594,N_20209,N_20268);
or U20595 (N_20595,N_20239,N_20260);
xor U20596 (N_20596,N_20395,N_20252);
nand U20597 (N_20597,N_20259,N_20298);
xnor U20598 (N_20598,N_20252,N_20287);
xnor U20599 (N_20599,N_20216,N_20368);
or U20600 (N_20600,N_20443,N_20439);
nand U20601 (N_20601,N_20404,N_20543);
xor U20602 (N_20602,N_20533,N_20497);
or U20603 (N_20603,N_20458,N_20590);
xnor U20604 (N_20604,N_20518,N_20504);
nor U20605 (N_20605,N_20547,N_20414);
xnor U20606 (N_20606,N_20452,N_20594);
xor U20607 (N_20607,N_20586,N_20446);
or U20608 (N_20608,N_20480,N_20516);
and U20609 (N_20609,N_20569,N_20402);
nor U20610 (N_20610,N_20420,N_20463);
xor U20611 (N_20611,N_20496,N_20401);
or U20612 (N_20612,N_20503,N_20418);
nand U20613 (N_20613,N_20588,N_20406);
and U20614 (N_20614,N_20474,N_20537);
xnor U20615 (N_20615,N_20527,N_20583);
nand U20616 (N_20616,N_20515,N_20502);
and U20617 (N_20617,N_20541,N_20506);
xor U20618 (N_20618,N_20529,N_20449);
xor U20619 (N_20619,N_20400,N_20520);
and U20620 (N_20620,N_20558,N_20486);
nor U20621 (N_20621,N_20511,N_20563);
and U20622 (N_20622,N_20560,N_20552);
xnor U20623 (N_20623,N_20495,N_20582);
xnor U20624 (N_20624,N_20479,N_20556);
or U20625 (N_20625,N_20501,N_20572);
or U20626 (N_20626,N_20465,N_20491);
nor U20627 (N_20627,N_20514,N_20448);
or U20628 (N_20628,N_20576,N_20468);
or U20629 (N_20629,N_20567,N_20461);
or U20630 (N_20630,N_20460,N_20485);
or U20631 (N_20631,N_20444,N_20554);
nor U20632 (N_20632,N_20492,N_20459);
nor U20633 (N_20633,N_20415,N_20548);
nand U20634 (N_20634,N_20538,N_20507);
nand U20635 (N_20635,N_20544,N_20477);
and U20636 (N_20636,N_20530,N_20573);
nand U20637 (N_20637,N_20591,N_20416);
xor U20638 (N_20638,N_20435,N_20475);
and U20639 (N_20639,N_20542,N_20429);
and U20640 (N_20640,N_20499,N_20578);
xnor U20641 (N_20641,N_20467,N_20412);
or U20642 (N_20642,N_20577,N_20551);
nand U20643 (N_20643,N_20453,N_20483);
and U20644 (N_20644,N_20505,N_20431);
nand U20645 (N_20645,N_20462,N_20419);
xor U20646 (N_20646,N_20596,N_20592);
and U20647 (N_20647,N_20476,N_20433);
nand U20648 (N_20648,N_20424,N_20469);
nand U20649 (N_20649,N_20488,N_20535);
or U20650 (N_20650,N_20528,N_20545);
xor U20651 (N_20651,N_20598,N_20571);
and U20652 (N_20652,N_20482,N_20473);
and U20653 (N_20653,N_20472,N_20490);
or U20654 (N_20654,N_20489,N_20428);
xnor U20655 (N_20655,N_20405,N_20432);
and U20656 (N_20656,N_20534,N_20559);
nand U20657 (N_20657,N_20484,N_20561);
nor U20658 (N_20658,N_20536,N_20539);
xor U20659 (N_20659,N_20442,N_20454);
or U20660 (N_20660,N_20589,N_20521);
xnor U20661 (N_20661,N_20438,N_20456);
nor U20662 (N_20662,N_20519,N_20526);
or U20663 (N_20663,N_20512,N_20427);
nand U20664 (N_20664,N_20532,N_20466);
nor U20665 (N_20665,N_20597,N_20562);
xnor U20666 (N_20666,N_20531,N_20555);
and U20667 (N_20667,N_20430,N_20549);
xor U20668 (N_20668,N_20557,N_20585);
or U20669 (N_20669,N_20524,N_20437);
and U20670 (N_20670,N_20464,N_20426);
nand U20671 (N_20671,N_20408,N_20566);
nand U20672 (N_20672,N_20575,N_20481);
xor U20673 (N_20673,N_20540,N_20421);
and U20674 (N_20674,N_20493,N_20546);
nor U20675 (N_20675,N_20574,N_20525);
xor U20676 (N_20676,N_20471,N_20595);
or U20677 (N_20677,N_20564,N_20593);
nor U20678 (N_20678,N_20550,N_20450);
nand U20679 (N_20679,N_20494,N_20411);
and U20680 (N_20680,N_20510,N_20440);
xor U20681 (N_20681,N_20565,N_20457);
nand U20682 (N_20682,N_20498,N_20425);
nor U20683 (N_20683,N_20417,N_20570);
nand U20684 (N_20684,N_20413,N_20584);
nand U20685 (N_20685,N_20409,N_20423);
or U20686 (N_20686,N_20447,N_20599);
and U20687 (N_20687,N_20522,N_20509);
or U20688 (N_20688,N_20436,N_20434);
or U20689 (N_20689,N_20441,N_20410);
nand U20690 (N_20690,N_20478,N_20451);
nor U20691 (N_20691,N_20422,N_20403);
nand U20692 (N_20692,N_20587,N_20568);
and U20693 (N_20693,N_20470,N_20523);
xnor U20694 (N_20694,N_20553,N_20407);
nor U20695 (N_20695,N_20581,N_20513);
and U20696 (N_20696,N_20500,N_20517);
nor U20697 (N_20697,N_20579,N_20445);
and U20698 (N_20698,N_20580,N_20487);
or U20699 (N_20699,N_20455,N_20508);
and U20700 (N_20700,N_20417,N_20584);
nand U20701 (N_20701,N_20491,N_20576);
and U20702 (N_20702,N_20599,N_20570);
and U20703 (N_20703,N_20583,N_20483);
and U20704 (N_20704,N_20409,N_20541);
nand U20705 (N_20705,N_20401,N_20470);
nor U20706 (N_20706,N_20594,N_20570);
or U20707 (N_20707,N_20565,N_20524);
nand U20708 (N_20708,N_20494,N_20527);
and U20709 (N_20709,N_20555,N_20529);
nor U20710 (N_20710,N_20442,N_20439);
nor U20711 (N_20711,N_20469,N_20479);
or U20712 (N_20712,N_20480,N_20449);
xnor U20713 (N_20713,N_20499,N_20471);
nor U20714 (N_20714,N_20536,N_20572);
or U20715 (N_20715,N_20418,N_20530);
nand U20716 (N_20716,N_20429,N_20482);
nor U20717 (N_20717,N_20493,N_20532);
xor U20718 (N_20718,N_20536,N_20560);
and U20719 (N_20719,N_20527,N_20523);
nor U20720 (N_20720,N_20536,N_20451);
nor U20721 (N_20721,N_20514,N_20443);
nor U20722 (N_20722,N_20588,N_20462);
nor U20723 (N_20723,N_20540,N_20428);
nand U20724 (N_20724,N_20484,N_20512);
nand U20725 (N_20725,N_20487,N_20445);
or U20726 (N_20726,N_20557,N_20412);
nor U20727 (N_20727,N_20501,N_20508);
xnor U20728 (N_20728,N_20483,N_20588);
xor U20729 (N_20729,N_20421,N_20444);
or U20730 (N_20730,N_20460,N_20411);
and U20731 (N_20731,N_20569,N_20479);
or U20732 (N_20732,N_20431,N_20578);
and U20733 (N_20733,N_20449,N_20445);
and U20734 (N_20734,N_20556,N_20568);
xor U20735 (N_20735,N_20409,N_20579);
nand U20736 (N_20736,N_20503,N_20493);
or U20737 (N_20737,N_20472,N_20546);
xnor U20738 (N_20738,N_20531,N_20487);
nor U20739 (N_20739,N_20535,N_20527);
nor U20740 (N_20740,N_20512,N_20522);
or U20741 (N_20741,N_20575,N_20597);
or U20742 (N_20742,N_20508,N_20559);
nand U20743 (N_20743,N_20552,N_20477);
or U20744 (N_20744,N_20491,N_20545);
xor U20745 (N_20745,N_20522,N_20486);
and U20746 (N_20746,N_20546,N_20435);
and U20747 (N_20747,N_20449,N_20538);
and U20748 (N_20748,N_20486,N_20473);
nor U20749 (N_20749,N_20432,N_20551);
or U20750 (N_20750,N_20527,N_20465);
nor U20751 (N_20751,N_20441,N_20455);
nand U20752 (N_20752,N_20488,N_20563);
nand U20753 (N_20753,N_20587,N_20502);
nand U20754 (N_20754,N_20589,N_20572);
and U20755 (N_20755,N_20449,N_20558);
nand U20756 (N_20756,N_20436,N_20451);
nand U20757 (N_20757,N_20589,N_20573);
or U20758 (N_20758,N_20458,N_20485);
nor U20759 (N_20759,N_20551,N_20541);
and U20760 (N_20760,N_20505,N_20443);
or U20761 (N_20761,N_20582,N_20425);
or U20762 (N_20762,N_20582,N_20537);
nor U20763 (N_20763,N_20582,N_20517);
xor U20764 (N_20764,N_20402,N_20465);
xor U20765 (N_20765,N_20533,N_20553);
and U20766 (N_20766,N_20574,N_20470);
nand U20767 (N_20767,N_20425,N_20452);
and U20768 (N_20768,N_20466,N_20562);
nor U20769 (N_20769,N_20452,N_20556);
or U20770 (N_20770,N_20468,N_20401);
nand U20771 (N_20771,N_20571,N_20515);
nand U20772 (N_20772,N_20442,N_20504);
or U20773 (N_20773,N_20451,N_20577);
and U20774 (N_20774,N_20482,N_20460);
nor U20775 (N_20775,N_20420,N_20413);
nor U20776 (N_20776,N_20438,N_20507);
and U20777 (N_20777,N_20415,N_20561);
or U20778 (N_20778,N_20537,N_20465);
xor U20779 (N_20779,N_20496,N_20554);
xor U20780 (N_20780,N_20437,N_20479);
or U20781 (N_20781,N_20523,N_20530);
and U20782 (N_20782,N_20460,N_20586);
or U20783 (N_20783,N_20461,N_20575);
and U20784 (N_20784,N_20465,N_20571);
nor U20785 (N_20785,N_20498,N_20559);
xnor U20786 (N_20786,N_20435,N_20473);
or U20787 (N_20787,N_20417,N_20573);
nor U20788 (N_20788,N_20527,N_20512);
nor U20789 (N_20789,N_20409,N_20470);
and U20790 (N_20790,N_20495,N_20542);
and U20791 (N_20791,N_20498,N_20551);
and U20792 (N_20792,N_20494,N_20534);
xnor U20793 (N_20793,N_20444,N_20437);
xnor U20794 (N_20794,N_20574,N_20469);
nand U20795 (N_20795,N_20403,N_20517);
and U20796 (N_20796,N_20557,N_20492);
nand U20797 (N_20797,N_20402,N_20520);
nand U20798 (N_20798,N_20402,N_20556);
or U20799 (N_20799,N_20454,N_20531);
or U20800 (N_20800,N_20773,N_20689);
or U20801 (N_20801,N_20648,N_20684);
and U20802 (N_20802,N_20683,N_20762);
and U20803 (N_20803,N_20605,N_20701);
nand U20804 (N_20804,N_20677,N_20670);
nand U20805 (N_20805,N_20797,N_20758);
nand U20806 (N_20806,N_20618,N_20766);
nand U20807 (N_20807,N_20749,N_20641);
and U20808 (N_20808,N_20671,N_20777);
or U20809 (N_20809,N_20616,N_20622);
and U20810 (N_20810,N_20698,N_20752);
or U20811 (N_20811,N_20717,N_20647);
nor U20812 (N_20812,N_20632,N_20775);
and U20813 (N_20813,N_20644,N_20761);
xnor U20814 (N_20814,N_20627,N_20780);
or U20815 (N_20815,N_20654,N_20636);
xnor U20816 (N_20816,N_20601,N_20700);
or U20817 (N_20817,N_20722,N_20739);
xnor U20818 (N_20818,N_20721,N_20709);
nand U20819 (N_20819,N_20609,N_20748);
or U20820 (N_20820,N_20634,N_20687);
nor U20821 (N_20821,N_20665,N_20741);
nand U20822 (N_20822,N_20705,N_20681);
nor U20823 (N_20823,N_20637,N_20682);
or U20824 (N_20824,N_20765,N_20695);
and U20825 (N_20825,N_20633,N_20646);
and U20826 (N_20826,N_20694,N_20640);
xor U20827 (N_20827,N_20734,N_20613);
and U20828 (N_20828,N_20661,N_20679);
or U20829 (N_20829,N_20785,N_20638);
nor U20830 (N_20830,N_20685,N_20787);
or U20831 (N_20831,N_20602,N_20617);
and U20832 (N_20832,N_20628,N_20639);
or U20833 (N_20833,N_20743,N_20727);
nand U20834 (N_20834,N_20611,N_20651);
or U20835 (N_20835,N_20754,N_20759);
nand U20836 (N_20836,N_20790,N_20673);
xnor U20837 (N_20837,N_20623,N_20652);
xnor U20838 (N_20838,N_20686,N_20629);
nand U20839 (N_20839,N_20764,N_20658);
nor U20840 (N_20840,N_20799,N_20619);
or U20841 (N_20841,N_20726,N_20653);
or U20842 (N_20842,N_20635,N_20669);
nor U20843 (N_20843,N_20772,N_20767);
xor U20844 (N_20844,N_20704,N_20630);
and U20845 (N_20845,N_20750,N_20776);
nor U20846 (N_20846,N_20731,N_20668);
nor U20847 (N_20847,N_20782,N_20608);
xnor U20848 (N_20848,N_20793,N_20699);
xnor U20849 (N_20849,N_20600,N_20763);
and U20850 (N_20850,N_20707,N_20626);
nand U20851 (N_20851,N_20604,N_20738);
and U20852 (N_20852,N_20783,N_20789);
xnor U20853 (N_20853,N_20737,N_20672);
or U20854 (N_20854,N_20674,N_20693);
nor U20855 (N_20855,N_20794,N_20740);
nand U20856 (N_20856,N_20696,N_20614);
or U20857 (N_20857,N_20656,N_20728);
nor U20858 (N_20858,N_20755,N_20712);
and U20859 (N_20859,N_20798,N_20603);
nand U20860 (N_20860,N_20702,N_20650);
nand U20861 (N_20861,N_20708,N_20713);
or U20862 (N_20862,N_20744,N_20621);
xnor U20863 (N_20863,N_20676,N_20659);
or U20864 (N_20864,N_20706,N_20688);
nor U20865 (N_20865,N_20649,N_20742);
nor U20866 (N_20866,N_20757,N_20725);
xor U20867 (N_20867,N_20723,N_20786);
and U20868 (N_20868,N_20666,N_20733);
nand U20869 (N_20869,N_20747,N_20732);
and U20870 (N_20870,N_20680,N_20642);
xnor U20871 (N_20871,N_20662,N_20664);
xor U20872 (N_20872,N_20631,N_20692);
nor U20873 (N_20873,N_20792,N_20657);
and U20874 (N_20874,N_20612,N_20795);
xnor U20875 (N_20875,N_20730,N_20615);
and U20876 (N_20876,N_20714,N_20751);
nand U20877 (N_20877,N_20796,N_20645);
xnor U20878 (N_20878,N_20724,N_20678);
or U20879 (N_20879,N_20720,N_20655);
xnor U20880 (N_20880,N_20675,N_20756);
nor U20881 (N_20881,N_20778,N_20610);
or U20882 (N_20882,N_20729,N_20736);
nand U20883 (N_20883,N_20769,N_20625);
or U20884 (N_20884,N_20760,N_20753);
and U20885 (N_20885,N_20703,N_20715);
nand U20886 (N_20886,N_20779,N_20768);
and U20887 (N_20887,N_20711,N_20771);
or U20888 (N_20888,N_20774,N_20784);
nand U20889 (N_20889,N_20607,N_20606);
or U20890 (N_20890,N_20745,N_20690);
nand U20891 (N_20891,N_20667,N_20620);
nand U20892 (N_20892,N_20624,N_20781);
nor U20893 (N_20893,N_20710,N_20716);
nor U20894 (N_20894,N_20746,N_20691);
and U20895 (N_20895,N_20791,N_20719);
nand U20896 (N_20896,N_20788,N_20735);
and U20897 (N_20897,N_20718,N_20697);
nand U20898 (N_20898,N_20643,N_20770);
or U20899 (N_20899,N_20663,N_20660);
xnor U20900 (N_20900,N_20730,N_20629);
and U20901 (N_20901,N_20603,N_20700);
or U20902 (N_20902,N_20613,N_20624);
xor U20903 (N_20903,N_20640,N_20765);
and U20904 (N_20904,N_20656,N_20622);
xor U20905 (N_20905,N_20642,N_20643);
and U20906 (N_20906,N_20701,N_20668);
nand U20907 (N_20907,N_20702,N_20645);
nor U20908 (N_20908,N_20734,N_20751);
nand U20909 (N_20909,N_20740,N_20736);
nor U20910 (N_20910,N_20671,N_20775);
nand U20911 (N_20911,N_20768,N_20707);
and U20912 (N_20912,N_20644,N_20777);
nor U20913 (N_20913,N_20647,N_20778);
nor U20914 (N_20914,N_20799,N_20622);
nand U20915 (N_20915,N_20678,N_20778);
xnor U20916 (N_20916,N_20699,N_20605);
nand U20917 (N_20917,N_20789,N_20669);
nor U20918 (N_20918,N_20730,N_20610);
xor U20919 (N_20919,N_20796,N_20683);
and U20920 (N_20920,N_20683,N_20695);
and U20921 (N_20921,N_20650,N_20681);
nor U20922 (N_20922,N_20688,N_20709);
or U20923 (N_20923,N_20607,N_20716);
nand U20924 (N_20924,N_20616,N_20712);
xnor U20925 (N_20925,N_20752,N_20663);
nand U20926 (N_20926,N_20727,N_20720);
nor U20927 (N_20927,N_20652,N_20607);
nand U20928 (N_20928,N_20730,N_20613);
xor U20929 (N_20929,N_20703,N_20716);
xor U20930 (N_20930,N_20616,N_20611);
xnor U20931 (N_20931,N_20625,N_20799);
xnor U20932 (N_20932,N_20688,N_20725);
or U20933 (N_20933,N_20722,N_20737);
nand U20934 (N_20934,N_20764,N_20632);
xor U20935 (N_20935,N_20685,N_20620);
and U20936 (N_20936,N_20691,N_20630);
nand U20937 (N_20937,N_20739,N_20643);
nand U20938 (N_20938,N_20601,N_20733);
nor U20939 (N_20939,N_20688,N_20601);
and U20940 (N_20940,N_20788,N_20638);
and U20941 (N_20941,N_20711,N_20617);
and U20942 (N_20942,N_20754,N_20652);
and U20943 (N_20943,N_20737,N_20723);
xor U20944 (N_20944,N_20667,N_20721);
nand U20945 (N_20945,N_20600,N_20777);
nand U20946 (N_20946,N_20607,N_20661);
nor U20947 (N_20947,N_20760,N_20711);
xor U20948 (N_20948,N_20717,N_20664);
nor U20949 (N_20949,N_20766,N_20702);
or U20950 (N_20950,N_20716,N_20679);
xor U20951 (N_20951,N_20758,N_20743);
xnor U20952 (N_20952,N_20790,N_20728);
and U20953 (N_20953,N_20760,N_20663);
nor U20954 (N_20954,N_20749,N_20704);
nand U20955 (N_20955,N_20774,N_20626);
or U20956 (N_20956,N_20754,N_20628);
nand U20957 (N_20957,N_20670,N_20613);
and U20958 (N_20958,N_20676,N_20724);
or U20959 (N_20959,N_20697,N_20773);
and U20960 (N_20960,N_20735,N_20644);
nor U20961 (N_20961,N_20721,N_20701);
xor U20962 (N_20962,N_20733,N_20614);
nand U20963 (N_20963,N_20625,N_20659);
nand U20964 (N_20964,N_20605,N_20781);
xnor U20965 (N_20965,N_20668,N_20789);
and U20966 (N_20966,N_20704,N_20696);
nor U20967 (N_20967,N_20650,N_20673);
and U20968 (N_20968,N_20747,N_20614);
nor U20969 (N_20969,N_20678,N_20791);
nor U20970 (N_20970,N_20777,N_20676);
xnor U20971 (N_20971,N_20742,N_20743);
and U20972 (N_20972,N_20790,N_20747);
or U20973 (N_20973,N_20751,N_20776);
and U20974 (N_20974,N_20738,N_20633);
and U20975 (N_20975,N_20670,N_20774);
xor U20976 (N_20976,N_20677,N_20767);
nor U20977 (N_20977,N_20780,N_20636);
and U20978 (N_20978,N_20605,N_20686);
nor U20979 (N_20979,N_20624,N_20766);
and U20980 (N_20980,N_20714,N_20788);
nand U20981 (N_20981,N_20784,N_20699);
xor U20982 (N_20982,N_20762,N_20695);
and U20983 (N_20983,N_20679,N_20748);
or U20984 (N_20984,N_20787,N_20762);
and U20985 (N_20985,N_20679,N_20729);
nor U20986 (N_20986,N_20623,N_20665);
or U20987 (N_20987,N_20633,N_20634);
and U20988 (N_20988,N_20769,N_20725);
xor U20989 (N_20989,N_20630,N_20746);
nand U20990 (N_20990,N_20692,N_20610);
xnor U20991 (N_20991,N_20611,N_20708);
nand U20992 (N_20992,N_20707,N_20721);
nand U20993 (N_20993,N_20650,N_20675);
nor U20994 (N_20994,N_20630,N_20780);
and U20995 (N_20995,N_20746,N_20685);
nand U20996 (N_20996,N_20791,N_20619);
nor U20997 (N_20997,N_20652,N_20644);
and U20998 (N_20998,N_20685,N_20674);
xor U20999 (N_20999,N_20745,N_20694);
nor U21000 (N_21000,N_20966,N_20886);
nand U21001 (N_21001,N_20950,N_20839);
xor U21002 (N_21002,N_20980,N_20864);
and U21003 (N_21003,N_20938,N_20865);
nand U21004 (N_21004,N_20885,N_20947);
nand U21005 (N_21005,N_20835,N_20841);
or U21006 (N_21006,N_20853,N_20939);
xnor U21007 (N_21007,N_20895,N_20802);
and U21008 (N_21008,N_20911,N_20876);
nor U21009 (N_21009,N_20951,N_20908);
nor U21010 (N_21010,N_20971,N_20827);
and U21011 (N_21011,N_20994,N_20846);
or U21012 (N_21012,N_20873,N_20910);
nand U21013 (N_21013,N_20817,N_20834);
nand U21014 (N_21014,N_20945,N_20807);
and U21015 (N_21015,N_20992,N_20915);
xor U21016 (N_21016,N_20958,N_20949);
xor U21017 (N_21017,N_20892,N_20869);
or U21018 (N_21018,N_20888,N_20926);
nor U21019 (N_21019,N_20859,N_20815);
and U21020 (N_21020,N_20850,N_20989);
xnor U21021 (N_21021,N_20882,N_20824);
nor U21022 (N_21022,N_20900,N_20964);
or U21023 (N_21023,N_20973,N_20872);
nor U21024 (N_21024,N_20984,N_20821);
xnor U21025 (N_21025,N_20961,N_20906);
nor U21026 (N_21026,N_20852,N_20977);
nand U21027 (N_21027,N_20962,N_20995);
and U21028 (N_21028,N_20952,N_20975);
or U21029 (N_21029,N_20935,N_20828);
or U21030 (N_21030,N_20967,N_20981);
and U21031 (N_21031,N_20861,N_20810);
or U21032 (N_21032,N_20880,N_20940);
nor U21033 (N_21033,N_20843,N_20884);
nor U21034 (N_21034,N_20899,N_20965);
nand U21035 (N_21035,N_20857,N_20878);
xor U21036 (N_21036,N_20946,N_20918);
nand U21037 (N_21037,N_20890,N_20909);
nor U21038 (N_21038,N_20932,N_20806);
nand U21039 (N_21039,N_20985,N_20803);
nand U21040 (N_21040,N_20879,N_20830);
xnor U21041 (N_21041,N_20875,N_20976);
nor U21042 (N_21042,N_20953,N_20905);
and U21043 (N_21043,N_20931,N_20874);
or U21044 (N_21044,N_20826,N_20963);
or U21045 (N_21045,N_20948,N_20901);
or U21046 (N_21046,N_20896,N_20928);
nor U21047 (N_21047,N_20955,N_20829);
xor U21048 (N_21048,N_20999,N_20837);
xor U21049 (N_21049,N_20968,N_20930);
nand U21050 (N_21050,N_20856,N_20912);
xnor U21051 (N_21051,N_20867,N_20816);
and U21052 (N_21052,N_20897,N_20917);
nand U21053 (N_21053,N_20820,N_20929);
xnor U21054 (N_21054,N_20990,N_20954);
xnor U21055 (N_21055,N_20956,N_20972);
nand U21056 (N_21056,N_20894,N_20851);
or U21057 (N_21057,N_20840,N_20836);
or U21058 (N_21058,N_20922,N_20871);
and U21059 (N_21059,N_20848,N_20822);
xor U21060 (N_21060,N_20889,N_20898);
and U21061 (N_21061,N_20914,N_20814);
xor U21062 (N_21062,N_20979,N_20927);
nor U21063 (N_21063,N_20811,N_20863);
or U21064 (N_21064,N_20924,N_20937);
or U21065 (N_21065,N_20855,N_20960);
and U21066 (N_21066,N_20877,N_20969);
and U21067 (N_21067,N_20891,N_20804);
or U21068 (N_21068,N_20903,N_20933);
or U21069 (N_21069,N_20893,N_20832);
xnor U21070 (N_21070,N_20902,N_20849);
xor U21071 (N_21071,N_20854,N_20808);
nor U21072 (N_21072,N_20904,N_20805);
nand U21073 (N_21073,N_20957,N_20858);
or U21074 (N_21074,N_20862,N_20813);
or U21075 (N_21075,N_20988,N_20943);
or U21076 (N_21076,N_20801,N_20860);
nand U21077 (N_21077,N_20818,N_20845);
or U21078 (N_21078,N_20831,N_20944);
nor U21079 (N_21079,N_20998,N_20825);
or U21080 (N_21080,N_20838,N_20983);
nand U21081 (N_21081,N_20974,N_20987);
or U21082 (N_21082,N_20913,N_20833);
xor U21083 (N_21083,N_20934,N_20842);
and U21084 (N_21084,N_20942,N_20916);
nor U21085 (N_21085,N_20887,N_20809);
or U21086 (N_21086,N_20883,N_20978);
or U21087 (N_21087,N_20881,N_20923);
nor U21088 (N_21088,N_20920,N_20907);
and U21089 (N_21089,N_20993,N_20921);
or U21090 (N_21090,N_20996,N_20819);
xnor U21091 (N_21091,N_20866,N_20823);
xor U21092 (N_21092,N_20991,N_20844);
nor U21093 (N_21093,N_20982,N_20986);
xor U21094 (N_21094,N_20868,N_20847);
and U21095 (N_21095,N_20925,N_20800);
and U21096 (N_21096,N_20997,N_20970);
nor U21097 (N_21097,N_20941,N_20959);
or U21098 (N_21098,N_20936,N_20812);
xnor U21099 (N_21099,N_20870,N_20919);
nor U21100 (N_21100,N_20989,N_20846);
nand U21101 (N_21101,N_20977,N_20952);
nand U21102 (N_21102,N_20865,N_20856);
nand U21103 (N_21103,N_20932,N_20984);
nand U21104 (N_21104,N_20968,N_20810);
or U21105 (N_21105,N_20816,N_20931);
xnor U21106 (N_21106,N_20873,N_20935);
or U21107 (N_21107,N_20826,N_20986);
nand U21108 (N_21108,N_20913,N_20995);
xnor U21109 (N_21109,N_20986,N_20856);
nor U21110 (N_21110,N_20958,N_20972);
xor U21111 (N_21111,N_20908,N_20845);
nand U21112 (N_21112,N_20820,N_20914);
nor U21113 (N_21113,N_20876,N_20919);
or U21114 (N_21114,N_20935,N_20926);
and U21115 (N_21115,N_20895,N_20916);
and U21116 (N_21116,N_20973,N_20830);
or U21117 (N_21117,N_20922,N_20943);
and U21118 (N_21118,N_20919,N_20807);
or U21119 (N_21119,N_20895,N_20922);
nor U21120 (N_21120,N_20985,N_20922);
nor U21121 (N_21121,N_20958,N_20861);
nor U21122 (N_21122,N_20980,N_20853);
xnor U21123 (N_21123,N_20952,N_20862);
nor U21124 (N_21124,N_20922,N_20935);
nor U21125 (N_21125,N_20962,N_20887);
nor U21126 (N_21126,N_20908,N_20843);
nor U21127 (N_21127,N_20811,N_20821);
nor U21128 (N_21128,N_20862,N_20979);
and U21129 (N_21129,N_20994,N_20938);
nor U21130 (N_21130,N_20898,N_20864);
nand U21131 (N_21131,N_20800,N_20872);
xor U21132 (N_21132,N_20947,N_20892);
nor U21133 (N_21133,N_20887,N_20831);
nor U21134 (N_21134,N_20859,N_20860);
and U21135 (N_21135,N_20835,N_20964);
or U21136 (N_21136,N_20819,N_20961);
xor U21137 (N_21137,N_20977,N_20916);
xnor U21138 (N_21138,N_20887,N_20942);
nor U21139 (N_21139,N_20975,N_20915);
nor U21140 (N_21140,N_20933,N_20883);
xor U21141 (N_21141,N_20902,N_20955);
nor U21142 (N_21142,N_20986,N_20897);
nor U21143 (N_21143,N_20893,N_20903);
nand U21144 (N_21144,N_20891,N_20862);
nand U21145 (N_21145,N_20985,N_20970);
nand U21146 (N_21146,N_20997,N_20896);
or U21147 (N_21147,N_20999,N_20899);
and U21148 (N_21148,N_20882,N_20931);
nand U21149 (N_21149,N_20826,N_20910);
xor U21150 (N_21150,N_20817,N_20952);
nor U21151 (N_21151,N_20988,N_20992);
nand U21152 (N_21152,N_20998,N_20874);
or U21153 (N_21153,N_20950,N_20967);
nor U21154 (N_21154,N_20903,N_20830);
xnor U21155 (N_21155,N_20877,N_20886);
or U21156 (N_21156,N_20877,N_20912);
and U21157 (N_21157,N_20948,N_20964);
nor U21158 (N_21158,N_20893,N_20840);
xor U21159 (N_21159,N_20923,N_20862);
nor U21160 (N_21160,N_20873,N_20991);
or U21161 (N_21161,N_20989,N_20958);
nand U21162 (N_21162,N_20985,N_20829);
nand U21163 (N_21163,N_20921,N_20932);
or U21164 (N_21164,N_20911,N_20890);
xor U21165 (N_21165,N_20971,N_20958);
or U21166 (N_21166,N_20861,N_20966);
or U21167 (N_21167,N_20812,N_20885);
and U21168 (N_21168,N_20825,N_20970);
and U21169 (N_21169,N_20964,N_20879);
and U21170 (N_21170,N_20991,N_20939);
or U21171 (N_21171,N_20979,N_20958);
or U21172 (N_21172,N_20868,N_20921);
nand U21173 (N_21173,N_20918,N_20915);
xor U21174 (N_21174,N_20819,N_20922);
and U21175 (N_21175,N_20854,N_20983);
nand U21176 (N_21176,N_20893,N_20830);
xnor U21177 (N_21177,N_20989,N_20880);
xor U21178 (N_21178,N_20942,N_20861);
or U21179 (N_21179,N_20874,N_20916);
nor U21180 (N_21180,N_20909,N_20901);
or U21181 (N_21181,N_20808,N_20871);
nor U21182 (N_21182,N_20880,N_20874);
and U21183 (N_21183,N_20906,N_20902);
or U21184 (N_21184,N_20956,N_20902);
nand U21185 (N_21185,N_20978,N_20974);
nand U21186 (N_21186,N_20912,N_20954);
nor U21187 (N_21187,N_20956,N_20927);
nand U21188 (N_21188,N_20861,N_20866);
or U21189 (N_21189,N_20930,N_20956);
nor U21190 (N_21190,N_20871,N_20960);
xor U21191 (N_21191,N_20926,N_20991);
and U21192 (N_21192,N_20844,N_20914);
nor U21193 (N_21193,N_20944,N_20807);
xnor U21194 (N_21194,N_20915,N_20800);
nand U21195 (N_21195,N_20947,N_20845);
nand U21196 (N_21196,N_20888,N_20865);
and U21197 (N_21197,N_20987,N_20964);
and U21198 (N_21198,N_20949,N_20860);
nor U21199 (N_21199,N_20842,N_20880);
nand U21200 (N_21200,N_21147,N_21191);
xnor U21201 (N_21201,N_21032,N_21042);
xnor U21202 (N_21202,N_21016,N_21010);
nor U21203 (N_21203,N_21188,N_21176);
or U21204 (N_21204,N_21094,N_21174);
nor U21205 (N_21205,N_21080,N_21001);
nor U21206 (N_21206,N_21169,N_21096);
nand U21207 (N_21207,N_21167,N_21054);
and U21208 (N_21208,N_21002,N_21053);
nand U21209 (N_21209,N_21089,N_21051);
or U21210 (N_21210,N_21012,N_21024);
nor U21211 (N_21211,N_21112,N_21099);
nor U21212 (N_21212,N_21159,N_21045);
nand U21213 (N_21213,N_21057,N_21088);
and U21214 (N_21214,N_21157,N_21034);
nand U21215 (N_21215,N_21066,N_21003);
or U21216 (N_21216,N_21052,N_21173);
xor U21217 (N_21217,N_21067,N_21150);
nor U21218 (N_21218,N_21193,N_21126);
and U21219 (N_21219,N_21113,N_21171);
nand U21220 (N_21220,N_21058,N_21175);
or U21221 (N_21221,N_21102,N_21185);
nor U21222 (N_21222,N_21164,N_21049);
nor U21223 (N_21223,N_21129,N_21161);
or U21224 (N_21224,N_21124,N_21040);
xnor U21225 (N_21225,N_21120,N_21144);
nor U21226 (N_21226,N_21118,N_21139);
xor U21227 (N_21227,N_21141,N_21026);
nor U21228 (N_21228,N_21182,N_21004);
nand U21229 (N_21229,N_21046,N_21184);
and U21230 (N_21230,N_21162,N_21149);
xnor U21231 (N_21231,N_21166,N_21109);
xor U21232 (N_21232,N_21130,N_21189);
nand U21233 (N_21233,N_21105,N_21068);
and U21234 (N_21234,N_21019,N_21095);
xor U21235 (N_21235,N_21092,N_21047);
or U21236 (N_21236,N_21014,N_21060);
xor U21237 (N_21237,N_21145,N_21000);
xnor U21238 (N_21238,N_21069,N_21114);
or U21239 (N_21239,N_21165,N_21005);
and U21240 (N_21240,N_21097,N_21017);
nand U21241 (N_21241,N_21084,N_21143);
and U21242 (N_21242,N_21076,N_21106);
nand U21243 (N_21243,N_21059,N_21151);
or U21244 (N_21244,N_21025,N_21107);
nor U21245 (N_21245,N_21125,N_21136);
or U21246 (N_21246,N_21072,N_21163);
or U21247 (N_21247,N_21071,N_21091);
and U21248 (N_21248,N_21074,N_21056);
xnor U21249 (N_21249,N_21198,N_21160);
and U21250 (N_21250,N_21044,N_21197);
xor U21251 (N_21251,N_21038,N_21108);
or U21252 (N_21252,N_21152,N_21153);
xnor U21253 (N_21253,N_21148,N_21128);
nand U21254 (N_21254,N_21075,N_21022);
nand U21255 (N_21255,N_21154,N_21135);
and U21256 (N_21256,N_21179,N_21020);
nand U21257 (N_21257,N_21006,N_21023);
or U21258 (N_21258,N_21127,N_21156);
nand U21259 (N_21259,N_21083,N_21008);
xor U21260 (N_21260,N_21142,N_21041);
nand U21261 (N_21261,N_21086,N_21186);
xor U21262 (N_21262,N_21050,N_21085);
nor U21263 (N_21263,N_21048,N_21077);
xnor U21264 (N_21264,N_21015,N_21177);
or U21265 (N_21265,N_21104,N_21007);
and U21266 (N_21266,N_21180,N_21055);
nand U21267 (N_21267,N_21122,N_21115);
nor U21268 (N_21268,N_21009,N_21181);
or U21269 (N_21269,N_21187,N_21013);
or U21270 (N_21270,N_21039,N_21110);
nor U21271 (N_21271,N_21064,N_21146);
xnor U21272 (N_21272,N_21199,N_21100);
xnor U21273 (N_21273,N_21021,N_21116);
or U21274 (N_21274,N_21101,N_21103);
or U21275 (N_21275,N_21037,N_21028);
xor U21276 (N_21276,N_21029,N_21178);
or U21277 (N_21277,N_21192,N_21196);
or U21278 (N_21278,N_21117,N_21168);
nor U21279 (N_21279,N_21121,N_21111);
xnor U21280 (N_21280,N_21081,N_21131);
xor U21281 (N_21281,N_21027,N_21155);
nand U21282 (N_21282,N_21079,N_21030);
nor U21283 (N_21283,N_21158,N_21138);
and U21284 (N_21284,N_21082,N_21035);
xnor U21285 (N_21285,N_21087,N_21033);
nand U21286 (N_21286,N_21093,N_21098);
xor U21287 (N_21287,N_21170,N_21190);
nor U21288 (N_21288,N_21036,N_21070);
nor U21289 (N_21289,N_21133,N_21061);
nand U21290 (N_21290,N_21090,N_21065);
xor U21291 (N_21291,N_21063,N_21018);
nor U21292 (N_21292,N_21183,N_21137);
or U21293 (N_21293,N_21062,N_21172);
or U21294 (N_21294,N_21011,N_21194);
nor U21295 (N_21295,N_21043,N_21031);
or U21296 (N_21296,N_21078,N_21134);
and U21297 (N_21297,N_21195,N_21073);
or U21298 (N_21298,N_21132,N_21119);
and U21299 (N_21299,N_21123,N_21140);
nor U21300 (N_21300,N_21158,N_21187);
and U21301 (N_21301,N_21096,N_21163);
nand U21302 (N_21302,N_21139,N_21077);
nor U21303 (N_21303,N_21146,N_21046);
xnor U21304 (N_21304,N_21075,N_21190);
nor U21305 (N_21305,N_21068,N_21038);
nand U21306 (N_21306,N_21126,N_21097);
nand U21307 (N_21307,N_21061,N_21034);
nor U21308 (N_21308,N_21098,N_21162);
nand U21309 (N_21309,N_21198,N_21029);
and U21310 (N_21310,N_21197,N_21156);
nor U21311 (N_21311,N_21103,N_21086);
and U21312 (N_21312,N_21032,N_21071);
nand U21313 (N_21313,N_21119,N_21189);
or U21314 (N_21314,N_21007,N_21054);
or U21315 (N_21315,N_21186,N_21078);
nor U21316 (N_21316,N_21178,N_21120);
nor U21317 (N_21317,N_21011,N_21141);
or U21318 (N_21318,N_21157,N_21162);
or U21319 (N_21319,N_21133,N_21198);
or U21320 (N_21320,N_21091,N_21144);
xnor U21321 (N_21321,N_21149,N_21159);
or U21322 (N_21322,N_21178,N_21108);
and U21323 (N_21323,N_21056,N_21086);
nand U21324 (N_21324,N_21010,N_21127);
and U21325 (N_21325,N_21186,N_21112);
and U21326 (N_21326,N_21040,N_21047);
and U21327 (N_21327,N_21032,N_21077);
xnor U21328 (N_21328,N_21177,N_21178);
and U21329 (N_21329,N_21044,N_21031);
nor U21330 (N_21330,N_21099,N_21040);
nand U21331 (N_21331,N_21101,N_21097);
xnor U21332 (N_21332,N_21196,N_21082);
nor U21333 (N_21333,N_21157,N_21177);
nor U21334 (N_21334,N_21166,N_21082);
or U21335 (N_21335,N_21183,N_21068);
nand U21336 (N_21336,N_21138,N_21074);
and U21337 (N_21337,N_21125,N_21191);
nand U21338 (N_21338,N_21095,N_21027);
and U21339 (N_21339,N_21177,N_21084);
and U21340 (N_21340,N_21130,N_21158);
or U21341 (N_21341,N_21042,N_21146);
nand U21342 (N_21342,N_21146,N_21126);
nand U21343 (N_21343,N_21118,N_21066);
nand U21344 (N_21344,N_21051,N_21075);
nand U21345 (N_21345,N_21080,N_21020);
or U21346 (N_21346,N_21007,N_21160);
nor U21347 (N_21347,N_21183,N_21096);
nor U21348 (N_21348,N_21118,N_21059);
xor U21349 (N_21349,N_21101,N_21096);
nand U21350 (N_21350,N_21190,N_21150);
nand U21351 (N_21351,N_21082,N_21078);
nand U21352 (N_21352,N_21020,N_21105);
nor U21353 (N_21353,N_21126,N_21076);
and U21354 (N_21354,N_21121,N_21181);
nand U21355 (N_21355,N_21135,N_21169);
nor U21356 (N_21356,N_21187,N_21156);
nor U21357 (N_21357,N_21192,N_21122);
nor U21358 (N_21358,N_21138,N_21160);
nand U21359 (N_21359,N_21103,N_21193);
nand U21360 (N_21360,N_21144,N_21049);
nand U21361 (N_21361,N_21135,N_21012);
nor U21362 (N_21362,N_21099,N_21124);
and U21363 (N_21363,N_21110,N_21123);
xnor U21364 (N_21364,N_21029,N_21031);
and U21365 (N_21365,N_21032,N_21018);
or U21366 (N_21366,N_21068,N_21147);
or U21367 (N_21367,N_21169,N_21065);
and U21368 (N_21368,N_21173,N_21033);
or U21369 (N_21369,N_21176,N_21071);
or U21370 (N_21370,N_21182,N_21184);
nand U21371 (N_21371,N_21067,N_21016);
and U21372 (N_21372,N_21115,N_21119);
or U21373 (N_21373,N_21113,N_21042);
or U21374 (N_21374,N_21023,N_21037);
xnor U21375 (N_21375,N_21123,N_21080);
xor U21376 (N_21376,N_21085,N_21029);
and U21377 (N_21377,N_21189,N_21060);
or U21378 (N_21378,N_21180,N_21116);
or U21379 (N_21379,N_21188,N_21180);
nand U21380 (N_21380,N_21067,N_21095);
nor U21381 (N_21381,N_21120,N_21170);
xor U21382 (N_21382,N_21062,N_21088);
xnor U21383 (N_21383,N_21079,N_21037);
nor U21384 (N_21384,N_21148,N_21055);
nand U21385 (N_21385,N_21167,N_21035);
nand U21386 (N_21386,N_21149,N_21061);
nand U21387 (N_21387,N_21049,N_21186);
or U21388 (N_21388,N_21045,N_21044);
xor U21389 (N_21389,N_21075,N_21045);
and U21390 (N_21390,N_21018,N_21061);
nand U21391 (N_21391,N_21041,N_21068);
nor U21392 (N_21392,N_21092,N_21056);
and U21393 (N_21393,N_21177,N_21075);
nand U21394 (N_21394,N_21000,N_21022);
nand U21395 (N_21395,N_21185,N_21175);
xnor U21396 (N_21396,N_21124,N_21045);
nand U21397 (N_21397,N_21197,N_21126);
and U21398 (N_21398,N_21033,N_21110);
or U21399 (N_21399,N_21003,N_21156);
nand U21400 (N_21400,N_21223,N_21222);
nor U21401 (N_21401,N_21368,N_21208);
nor U21402 (N_21402,N_21270,N_21246);
nand U21403 (N_21403,N_21260,N_21317);
or U21404 (N_21404,N_21243,N_21337);
nor U21405 (N_21405,N_21296,N_21325);
xor U21406 (N_21406,N_21326,N_21218);
nor U21407 (N_21407,N_21248,N_21363);
and U21408 (N_21408,N_21366,N_21341);
or U21409 (N_21409,N_21261,N_21256);
xnor U21410 (N_21410,N_21230,N_21344);
nand U21411 (N_21411,N_21315,N_21276);
or U21412 (N_21412,N_21233,N_21357);
nand U21413 (N_21413,N_21227,N_21397);
nor U21414 (N_21414,N_21356,N_21288);
or U21415 (N_21415,N_21214,N_21347);
and U21416 (N_21416,N_21345,N_21232);
or U21417 (N_21417,N_21310,N_21299);
or U21418 (N_21418,N_21300,N_21352);
nor U21419 (N_21419,N_21239,N_21219);
and U21420 (N_21420,N_21376,N_21245);
nor U21421 (N_21421,N_21302,N_21367);
xor U21422 (N_21422,N_21285,N_21396);
and U21423 (N_21423,N_21277,N_21254);
or U21424 (N_21424,N_21379,N_21200);
nand U21425 (N_21425,N_21330,N_21321);
nor U21426 (N_21426,N_21263,N_21203);
or U21427 (N_21427,N_21377,N_21272);
or U21428 (N_21428,N_21361,N_21206);
xnor U21429 (N_21429,N_21250,N_21381);
or U21430 (N_21430,N_21311,N_21336);
nor U21431 (N_21431,N_21384,N_21268);
and U21432 (N_21432,N_21283,N_21202);
xnor U21433 (N_21433,N_21327,N_21294);
nor U21434 (N_21434,N_21224,N_21324);
xnor U21435 (N_21435,N_21314,N_21213);
nand U21436 (N_21436,N_21284,N_21318);
and U21437 (N_21437,N_21390,N_21343);
nand U21438 (N_21438,N_21398,N_21255);
xnor U21439 (N_21439,N_21328,N_21238);
nor U21440 (N_21440,N_21372,N_21215);
nor U21441 (N_21441,N_21228,N_21333);
nor U21442 (N_21442,N_21349,N_21395);
or U21443 (N_21443,N_21266,N_21293);
or U21444 (N_21444,N_21348,N_21249);
nor U21445 (N_21445,N_21399,N_21295);
nand U21446 (N_21446,N_21275,N_21291);
nor U21447 (N_21447,N_21359,N_21267);
and U21448 (N_21448,N_21350,N_21216);
nor U21449 (N_21449,N_21375,N_21307);
xnor U21450 (N_21450,N_21305,N_21335);
or U21451 (N_21451,N_21242,N_21229);
and U21452 (N_21452,N_21386,N_21286);
and U21453 (N_21453,N_21393,N_21209);
or U21454 (N_21454,N_21306,N_21225);
and U21455 (N_21455,N_21259,N_21378);
xor U21456 (N_21456,N_21388,N_21211);
and U21457 (N_21457,N_21385,N_21308);
xnor U21458 (N_21458,N_21240,N_21370);
nand U21459 (N_21459,N_21226,N_21252);
nand U21460 (N_21460,N_21303,N_21304);
nand U21461 (N_21461,N_21360,N_21392);
nor U21462 (N_21462,N_21292,N_21319);
or U21463 (N_21463,N_21364,N_21323);
xor U21464 (N_21464,N_21358,N_21247);
nand U21465 (N_21465,N_21329,N_21221);
nor U21466 (N_21466,N_21374,N_21234);
xor U21467 (N_21467,N_21301,N_21340);
and U21468 (N_21468,N_21236,N_21281);
and U21469 (N_21469,N_21369,N_21264);
nor U21470 (N_21470,N_21298,N_21273);
or U21471 (N_21471,N_21353,N_21383);
nand U21472 (N_21472,N_21365,N_21237);
nor U21473 (N_21473,N_21279,N_21262);
xor U21474 (N_21474,N_21204,N_21201);
nand U21475 (N_21475,N_21217,N_21338);
nor U21476 (N_21476,N_21331,N_21251);
or U21477 (N_21477,N_21351,N_21362);
and U21478 (N_21478,N_21354,N_21355);
and U21479 (N_21479,N_21282,N_21271);
or U21480 (N_21480,N_21253,N_21207);
nand U21481 (N_21481,N_21231,N_21309);
or U21482 (N_21482,N_21290,N_21339);
or U21483 (N_21483,N_21297,N_21265);
nor U21484 (N_21484,N_21391,N_21320);
or U21485 (N_21485,N_21244,N_21205);
and U21486 (N_21486,N_21235,N_21382);
nor U21487 (N_21487,N_21313,N_21373);
xor U21488 (N_21488,N_21394,N_21278);
or U21489 (N_21489,N_21210,N_21334);
and U21490 (N_21490,N_21322,N_21269);
nand U21491 (N_21491,N_21289,N_21346);
and U21492 (N_21492,N_21387,N_21212);
xnor U21493 (N_21493,N_21274,N_21241);
nor U21494 (N_21494,N_21316,N_21371);
and U21495 (N_21495,N_21389,N_21258);
xor U21496 (N_21496,N_21257,N_21287);
xor U21497 (N_21497,N_21312,N_21220);
or U21498 (N_21498,N_21380,N_21342);
xnor U21499 (N_21499,N_21280,N_21332);
and U21500 (N_21500,N_21205,N_21223);
and U21501 (N_21501,N_21256,N_21303);
or U21502 (N_21502,N_21223,N_21329);
xnor U21503 (N_21503,N_21257,N_21251);
and U21504 (N_21504,N_21291,N_21242);
xnor U21505 (N_21505,N_21365,N_21230);
nand U21506 (N_21506,N_21366,N_21354);
nor U21507 (N_21507,N_21278,N_21241);
nor U21508 (N_21508,N_21337,N_21386);
nand U21509 (N_21509,N_21359,N_21369);
nor U21510 (N_21510,N_21211,N_21265);
nor U21511 (N_21511,N_21244,N_21271);
xnor U21512 (N_21512,N_21369,N_21238);
and U21513 (N_21513,N_21372,N_21274);
nand U21514 (N_21514,N_21354,N_21258);
xor U21515 (N_21515,N_21378,N_21283);
and U21516 (N_21516,N_21268,N_21293);
or U21517 (N_21517,N_21269,N_21214);
and U21518 (N_21518,N_21266,N_21367);
or U21519 (N_21519,N_21289,N_21293);
xor U21520 (N_21520,N_21391,N_21389);
nor U21521 (N_21521,N_21207,N_21209);
xnor U21522 (N_21522,N_21376,N_21346);
or U21523 (N_21523,N_21362,N_21261);
nand U21524 (N_21524,N_21247,N_21291);
xor U21525 (N_21525,N_21349,N_21374);
xnor U21526 (N_21526,N_21218,N_21237);
xor U21527 (N_21527,N_21241,N_21228);
nor U21528 (N_21528,N_21266,N_21256);
or U21529 (N_21529,N_21329,N_21280);
and U21530 (N_21530,N_21365,N_21346);
or U21531 (N_21531,N_21391,N_21250);
nor U21532 (N_21532,N_21243,N_21320);
nand U21533 (N_21533,N_21276,N_21373);
nor U21534 (N_21534,N_21297,N_21347);
or U21535 (N_21535,N_21252,N_21280);
xor U21536 (N_21536,N_21203,N_21239);
nor U21537 (N_21537,N_21257,N_21262);
xor U21538 (N_21538,N_21397,N_21267);
or U21539 (N_21539,N_21201,N_21327);
or U21540 (N_21540,N_21235,N_21259);
xor U21541 (N_21541,N_21303,N_21228);
nand U21542 (N_21542,N_21205,N_21385);
nor U21543 (N_21543,N_21209,N_21208);
or U21544 (N_21544,N_21252,N_21314);
nor U21545 (N_21545,N_21262,N_21204);
and U21546 (N_21546,N_21259,N_21373);
nor U21547 (N_21547,N_21201,N_21371);
xor U21548 (N_21548,N_21245,N_21303);
xnor U21549 (N_21549,N_21237,N_21267);
or U21550 (N_21550,N_21304,N_21368);
nor U21551 (N_21551,N_21394,N_21254);
xnor U21552 (N_21552,N_21201,N_21346);
nor U21553 (N_21553,N_21266,N_21316);
nor U21554 (N_21554,N_21260,N_21202);
or U21555 (N_21555,N_21393,N_21392);
xnor U21556 (N_21556,N_21246,N_21220);
xnor U21557 (N_21557,N_21297,N_21387);
or U21558 (N_21558,N_21301,N_21206);
and U21559 (N_21559,N_21240,N_21342);
and U21560 (N_21560,N_21281,N_21370);
and U21561 (N_21561,N_21271,N_21259);
xor U21562 (N_21562,N_21293,N_21238);
nand U21563 (N_21563,N_21339,N_21298);
or U21564 (N_21564,N_21394,N_21216);
or U21565 (N_21565,N_21205,N_21340);
xnor U21566 (N_21566,N_21286,N_21355);
xnor U21567 (N_21567,N_21272,N_21273);
and U21568 (N_21568,N_21202,N_21324);
xnor U21569 (N_21569,N_21377,N_21311);
nor U21570 (N_21570,N_21322,N_21284);
and U21571 (N_21571,N_21340,N_21203);
nor U21572 (N_21572,N_21306,N_21282);
and U21573 (N_21573,N_21287,N_21211);
nor U21574 (N_21574,N_21283,N_21350);
and U21575 (N_21575,N_21264,N_21331);
and U21576 (N_21576,N_21231,N_21371);
nor U21577 (N_21577,N_21229,N_21237);
nor U21578 (N_21578,N_21398,N_21278);
nor U21579 (N_21579,N_21268,N_21223);
or U21580 (N_21580,N_21371,N_21293);
or U21581 (N_21581,N_21204,N_21295);
or U21582 (N_21582,N_21283,N_21252);
nand U21583 (N_21583,N_21225,N_21325);
and U21584 (N_21584,N_21238,N_21397);
xor U21585 (N_21585,N_21222,N_21332);
xor U21586 (N_21586,N_21397,N_21269);
nor U21587 (N_21587,N_21303,N_21365);
and U21588 (N_21588,N_21206,N_21213);
nand U21589 (N_21589,N_21362,N_21379);
xor U21590 (N_21590,N_21277,N_21342);
or U21591 (N_21591,N_21251,N_21273);
and U21592 (N_21592,N_21299,N_21263);
nor U21593 (N_21593,N_21297,N_21291);
nor U21594 (N_21594,N_21361,N_21372);
nand U21595 (N_21595,N_21369,N_21390);
nand U21596 (N_21596,N_21284,N_21301);
nand U21597 (N_21597,N_21376,N_21285);
nand U21598 (N_21598,N_21304,N_21230);
and U21599 (N_21599,N_21217,N_21254);
nor U21600 (N_21600,N_21486,N_21570);
or U21601 (N_21601,N_21495,N_21494);
or U21602 (N_21602,N_21471,N_21561);
or U21603 (N_21603,N_21594,N_21473);
xnor U21604 (N_21604,N_21425,N_21453);
and U21605 (N_21605,N_21408,N_21563);
nor U21606 (N_21606,N_21510,N_21566);
nor U21607 (N_21607,N_21491,N_21543);
nor U21608 (N_21608,N_21518,N_21550);
nand U21609 (N_21609,N_21411,N_21447);
and U21610 (N_21610,N_21466,N_21525);
and U21611 (N_21611,N_21546,N_21520);
and U21612 (N_21612,N_21435,N_21428);
nand U21613 (N_21613,N_21412,N_21487);
nor U21614 (N_21614,N_21501,N_21574);
and U21615 (N_21615,N_21476,N_21555);
or U21616 (N_21616,N_21492,N_21457);
nor U21617 (N_21617,N_21438,N_21537);
nand U21618 (N_21618,N_21405,N_21461);
nand U21619 (N_21619,N_21533,N_21404);
nor U21620 (N_21620,N_21400,N_21474);
nand U21621 (N_21621,N_21549,N_21464);
nand U21622 (N_21622,N_21415,N_21540);
or U21623 (N_21623,N_21512,N_21436);
nand U21624 (N_21624,N_21517,N_21579);
and U21625 (N_21625,N_21527,N_21523);
nand U21626 (N_21626,N_21449,N_21547);
and U21627 (N_21627,N_21552,N_21452);
nand U21628 (N_21628,N_21556,N_21529);
xor U21629 (N_21629,N_21554,N_21432);
nor U21630 (N_21630,N_21427,N_21401);
xor U21631 (N_21631,N_21562,N_21524);
xor U21632 (N_21632,N_21542,N_21481);
and U21633 (N_21633,N_21541,N_21505);
or U21634 (N_21634,N_21448,N_21484);
xnor U21635 (N_21635,N_21446,N_21493);
nor U21636 (N_21636,N_21515,N_21407);
nor U21637 (N_21637,N_21508,N_21587);
xnor U21638 (N_21638,N_21430,N_21565);
nand U21639 (N_21639,N_21509,N_21483);
or U21640 (N_21640,N_21419,N_21567);
and U21641 (N_21641,N_21409,N_21599);
or U21642 (N_21642,N_21584,N_21454);
nor U21643 (N_21643,N_21580,N_21459);
nor U21644 (N_21644,N_21530,N_21433);
nand U21645 (N_21645,N_21465,N_21504);
or U21646 (N_21646,N_21500,N_21478);
or U21647 (N_21647,N_21536,N_21485);
xnor U21648 (N_21648,N_21531,N_21444);
xnor U21649 (N_21649,N_21560,N_21519);
nand U21650 (N_21650,N_21539,N_21422);
or U21651 (N_21651,N_21403,N_21548);
and U21652 (N_21652,N_21462,N_21467);
and U21653 (N_21653,N_21434,N_21414);
and U21654 (N_21654,N_21589,N_21581);
xor U21655 (N_21655,N_21431,N_21455);
or U21656 (N_21656,N_21424,N_21406);
xnor U21657 (N_21657,N_21490,N_21417);
nor U21658 (N_21658,N_21445,N_21437);
nor U21659 (N_21659,N_21402,N_21586);
nand U21660 (N_21660,N_21582,N_21470);
xnor U21661 (N_21661,N_21513,N_21583);
and U21662 (N_21662,N_21507,N_21571);
xor U21663 (N_21663,N_21469,N_21553);
nor U21664 (N_21664,N_21576,N_21440);
xor U21665 (N_21665,N_21410,N_21593);
and U21666 (N_21666,N_21468,N_21573);
nand U21667 (N_21667,N_21488,N_21585);
xnor U21668 (N_21668,N_21418,N_21559);
xor U21669 (N_21669,N_21456,N_21522);
nand U21670 (N_21670,N_21429,N_21480);
xor U21671 (N_21671,N_21569,N_21572);
and U21672 (N_21672,N_21477,N_21506);
xor U21673 (N_21673,N_21458,N_21597);
and U21674 (N_21674,N_21516,N_21545);
and U21675 (N_21675,N_21590,N_21595);
and U21676 (N_21676,N_21496,N_21578);
nand U21677 (N_21677,N_21534,N_21475);
nand U21678 (N_21678,N_21463,N_21568);
xnor U21679 (N_21679,N_21443,N_21511);
or U21680 (N_21680,N_21538,N_21502);
and U21681 (N_21681,N_21558,N_21420);
or U21682 (N_21682,N_21423,N_21577);
and U21683 (N_21683,N_21441,N_21528);
and U21684 (N_21684,N_21439,N_21551);
or U21685 (N_21685,N_21426,N_21413);
and U21686 (N_21686,N_21575,N_21472);
xnor U21687 (N_21687,N_21588,N_21498);
xnor U21688 (N_21688,N_21526,N_21532);
xnor U21689 (N_21689,N_21499,N_21497);
nor U21690 (N_21690,N_21450,N_21442);
xor U21691 (N_21691,N_21460,N_21479);
and U21692 (N_21692,N_21489,N_21535);
nor U21693 (N_21693,N_21421,N_21592);
xor U21694 (N_21694,N_21544,N_21514);
xor U21695 (N_21695,N_21482,N_21596);
nor U21696 (N_21696,N_21503,N_21564);
and U21697 (N_21697,N_21451,N_21598);
nand U21698 (N_21698,N_21591,N_21521);
nor U21699 (N_21699,N_21416,N_21557);
xnor U21700 (N_21700,N_21590,N_21550);
and U21701 (N_21701,N_21422,N_21467);
or U21702 (N_21702,N_21434,N_21407);
nand U21703 (N_21703,N_21526,N_21454);
or U21704 (N_21704,N_21404,N_21422);
or U21705 (N_21705,N_21495,N_21524);
nor U21706 (N_21706,N_21433,N_21522);
xnor U21707 (N_21707,N_21454,N_21544);
and U21708 (N_21708,N_21540,N_21451);
xnor U21709 (N_21709,N_21574,N_21407);
xnor U21710 (N_21710,N_21422,N_21524);
nor U21711 (N_21711,N_21434,N_21480);
or U21712 (N_21712,N_21405,N_21565);
and U21713 (N_21713,N_21433,N_21540);
nand U21714 (N_21714,N_21536,N_21475);
and U21715 (N_21715,N_21536,N_21505);
and U21716 (N_21716,N_21540,N_21571);
xor U21717 (N_21717,N_21551,N_21544);
nand U21718 (N_21718,N_21437,N_21490);
and U21719 (N_21719,N_21593,N_21482);
xnor U21720 (N_21720,N_21406,N_21551);
nor U21721 (N_21721,N_21592,N_21591);
nand U21722 (N_21722,N_21435,N_21423);
nand U21723 (N_21723,N_21447,N_21517);
and U21724 (N_21724,N_21413,N_21431);
or U21725 (N_21725,N_21429,N_21477);
nand U21726 (N_21726,N_21403,N_21407);
nand U21727 (N_21727,N_21455,N_21402);
nor U21728 (N_21728,N_21436,N_21473);
xor U21729 (N_21729,N_21575,N_21425);
xnor U21730 (N_21730,N_21578,N_21491);
or U21731 (N_21731,N_21418,N_21580);
nor U21732 (N_21732,N_21448,N_21561);
and U21733 (N_21733,N_21520,N_21440);
xor U21734 (N_21734,N_21563,N_21435);
or U21735 (N_21735,N_21475,N_21470);
nor U21736 (N_21736,N_21578,N_21521);
nand U21737 (N_21737,N_21454,N_21561);
and U21738 (N_21738,N_21429,N_21474);
nand U21739 (N_21739,N_21587,N_21535);
xor U21740 (N_21740,N_21590,N_21419);
and U21741 (N_21741,N_21481,N_21419);
and U21742 (N_21742,N_21455,N_21446);
nand U21743 (N_21743,N_21531,N_21540);
nor U21744 (N_21744,N_21522,N_21427);
and U21745 (N_21745,N_21432,N_21461);
xor U21746 (N_21746,N_21407,N_21405);
and U21747 (N_21747,N_21513,N_21501);
nand U21748 (N_21748,N_21466,N_21553);
and U21749 (N_21749,N_21557,N_21587);
nand U21750 (N_21750,N_21457,N_21548);
nand U21751 (N_21751,N_21561,N_21512);
or U21752 (N_21752,N_21530,N_21553);
xnor U21753 (N_21753,N_21538,N_21485);
or U21754 (N_21754,N_21529,N_21548);
xor U21755 (N_21755,N_21438,N_21585);
nand U21756 (N_21756,N_21586,N_21419);
nand U21757 (N_21757,N_21491,N_21573);
or U21758 (N_21758,N_21520,N_21499);
and U21759 (N_21759,N_21439,N_21468);
nand U21760 (N_21760,N_21435,N_21561);
nand U21761 (N_21761,N_21570,N_21537);
or U21762 (N_21762,N_21416,N_21432);
and U21763 (N_21763,N_21471,N_21489);
xnor U21764 (N_21764,N_21573,N_21503);
xor U21765 (N_21765,N_21466,N_21430);
or U21766 (N_21766,N_21578,N_21526);
xor U21767 (N_21767,N_21410,N_21457);
and U21768 (N_21768,N_21550,N_21493);
xnor U21769 (N_21769,N_21421,N_21471);
nand U21770 (N_21770,N_21415,N_21416);
and U21771 (N_21771,N_21534,N_21413);
and U21772 (N_21772,N_21452,N_21523);
nor U21773 (N_21773,N_21572,N_21476);
nand U21774 (N_21774,N_21414,N_21491);
nor U21775 (N_21775,N_21456,N_21532);
nor U21776 (N_21776,N_21484,N_21410);
nand U21777 (N_21777,N_21459,N_21446);
and U21778 (N_21778,N_21434,N_21445);
nor U21779 (N_21779,N_21546,N_21526);
and U21780 (N_21780,N_21579,N_21421);
nand U21781 (N_21781,N_21598,N_21437);
and U21782 (N_21782,N_21428,N_21493);
and U21783 (N_21783,N_21469,N_21547);
nor U21784 (N_21784,N_21418,N_21541);
and U21785 (N_21785,N_21588,N_21471);
nand U21786 (N_21786,N_21413,N_21485);
xor U21787 (N_21787,N_21546,N_21588);
xor U21788 (N_21788,N_21579,N_21401);
or U21789 (N_21789,N_21499,N_21445);
nor U21790 (N_21790,N_21415,N_21446);
xor U21791 (N_21791,N_21561,N_21525);
or U21792 (N_21792,N_21487,N_21420);
or U21793 (N_21793,N_21563,N_21523);
and U21794 (N_21794,N_21581,N_21582);
nand U21795 (N_21795,N_21524,N_21475);
and U21796 (N_21796,N_21400,N_21576);
or U21797 (N_21797,N_21429,N_21440);
and U21798 (N_21798,N_21498,N_21560);
nand U21799 (N_21799,N_21469,N_21419);
and U21800 (N_21800,N_21694,N_21783);
xor U21801 (N_21801,N_21661,N_21691);
and U21802 (N_21802,N_21678,N_21746);
nand U21803 (N_21803,N_21726,N_21735);
nor U21804 (N_21804,N_21625,N_21713);
and U21805 (N_21805,N_21685,N_21698);
and U21806 (N_21806,N_21629,N_21706);
nand U21807 (N_21807,N_21667,N_21631);
nand U21808 (N_21808,N_21637,N_21788);
or U21809 (N_21809,N_21703,N_21708);
xor U21810 (N_21810,N_21707,N_21765);
nand U21811 (N_21811,N_21657,N_21680);
nor U21812 (N_21812,N_21687,N_21797);
nor U21813 (N_21813,N_21792,N_21686);
xnor U21814 (N_21814,N_21697,N_21612);
and U21815 (N_21815,N_21767,N_21776);
nand U21816 (N_21816,N_21790,N_21604);
and U21817 (N_21817,N_21620,N_21681);
xor U21818 (N_21818,N_21768,N_21761);
nor U21819 (N_21819,N_21745,N_21764);
and U21820 (N_21820,N_21702,N_21756);
nand U21821 (N_21821,N_21605,N_21696);
xnor U21822 (N_21822,N_21688,N_21608);
nor U21823 (N_21823,N_21627,N_21616);
and U21824 (N_21824,N_21738,N_21695);
xor U21825 (N_21825,N_21643,N_21613);
nand U21826 (N_21826,N_21789,N_21791);
nor U21827 (N_21827,N_21712,N_21699);
and U21828 (N_21828,N_21720,N_21650);
xor U21829 (N_21829,N_21781,N_21648);
nand U21830 (N_21830,N_21622,N_21607);
nor U21831 (N_21831,N_21749,N_21773);
nand U21832 (N_21832,N_21645,N_21711);
xor U21833 (N_21833,N_21611,N_21615);
or U21834 (N_21834,N_21652,N_21653);
and U21835 (N_21835,N_21617,N_21601);
xor U21836 (N_21836,N_21772,N_21618);
xnor U21837 (N_21837,N_21673,N_21717);
and U21838 (N_21838,N_21668,N_21600);
and U21839 (N_21839,N_21741,N_21744);
nand U21840 (N_21840,N_21610,N_21742);
xor U21841 (N_21841,N_21676,N_21621);
nor U21842 (N_21842,N_21795,N_21736);
nand U21843 (N_21843,N_21662,N_21692);
nor U21844 (N_21844,N_21710,N_21731);
and U21845 (N_21845,N_21727,N_21778);
and U21846 (N_21846,N_21669,N_21665);
or U21847 (N_21847,N_21759,N_21739);
xnor U21848 (N_21848,N_21655,N_21671);
xnor U21849 (N_21849,N_21635,N_21656);
or U21850 (N_21850,N_21684,N_21641);
nor U21851 (N_21851,N_21649,N_21777);
or U21852 (N_21852,N_21628,N_21754);
nand U21853 (N_21853,N_21704,N_21647);
and U21854 (N_21854,N_21760,N_21798);
nand U21855 (N_21855,N_21782,N_21701);
nor U21856 (N_21856,N_21677,N_21624);
nand U21857 (N_21857,N_21793,N_21670);
nand U21858 (N_21858,N_21651,N_21603);
nor U21859 (N_21859,N_21715,N_21762);
xnor U21860 (N_21860,N_21658,N_21747);
nor U21861 (N_21861,N_21728,N_21619);
or U21862 (N_21862,N_21682,N_21757);
nor U21863 (N_21863,N_21716,N_21639);
xnor U21864 (N_21864,N_21733,N_21638);
and U21865 (N_21865,N_21636,N_21700);
or U21866 (N_21866,N_21780,N_21799);
or U21867 (N_21867,N_21609,N_21771);
nand U21868 (N_21868,N_21659,N_21654);
xor U21869 (N_21869,N_21779,N_21614);
nand U21870 (N_21870,N_21748,N_21606);
nand U21871 (N_21871,N_21642,N_21626);
or U21872 (N_21872,N_21689,N_21758);
nand U21873 (N_21873,N_21722,N_21623);
xor U21874 (N_21874,N_21719,N_21709);
xor U21875 (N_21875,N_21725,N_21690);
xor U21876 (N_21876,N_21769,N_21633);
xnor U21877 (N_21877,N_21723,N_21674);
and U21878 (N_21878,N_21786,N_21718);
or U21879 (N_21879,N_21714,N_21740);
xnor U21880 (N_21880,N_21672,N_21660);
and U21881 (N_21881,N_21763,N_21646);
xnor U21882 (N_21882,N_21737,N_21775);
nor U21883 (N_21883,N_21683,N_21732);
and U21884 (N_21884,N_21664,N_21724);
nor U21885 (N_21885,N_21679,N_21785);
xor U21886 (N_21886,N_21634,N_21663);
xnor U21887 (N_21887,N_21766,N_21705);
nand U21888 (N_21888,N_21770,N_21751);
nor U21889 (N_21889,N_21743,N_21729);
and U21890 (N_21890,N_21774,N_21630);
or U21891 (N_21891,N_21794,N_21640);
nor U21892 (N_21892,N_21666,N_21730);
nand U21893 (N_21893,N_21787,N_21632);
xnor U21894 (N_21894,N_21784,N_21752);
or U21895 (N_21895,N_21602,N_21753);
nand U21896 (N_21896,N_21734,N_21644);
and U21897 (N_21897,N_21755,N_21750);
and U21898 (N_21898,N_21721,N_21693);
and U21899 (N_21899,N_21675,N_21796);
xnor U21900 (N_21900,N_21784,N_21602);
or U21901 (N_21901,N_21702,N_21696);
and U21902 (N_21902,N_21638,N_21674);
or U21903 (N_21903,N_21604,N_21642);
or U21904 (N_21904,N_21696,N_21668);
nor U21905 (N_21905,N_21776,N_21746);
xor U21906 (N_21906,N_21679,N_21623);
nand U21907 (N_21907,N_21765,N_21722);
nand U21908 (N_21908,N_21741,N_21757);
nor U21909 (N_21909,N_21700,N_21624);
nor U21910 (N_21910,N_21653,N_21703);
nand U21911 (N_21911,N_21776,N_21690);
nand U21912 (N_21912,N_21700,N_21784);
xor U21913 (N_21913,N_21721,N_21744);
nor U21914 (N_21914,N_21748,N_21613);
and U21915 (N_21915,N_21795,N_21650);
or U21916 (N_21916,N_21779,N_21690);
xor U21917 (N_21917,N_21667,N_21670);
xor U21918 (N_21918,N_21607,N_21782);
nor U21919 (N_21919,N_21668,N_21726);
or U21920 (N_21920,N_21745,N_21677);
xor U21921 (N_21921,N_21658,N_21724);
or U21922 (N_21922,N_21625,N_21768);
xnor U21923 (N_21923,N_21726,N_21643);
xnor U21924 (N_21924,N_21779,N_21731);
or U21925 (N_21925,N_21605,N_21694);
nor U21926 (N_21926,N_21699,N_21713);
or U21927 (N_21927,N_21692,N_21621);
and U21928 (N_21928,N_21656,N_21666);
nor U21929 (N_21929,N_21719,N_21741);
and U21930 (N_21930,N_21744,N_21652);
nand U21931 (N_21931,N_21627,N_21775);
nand U21932 (N_21932,N_21681,N_21708);
xnor U21933 (N_21933,N_21761,N_21626);
xor U21934 (N_21934,N_21767,N_21703);
and U21935 (N_21935,N_21664,N_21624);
nor U21936 (N_21936,N_21768,N_21712);
xor U21937 (N_21937,N_21720,N_21643);
and U21938 (N_21938,N_21792,N_21765);
nand U21939 (N_21939,N_21717,N_21680);
nand U21940 (N_21940,N_21739,N_21681);
nand U21941 (N_21941,N_21692,N_21618);
or U21942 (N_21942,N_21608,N_21709);
and U21943 (N_21943,N_21606,N_21696);
or U21944 (N_21944,N_21746,N_21695);
or U21945 (N_21945,N_21632,N_21739);
or U21946 (N_21946,N_21613,N_21736);
xnor U21947 (N_21947,N_21711,N_21792);
xnor U21948 (N_21948,N_21696,N_21670);
nand U21949 (N_21949,N_21634,N_21717);
xnor U21950 (N_21950,N_21696,N_21763);
or U21951 (N_21951,N_21633,N_21648);
nand U21952 (N_21952,N_21647,N_21670);
or U21953 (N_21953,N_21764,N_21602);
xor U21954 (N_21954,N_21615,N_21640);
xnor U21955 (N_21955,N_21609,N_21781);
nor U21956 (N_21956,N_21733,N_21747);
xnor U21957 (N_21957,N_21740,N_21754);
nand U21958 (N_21958,N_21706,N_21730);
or U21959 (N_21959,N_21766,N_21680);
nor U21960 (N_21960,N_21757,N_21729);
xnor U21961 (N_21961,N_21723,N_21773);
nand U21962 (N_21962,N_21677,N_21714);
and U21963 (N_21963,N_21709,N_21769);
and U21964 (N_21964,N_21605,N_21689);
or U21965 (N_21965,N_21619,N_21675);
and U21966 (N_21966,N_21624,N_21679);
xnor U21967 (N_21967,N_21600,N_21772);
and U21968 (N_21968,N_21628,N_21785);
xor U21969 (N_21969,N_21792,N_21782);
nand U21970 (N_21970,N_21706,N_21788);
or U21971 (N_21971,N_21776,N_21757);
xnor U21972 (N_21972,N_21737,N_21683);
or U21973 (N_21973,N_21786,N_21633);
xnor U21974 (N_21974,N_21692,N_21601);
or U21975 (N_21975,N_21653,N_21776);
xnor U21976 (N_21976,N_21771,N_21766);
and U21977 (N_21977,N_21721,N_21644);
and U21978 (N_21978,N_21743,N_21659);
nor U21979 (N_21979,N_21781,N_21711);
or U21980 (N_21980,N_21634,N_21688);
nor U21981 (N_21981,N_21719,N_21662);
nor U21982 (N_21982,N_21653,N_21637);
xor U21983 (N_21983,N_21761,N_21652);
nand U21984 (N_21984,N_21634,N_21711);
and U21985 (N_21985,N_21689,N_21784);
nand U21986 (N_21986,N_21775,N_21636);
nand U21987 (N_21987,N_21694,N_21657);
or U21988 (N_21988,N_21753,N_21733);
xnor U21989 (N_21989,N_21753,N_21766);
xnor U21990 (N_21990,N_21778,N_21643);
nand U21991 (N_21991,N_21795,N_21622);
xor U21992 (N_21992,N_21610,N_21712);
nor U21993 (N_21993,N_21657,N_21617);
and U21994 (N_21994,N_21648,N_21641);
and U21995 (N_21995,N_21616,N_21770);
and U21996 (N_21996,N_21766,N_21671);
or U21997 (N_21997,N_21726,N_21774);
nand U21998 (N_21998,N_21674,N_21759);
nand U21999 (N_21999,N_21712,N_21640);
and U22000 (N_22000,N_21899,N_21850);
or U22001 (N_22001,N_21979,N_21837);
nor U22002 (N_22002,N_21905,N_21940);
nor U22003 (N_22003,N_21948,N_21961);
and U22004 (N_22004,N_21885,N_21896);
nor U22005 (N_22005,N_21897,N_21879);
xnor U22006 (N_22006,N_21802,N_21860);
and U22007 (N_22007,N_21864,N_21811);
and U22008 (N_22008,N_21992,N_21941);
nor U22009 (N_22009,N_21924,N_21804);
nand U22010 (N_22010,N_21916,N_21982);
or U22011 (N_22011,N_21970,N_21815);
nor U22012 (N_22012,N_21945,N_21892);
nor U22013 (N_22013,N_21848,N_21950);
or U22014 (N_22014,N_21859,N_21981);
and U22015 (N_22015,N_21920,N_21898);
xnor U22016 (N_22016,N_21833,N_21816);
and U22017 (N_22017,N_21968,N_21978);
nand U22018 (N_22018,N_21937,N_21953);
and U22019 (N_22019,N_21952,N_21831);
nor U22020 (N_22020,N_21801,N_21889);
xnor U22021 (N_22021,N_21954,N_21972);
nand U22022 (N_22022,N_21977,N_21825);
and U22023 (N_22023,N_21999,N_21980);
or U22024 (N_22024,N_21910,N_21949);
and U22025 (N_22025,N_21932,N_21975);
and U22026 (N_22026,N_21836,N_21988);
nor U22027 (N_22027,N_21915,N_21935);
or U22028 (N_22028,N_21857,N_21925);
or U22029 (N_22029,N_21913,N_21820);
or U22030 (N_22030,N_21921,N_21883);
nor U22031 (N_22031,N_21822,N_21803);
xnor U22032 (N_22032,N_21839,N_21844);
xor U22033 (N_22033,N_21873,N_21823);
nor U22034 (N_22034,N_21914,N_21918);
or U22035 (N_22035,N_21967,N_21923);
xnor U22036 (N_22036,N_21929,N_21829);
nand U22037 (N_22037,N_21909,N_21907);
and U22038 (N_22038,N_21955,N_21934);
xor U22039 (N_22039,N_21863,N_21989);
or U22040 (N_22040,N_21881,N_21947);
or U22041 (N_22041,N_21997,N_21986);
nand U22042 (N_22042,N_21966,N_21854);
nor U22043 (N_22043,N_21998,N_21846);
and U22044 (N_22044,N_21842,N_21878);
nand U22045 (N_22045,N_21819,N_21812);
and U22046 (N_22046,N_21900,N_21991);
nor U22047 (N_22047,N_21888,N_21845);
and U22048 (N_22048,N_21813,N_21926);
xor U22049 (N_22049,N_21886,N_21867);
xnor U22050 (N_22050,N_21862,N_21903);
and U22051 (N_22051,N_21834,N_21922);
nor U22052 (N_22052,N_21853,N_21957);
xor U22053 (N_22053,N_21895,N_21874);
or U22054 (N_22054,N_21987,N_21818);
nand U22055 (N_22055,N_21993,N_21984);
or U22056 (N_22056,N_21858,N_21866);
nor U22057 (N_22057,N_21884,N_21835);
xor U22058 (N_22058,N_21944,N_21906);
xor U22059 (N_22059,N_21814,N_21958);
xor U22060 (N_22060,N_21807,N_21827);
xnor U22061 (N_22061,N_21928,N_21962);
nand U22062 (N_22062,N_21855,N_21868);
nand U22063 (N_22063,N_21840,N_21865);
nor U22064 (N_22064,N_21927,N_21936);
and U22065 (N_22065,N_21951,N_21912);
nand U22066 (N_22066,N_21956,N_21843);
or U22067 (N_22067,N_21869,N_21974);
nor U22068 (N_22068,N_21852,N_21917);
nor U22069 (N_22069,N_21875,N_21861);
nor U22070 (N_22070,N_21838,N_21849);
nand U22071 (N_22071,N_21938,N_21876);
and U22072 (N_22072,N_21809,N_21810);
xor U22073 (N_22073,N_21805,N_21800);
and U22074 (N_22074,N_21990,N_21960);
and U22075 (N_22075,N_21901,N_21817);
or U22076 (N_22076,N_21872,N_21943);
nand U22077 (N_22077,N_21996,N_21904);
and U22078 (N_22078,N_21902,N_21826);
xor U22079 (N_22079,N_21806,N_21847);
and U22080 (N_22080,N_21891,N_21824);
or U22081 (N_22081,N_21911,N_21828);
and U22082 (N_22082,N_21856,N_21994);
xnor U22083 (N_22083,N_21976,N_21894);
and U22084 (N_22084,N_21851,N_21963);
or U22085 (N_22085,N_21939,N_21882);
and U22086 (N_22086,N_21893,N_21933);
xnor U22087 (N_22087,N_21841,N_21880);
or U22088 (N_22088,N_21871,N_21887);
xnor U22089 (N_22089,N_21890,N_21969);
nor U22090 (N_22090,N_21908,N_21931);
and U22091 (N_22091,N_21946,N_21959);
nand U22092 (N_22092,N_21870,N_21995);
or U22093 (N_22093,N_21919,N_21971);
nand U22094 (N_22094,N_21983,N_21821);
or U22095 (N_22095,N_21808,N_21830);
or U22096 (N_22096,N_21877,N_21973);
or U22097 (N_22097,N_21832,N_21964);
nor U22098 (N_22098,N_21965,N_21985);
nor U22099 (N_22099,N_21930,N_21942);
xor U22100 (N_22100,N_21851,N_21938);
nor U22101 (N_22101,N_21944,N_21876);
nor U22102 (N_22102,N_21941,N_21815);
xnor U22103 (N_22103,N_21949,N_21838);
xor U22104 (N_22104,N_21809,N_21883);
and U22105 (N_22105,N_21942,N_21800);
and U22106 (N_22106,N_21863,N_21876);
and U22107 (N_22107,N_21854,N_21920);
and U22108 (N_22108,N_21956,N_21987);
xnor U22109 (N_22109,N_21849,N_21828);
or U22110 (N_22110,N_21872,N_21880);
and U22111 (N_22111,N_21940,N_21906);
nor U22112 (N_22112,N_21896,N_21838);
or U22113 (N_22113,N_21959,N_21827);
and U22114 (N_22114,N_21856,N_21802);
and U22115 (N_22115,N_21972,N_21812);
or U22116 (N_22116,N_21843,N_21837);
and U22117 (N_22117,N_21813,N_21965);
or U22118 (N_22118,N_21814,N_21807);
nor U22119 (N_22119,N_21824,N_21905);
and U22120 (N_22120,N_21846,N_21949);
and U22121 (N_22121,N_21987,N_21896);
nor U22122 (N_22122,N_21857,N_21801);
nand U22123 (N_22123,N_21802,N_21826);
and U22124 (N_22124,N_21813,N_21838);
nor U22125 (N_22125,N_21997,N_21828);
and U22126 (N_22126,N_21827,N_21900);
or U22127 (N_22127,N_21989,N_21834);
and U22128 (N_22128,N_21879,N_21820);
xnor U22129 (N_22129,N_21925,N_21904);
and U22130 (N_22130,N_21888,N_21934);
xor U22131 (N_22131,N_21938,N_21836);
and U22132 (N_22132,N_21957,N_21955);
or U22133 (N_22133,N_21806,N_21986);
nor U22134 (N_22134,N_21937,N_21988);
nand U22135 (N_22135,N_21929,N_21972);
or U22136 (N_22136,N_21868,N_21938);
nor U22137 (N_22137,N_21900,N_21990);
nand U22138 (N_22138,N_21914,N_21900);
xor U22139 (N_22139,N_21828,N_21921);
or U22140 (N_22140,N_21917,N_21887);
or U22141 (N_22141,N_21811,N_21889);
nand U22142 (N_22142,N_21985,N_21931);
and U22143 (N_22143,N_21951,N_21876);
xnor U22144 (N_22144,N_21925,N_21994);
nand U22145 (N_22145,N_21942,N_21803);
nor U22146 (N_22146,N_21932,N_21858);
nand U22147 (N_22147,N_21988,N_21965);
xor U22148 (N_22148,N_21952,N_21889);
and U22149 (N_22149,N_21837,N_21944);
or U22150 (N_22150,N_21833,N_21805);
xor U22151 (N_22151,N_21932,N_21804);
nand U22152 (N_22152,N_21993,N_21805);
nand U22153 (N_22153,N_21821,N_21930);
nor U22154 (N_22154,N_21997,N_21870);
xnor U22155 (N_22155,N_21972,N_21840);
and U22156 (N_22156,N_21831,N_21809);
and U22157 (N_22157,N_21895,N_21889);
nand U22158 (N_22158,N_21861,N_21847);
xor U22159 (N_22159,N_21975,N_21938);
and U22160 (N_22160,N_21900,N_21956);
nor U22161 (N_22161,N_21915,N_21870);
nand U22162 (N_22162,N_21803,N_21926);
nand U22163 (N_22163,N_21930,N_21972);
nand U22164 (N_22164,N_21807,N_21970);
xor U22165 (N_22165,N_21990,N_21893);
and U22166 (N_22166,N_21903,N_21993);
and U22167 (N_22167,N_21980,N_21928);
xor U22168 (N_22168,N_21932,N_21977);
and U22169 (N_22169,N_21857,N_21949);
and U22170 (N_22170,N_21968,N_21998);
nand U22171 (N_22171,N_21830,N_21990);
xor U22172 (N_22172,N_21903,N_21933);
and U22173 (N_22173,N_21804,N_21898);
or U22174 (N_22174,N_21977,N_21981);
nor U22175 (N_22175,N_21828,N_21978);
nand U22176 (N_22176,N_21823,N_21974);
nor U22177 (N_22177,N_21963,N_21994);
and U22178 (N_22178,N_21815,N_21991);
nor U22179 (N_22179,N_21943,N_21865);
or U22180 (N_22180,N_21903,N_21871);
nand U22181 (N_22181,N_21875,N_21821);
nor U22182 (N_22182,N_21898,N_21826);
xor U22183 (N_22183,N_21820,N_21852);
or U22184 (N_22184,N_21974,N_21906);
xor U22185 (N_22185,N_21820,N_21993);
nor U22186 (N_22186,N_21826,N_21946);
nand U22187 (N_22187,N_21827,N_21902);
or U22188 (N_22188,N_21962,N_21997);
nand U22189 (N_22189,N_21879,N_21885);
and U22190 (N_22190,N_21860,N_21909);
nand U22191 (N_22191,N_21909,N_21984);
xor U22192 (N_22192,N_21901,N_21845);
nor U22193 (N_22193,N_21966,N_21822);
and U22194 (N_22194,N_21867,N_21835);
or U22195 (N_22195,N_21829,N_21946);
and U22196 (N_22196,N_21980,N_21962);
xnor U22197 (N_22197,N_21995,N_21897);
xor U22198 (N_22198,N_21932,N_21829);
nand U22199 (N_22199,N_21907,N_21849);
or U22200 (N_22200,N_22184,N_22065);
nand U22201 (N_22201,N_22025,N_22187);
and U22202 (N_22202,N_22029,N_22108);
and U22203 (N_22203,N_22146,N_22079);
or U22204 (N_22204,N_22027,N_22170);
and U22205 (N_22205,N_22034,N_22111);
or U22206 (N_22206,N_22126,N_22199);
xor U22207 (N_22207,N_22157,N_22072);
xnor U22208 (N_22208,N_22061,N_22008);
nand U22209 (N_22209,N_22002,N_22055);
or U22210 (N_22210,N_22168,N_22054);
xor U22211 (N_22211,N_22151,N_22016);
xnor U22212 (N_22212,N_22032,N_22062);
xnor U22213 (N_22213,N_22039,N_22124);
xor U22214 (N_22214,N_22183,N_22022);
nor U22215 (N_22215,N_22192,N_22005);
nand U22216 (N_22216,N_22070,N_22119);
or U22217 (N_22217,N_22095,N_22182);
xnor U22218 (N_22218,N_22020,N_22118);
or U22219 (N_22219,N_22035,N_22149);
nand U22220 (N_22220,N_22051,N_22046);
or U22221 (N_22221,N_22080,N_22147);
nand U22222 (N_22222,N_22144,N_22197);
and U22223 (N_22223,N_22037,N_22106);
and U22224 (N_22224,N_22099,N_22090);
nand U22225 (N_22225,N_22148,N_22089);
and U22226 (N_22226,N_22073,N_22077);
or U22227 (N_22227,N_22033,N_22057);
or U22228 (N_22228,N_22173,N_22024);
xor U22229 (N_22229,N_22010,N_22139);
nor U22230 (N_22230,N_22094,N_22038);
nor U22231 (N_22231,N_22086,N_22013);
and U22232 (N_22232,N_22175,N_22190);
and U22233 (N_22233,N_22009,N_22114);
and U22234 (N_22234,N_22128,N_22116);
or U22235 (N_22235,N_22004,N_22142);
nor U22236 (N_22236,N_22076,N_22195);
and U22237 (N_22237,N_22171,N_22044);
nand U22238 (N_22238,N_22117,N_22121);
or U22239 (N_22239,N_22011,N_22085);
xnor U22240 (N_22240,N_22166,N_22049);
or U22241 (N_22241,N_22067,N_22075);
or U22242 (N_22242,N_22040,N_22015);
and U22243 (N_22243,N_22084,N_22036);
xnor U22244 (N_22244,N_22135,N_22069);
nand U22245 (N_22245,N_22134,N_22019);
or U22246 (N_22246,N_22056,N_22141);
and U22247 (N_22247,N_22179,N_22045);
or U22248 (N_22248,N_22127,N_22165);
or U22249 (N_22249,N_22007,N_22154);
nor U22250 (N_22250,N_22000,N_22105);
and U22251 (N_22251,N_22041,N_22050);
and U22252 (N_22252,N_22176,N_22001);
nor U22253 (N_22253,N_22006,N_22059);
nor U22254 (N_22254,N_22178,N_22028);
xnor U22255 (N_22255,N_22185,N_22196);
nand U22256 (N_22256,N_22125,N_22091);
xor U22257 (N_22257,N_22064,N_22043);
nor U22258 (N_22258,N_22103,N_22169);
nor U22259 (N_22259,N_22181,N_22058);
and U22260 (N_22260,N_22053,N_22177);
and U22261 (N_22261,N_22145,N_22186);
or U22262 (N_22262,N_22048,N_22140);
nand U22263 (N_22263,N_22068,N_22153);
xor U22264 (N_22264,N_22189,N_22074);
and U22265 (N_22265,N_22021,N_22122);
nor U22266 (N_22266,N_22167,N_22156);
nand U22267 (N_22267,N_22042,N_22012);
xor U22268 (N_22268,N_22123,N_22030);
and U22269 (N_22269,N_22138,N_22160);
nand U22270 (N_22270,N_22152,N_22172);
and U22271 (N_22271,N_22180,N_22096);
and U22272 (N_22272,N_22097,N_22112);
nor U22273 (N_22273,N_22133,N_22159);
and U22274 (N_22274,N_22063,N_22102);
nand U22275 (N_22275,N_22017,N_22081);
and U22276 (N_22276,N_22066,N_22018);
or U22277 (N_22277,N_22060,N_22023);
nand U22278 (N_22278,N_22191,N_22158);
or U22279 (N_22279,N_22143,N_22155);
xnor U22280 (N_22280,N_22164,N_22052);
and U22281 (N_22281,N_22198,N_22193);
nor U22282 (N_22282,N_22078,N_22098);
and U22283 (N_22283,N_22104,N_22188);
nand U22284 (N_22284,N_22163,N_22100);
nand U22285 (N_22285,N_22088,N_22136);
and U22286 (N_22286,N_22101,N_22092);
xor U22287 (N_22287,N_22014,N_22130);
xor U22288 (N_22288,N_22174,N_22132);
and U22289 (N_22289,N_22093,N_22109);
and U22290 (N_22290,N_22162,N_22047);
or U22291 (N_22291,N_22137,N_22131);
nor U22292 (N_22292,N_22026,N_22110);
nand U22293 (N_22293,N_22150,N_22031);
xor U22294 (N_22294,N_22115,N_22003);
or U22295 (N_22295,N_22161,N_22120);
nand U22296 (N_22296,N_22129,N_22082);
or U22297 (N_22297,N_22113,N_22194);
or U22298 (N_22298,N_22071,N_22107);
or U22299 (N_22299,N_22087,N_22083);
nor U22300 (N_22300,N_22104,N_22013);
nor U22301 (N_22301,N_22029,N_22159);
xnor U22302 (N_22302,N_22008,N_22184);
nor U22303 (N_22303,N_22160,N_22145);
or U22304 (N_22304,N_22081,N_22159);
and U22305 (N_22305,N_22101,N_22107);
nand U22306 (N_22306,N_22112,N_22117);
and U22307 (N_22307,N_22068,N_22092);
or U22308 (N_22308,N_22198,N_22178);
nor U22309 (N_22309,N_22028,N_22118);
nand U22310 (N_22310,N_22081,N_22070);
and U22311 (N_22311,N_22180,N_22091);
nor U22312 (N_22312,N_22023,N_22000);
nand U22313 (N_22313,N_22166,N_22188);
nand U22314 (N_22314,N_22170,N_22100);
nor U22315 (N_22315,N_22088,N_22005);
nor U22316 (N_22316,N_22058,N_22143);
or U22317 (N_22317,N_22027,N_22051);
and U22318 (N_22318,N_22148,N_22114);
nand U22319 (N_22319,N_22119,N_22010);
nand U22320 (N_22320,N_22006,N_22069);
and U22321 (N_22321,N_22147,N_22172);
or U22322 (N_22322,N_22019,N_22074);
and U22323 (N_22323,N_22156,N_22161);
or U22324 (N_22324,N_22194,N_22114);
nor U22325 (N_22325,N_22186,N_22106);
and U22326 (N_22326,N_22046,N_22104);
nor U22327 (N_22327,N_22103,N_22032);
nand U22328 (N_22328,N_22118,N_22132);
or U22329 (N_22329,N_22000,N_22135);
or U22330 (N_22330,N_22109,N_22154);
xor U22331 (N_22331,N_22030,N_22067);
and U22332 (N_22332,N_22047,N_22065);
xor U22333 (N_22333,N_22050,N_22140);
or U22334 (N_22334,N_22102,N_22132);
or U22335 (N_22335,N_22106,N_22174);
or U22336 (N_22336,N_22162,N_22006);
and U22337 (N_22337,N_22157,N_22144);
or U22338 (N_22338,N_22075,N_22000);
nor U22339 (N_22339,N_22193,N_22019);
xnor U22340 (N_22340,N_22177,N_22000);
xnor U22341 (N_22341,N_22031,N_22125);
xor U22342 (N_22342,N_22004,N_22199);
and U22343 (N_22343,N_22110,N_22021);
xnor U22344 (N_22344,N_22155,N_22091);
and U22345 (N_22345,N_22185,N_22080);
nand U22346 (N_22346,N_22101,N_22122);
xor U22347 (N_22347,N_22108,N_22175);
nor U22348 (N_22348,N_22124,N_22020);
nor U22349 (N_22349,N_22131,N_22010);
nand U22350 (N_22350,N_22055,N_22030);
and U22351 (N_22351,N_22050,N_22143);
nand U22352 (N_22352,N_22048,N_22155);
nor U22353 (N_22353,N_22120,N_22166);
xnor U22354 (N_22354,N_22113,N_22115);
xor U22355 (N_22355,N_22062,N_22036);
nand U22356 (N_22356,N_22187,N_22012);
nor U22357 (N_22357,N_22130,N_22107);
nor U22358 (N_22358,N_22175,N_22166);
nor U22359 (N_22359,N_22120,N_22104);
and U22360 (N_22360,N_22040,N_22101);
nand U22361 (N_22361,N_22148,N_22122);
nor U22362 (N_22362,N_22050,N_22153);
and U22363 (N_22363,N_22149,N_22033);
and U22364 (N_22364,N_22104,N_22124);
nand U22365 (N_22365,N_22166,N_22131);
xnor U22366 (N_22366,N_22022,N_22075);
or U22367 (N_22367,N_22029,N_22155);
nor U22368 (N_22368,N_22129,N_22111);
xor U22369 (N_22369,N_22007,N_22006);
and U22370 (N_22370,N_22016,N_22013);
and U22371 (N_22371,N_22131,N_22022);
nand U22372 (N_22372,N_22199,N_22081);
nor U22373 (N_22373,N_22183,N_22001);
nand U22374 (N_22374,N_22101,N_22162);
or U22375 (N_22375,N_22091,N_22183);
and U22376 (N_22376,N_22191,N_22155);
nand U22377 (N_22377,N_22194,N_22122);
xor U22378 (N_22378,N_22097,N_22198);
nor U22379 (N_22379,N_22033,N_22056);
and U22380 (N_22380,N_22164,N_22160);
nand U22381 (N_22381,N_22003,N_22051);
and U22382 (N_22382,N_22157,N_22192);
nand U22383 (N_22383,N_22165,N_22020);
xnor U22384 (N_22384,N_22169,N_22137);
and U22385 (N_22385,N_22129,N_22091);
nand U22386 (N_22386,N_22101,N_22064);
nor U22387 (N_22387,N_22048,N_22037);
nand U22388 (N_22388,N_22161,N_22183);
nor U22389 (N_22389,N_22077,N_22184);
and U22390 (N_22390,N_22032,N_22061);
xnor U22391 (N_22391,N_22028,N_22085);
and U22392 (N_22392,N_22195,N_22074);
or U22393 (N_22393,N_22063,N_22025);
nand U22394 (N_22394,N_22145,N_22182);
nand U22395 (N_22395,N_22029,N_22003);
nor U22396 (N_22396,N_22162,N_22089);
xnor U22397 (N_22397,N_22098,N_22008);
nand U22398 (N_22398,N_22125,N_22081);
nor U22399 (N_22399,N_22184,N_22179);
or U22400 (N_22400,N_22217,N_22322);
nand U22401 (N_22401,N_22264,N_22346);
nand U22402 (N_22402,N_22309,N_22221);
or U22403 (N_22403,N_22363,N_22307);
xnor U22404 (N_22404,N_22371,N_22200);
nor U22405 (N_22405,N_22288,N_22302);
nor U22406 (N_22406,N_22215,N_22291);
xor U22407 (N_22407,N_22209,N_22367);
xor U22408 (N_22408,N_22321,N_22252);
xor U22409 (N_22409,N_22207,N_22331);
or U22410 (N_22410,N_22384,N_22206);
xnor U22411 (N_22411,N_22202,N_22389);
xnor U22412 (N_22412,N_22328,N_22324);
xnor U22413 (N_22413,N_22332,N_22292);
and U22414 (N_22414,N_22250,N_22255);
and U22415 (N_22415,N_22240,N_22232);
xnor U22416 (N_22416,N_22238,N_22356);
or U22417 (N_22417,N_22313,N_22201);
xnor U22418 (N_22418,N_22341,N_22380);
nor U22419 (N_22419,N_22224,N_22257);
or U22420 (N_22420,N_22253,N_22355);
nor U22421 (N_22421,N_22325,N_22266);
nand U22422 (N_22422,N_22226,N_22228);
and U22423 (N_22423,N_22282,N_22391);
nand U22424 (N_22424,N_22392,N_22305);
and U22425 (N_22425,N_22373,N_22233);
nor U22426 (N_22426,N_22345,N_22340);
nor U22427 (N_22427,N_22388,N_22230);
nor U22428 (N_22428,N_22204,N_22294);
xor U22429 (N_22429,N_22268,N_22376);
and U22430 (N_22430,N_22378,N_22258);
and U22431 (N_22431,N_22245,N_22386);
or U22432 (N_22432,N_22320,N_22285);
nor U22433 (N_22433,N_22352,N_22335);
nor U22434 (N_22434,N_22286,N_22212);
xor U22435 (N_22435,N_22281,N_22234);
or U22436 (N_22436,N_22348,N_22377);
or U22437 (N_22437,N_22396,N_22398);
xor U22438 (N_22438,N_22360,N_22299);
and U22439 (N_22439,N_22385,N_22354);
xor U22440 (N_22440,N_22370,N_22369);
nor U22441 (N_22441,N_22342,N_22297);
nor U22442 (N_22442,N_22219,N_22275);
nor U22443 (N_22443,N_22210,N_22382);
and U22444 (N_22444,N_22394,N_22225);
xnor U22445 (N_22445,N_22337,N_22277);
and U22446 (N_22446,N_22243,N_22269);
nand U22447 (N_22447,N_22251,N_22375);
or U22448 (N_22448,N_22308,N_22280);
nand U22449 (N_22449,N_22247,N_22312);
xnor U22450 (N_22450,N_22214,N_22372);
and U22451 (N_22451,N_22241,N_22289);
and U22452 (N_22452,N_22290,N_22301);
and U22453 (N_22453,N_22284,N_22274);
or U22454 (N_22454,N_22229,N_22242);
xnor U22455 (N_22455,N_22351,N_22390);
nor U22456 (N_22456,N_22362,N_22383);
or U22457 (N_22457,N_22316,N_22248);
or U22458 (N_22458,N_22237,N_22236);
or U22459 (N_22459,N_22261,N_22319);
xor U22460 (N_22460,N_22374,N_22353);
nor U22461 (N_22461,N_22333,N_22218);
and U22462 (N_22462,N_22216,N_22263);
nor U22463 (N_22463,N_22296,N_22279);
nor U22464 (N_22464,N_22399,N_22349);
and U22465 (N_22465,N_22361,N_22379);
nor U22466 (N_22466,N_22272,N_22256);
and U22467 (N_22467,N_22278,N_22259);
xor U22468 (N_22468,N_22350,N_22213);
xnor U22469 (N_22469,N_22300,N_22395);
and U22470 (N_22470,N_22317,N_22311);
or U22471 (N_22471,N_22271,N_22347);
and U22472 (N_22472,N_22336,N_22323);
nand U22473 (N_22473,N_22365,N_22246);
xnor U22474 (N_22474,N_22303,N_22270);
xnor U22475 (N_22475,N_22273,N_22344);
or U22476 (N_22476,N_22298,N_22220);
and U22477 (N_22477,N_22326,N_22387);
xor U22478 (N_22478,N_22262,N_22235);
nor U22479 (N_22479,N_22358,N_22223);
nand U22480 (N_22480,N_22304,N_22364);
xnor U22481 (N_22481,N_22339,N_22283);
nand U22482 (N_22482,N_22338,N_22276);
nand U22483 (N_22483,N_22295,N_22231);
and U22484 (N_22484,N_22393,N_22310);
nor U22485 (N_22485,N_22357,N_22359);
nand U22486 (N_22486,N_22329,N_22318);
or U22487 (N_22487,N_22287,N_22315);
nand U22488 (N_22488,N_22381,N_22205);
and U22489 (N_22489,N_22249,N_22327);
xor U22490 (N_22490,N_22306,N_22343);
or U22491 (N_22491,N_22265,N_22368);
xor U22492 (N_22492,N_22260,N_22397);
xor U22493 (N_22493,N_22330,N_22222);
or U22494 (N_22494,N_22208,N_22227);
and U22495 (N_22495,N_22267,N_22244);
and U22496 (N_22496,N_22293,N_22334);
nor U22497 (N_22497,N_22254,N_22314);
nor U22498 (N_22498,N_22366,N_22211);
nand U22499 (N_22499,N_22239,N_22203);
xnor U22500 (N_22500,N_22254,N_22258);
nand U22501 (N_22501,N_22274,N_22302);
xnor U22502 (N_22502,N_22254,N_22338);
or U22503 (N_22503,N_22367,N_22370);
and U22504 (N_22504,N_22290,N_22207);
xor U22505 (N_22505,N_22252,N_22308);
or U22506 (N_22506,N_22351,N_22213);
or U22507 (N_22507,N_22364,N_22258);
and U22508 (N_22508,N_22319,N_22386);
nor U22509 (N_22509,N_22243,N_22302);
xnor U22510 (N_22510,N_22321,N_22309);
nor U22511 (N_22511,N_22210,N_22261);
xor U22512 (N_22512,N_22256,N_22209);
nand U22513 (N_22513,N_22283,N_22338);
nand U22514 (N_22514,N_22209,N_22265);
xnor U22515 (N_22515,N_22292,N_22339);
nand U22516 (N_22516,N_22283,N_22368);
nand U22517 (N_22517,N_22207,N_22347);
nor U22518 (N_22518,N_22316,N_22302);
xor U22519 (N_22519,N_22271,N_22358);
xnor U22520 (N_22520,N_22237,N_22365);
nor U22521 (N_22521,N_22357,N_22306);
nor U22522 (N_22522,N_22213,N_22397);
nand U22523 (N_22523,N_22337,N_22363);
nor U22524 (N_22524,N_22260,N_22222);
and U22525 (N_22525,N_22302,N_22371);
nand U22526 (N_22526,N_22269,N_22249);
xor U22527 (N_22527,N_22235,N_22202);
nor U22528 (N_22528,N_22309,N_22357);
xnor U22529 (N_22529,N_22260,N_22327);
nand U22530 (N_22530,N_22272,N_22303);
and U22531 (N_22531,N_22383,N_22254);
or U22532 (N_22532,N_22222,N_22240);
nor U22533 (N_22533,N_22392,N_22205);
nor U22534 (N_22534,N_22329,N_22240);
nand U22535 (N_22535,N_22227,N_22380);
and U22536 (N_22536,N_22226,N_22243);
nand U22537 (N_22537,N_22279,N_22396);
xor U22538 (N_22538,N_22382,N_22365);
xor U22539 (N_22539,N_22357,N_22380);
or U22540 (N_22540,N_22267,N_22264);
or U22541 (N_22541,N_22354,N_22329);
nor U22542 (N_22542,N_22346,N_22331);
and U22543 (N_22543,N_22367,N_22371);
and U22544 (N_22544,N_22275,N_22242);
nor U22545 (N_22545,N_22326,N_22301);
nand U22546 (N_22546,N_22367,N_22294);
nand U22547 (N_22547,N_22251,N_22370);
nand U22548 (N_22548,N_22315,N_22225);
nand U22549 (N_22549,N_22263,N_22341);
xnor U22550 (N_22550,N_22216,N_22328);
or U22551 (N_22551,N_22323,N_22230);
and U22552 (N_22552,N_22367,N_22368);
nand U22553 (N_22553,N_22269,N_22299);
nor U22554 (N_22554,N_22376,N_22365);
and U22555 (N_22555,N_22355,N_22286);
xor U22556 (N_22556,N_22380,N_22368);
xnor U22557 (N_22557,N_22248,N_22300);
or U22558 (N_22558,N_22294,N_22356);
nand U22559 (N_22559,N_22298,N_22247);
nand U22560 (N_22560,N_22396,N_22395);
and U22561 (N_22561,N_22363,N_22259);
xor U22562 (N_22562,N_22212,N_22255);
nor U22563 (N_22563,N_22314,N_22307);
or U22564 (N_22564,N_22208,N_22216);
nand U22565 (N_22565,N_22259,N_22354);
nor U22566 (N_22566,N_22328,N_22268);
nand U22567 (N_22567,N_22386,N_22343);
nor U22568 (N_22568,N_22337,N_22350);
xnor U22569 (N_22569,N_22374,N_22388);
nand U22570 (N_22570,N_22360,N_22206);
xnor U22571 (N_22571,N_22394,N_22329);
and U22572 (N_22572,N_22381,N_22306);
and U22573 (N_22573,N_22307,N_22217);
nand U22574 (N_22574,N_22226,N_22260);
and U22575 (N_22575,N_22265,N_22260);
nand U22576 (N_22576,N_22372,N_22235);
and U22577 (N_22577,N_22330,N_22317);
or U22578 (N_22578,N_22359,N_22324);
or U22579 (N_22579,N_22215,N_22294);
and U22580 (N_22580,N_22250,N_22301);
or U22581 (N_22581,N_22230,N_22215);
nand U22582 (N_22582,N_22251,N_22207);
nor U22583 (N_22583,N_22263,N_22323);
nor U22584 (N_22584,N_22268,N_22339);
and U22585 (N_22585,N_22338,N_22343);
and U22586 (N_22586,N_22332,N_22320);
nor U22587 (N_22587,N_22354,N_22363);
and U22588 (N_22588,N_22395,N_22317);
or U22589 (N_22589,N_22216,N_22237);
or U22590 (N_22590,N_22332,N_22263);
nand U22591 (N_22591,N_22306,N_22211);
nand U22592 (N_22592,N_22381,N_22395);
xnor U22593 (N_22593,N_22239,N_22240);
nor U22594 (N_22594,N_22254,N_22362);
nand U22595 (N_22595,N_22307,N_22341);
and U22596 (N_22596,N_22395,N_22252);
xor U22597 (N_22597,N_22347,N_22300);
and U22598 (N_22598,N_22290,N_22361);
xnor U22599 (N_22599,N_22392,N_22309);
nor U22600 (N_22600,N_22404,N_22489);
nor U22601 (N_22601,N_22565,N_22571);
nor U22602 (N_22602,N_22563,N_22487);
nand U22603 (N_22603,N_22468,N_22510);
xor U22604 (N_22604,N_22409,N_22435);
or U22605 (N_22605,N_22470,N_22538);
nor U22606 (N_22606,N_22588,N_22596);
or U22607 (N_22607,N_22570,N_22480);
or U22608 (N_22608,N_22533,N_22449);
nor U22609 (N_22609,N_22436,N_22530);
nand U22610 (N_22610,N_22467,N_22513);
nor U22611 (N_22611,N_22521,N_22502);
nand U22612 (N_22612,N_22592,N_22417);
and U22613 (N_22613,N_22434,N_22514);
nor U22614 (N_22614,N_22483,N_22526);
nand U22615 (N_22615,N_22549,N_22460);
nand U22616 (N_22616,N_22454,N_22472);
and U22617 (N_22617,N_22585,N_22474);
nor U22618 (N_22618,N_22567,N_22503);
nand U22619 (N_22619,N_22442,N_22437);
nor U22620 (N_22620,N_22402,N_22425);
and U22621 (N_22621,N_22481,N_22581);
nand U22622 (N_22622,N_22452,N_22583);
nor U22623 (N_22623,N_22555,N_22414);
and U22624 (N_22624,N_22426,N_22575);
or U22625 (N_22625,N_22457,N_22546);
nand U22626 (N_22626,N_22529,N_22589);
nand U22627 (N_22627,N_22462,N_22450);
nand U22628 (N_22628,N_22422,N_22443);
nand U22629 (N_22629,N_22445,N_22542);
and U22630 (N_22630,N_22478,N_22586);
nor U22631 (N_22631,N_22518,N_22578);
nor U22632 (N_22632,N_22593,N_22492);
xor U22633 (N_22633,N_22576,N_22441);
and U22634 (N_22634,N_22531,N_22459);
xnor U22635 (N_22635,N_22495,N_22523);
or U22636 (N_22636,N_22537,N_22559);
xor U22637 (N_22637,N_22562,N_22534);
xnor U22638 (N_22638,N_22564,N_22451);
or U22639 (N_22639,N_22488,N_22594);
xor U22640 (N_22640,N_22591,N_22477);
xor U22641 (N_22641,N_22572,N_22547);
and U22642 (N_22642,N_22541,N_22520);
nand U22643 (N_22643,N_22551,N_22558);
or U22644 (N_22644,N_22496,N_22515);
or U22645 (N_22645,N_22401,N_22427);
and U22646 (N_22646,N_22507,N_22482);
and U22647 (N_22647,N_22582,N_22550);
and U22648 (N_22648,N_22439,N_22506);
nand U22649 (N_22649,N_22539,N_22476);
nor U22650 (N_22650,N_22473,N_22519);
nor U22651 (N_22651,N_22509,N_22553);
or U22652 (N_22652,N_22556,N_22440);
or U22653 (N_22653,N_22577,N_22403);
or U22654 (N_22654,N_22433,N_22464);
xnor U22655 (N_22655,N_22566,N_22438);
xor U22656 (N_22656,N_22432,N_22552);
nor U22657 (N_22657,N_22536,N_22423);
xnor U22658 (N_22658,N_22497,N_22505);
nand U22659 (N_22659,N_22524,N_22516);
nor U22660 (N_22660,N_22499,N_22574);
xor U22661 (N_22661,N_22498,N_22557);
nand U22662 (N_22662,N_22418,N_22453);
nand U22663 (N_22663,N_22479,N_22421);
or U22664 (N_22664,N_22416,N_22508);
xor U22665 (N_22665,N_22579,N_22522);
and U22666 (N_22666,N_22599,N_22412);
xor U22667 (N_22667,N_22527,N_22517);
nor U22668 (N_22668,N_22420,N_22463);
nand U22669 (N_22669,N_22548,N_22466);
xnor U22670 (N_22670,N_22447,N_22590);
xor U22671 (N_22671,N_22587,N_22475);
and U22672 (N_22672,N_22573,N_22408);
or U22673 (N_22673,N_22569,N_22400);
or U22674 (N_22674,N_22428,N_22511);
or U22675 (N_22675,N_22544,N_22532);
xnor U22676 (N_22676,N_22410,N_22407);
nand U22677 (N_22677,N_22415,N_22484);
or U22678 (N_22678,N_22528,N_22561);
and U22679 (N_22679,N_22491,N_22545);
xor U22680 (N_22680,N_22455,N_22543);
nor U22681 (N_22681,N_22444,N_22456);
xor U22682 (N_22682,N_22448,N_22406);
nor U22683 (N_22683,N_22419,N_22430);
and U22684 (N_22684,N_22446,N_22525);
or U22685 (N_22685,N_22429,N_22431);
xor U22686 (N_22686,N_22512,N_22595);
nand U22687 (N_22687,N_22411,N_22493);
or U22688 (N_22688,N_22461,N_22405);
xor U22689 (N_22689,N_22597,N_22580);
xor U22690 (N_22690,N_22494,N_22535);
and U22691 (N_22691,N_22501,N_22554);
or U22692 (N_22692,N_22540,N_22584);
nor U22693 (N_22693,N_22458,N_22471);
nand U22694 (N_22694,N_22485,N_22413);
nand U22695 (N_22695,N_22490,N_22424);
nand U22696 (N_22696,N_22469,N_22598);
and U22697 (N_22697,N_22500,N_22504);
nor U22698 (N_22698,N_22465,N_22486);
nor U22699 (N_22699,N_22560,N_22568);
nor U22700 (N_22700,N_22593,N_22539);
and U22701 (N_22701,N_22498,N_22534);
xnor U22702 (N_22702,N_22425,N_22429);
nor U22703 (N_22703,N_22534,N_22568);
nand U22704 (N_22704,N_22568,N_22574);
nand U22705 (N_22705,N_22452,N_22438);
and U22706 (N_22706,N_22553,N_22457);
nor U22707 (N_22707,N_22506,N_22509);
nand U22708 (N_22708,N_22434,N_22485);
nor U22709 (N_22709,N_22529,N_22535);
xor U22710 (N_22710,N_22466,N_22546);
nand U22711 (N_22711,N_22528,N_22511);
xnor U22712 (N_22712,N_22548,N_22589);
and U22713 (N_22713,N_22598,N_22459);
and U22714 (N_22714,N_22585,N_22406);
xnor U22715 (N_22715,N_22463,N_22413);
xor U22716 (N_22716,N_22563,N_22585);
nand U22717 (N_22717,N_22492,N_22468);
and U22718 (N_22718,N_22550,N_22421);
or U22719 (N_22719,N_22592,N_22476);
nand U22720 (N_22720,N_22575,N_22480);
and U22721 (N_22721,N_22458,N_22526);
xor U22722 (N_22722,N_22499,N_22409);
and U22723 (N_22723,N_22440,N_22489);
xnor U22724 (N_22724,N_22551,N_22423);
or U22725 (N_22725,N_22532,N_22414);
nand U22726 (N_22726,N_22408,N_22516);
and U22727 (N_22727,N_22504,N_22573);
nor U22728 (N_22728,N_22468,N_22454);
and U22729 (N_22729,N_22596,N_22501);
or U22730 (N_22730,N_22582,N_22518);
nor U22731 (N_22731,N_22440,N_22414);
nand U22732 (N_22732,N_22434,N_22551);
and U22733 (N_22733,N_22494,N_22538);
xor U22734 (N_22734,N_22447,N_22473);
xor U22735 (N_22735,N_22581,N_22439);
nand U22736 (N_22736,N_22598,N_22512);
nor U22737 (N_22737,N_22404,N_22518);
nand U22738 (N_22738,N_22517,N_22553);
xnor U22739 (N_22739,N_22509,N_22590);
nand U22740 (N_22740,N_22597,N_22401);
and U22741 (N_22741,N_22578,N_22408);
and U22742 (N_22742,N_22462,N_22503);
nor U22743 (N_22743,N_22522,N_22598);
xnor U22744 (N_22744,N_22438,N_22561);
nand U22745 (N_22745,N_22523,N_22580);
nor U22746 (N_22746,N_22520,N_22461);
xnor U22747 (N_22747,N_22505,N_22424);
nand U22748 (N_22748,N_22535,N_22584);
xnor U22749 (N_22749,N_22446,N_22465);
nand U22750 (N_22750,N_22505,N_22487);
nor U22751 (N_22751,N_22465,N_22440);
nand U22752 (N_22752,N_22559,N_22567);
or U22753 (N_22753,N_22535,N_22590);
or U22754 (N_22754,N_22488,N_22521);
nand U22755 (N_22755,N_22543,N_22528);
or U22756 (N_22756,N_22476,N_22434);
nor U22757 (N_22757,N_22596,N_22493);
xnor U22758 (N_22758,N_22499,N_22406);
nor U22759 (N_22759,N_22554,N_22429);
or U22760 (N_22760,N_22488,N_22575);
xor U22761 (N_22761,N_22525,N_22476);
xnor U22762 (N_22762,N_22435,N_22438);
and U22763 (N_22763,N_22592,N_22461);
xor U22764 (N_22764,N_22529,N_22519);
or U22765 (N_22765,N_22561,N_22475);
and U22766 (N_22766,N_22515,N_22516);
or U22767 (N_22767,N_22595,N_22467);
xor U22768 (N_22768,N_22475,N_22541);
xnor U22769 (N_22769,N_22483,N_22480);
nand U22770 (N_22770,N_22403,N_22472);
nor U22771 (N_22771,N_22518,N_22510);
xor U22772 (N_22772,N_22430,N_22411);
nor U22773 (N_22773,N_22517,N_22409);
and U22774 (N_22774,N_22569,N_22490);
xnor U22775 (N_22775,N_22538,N_22439);
nor U22776 (N_22776,N_22403,N_22412);
or U22777 (N_22777,N_22532,N_22599);
and U22778 (N_22778,N_22413,N_22570);
nand U22779 (N_22779,N_22421,N_22405);
or U22780 (N_22780,N_22443,N_22475);
xnor U22781 (N_22781,N_22474,N_22524);
and U22782 (N_22782,N_22516,N_22534);
and U22783 (N_22783,N_22494,N_22482);
or U22784 (N_22784,N_22509,N_22558);
or U22785 (N_22785,N_22571,N_22414);
nor U22786 (N_22786,N_22430,N_22493);
or U22787 (N_22787,N_22511,N_22446);
xor U22788 (N_22788,N_22551,N_22413);
nand U22789 (N_22789,N_22468,N_22509);
or U22790 (N_22790,N_22485,N_22565);
nor U22791 (N_22791,N_22569,N_22501);
and U22792 (N_22792,N_22482,N_22510);
and U22793 (N_22793,N_22528,N_22404);
xor U22794 (N_22794,N_22414,N_22591);
or U22795 (N_22795,N_22578,N_22562);
xnor U22796 (N_22796,N_22401,N_22469);
or U22797 (N_22797,N_22534,N_22514);
nor U22798 (N_22798,N_22531,N_22574);
nor U22799 (N_22799,N_22426,N_22401);
nand U22800 (N_22800,N_22743,N_22710);
nand U22801 (N_22801,N_22745,N_22796);
xor U22802 (N_22802,N_22618,N_22721);
or U22803 (N_22803,N_22601,N_22769);
nand U22804 (N_22804,N_22623,N_22643);
or U22805 (N_22805,N_22685,N_22666);
and U22806 (N_22806,N_22770,N_22642);
nor U22807 (N_22807,N_22787,N_22621);
nor U22808 (N_22808,N_22698,N_22789);
xnor U22809 (N_22809,N_22764,N_22793);
and U22810 (N_22810,N_22779,N_22727);
nand U22811 (N_22811,N_22628,N_22708);
nor U22812 (N_22812,N_22772,N_22794);
nand U22813 (N_22813,N_22672,N_22693);
nand U22814 (N_22814,N_22649,N_22695);
nand U22815 (N_22815,N_22748,N_22603);
or U22816 (N_22816,N_22783,N_22722);
nor U22817 (N_22817,N_22737,N_22647);
or U22818 (N_22818,N_22690,N_22646);
or U22819 (N_22819,N_22637,N_22683);
nand U22820 (N_22820,N_22633,N_22746);
nand U22821 (N_22821,N_22624,N_22765);
and U22822 (N_22822,N_22723,N_22728);
or U22823 (N_22823,N_22788,N_22679);
or U22824 (N_22824,N_22711,N_22687);
or U22825 (N_22825,N_22724,N_22717);
and U22826 (N_22826,N_22620,N_22701);
xnor U22827 (N_22827,N_22634,N_22671);
or U22828 (N_22828,N_22640,N_22712);
nor U22829 (N_22829,N_22753,N_22689);
xnor U22830 (N_22830,N_22656,N_22664);
or U22831 (N_22831,N_22696,N_22714);
nand U22832 (N_22832,N_22617,N_22715);
xor U22833 (N_22833,N_22631,N_22729);
nor U22834 (N_22834,N_22720,N_22627);
nor U22835 (N_22835,N_22704,N_22638);
xnor U22836 (N_22836,N_22738,N_22609);
and U22837 (N_22837,N_22659,N_22725);
xor U22838 (N_22838,N_22706,N_22673);
nand U22839 (N_22839,N_22686,N_22670);
xnor U22840 (N_22840,N_22692,N_22668);
or U22841 (N_22841,N_22739,N_22755);
or U22842 (N_22842,N_22660,N_22699);
nand U22843 (N_22843,N_22632,N_22775);
or U22844 (N_22844,N_22785,N_22616);
nor U22845 (N_22845,N_22709,N_22636);
nand U22846 (N_22846,N_22754,N_22655);
and U22847 (N_22847,N_22726,N_22758);
nor U22848 (N_22848,N_22768,N_22602);
and U22849 (N_22849,N_22781,N_22639);
nand U22850 (N_22850,N_22661,N_22719);
nand U22851 (N_22851,N_22799,N_22736);
or U22852 (N_22852,N_22644,N_22707);
nand U22853 (N_22853,N_22742,N_22676);
or U22854 (N_22854,N_22648,N_22763);
and U22855 (N_22855,N_22607,N_22650);
nand U22856 (N_22856,N_22790,N_22741);
and U22857 (N_22857,N_22751,N_22777);
nand U22858 (N_22858,N_22713,N_22730);
nor U22859 (N_22859,N_22611,N_22675);
nor U22860 (N_22860,N_22606,N_22749);
and U22861 (N_22861,N_22688,N_22798);
or U22862 (N_22862,N_22733,N_22629);
xor U22863 (N_22863,N_22776,N_22716);
and U22864 (N_22864,N_22731,N_22780);
and U22865 (N_22865,N_22625,N_22635);
xor U22866 (N_22866,N_22612,N_22734);
nor U22867 (N_22867,N_22757,N_22651);
and U22868 (N_22868,N_22681,N_22604);
or U22869 (N_22869,N_22740,N_22663);
nor U22870 (N_22870,N_22784,N_22684);
xnor U22871 (N_22871,N_22680,N_22662);
xnor U22872 (N_22872,N_22792,N_22702);
nand U22873 (N_22873,N_22600,N_22771);
xor U22874 (N_22874,N_22752,N_22700);
or U22875 (N_22875,N_22667,N_22762);
and U22876 (N_22876,N_22760,N_22732);
nand U22877 (N_22877,N_22678,N_22605);
xor U22878 (N_22878,N_22615,N_22744);
or U22879 (N_22879,N_22645,N_22791);
nand U22880 (N_22880,N_22759,N_22703);
nor U22881 (N_22881,N_22622,N_22761);
xnor U22882 (N_22882,N_22782,N_22665);
nor U22883 (N_22883,N_22654,N_22608);
xnor U22884 (N_22884,N_22652,N_22657);
xor U22885 (N_22885,N_22613,N_22674);
or U22886 (N_22886,N_22677,N_22619);
nor U22887 (N_22887,N_22682,N_22756);
or U22888 (N_22888,N_22630,N_22641);
xor U22889 (N_22889,N_22766,N_22614);
xor U22890 (N_22890,N_22718,N_22735);
or U22891 (N_22891,N_22750,N_22767);
nor U22892 (N_22892,N_22694,N_22669);
nand U22893 (N_22893,N_22697,N_22610);
or U22894 (N_22894,N_22747,N_22786);
nand U22895 (N_22895,N_22778,N_22626);
xnor U22896 (N_22896,N_22653,N_22797);
or U22897 (N_22897,N_22658,N_22773);
xor U22898 (N_22898,N_22691,N_22774);
nor U22899 (N_22899,N_22795,N_22705);
nor U22900 (N_22900,N_22722,N_22645);
xor U22901 (N_22901,N_22721,N_22630);
or U22902 (N_22902,N_22756,N_22651);
and U22903 (N_22903,N_22639,N_22672);
nor U22904 (N_22904,N_22608,N_22603);
nor U22905 (N_22905,N_22657,N_22734);
or U22906 (N_22906,N_22751,N_22611);
nor U22907 (N_22907,N_22611,N_22699);
xnor U22908 (N_22908,N_22677,N_22759);
xnor U22909 (N_22909,N_22787,N_22657);
or U22910 (N_22910,N_22754,N_22701);
xor U22911 (N_22911,N_22770,N_22662);
xor U22912 (N_22912,N_22665,N_22789);
or U22913 (N_22913,N_22663,N_22602);
xnor U22914 (N_22914,N_22663,N_22680);
nand U22915 (N_22915,N_22615,N_22775);
or U22916 (N_22916,N_22681,N_22772);
xor U22917 (N_22917,N_22691,N_22756);
and U22918 (N_22918,N_22759,N_22784);
or U22919 (N_22919,N_22717,N_22626);
and U22920 (N_22920,N_22601,N_22741);
xnor U22921 (N_22921,N_22653,N_22695);
and U22922 (N_22922,N_22737,N_22685);
nor U22923 (N_22923,N_22660,N_22755);
and U22924 (N_22924,N_22797,N_22627);
or U22925 (N_22925,N_22791,N_22736);
and U22926 (N_22926,N_22782,N_22798);
or U22927 (N_22927,N_22711,N_22628);
nor U22928 (N_22928,N_22768,N_22648);
xor U22929 (N_22929,N_22794,N_22771);
and U22930 (N_22930,N_22606,N_22731);
nor U22931 (N_22931,N_22678,N_22736);
and U22932 (N_22932,N_22610,N_22675);
nor U22933 (N_22933,N_22698,N_22774);
xnor U22934 (N_22934,N_22783,N_22673);
xor U22935 (N_22935,N_22695,N_22717);
or U22936 (N_22936,N_22745,N_22712);
or U22937 (N_22937,N_22694,N_22748);
nor U22938 (N_22938,N_22606,N_22698);
or U22939 (N_22939,N_22669,N_22763);
and U22940 (N_22940,N_22783,N_22753);
nor U22941 (N_22941,N_22779,N_22721);
nor U22942 (N_22942,N_22706,N_22665);
nor U22943 (N_22943,N_22691,N_22617);
nand U22944 (N_22944,N_22770,N_22740);
and U22945 (N_22945,N_22642,N_22634);
and U22946 (N_22946,N_22629,N_22689);
or U22947 (N_22947,N_22696,N_22731);
nand U22948 (N_22948,N_22659,N_22781);
nand U22949 (N_22949,N_22657,N_22696);
xnor U22950 (N_22950,N_22617,N_22776);
nand U22951 (N_22951,N_22633,N_22726);
nor U22952 (N_22952,N_22694,N_22766);
or U22953 (N_22953,N_22662,N_22743);
and U22954 (N_22954,N_22794,N_22741);
and U22955 (N_22955,N_22708,N_22700);
nor U22956 (N_22956,N_22729,N_22604);
xnor U22957 (N_22957,N_22764,N_22690);
nor U22958 (N_22958,N_22743,N_22761);
xor U22959 (N_22959,N_22680,N_22698);
xnor U22960 (N_22960,N_22758,N_22681);
xor U22961 (N_22961,N_22760,N_22724);
xnor U22962 (N_22962,N_22613,N_22675);
nor U22963 (N_22963,N_22738,N_22699);
nor U22964 (N_22964,N_22793,N_22618);
and U22965 (N_22965,N_22762,N_22771);
nor U22966 (N_22966,N_22759,N_22681);
or U22967 (N_22967,N_22618,N_22727);
xnor U22968 (N_22968,N_22626,N_22793);
nor U22969 (N_22969,N_22719,N_22630);
and U22970 (N_22970,N_22796,N_22650);
xnor U22971 (N_22971,N_22706,N_22799);
or U22972 (N_22972,N_22765,N_22658);
or U22973 (N_22973,N_22799,N_22777);
and U22974 (N_22974,N_22648,N_22652);
and U22975 (N_22975,N_22756,N_22749);
xnor U22976 (N_22976,N_22724,N_22751);
nand U22977 (N_22977,N_22765,N_22676);
and U22978 (N_22978,N_22755,N_22648);
nand U22979 (N_22979,N_22605,N_22704);
nand U22980 (N_22980,N_22601,N_22740);
nor U22981 (N_22981,N_22637,N_22784);
or U22982 (N_22982,N_22631,N_22760);
nand U22983 (N_22983,N_22618,N_22716);
and U22984 (N_22984,N_22791,N_22737);
or U22985 (N_22985,N_22779,N_22739);
xor U22986 (N_22986,N_22707,N_22794);
xor U22987 (N_22987,N_22719,N_22756);
nor U22988 (N_22988,N_22683,N_22706);
nor U22989 (N_22989,N_22789,N_22774);
or U22990 (N_22990,N_22775,N_22635);
nand U22991 (N_22991,N_22676,N_22795);
nand U22992 (N_22992,N_22747,N_22613);
and U22993 (N_22993,N_22659,N_22733);
nor U22994 (N_22994,N_22717,N_22748);
and U22995 (N_22995,N_22664,N_22740);
and U22996 (N_22996,N_22604,N_22790);
nor U22997 (N_22997,N_22746,N_22686);
nand U22998 (N_22998,N_22615,N_22712);
and U22999 (N_22999,N_22730,N_22780);
nand U23000 (N_23000,N_22965,N_22955);
and U23001 (N_23001,N_22908,N_22966);
nor U23002 (N_23002,N_22812,N_22915);
xnor U23003 (N_23003,N_22942,N_22933);
and U23004 (N_23004,N_22929,N_22880);
or U23005 (N_23005,N_22995,N_22868);
xnor U23006 (N_23006,N_22870,N_22976);
nand U23007 (N_23007,N_22846,N_22820);
xnor U23008 (N_23008,N_22991,N_22875);
xor U23009 (N_23009,N_22809,N_22824);
or U23010 (N_23010,N_22849,N_22805);
and U23011 (N_23011,N_22927,N_22903);
xor U23012 (N_23012,N_22997,N_22877);
and U23013 (N_23013,N_22807,N_22811);
nand U23014 (N_23014,N_22937,N_22922);
xor U23015 (N_23015,N_22825,N_22841);
and U23016 (N_23016,N_22934,N_22860);
or U23017 (N_23017,N_22885,N_22948);
xor U23018 (N_23018,N_22823,N_22980);
nor U23019 (N_23019,N_22891,N_22884);
nor U23020 (N_23020,N_22800,N_22900);
nand U23021 (N_23021,N_22837,N_22974);
or U23022 (N_23022,N_22847,N_22897);
nand U23023 (N_23023,N_22865,N_22913);
xnor U23024 (N_23024,N_22834,N_22852);
nand U23025 (N_23025,N_22986,N_22924);
nand U23026 (N_23026,N_22866,N_22818);
or U23027 (N_23027,N_22972,N_22964);
or U23028 (N_23028,N_22882,N_22978);
and U23029 (N_23029,N_22961,N_22916);
and U23030 (N_23030,N_22968,N_22926);
xor U23031 (N_23031,N_22979,N_22804);
nand U23032 (N_23032,N_22844,N_22993);
nand U23033 (N_23033,N_22887,N_22826);
and U23034 (N_23034,N_22985,N_22821);
nor U23035 (N_23035,N_22902,N_22911);
or U23036 (N_23036,N_22836,N_22827);
nand U23037 (N_23037,N_22910,N_22975);
nand U23038 (N_23038,N_22947,N_22905);
xnor U23039 (N_23039,N_22919,N_22973);
nand U23040 (N_23040,N_22958,N_22944);
nand U23041 (N_23041,N_22989,N_22918);
nand U23042 (N_23042,N_22940,N_22938);
nor U23043 (N_23043,N_22803,N_22856);
xnor U23044 (N_23044,N_22983,N_22894);
and U23045 (N_23045,N_22822,N_22967);
xor U23046 (N_23046,N_22899,N_22838);
nor U23047 (N_23047,N_22878,N_22890);
nand U23048 (N_23048,N_22867,N_22923);
xnor U23049 (N_23049,N_22906,N_22828);
nand U23050 (N_23050,N_22941,N_22802);
or U23051 (N_23051,N_22872,N_22896);
and U23052 (N_23052,N_22883,N_22801);
and U23053 (N_23053,N_22859,N_22831);
and U23054 (N_23054,N_22829,N_22932);
nor U23055 (N_23055,N_22998,N_22819);
xor U23056 (N_23056,N_22851,N_22814);
and U23057 (N_23057,N_22842,N_22839);
xnor U23058 (N_23058,N_22898,N_22833);
nand U23059 (N_23059,N_22850,N_22871);
or U23060 (N_23060,N_22949,N_22810);
or U23061 (N_23061,N_22914,N_22858);
xnor U23062 (N_23062,N_22892,N_22853);
xnor U23063 (N_23063,N_22854,N_22888);
xor U23064 (N_23064,N_22953,N_22988);
or U23065 (N_23065,N_22943,N_22909);
and U23066 (N_23066,N_22996,N_22904);
nor U23067 (N_23067,N_22928,N_22845);
xor U23068 (N_23068,N_22963,N_22879);
nand U23069 (N_23069,N_22984,N_22855);
xor U23070 (N_23070,N_22864,N_22840);
or U23071 (N_23071,N_22925,N_22889);
xor U23072 (N_23072,N_22990,N_22936);
nand U23073 (N_23073,N_22806,N_22946);
nor U23074 (N_23074,N_22969,N_22962);
xor U23075 (N_23075,N_22999,N_22920);
and U23076 (N_23076,N_22876,N_22817);
nor U23077 (N_23077,N_22815,N_22931);
nand U23078 (N_23078,N_22808,N_22954);
nor U23079 (N_23079,N_22901,N_22862);
nor U23080 (N_23080,N_22950,N_22895);
and U23081 (N_23081,N_22956,N_22912);
and U23082 (N_23082,N_22874,N_22970);
xnor U23083 (N_23083,N_22971,N_22816);
or U23084 (N_23084,N_22959,N_22848);
nor U23085 (N_23085,N_22977,N_22857);
nor U23086 (N_23086,N_22930,N_22830);
nor U23087 (N_23087,N_22869,N_22957);
and U23088 (N_23088,N_22981,N_22935);
nand U23089 (N_23089,N_22921,N_22994);
and U23090 (N_23090,N_22952,N_22886);
xor U23091 (N_23091,N_22843,N_22939);
xnor U23092 (N_23092,N_22992,N_22960);
and U23093 (N_23093,N_22907,N_22951);
or U23094 (N_23094,N_22917,N_22813);
or U23095 (N_23095,N_22835,N_22832);
nand U23096 (N_23096,N_22861,N_22881);
nand U23097 (N_23097,N_22982,N_22893);
nor U23098 (N_23098,N_22987,N_22945);
nand U23099 (N_23099,N_22873,N_22863);
nor U23100 (N_23100,N_22804,N_22826);
nand U23101 (N_23101,N_22996,N_22971);
and U23102 (N_23102,N_22984,N_22912);
and U23103 (N_23103,N_22891,N_22860);
xor U23104 (N_23104,N_22885,N_22910);
nor U23105 (N_23105,N_22868,N_22870);
or U23106 (N_23106,N_22897,N_22890);
or U23107 (N_23107,N_22846,N_22915);
nor U23108 (N_23108,N_22804,N_22998);
and U23109 (N_23109,N_22801,N_22829);
nor U23110 (N_23110,N_22871,N_22986);
nand U23111 (N_23111,N_22899,N_22992);
nand U23112 (N_23112,N_22999,N_22936);
xor U23113 (N_23113,N_22972,N_22802);
xnor U23114 (N_23114,N_22884,N_22839);
nand U23115 (N_23115,N_22893,N_22868);
or U23116 (N_23116,N_22835,N_22913);
and U23117 (N_23117,N_22977,N_22844);
nor U23118 (N_23118,N_22896,N_22863);
xor U23119 (N_23119,N_22990,N_22842);
xor U23120 (N_23120,N_22912,N_22844);
or U23121 (N_23121,N_22985,N_22931);
and U23122 (N_23122,N_22933,N_22810);
xor U23123 (N_23123,N_22938,N_22980);
nand U23124 (N_23124,N_22887,N_22853);
and U23125 (N_23125,N_22828,N_22930);
nor U23126 (N_23126,N_22899,N_22916);
and U23127 (N_23127,N_22910,N_22992);
xnor U23128 (N_23128,N_22927,N_22916);
nand U23129 (N_23129,N_22912,N_22990);
nand U23130 (N_23130,N_22987,N_22838);
or U23131 (N_23131,N_22998,N_22840);
nand U23132 (N_23132,N_22830,N_22945);
xor U23133 (N_23133,N_22815,N_22986);
nand U23134 (N_23134,N_22978,N_22921);
nor U23135 (N_23135,N_22909,N_22889);
or U23136 (N_23136,N_22847,N_22931);
or U23137 (N_23137,N_22895,N_22908);
and U23138 (N_23138,N_22842,N_22871);
or U23139 (N_23139,N_22909,N_22877);
xor U23140 (N_23140,N_22958,N_22952);
xnor U23141 (N_23141,N_22828,N_22870);
or U23142 (N_23142,N_22960,N_22801);
or U23143 (N_23143,N_22803,N_22870);
nor U23144 (N_23144,N_22911,N_22865);
or U23145 (N_23145,N_22918,N_22853);
nand U23146 (N_23146,N_22963,N_22914);
xnor U23147 (N_23147,N_22801,N_22877);
xor U23148 (N_23148,N_22812,N_22950);
nor U23149 (N_23149,N_22872,N_22841);
xor U23150 (N_23150,N_22870,N_22890);
nand U23151 (N_23151,N_22816,N_22926);
or U23152 (N_23152,N_22807,N_22835);
nand U23153 (N_23153,N_22973,N_22953);
xor U23154 (N_23154,N_22831,N_22993);
nor U23155 (N_23155,N_22975,N_22938);
or U23156 (N_23156,N_22918,N_22815);
nand U23157 (N_23157,N_22840,N_22845);
nand U23158 (N_23158,N_22837,N_22937);
and U23159 (N_23159,N_22856,N_22995);
and U23160 (N_23160,N_22837,N_22822);
nor U23161 (N_23161,N_22961,N_22856);
or U23162 (N_23162,N_22816,N_22802);
nor U23163 (N_23163,N_22906,N_22806);
or U23164 (N_23164,N_22929,N_22978);
or U23165 (N_23165,N_22876,N_22906);
and U23166 (N_23166,N_22834,N_22952);
xor U23167 (N_23167,N_22949,N_22947);
and U23168 (N_23168,N_22882,N_22865);
xor U23169 (N_23169,N_22902,N_22948);
or U23170 (N_23170,N_22873,N_22841);
nand U23171 (N_23171,N_22918,N_22890);
and U23172 (N_23172,N_22872,N_22912);
xor U23173 (N_23173,N_22894,N_22829);
or U23174 (N_23174,N_22995,N_22961);
nand U23175 (N_23175,N_22903,N_22809);
or U23176 (N_23176,N_22883,N_22964);
and U23177 (N_23177,N_22855,N_22870);
xnor U23178 (N_23178,N_22845,N_22863);
nor U23179 (N_23179,N_22973,N_22898);
and U23180 (N_23180,N_22895,N_22916);
nor U23181 (N_23181,N_22845,N_22917);
and U23182 (N_23182,N_22914,N_22926);
and U23183 (N_23183,N_22839,N_22852);
xor U23184 (N_23184,N_22973,N_22878);
nand U23185 (N_23185,N_22892,N_22894);
or U23186 (N_23186,N_22897,N_22975);
nor U23187 (N_23187,N_22868,N_22882);
nor U23188 (N_23188,N_22820,N_22981);
and U23189 (N_23189,N_22957,N_22895);
nand U23190 (N_23190,N_22986,N_22994);
xor U23191 (N_23191,N_22841,N_22845);
and U23192 (N_23192,N_22940,N_22971);
and U23193 (N_23193,N_22947,N_22891);
xor U23194 (N_23194,N_22928,N_22955);
or U23195 (N_23195,N_22940,N_22858);
and U23196 (N_23196,N_22867,N_22857);
nor U23197 (N_23197,N_22829,N_22976);
or U23198 (N_23198,N_22940,N_22879);
nand U23199 (N_23199,N_22859,N_22908);
or U23200 (N_23200,N_23114,N_23111);
and U23201 (N_23201,N_23040,N_23179);
or U23202 (N_23202,N_23047,N_23096);
xor U23203 (N_23203,N_23050,N_23084);
nor U23204 (N_23204,N_23000,N_23070);
xor U23205 (N_23205,N_23154,N_23128);
or U23206 (N_23206,N_23081,N_23143);
nand U23207 (N_23207,N_23086,N_23164);
nor U23208 (N_23208,N_23008,N_23026);
nand U23209 (N_23209,N_23137,N_23094);
and U23210 (N_23210,N_23069,N_23056);
and U23211 (N_23211,N_23105,N_23109);
or U23212 (N_23212,N_23065,N_23034);
nand U23213 (N_23213,N_23108,N_23027);
or U23214 (N_23214,N_23018,N_23068);
or U23215 (N_23215,N_23085,N_23103);
and U23216 (N_23216,N_23054,N_23199);
or U23217 (N_23217,N_23042,N_23005);
nor U23218 (N_23218,N_23122,N_23064);
and U23219 (N_23219,N_23171,N_23090);
nor U23220 (N_23220,N_23145,N_23093);
nand U23221 (N_23221,N_23112,N_23038);
nor U23222 (N_23222,N_23131,N_23014);
and U23223 (N_23223,N_23148,N_23039);
nor U23224 (N_23224,N_23023,N_23155);
nor U23225 (N_23225,N_23049,N_23072);
nand U23226 (N_23226,N_23033,N_23187);
xor U23227 (N_23227,N_23170,N_23194);
xnor U23228 (N_23228,N_23101,N_23166);
xnor U23229 (N_23229,N_23041,N_23120);
nand U23230 (N_23230,N_23193,N_23097);
or U23231 (N_23231,N_23123,N_23061);
or U23232 (N_23232,N_23019,N_23010);
nand U23233 (N_23233,N_23020,N_23104);
xor U23234 (N_23234,N_23058,N_23102);
nand U23235 (N_23235,N_23035,N_23092);
nor U23236 (N_23236,N_23172,N_23181);
or U23237 (N_23237,N_23012,N_23059);
nor U23238 (N_23238,N_23141,N_23075);
xor U23239 (N_23239,N_23060,N_23133);
and U23240 (N_23240,N_23195,N_23198);
nand U23241 (N_23241,N_23189,N_23029);
nor U23242 (N_23242,N_23046,N_23113);
and U23243 (N_23243,N_23186,N_23134);
or U23244 (N_23244,N_23175,N_23051);
and U23245 (N_23245,N_23159,N_23074);
nor U23246 (N_23246,N_23173,N_23140);
and U23247 (N_23247,N_23174,N_23160);
xnor U23248 (N_23248,N_23052,N_23153);
and U23249 (N_23249,N_23004,N_23163);
or U23250 (N_23250,N_23138,N_23150);
and U23251 (N_23251,N_23082,N_23165);
and U23252 (N_23252,N_23188,N_23158);
nand U23253 (N_23253,N_23191,N_23146);
and U23254 (N_23254,N_23157,N_23037);
nor U23255 (N_23255,N_23182,N_23073);
xnor U23256 (N_23256,N_23169,N_23080);
nand U23257 (N_23257,N_23192,N_23045);
or U23258 (N_23258,N_23127,N_23190);
nand U23259 (N_23259,N_23017,N_23151);
nand U23260 (N_23260,N_23178,N_23129);
nand U23261 (N_23261,N_23006,N_23067);
or U23262 (N_23262,N_23149,N_23001);
and U23263 (N_23263,N_23055,N_23197);
nor U23264 (N_23264,N_23044,N_23142);
nand U23265 (N_23265,N_23036,N_23062);
and U23266 (N_23266,N_23088,N_23007);
or U23267 (N_23267,N_23136,N_23098);
nand U23268 (N_23268,N_23078,N_23196);
nor U23269 (N_23269,N_23162,N_23025);
and U23270 (N_23270,N_23022,N_23013);
xnor U23271 (N_23271,N_23021,N_23002);
nor U23272 (N_23272,N_23144,N_23126);
and U23273 (N_23273,N_23183,N_23016);
xor U23274 (N_23274,N_23115,N_23135);
or U23275 (N_23275,N_23076,N_23066);
or U23276 (N_23276,N_23139,N_23130);
or U23277 (N_23277,N_23156,N_23168);
xnor U23278 (N_23278,N_23089,N_23106);
xor U23279 (N_23279,N_23161,N_23167);
and U23280 (N_23280,N_23077,N_23185);
xnor U23281 (N_23281,N_23124,N_23087);
nand U23282 (N_23282,N_23121,N_23095);
and U23283 (N_23283,N_23043,N_23118);
or U23284 (N_23284,N_23177,N_23119);
and U23285 (N_23285,N_23125,N_23003);
nor U23286 (N_23286,N_23009,N_23107);
nand U23287 (N_23287,N_23083,N_23099);
or U23288 (N_23288,N_23176,N_23071);
or U23289 (N_23289,N_23015,N_23152);
nand U23290 (N_23290,N_23057,N_23117);
and U23291 (N_23291,N_23053,N_23132);
or U23292 (N_23292,N_23030,N_23180);
nand U23293 (N_23293,N_23032,N_23024);
xnor U23294 (N_23294,N_23028,N_23079);
xor U23295 (N_23295,N_23116,N_23100);
and U23296 (N_23296,N_23091,N_23048);
xor U23297 (N_23297,N_23011,N_23063);
nand U23298 (N_23298,N_23031,N_23110);
or U23299 (N_23299,N_23147,N_23184);
nor U23300 (N_23300,N_23173,N_23086);
and U23301 (N_23301,N_23071,N_23014);
and U23302 (N_23302,N_23163,N_23056);
and U23303 (N_23303,N_23117,N_23073);
and U23304 (N_23304,N_23117,N_23021);
nand U23305 (N_23305,N_23178,N_23159);
xnor U23306 (N_23306,N_23097,N_23153);
xor U23307 (N_23307,N_23065,N_23106);
nand U23308 (N_23308,N_23020,N_23193);
or U23309 (N_23309,N_23131,N_23026);
and U23310 (N_23310,N_23010,N_23046);
or U23311 (N_23311,N_23192,N_23140);
xnor U23312 (N_23312,N_23135,N_23110);
and U23313 (N_23313,N_23195,N_23051);
nand U23314 (N_23314,N_23074,N_23143);
or U23315 (N_23315,N_23172,N_23182);
xor U23316 (N_23316,N_23179,N_23001);
xor U23317 (N_23317,N_23065,N_23155);
nor U23318 (N_23318,N_23017,N_23003);
nor U23319 (N_23319,N_23029,N_23129);
or U23320 (N_23320,N_23178,N_23147);
nand U23321 (N_23321,N_23087,N_23090);
xor U23322 (N_23322,N_23105,N_23038);
or U23323 (N_23323,N_23083,N_23065);
and U23324 (N_23324,N_23128,N_23185);
and U23325 (N_23325,N_23175,N_23141);
or U23326 (N_23326,N_23014,N_23103);
nor U23327 (N_23327,N_23161,N_23037);
nand U23328 (N_23328,N_23030,N_23047);
nor U23329 (N_23329,N_23122,N_23183);
and U23330 (N_23330,N_23172,N_23085);
nand U23331 (N_23331,N_23091,N_23107);
xnor U23332 (N_23332,N_23114,N_23012);
nand U23333 (N_23333,N_23117,N_23131);
xor U23334 (N_23334,N_23199,N_23163);
xnor U23335 (N_23335,N_23100,N_23181);
xor U23336 (N_23336,N_23031,N_23190);
and U23337 (N_23337,N_23131,N_23016);
or U23338 (N_23338,N_23102,N_23052);
and U23339 (N_23339,N_23195,N_23076);
and U23340 (N_23340,N_23096,N_23183);
xor U23341 (N_23341,N_23111,N_23142);
and U23342 (N_23342,N_23152,N_23116);
or U23343 (N_23343,N_23025,N_23014);
nor U23344 (N_23344,N_23072,N_23192);
and U23345 (N_23345,N_23104,N_23044);
nand U23346 (N_23346,N_23043,N_23042);
or U23347 (N_23347,N_23098,N_23017);
or U23348 (N_23348,N_23174,N_23102);
and U23349 (N_23349,N_23057,N_23176);
nor U23350 (N_23350,N_23150,N_23014);
nand U23351 (N_23351,N_23035,N_23036);
nand U23352 (N_23352,N_23117,N_23072);
xor U23353 (N_23353,N_23108,N_23152);
nor U23354 (N_23354,N_23153,N_23002);
or U23355 (N_23355,N_23197,N_23063);
xor U23356 (N_23356,N_23163,N_23029);
nor U23357 (N_23357,N_23003,N_23140);
nor U23358 (N_23358,N_23097,N_23062);
nand U23359 (N_23359,N_23080,N_23175);
nor U23360 (N_23360,N_23045,N_23025);
nand U23361 (N_23361,N_23011,N_23123);
xnor U23362 (N_23362,N_23033,N_23180);
nand U23363 (N_23363,N_23165,N_23006);
nor U23364 (N_23364,N_23063,N_23062);
xnor U23365 (N_23365,N_23073,N_23168);
nor U23366 (N_23366,N_23014,N_23089);
nand U23367 (N_23367,N_23106,N_23108);
nor U23368 (N_23368,N_23094,N_23101);
nand U23369 (N_23369,N_23097,N_23189);
or U23370 (N_23370,N_23073,N_23091);
nor U23371 (N_23371,N_23041,N_23005);
xor U23372 (N_23372,N_23196,N_23013);
or U23373 (N_23373,N_23106,N_23159);
or U23374 (N_23374,N_23093,N_23002);
xnor U23375 (N_23375,N_23097,N_23020);
or U23376 (N_23376,N_23041,N_23172);
nor U23377 (N_23377,N_23100,N_23044);
nor U23378 (N_23378,N_23003,N_23028);
nor U23379 (N_23379,N_23132,N_23020);
nor U23380 (N_23380,N_23186,N_23187);
xor U23381 (N_23381,N_23183,N_23135);
xnor U23382 (N_23382,N_23135,N_23178);
or U23383 (N_23383,N_23145,N_23188);
or U23384 (N_23384,N_23007,N_23038);
or U23385 (N_23385,N_23027,N_23016);
and U23386 (N_23386,N_23041,N_23012);
nand U23387 (N_23387,N_23155,N_23169);
xnor U23388 (N_23388,N_23052,N_23146);
or U23389 (N_23389,N_23101,N_23087);
nor U23390 (N_23390,N_23152,N_23090);
nor U23391 (N_23391,N_23089,N_23048);
nor U23392 (N_23392,N_23031,N_23154);
and U23393 (N_23393,N_23033,N_23087);
nand U23394 (N_23394,N_23069,N_23062);
or U23395 (N_23395,N_23129,N_23135);
or U23396 (N_23396,N_23135,N_23117);
xnor U23397 (N_23397,N_23173,N_23161);
xnor U23398 (N_23398,N_23103,N_23119);
xor U23399 (N_23399,N_23037,N_23112);
nor U23400 (N_23400,N_23324,N_23238);
or U23401 (N_23401,N_23354,N_23387);
or U23402 (N_23402,N_23297,N_23374);
and U23403 (N_23403,N_23385,N_23283);
or U23404 (N_23404,N_23351,N_23355);
and U23405 (N_23405,N_23392,N_23276);
xor U23406 (N_23406,N_23240,N_23350);
or U23407 (N_23407,N_23292,N_23341);
nand U23408 (N_23408,N_23223,N_23303);
and U23409 (N_23409,N_23313,N_23381);
and U23410 (N_23410,N_23259,N_23268);
xnor U23411 (N_23411,N_23291,N_23287);
nor U23412 (N_23412,N_23231,N_23304);
nor U23413 (N_23413,N_23256,N_23221);
xnor U23414 (N_23414,N_23378,N_23248);
xnor U23415 (N_23415,N_23266,N_23214);
nand U23416 (N_23416,N_23315,N_23247);
xnor U23417 (N_23417,N_23229,N_23284);
xor U23418 (N_23418,N_23302,N_23314);
xor U23419 (N_23419,N_23212,N_23220);
or U23420 (N_23420,N_23311,N_23294);
nand U23421 (N_23421,N_23343,N_23293);
xnor U23422 (N_23422,N_23368,N_23376);
and U23423 (N_23423,N_23389,N_23337);
nand U23424 (N_23424,N_23328,N_23242);
nor U23425 (N_23425,N_23280,N_23249);
nand U23426 (N_23426,N_23356,N_23241);
nand U23427 (N_23427,N_23218,N_23282);
nand U23428 (N_23428,N_23306,N_23252);
and U23429 (N_23429,N_23257,N_23342);
and U23430 (N_23430,N_23344,N_23271);
xnor U23431 (N_23431,N_23200,N_23396);
nand U23432 (N_23432,N_23377,N_23373);
nand U23433 (N_23433,N_23333,N_23394);
nand U23434 (N_23434,N_23393,N_23281);
and U23435 (N_23435,N_23228,N_23295);
nand U23436 (N_23436,N_23367,N_23202);
nor U23437 (N_23437,N_23275,N_23310);
or U23438 (N_23438,N_23213,N_23232);
nor U23439 (N_23439,N_23349,N_23346);
and U23440 (N_23440,N_23301,N_23335);
nand U23441 (N_23441,N_23325,N_23334);
xnor U23442 (N_23442,N_23206,N_23362);
nand U23443 (N_23443,N_23234,N_23299);
or U23444 (N_23444,N_23285,N_23320);
and U23445 (N_23445,N_23258,N_23336);
nand U23446 (N_23446,N_23398,N_23254);
xor U23447 (N_23447,N_23222,N_23375);
and U23448 (N_23448,N_23226,N_23270);
nand U23449 (N_23449,N_23331,N_23345);
xor U23450 (N_23450,N_23316,N_23359);
nor U23451 (N_23451,N_23321,N_23279);
and U23452 (N_23452,N_23219,N_23309);
or U23453 (N_23453,N_23322,N_23253);
nand U23454 (N_23454,N_23384,N_23263);
and U23455 (N_23455,N_23216,N_23370);
nand U23456 (N_23456,N_23286,N_23205);
or U23457 (N_23457,N_23358,N_23211);
or U23458 (N_23458,N_23289,N_23217);
nor U23459 (N_23459,N_23274,N_23361);
xor U23460 (N_23460,N_23357,N_23265);
xnor U23461 (N_23461,N_23319,N_23261);
or U23462 (N_23462,N_23353,N_23397);
or U23463 (N_23463,N_23307,N_23391);
nand U23464 (N_23464,N_23383,N_23347);
xor U23465 (N_23465,N_23204,N_23338);
nor U23466 (N_23466,N_23224,N_23300);
nand U23467 (N_23467,N_23382,N_23380);
and U23468 (N_23468,N_23239,N_23201);
or U23469 (N_23469,N_23371,N_23250);
xnor U23470 (N_23470,N_23262,N_23207);
and U23471 (N_23471,N_23277,N_23208);
or U23472 (N_23472,N_23244,N_23236);
and U23473 (N_23473,N_23233,N_23251);
or U23474 (N_23474,N_23372,N_23225);
xor U23475 (N_23475,N_23305,N_23326);
and U23476 (N_23476,N_23339,N_23369);
nor U23477 (N_23477,N_23332,N_23323);
and U23478 (N_23478,N_23210,N_23296);
xnor U23479 (N_23479,N_23235,N_23308);
nor U23480 (N_23480,N_23388,N_23288);
nor U23481 (N_23481,N_23267,N_23269);
or U23482 (N_23482,N_23340,N_23329);
nand U23483 (N_23483,N_23318,N_23264);
nand U23484 (N_23484,N_23290,N_23327);
and U23485 (N_23485,N_23298,N_23245);
or U23486 (N_23486,N_23330,N_23227);
and U23487 (N_23487,N_23230,N_23364);
or U23488 (N_23488,N_23366,N_23399);
nor U23489 (N_23489,N_23278,N_23390);
nor U23490 (N_23490,N_23348,N_23215);
and U23491 (N_23491,N_23237,N_23365);
xor U23492 (N_23492,N_23209,N_23260);
or U23493 (N_23493,N_23255,N_23386);
nand U23494 (N_23494,N_23312,N_23395);
xor U23495 (N_23495,N_23273,N_23352);
xor U23496 (N_23496,N_23243,N_23272);
or U23497 (N_23497,N_23360,N_23246);
nor U23498 (N_23498,N_23363,N_23379);
nor U23499 (N_23499,N_23317,N_23203);
or U23500 (N_23500,N_23371,N_23365);
xor U23501 (N_23501,N_23272,N_23200);
or U23502 (N_23502,N_23204,N_23355);
xor U23503 (N_23503,N_23377,N_23399);
nor U23504 (N_23504,N_23387,N_23206);
nor U23505 (N_23505,N_23396,N_23211);
or U23506 (N_23506,N_23361,N_23255);
nand U23507 (N_23507,N_23302,N_23345);
or U23508 (N_23508,N_23205,N_23340);
nand U23509 (N_23509,N_23257,N_23320);
nor U23510 (N_23510,N_23334,N_23281);
xor U23511 (N_23511,N_23238,N_23234);
or U23512 (N_23512,N_23269,N_23273);
and U23513 (N_23513,N_23358,N_23396);
xnor U23514 (N_23514,N_23391,N_23238);
or U23515 (N_23515,N_23369,N_23335);
or U23516 (N_23516,N_23279,N_23334);
nor U23517 (N_23517,N_23335,N_23312);
or U23518 (N_23518,N_23296,N_23386);
nor U23519 (N_23519,N_23201,N_23298);
nor U23520 (N_23520,N_23360,N_23377);
and U23521 (N_23521,N_23377,N_23387);
xor U23522 (N_23522,N_23251,N_23278);
nand U23523 (N_23523,N_23361,N_23283);
nor U23524 (N_23524,N_23262,N_23321);
and U23525 (N_23525,N_23300,N_23261);
xnor U23526 (N_23526,N_23376,N_23330);
nor U23527 (N_23527,N_23397,N_23245);
xnor U23528 (N_23528,N_23222,N_23347);
nand U23529 (N_23529,N_23221,N_23349);
xor U23530 (N_23530,N_23325,N_23322);
xor U23531 (N_23531,N_23271,N_23221);
and U23532 (N_23532,N_23219,N_23264);
xnor U23533 (N_23533,N_23214,N_23230);
nor U23534 (N_23534,N_23302,N_23214);
xor U23535 (N_23535,N_23385,N_23288);
and U23536 (N_23536,N_23302,N_23355);
nand U23537 (N_23537,N_23380,N_23359);
or U23538 (N_23538,N_23253,N_23241);
nand U23539 (N_23539,N_23256,N_23206);
xnor U23540 (N_23540,N_23243,N_23329);
and U23541 (N_23541,N_23389,N_23254);
xor U23542 (N_23542,N_23229,N_23395);
and U23543 (N_23543,N_23366,N_23281);
nand U23544 (N_23544,N_23394,N_23319);
xor U23545 (N_23545,N_23223,N_23391);
or U23546 (N_23546,N_23286,N_23278);
nor U23547 (N_23547,N_23263,N_23256);
xnor U23548 (N_23548,N_23207,N_23374);
nor U23549 (N_23549,N_23336,N_23282);
and U23550 (N_23550,N_23307,N_23326);
nand U23551 (N_23551,N_23262,N_23273);
nand U23552 (N_23552,N_23287,N_23320);
or U23553 (N_23553,N_23335,N_23228);
xor U23554 (N_23554,N_23303,N_23204);
nor U23555 (N_23555,N_23349,N_23294);
xnor U23556 (N_23556,N_23310,N_23233);
nand U23557 (N_23557,N_23201,N_23302);
nand U23558 (N_23558,N_23355,N_23206);
and U23559 (N_23559,N_23380,N_23207);
nand U23560 (N_23560,N_23241,N_23324);
xor U23561 (N_23561,N_23368,N_23330);
xor U23562 (N_23562,N_23261,N_23224);
xnor U23563 (N_23563,N_23269,N_23294);
xnor U23564 (N_23564,N_23269,N_23260);
nor U23565 (N_23565,N_23201,N_23281);
or U23566 (N_23566,N_23386,N_23297);
and U23567 (N_23567,N_23316,N_23261);
nor U23568 (N_23568,N_23225,N_23367);
and U23569 (N_23569,N_23238,N_23263);
nor U23570 (N_23570,N_23377,N_23337);
and U23571 (N_23571,N_23219,N_23376);
nor U23572 (N_23572,N_23231,N_23347);
nand U23573 (N_23573,N_23215,N_23238);
xor U23574 (N_23574,N_23224,N_23377);
or U23575 (N_23575,N_23207,N_23346);
nand U23576 (N_23576,N_23368,N_23225);
and U23577 (N_23577,N_23378,N_23306);
nand U23578 (N_23578,N_23395,N_23398);
nand U23579 (N_23579,N_23316,N_23291);
nor U23580 (N_23580,N_23292,N_23323);
nand U23581 (N_23581,N_23368,N_23363);
and U23582 (N_23582,N_23206,N_23334);
nand U23583 (N_23583,N_23224,N_23264);
nand U23584 (N_23584,N_23249,N_23381);
and U23585 (N_23585,N_23340,N_23349);
xnor U23586 (N_23586,N_23314,N_23266);
nand U23587 (N_23587,N_23299,N_23353);
or U23588 (N_23588,N_23323,N_23288);
and U23589 (N_23589,N_23210,N_23354);
and U23590 (N_23590,N_23273,N_23219);
xor U23591 (N_23591,N_23303,N_23310);
and U23592 (N_23592,N_23248,N_23339);
nor U23593 (N_23593,N_23214,N_23340);
or U23594 (N_23594,N_23366,N_23339);
and U23595 (N_23595,N_23309,N_23336);
xor U23596 (N_23596,N_23233,N_23374);
or U23597 (N_23597,N_23379,N_23245);
xor U23598 (N_23598,N_23227,N_23368);
nor U23599 (N_23599,N_23355,N_23340);
or U23600 (N_23600,N_23588,N_23413);
nor U23601 (N_23601,N_23490,N_23441);
and U23602 (N_23602,N_23498,N_23405);
and U23603 (N_23603,N_23469,N_23591);
or U23604 (N_23604,N_23541,N_23404);
nand U23605 (N_23605,N_23552,N_23432);
nand U23606 (N_23606,N_23503,N_23408);
xor U23607 (N_23607,N_23568,N_23590);
xor U23608 (N_23608,N_23522,N_23415);
nor U23609 (N_23609,N_23485,N_23480);
nand U23610 (N_23610,N_23573,N_23418);
nand U23611 (N_23611,N_23487,N_23453);
xor U23612 (N_23612,N_23467,N_23407);
and U23613 (N_23613,N_23563,N_23452);
and U23614 (N_23614,N_23439,N_23505);
nand U23615 (N_23615,N_23481,N_23474);
and U23616 (N_23616,N_23527,N_23537);
or U23617 (N_23617,N_23547,N_23400);
nand U23618 (N_23618,N_23442,N_23513);
nor U23619 (N_23619,N_23411,N_23545);
xnor U23620 (N_23620,N_23523,N_23465);
xor U23621 (N_23621,N_23497,N_23575);
nor U23622 (N_23622,N_23509,N_23462);
xnor U23623 (N_23623,N_23542,N_23529);
and U23624 (N_23624,N_23491,N_23538);
nor U23625 (N_23625,N_23524,N_23496);
or U23626 (N_23626,N_23543,N_23517);
and U23627 (N_23627,N_23549,N_23586);
and U23628 (N_23628,N_23594,N_23535);
and U23629 (N_23629,N_23426,N_23571);
or U23630 (N_23630,N_23419,N_23435);
xnor U23631 (N_23631,N_23471,N_23593);
nor U23632 (N_23632,N_23581,N_23585);
nor U23633 (N_23633,N_23569,N_23457);
and U23634 (N_23634,N_23558,N_23427);
xnor U23635 (N_23635,N_23406,N_23566);
xnor U23636 (N_23636,N_23466,N_23533);
and U23637 (N_23637,N_23401,N_23478);
or U23638 (N_23638,N_23564,N_23477);
and U23639 (N_23639,N_23499,N_23515);
or U23640 (N_23640,N_23501,N_23482);
nor U23641 (N_23641,N_23551,N_23483);
or U23642 (N_23642,N_23451,N_23472);
or U23643 (N_23643,N_23484,N_23447);
or U23644 (N_23644,N_23560,N_23429);
nor U23645 (N_23645,N_23511,N_23479);
nor U23646 (N_23646,N_23463,N_23492);
and U23647 (N_23647,N_23531,N_23598);
nor U23648 (N_23648,N_23544,N_23434);
nor U23649 (N_23649,N_23576,N_23579);
or U23650 (N_23650,N_23436,N_23540);
nor U23651 (N_23651,N_23596,N_23430);
or U23652 (N_23652,N_23417,N_23433);
or U23653 (N_23653,N_23494,N_23473);
and U23654 (N_23654,N_23459,N_23449);
or U23655 (N_23655,N_23504,N_23448);
nor U23656 (N_23656,N_23450,N_23592);
or U23657 (N_23657,N_23414,N_23587);
xnor U23658 (N_23658,N_23532,N_23582);
and U23659 (N_23659,N_23597,N_23510);
or U23660 (N_23660,N_23536,N_23409);
nor U23661 (N_23661,N_23556,N_23574);
xnor U23662 (N_23662,N_23495,N_23550);
xnor U23663 (N_23663,N_23562,N_23488);
xnor U23664 (N_23664,N_23502,N_23526);
xor U23665 (N_23665,N_23559,N_23455);
nand U23666 (N_23666,N_23425,N_23475);
nand U23667 (N_23667,N_23534,N_23595);
nor U23668 (N_23668,N_23577,N_23528);
nand U23669 (N_23669,N_23489,N_23437);
and U23670 (N_23670,N_23519,N_23461);
nand U23671 (N_23671,N_23546,N_23565);
xnor U23672 (N_23672,N_23476,N_23403);
and U23673 (N_23673,N_23423,N_23420);
nor U23674 (N_23674,N_23521,N_23567);
xnor U23675 (N_23675,N_23570,N_23506);
or U23676 (N_23676,N_23554,N_23578);
and U23677 (N_23677,N_23416,N_23440);
xor U23678 (N_23678,N_23572,N_23443);
or U23679 (N_23679,N_23468,N_23539);
nand U23680 (N_23680,N_23454,N_23584);
nand U23681 (N_23681,N_23557,N_23589);
or U23682 (N_23682,N_23548,N_23516);
xor U23683 (N_23683,N_23410,N_23580);
xnor U23684 (N_23684,N_23470,N_23555);
or U23685 (N_23685,N_23512,N_23514);
xnor U23686 (N_23686,N_23456,N_23444);
nand U23687 (N_23687,N_23518,N_23402);
xor U23688 (N_23688,N_23458,N_23464);
nand U23689 (N_23689,N_23460,N_23508);
and U23690 (N_23690,N_23525,N_23438);
nor U23691 (N_23691,N_23486,N_23493);
xnor U23692 (N_23692,N_23445,N_23412);
or U23693 (N_23693,N_23530,N_23431);
nand U23694 (N_23694,N_23421,N_23507);
xor U23695 (N_23695,N_23424,N_23446);
and U23696 (N_23696,N_23553,N_23422);
nand U23697 (N_23697,N_23520,N_23500);
and U23698 (N_23698,N_23599,N_23428);
xnor U23699 (N_23699,N_23561,N_23583);
nor U23700 (N_23700,N_23470,N_23487);
or U23701 (N_23701,N_23464,N_23540);
nand U23702 (N_23702,N_23509,N_23400);
and U23703 (N_23703,N_23468,N_23408);
xor U23704 (N_23704,N_23564,N_23423);
nand U23705 (N_23705,N_23562,N_23409);
nor U23706 (N_23706,N_23522,N_23553);
nor U23707 (N_23707,N_23556,N_23561);
nor U23708 (N_23708,N_23569,N_23529);
xor U23709 (N_23709,N_23446,N_23406);
and U23710 (N_23710,N_23473,N_23546);
xor U23711 (N_23711,N_23517,N_23449);
and U23712 (N_23712,N_23511,N_23553);
nand U23713 (N_23713,N_23583,N_23457);
and U23714 (N_23714,N_23414,N_23497);
nand U23715 (N_23715,N_23590,N_23559);
or U23716 (N_23716,N_23575,N_23406);
nand U23717 (N_23717,N_23591,N_23405);
nand U23718 (N_23718,N_23412,N_23586);
or U23719 (N_23719,N_23547,N_23435);
and U23720 (N_23720,N_23462,N_23447);
nor U23721 (N_23721,N_23541,N_23509);
nand U23722 (N_23722,N_23453,N_23559);
nand U23723 (N_23723,N_23492,N_23560);
nor U23724 (N_23724,N_23537,N_23415);
xor U23725 (N_23725,N_23487,N_23540);
or U23726 (N_23726,N_23429,N_23476);
nor U23727 (N_23727,N_23529,N_23541);
or U23728 (N_23728,N_23460,N_23520);
or U23729 (N_23729,N_23489,N_23565);
and U23730 (N_23730,N_23502,N_23406);
or U23731 (N_23731,N_23404,N_23508);
and U23732 (N_23732,N_23586,N_23533);
xor U23733 (N_23733,N_23409,N_23574);
xnor U23734 (N_23734,N_23408,N_23451);
and U23735 (N_23735,N_23508,N_23545);
and U23736 (N_23736,N_23524,N_23425);
nand U23737 (N_23737,N_23455,N_23549);
nor U23738 (N_23738,N_23435,N_23451);
nor U23739 (N_23739,N_23549,N_23593);
nand U23740 (N_23740,N_23552,N_23502);
nand U23741 (N_23741,N_23534,N_23476);
nand U23742 (N_23742,N_23491,N_23517);
nand U23743 (N_23743,N_23599,N_23400);
xnor U23744 (N_23744,N_23511,N_23561);
nand U23745 (N_23745,N_23512,N_23484);
nand U23746 (N_23746,N_23550,N_23428);
and U23747 (N_23747,N_23589,N_23439);
and U23748 (N_23748,N_23530,N_23567);
or U23749 (N_23749,N_23589,N_23435);
or U23750 (N_23750,N_23465,N_23400);
nand U23751 (N_23751,N_23500,N_23413);
xor U23752 (N_23752,N_23476,N_23488);
and U23753 (N_23753,N_23427,N_23413);
nor U23754 (N_23754,N_23405,N_23435);
xor U23755 (N_23755,N_23557,N_23478);
nand U23756 (N_23756,N_23468,N_23515);
nor U23757 (N_23757,N_23436,N_23445);
or U23758 (N_23758,N_23559,N_23533);
nor U23759 (N_23759,N_23533,N_23549);
nor U23760 (N_23760,N_23410,N_23457);
or U23761 (N_23761,N_23587,N_23553);
or U23762 (N_23762,N_23417,N_23514);
and U23763 (N_23763,N_23441,N_23518);
nand U23764 (N_23764,N_23548,N_23587);
xor U23765 (N_23765,N_23466,N_23565);
and U23766 (N_23766,N_23550,N_23544);
or U23767 (N_23767,N_23502,N_23534);
nand U23768 (N_23768,N_23439,N_23458);
and U23769 (N_23769,N_23441,N_23429);
xnor U23770 (N_23770,N_23474,N_23498);
nor U23771 (N_23771,N_23470,N_23449);
xor U23772 (N_23772,N_23524,N_23466);
nand U23773 (N_23773,N_23418,N_23572);
or U23774 (N_23774,N_23578,N_23403);
nor U23775 (N_23775,N_23508,N_23547);
nor U23776 (N_23776,N_23420,N_23588);
or U23777 (N_23777,N_23478,N_23598);
xnor U23778 (N_23778,N_23523,N_23501);
xnor U23779 (N_23779,N_23430,N_23553);
nor U23780 (N_23780,N_23493,N_23406);
and U23781 (N_23781,N_23508,N_23431);
and U23782 (N_23782,N_23534,N_23591);
or U23783 (N_23783,N_23463,N_23471);
nand U23784 (N_23784,N_23471,N_23482);
and U23785 (N_23785,N_23537,N_23486);
and U23786 (N_23786,N_23577,N_23554);
nor U23787 (N_23787,N_23501,N_23579);
and U23788 (N_23788,N_23475,N_23415);
and U23789 (N_23789,N_23410,N_23518);
nand U23790 (N_23790,N_23545,N_23405);
and U23791 (N_23791,N_23440,N_23431);
or U23792 (N_23792,N_23420,N_23449);
and U23793 (N_23793,N_23412,N_23571);
xor U23794 (N_23794,N_23493,N_23563);
or U23795 (N_23795,N_23447,N_23430);
or U23796 (N_23796,N_23534,N_23475);
xnor U23797 (N_23797,N_23548,N_23562);
xor U23798 (N_23798,N_23433,N_23423);
and U23799 (N_23799,N_23560,N_23479);
and U23800 (N_23800,N_23649,N_23755);
and U23801 (N_23801,N_23741,N_23607);
nor U23802 (N_23802,N_23639,N_23784);
nor U23803 (N_23803,N_23660,N_23656);
nand U23804 (N_23804,N_23621,N_23609);
or U23805 (N_23805,N_23731,N_23771);
nor U23806 (N_23806,N_23602,N_23791);
nor U23807 (N_23807,N_23624,N_23664);
or U23808 (N_23808,N_23620,N_23631);
nor U23809 (N_23809,N_23718,N_23799);
xor U23810 (N_23810,N_23666,N_23782);
nor U23811 (N_23811,N_23630,N_23764);
nand U23812 (N_23812,N_23767,N_23770);
nor U23813 (N_23813,N_23680,N_23787);
and U23814 (N_23814,N_23780,N_23678);
and U23815 (N_23815,N_23761,N_23778);
xor U23816 (N_23816,N_23659,N_23793);
and U23817 (N_23817,N_23712,N_23798);
nor U23818 (N_23818,N_23629,N_23733);
nor U23819 (N_23819,N_23773,N_23600);
or U23820 (N_23820,N_23704,N_23688);
and U23821 (N_23821,N_23622,N_23722);
nand U23822 (N_23822,N_23717,N_23737);
and U23823 (N_23823,N_23681,N_23640);
nand U23824 (N_23824,N_23667,N_23642);
nor U23825 (N_23825,N_23613,N_23719);
nor U23826 (N_23826,N_23651,N_23753);
or U23827 (N_23827,N_23687,N_23652);
nor U23828 (N_23828,N_23781,N_23635);
and U23829 (N_23829,N_23674,N_23625);
and U23830 (N_23830,N_23750,N_23686);
xnor U23831 (N_23831,N_23647,N_23616);
nand U23832 (N_23832,N_23745,N_23683);
or U23833 (N_23833,N_23601,N_23700);
or U23834 (N_23834,N_23614,N_23610);
xor U23835 (N_23835,N_23714,N_23633);
and U23836 (N_23836,N_23709,N_23792);
and U23837 (N_23837,N_23788,N_23776);
nand U23838 (N_23838,N_23627,N_23760);
xor U23839 (N_23839,N_23708,N_23691);
xnor U23840 (N_23840,N_23746,N_23749);
xnor U23841 (N_23841,N_23744,N_23730);
and U23842 (N_23842,N_23675,N_23653);
nor U23843 (N_23843,N_23693,N_23604);
and U23844 (N_23844,N_23735,N_23632);
and U23845 (N_23845,N_23732,N_23606);
nand U23846 (N_23846,N_23617,N_23692);
and U23847 (N_23847,N_23650,N_23796);
and U23848 (N_23848,N_23762,N_23715);
or U23849 (N_23849,N_23637,N_23711);
nor U23850 (N_23850,N_23724,N_23789);
and U23851 (N_23851,N_23672,N_23729);
xnor U23852 (N_23852,N_23742,N_23648);
xnor U23853 (N_23853,N_23702,N_23641);
or U23854 (N_23854,N_23668,N_23603);
and U23855 (N_23855,N_23747,N_23794);
or U23856 (N_23856,N_23670,N_23685);
or U23857 (N_23857,N_23676,N_23689);
nand U23858 (N_23858,N_23765,N_23766);
and U23859 (N_23859,N_23636,N_23615);
nor U23860 (N_23860,N_23677,N_23772);
nor U23861 (N_23861,N_23665,N_23669);
and U23862 (N_23862,N_23756,N_23655);
nand U23863 (N_23863,N_23769,N_23618);
and U23864 (N_23864,N_23725,N_23701);
nor U23865 (N_23865,N_23738,N_23723);
or U23866 (N_23866,N_23626,N_23710);
or U23867 (N_23867,N_23786,N_23608);
or U23868 (N_23868,N_23619,N_23654);
nor U23869 (N_23869,N_23697,N_23758);
and U23870 (N_23870,N_23706,N_23736);
xor U23871 (N_23871,N_23726,N_23751);
or U23872 (N_23872,N_23645,N_23661);
nand U23873 (N_23873,N_23790,N_23695);
nor U23874 (N_23874,N_23743,N_23757);
and U23875 (N_23875,N_23671,N_23673);
nand U23876 (N_23876,N_23779,N_23740);
nand U23877 (N_23877,N_23623,N_23774);
nor U23878 (N_23878,N_23682,N_23720);
nor U23879 (N_23879,N_23739,N_23759);
xnor U23880 (N_23880,N_23763,N_23663);
nand U23881 (N_23881,N_23707,N_23696);
or U23882 (N_23882,N_23605,N_23777);
and U23883 (N_23883,N_23728,N_23628);
or U23884 (N_23884,N_23611,N_23638);
nor U23885 (N_23885,N_23699,N_23679);
nand U23886 (N_23886,N_23684,N_23658);
nor U23887 (N_23887,N_23752,N_23716);
and U23888 (N_23888,N_23705,N_23657);
or U23889 (N_23889,N_23783,N_23646);
xnor U23890 (N_23890,N_23785,N_23662);
and U23891 (N_23891,N_23775,N_23644);
xnor U23892 (N_23892,N_23703,N_23698);
xor U23893 (N_23893,N_23734,N_23690);
xnor U23894 (N_23894,N_23694,N_23634);
xnor U23895 (N_23895,N_23713,N_23795);
or U23896 (N_23896,N_23797,N_23612);
and U23897 (N_23897,N_23727,N_23721);
or U23898 (N_23898,N_23643,N_23754);
and U23899 (N_23899,N_23768,N_23748);
nand U23900 (N_23900,N_23637,N_23751);
nand U23901 (N_23901,N_23612,N_23754);
nor U23902 (N_23902,N_23669,N_23761);
and U23903 (N_23903,N_23656,N_23665);
nor U23904 (N_23904,N_23751,N_23632);
xor U23905 (N_23905,N_23692,N_23774);
nor U23906 (N_23906,N_23735,N_23693);
nand U23907 (N_23907,N_23607,N_23753);
and U23908 (N_23908,N_23691,N_23731);
nand U23909 (N_23909,N_23790,N_23703);
and U23910 (N_23910,N_23655,N_23601);
or U23911 (N_23911,N_23653,N_23787);
xor U23912 (N_23912,N_23611,N_23775);
xor U23913 (N_23913,N_23734,N_23723);
or U23914 (N_23914,N_23694,N_23736);
nor U23915 (N_23915,N_23696,N_23688);
xor U23916 (N_23916,N_23642,N_23624);
or U23917 (N_23917,N_23637,N_23607);
xor U23918 (N_23918,N_23613,N_23733);
nor U23919 (N_23919,N_23784,N_23611);
or U23920 (N_23920,N_23744,N_23629);
and U23921 (N_23921,N_23798,N_23729);
and U23922 (N_23922,N_23714,N_23615);
xnor U23923 (N_23923,N_23712,N_23705);
or U23924 (N_23924,N_23662,N_23637);
or U23925 (N_23925,N_23639,N_23665);
xor U23926 (N_23926,N_23623,N_23726);
and U23927 (N_23927,N_23758,N_23712);
or U23928 (N_23928,N_23776,N_23704);
nand U23929 (N_23929,N_23622,N_23627);
nor U23930 (N_23930,N_23623,N_23748);
or U23931 (N_23931,N_23790,N_23731);
xor U23932 (N_23932,N_23645,N_23736);
xor U23933 (N_23933,N_23756,N_23636);
and U23934 (N_23934,N_23682,N_23725);
xor U23935 (N_23935,N_23606,N_23687);
xnor U23936 (N_23936,N_23682,N_23655);
xnor U23937 (N_23937,N_23775,N_23605);
and U23938 (N_23938,N_23740,N_23701);
and U23939 (N_23939,N_23687,N_23674);
and U23940 (N_23940,N_23668,N_23604);
nand U23941 (N_23941,N_23715,N_23778);
nand U23942 (N_23942,N_23611,N_23799);
nand U23943 (N_23943,N_23729,N_23701);
nor U23944 (N_23944,N_23608,N_23677);
or U23945 (N_23945,N_23619,N_23645);
nor U23946 (N_23946,N_23691,N_23678);
xnor U23947 (N_23947,N_23704,N_23623);
and U23948 (N_23948,N_23666,N_23628);
or U23949 (N_23949,N_23671,N_23741);
or U23950 (N_23950,N_23740,N_23637);
xor U23951 (N_23951,N_23733,N_23671);
or U23952 (N_23952,N_23717,N_23758);
nand U23953 (N_23953,N_23615,N_23774);
nor U23954 (N_23954,N_23743,N_23697);
and U23955 (N_23955,N_23650,N_23656);
xnor U23956 (N_23956,N_23779,N_23770);
xnor U23957 (N_23957,N_23706,N_23717);
or U23958 (N_23958,N_23621,N_23651);
nand U23959 (N_23959,N_23692,N_23702);
and U23960 (N_23960,N_23611,N_23616);
nor U23961 (N_23961,N_23760,N_23775);
xor U23962 (N_23962,N_23765,N_23650);
or U23963 (N_23963,N_23675,N_23716);
nor U23964 (N_23964,N_23711,N_23683);
xor U23965 (N_23965,N_23612,N_23712);
nand U23966 (N_23966,N_23789,N_23765);
or U23967 (N_23967,N_23611,N_23600);
and U23968 (N_23968,N_23718,N_23689);
or U23969 (N_23969,N_23769,N_23784);
nor U23970 (N_23970,N_23751,N_23782);
nand U23971 (N_23971,N_23769,N_23640);
xnor U23972 (N_23972,N_23611,N_23686);
xor U23973 (N_23973,N_23701,N_23611);
nor U23974 (N_23974,N_23608,N_23743);
xor U23975 (N_23975,N_23754,N_23699);
or U23976 (N_23976,N_23632,N_23727);
nor U23977 (N_23977,N_23633,N_23748);
nor U23978 (N_23978,N_23703,N_23710);
nor U23979 (N_23979,N_23703,N_23713);
xor U23980 (N_23980,N_23776,N_23631);
xnor U23981 (N_23981,N_23774,N_23755);
nor U23982 (N_23982,N_23704,N_23603);
nor U23983 (N_23983,N_23798,N_23768);
xnor U23984 (N_23984,N_23638,N_23799);
or U23985 (N_23985,N_23684,N_23755);
xnor U23986 (N_23986,N_23786,N_23645);
nand U23987 (N_23987,N_23772,N_23625);
or U23988 (N_23988,N_23630,N_23613);
nand U23989 (N_23989,N_23613,N_23796);
or U23990 (N_23990,N_23614,N_23756);
nand U23991 (N_23991,N_23662,N_23621);
nand U23992 (N_23992,N_23772,N_23692);
nand U23993 (N_23993,N_23768,N_23656);
nor U23994 (N_23994,N_23730,N_23610);
or U23995 (N_23995,N_23760,N_23670);
nor U23996 (N_23996,N_23723,N_23716);
or U23997 (N_23997,N_23612,N_23773);
and U23998 (N_23998,N_23629,N_23680);
nor U23999 (N_23999,N_23789,N_23791);
xor U24000 (N_24000,N_23909,N_23858);
or U24001 (N_24001,N_23806,N_23917);
or U24002 (N_24002,N_23944,N_23824);
xor U24003 (N_24003,N_23869,N_23991);
or U24004 (N_24004,N_23870,N_23812);
or U24005 (N_24005,N_23998,N_23995);
xnor U24006 (N_24006,N_23993,N_23839);
or U24007 (N_24007,N_23952,N_23897);
nand U24008 (N_24008,N_23846,N_23800);
and U24009 (N_24009,N_23890,N_23941);
nor U24010 (N_24010,N_23903,N_23937);
nor U24011 (N_24011,N_23916,N_23901);
xnor U24012 (N_24012,N_23826,N_23946);
xor U24013 (N_24013,N_23996,N_23934);
xor U24014 (N_24014,N_23954,N_23857);
or U24015 (N_24015,N_23853,N_23864);
xor U24016 (N_24016,N_23927,N_23809);
xor U24017 (N_24017,N_23841,N_23896);
nor U24018 (N_24018,N_23965,N_23992);
and U24019 (N_24019,N_23950,N_23891);
xnor U24020 (N_24020,N_23838,N_23945);
nand U24021 (N_24021,N_23908,N_23842);
nand U24022 (N_24022,N_23820,N_23818);
xnor U24023 (N_24023,N_23935,N_23966);
or U24024 (N_24024,N_23971,N_23884);
or U24025 (N_24025,N_23975,N_23999);
and U24026 (N_24026,N_23802,N_23981);
nand U24027 (N_24027,N_23960,N_23930);
xnor U24028 (N_24028,N_23883,N_23905);
and U24029 (N_24029,N_23902,N_23977);
xnor U24030 (N_24030,N_23859,N_23840);
and U24031 (N_24031,N_23911,N_23973);
or U24032 (N_24032,N_23880,N_23913);
nand U24033 (N_24033,N_23974,N_23821);
nand U24034 (N_24034,N_23878,N_23819);
nor U24035 (N_24035,N_23807,N_23823);
nand U24036 (N_24036,N_23942,N_23926);
or U24037 (N_24037,N_23976,N_23827);
nor U24038 (N_24038,N_23968,N_23874);
nand U24039 (N_24039,N_23843,N_23956);
xnor U24040 (N_24040,N_23972,N_23875);
and U24041 (N_24041,N_23805,N_23929);
and U24042 (N_24042,N_23987,N_23886);
and U24043 (N_24043,N_23922,N_23907);
or U24044 (N_24044,N_23964,N_23943);
or U24045 (N_24045,N_23888,N_23881);
nand U24046 (N_24046,N_23863,N_23948);
xor U24047 (N_24047,N_23967,N_23918);
and U24048 (N_24048,N_23914,N_23816);
nor U24049 (N_24049,N_23804,N_23962);
xor U24050 (N_24050,N_23982,N_23920);
xor U24051 (N_24051,N_23835,N_23895);
and U24052 (N_24052,N_23953,N_23844);
or U24053 (N_24053,N_23959,N_23808);
or U24054 (N_24054,N_23892,N_23851);
and U24055 (N_24055,N_23949,N_23947);
nand U24056 (N_24056,N_23983,N_23871);
nor U24057 (N_24057,N_23958,N_23814);
nor U24058 (N_24058,N_23848,N_23882);
nand U24059 (N_24059,N_23803,N_23955);
or U24060 (N_24060,N_23997,N_23872);
nand U24061 (N_24061,N_23822,N_23928);
and U24062 (N_24062,N_23919,N_23810);
nand U24063 (N_24063,N_23849,N_23988);
and U24064 (N_24064,N_23801,N_23963);
and U24065 (N_24065,N_23852,N_23847);
nand U24066 (N_24066,N_23862,N_23832);
or U24067 (N_24067,N_23861,N_23811);
and U24068 (N_24068,N_23989,N_23940);
xor U24069 (N_24069,N_23828,N_23885);
or U24070 (N_24070,N_23984,N_23893);
xnor U24071 (N_24071,N_23855,N_23866);
nor U24072 (N_24072,N_23990,N_23831);
or U24073 (N_24073,N_23898,N_23877);
nand U24074 (N_24074,N_23969,N_23889);
nor U24075 (N_24075,N_23994,N_23957);
and U24076 (N_24076,N_23900,N_23837);
xor U24077 (N_24077,N_23932,N_23865);
nor U24078 (N_24078,N_23939,N_23921);
and U24079 (N_24079,N_23867,N_23850);
nor U24080 (N_24080,N_23815,N_23986);
nor U24081 (N_24081,N_23978,N_23834);
nand U24082 (N_24082,N_23951,N_23923);
or U24083 (N_24083,N_23931,N_23980);
and U24084 (N_24084,N_23873,N_23887);
xnor U24085 (N_24085,N_23899,N_23915);
nor U24086 (N_24086,N_23860,N_23933);
and U24087 (N_24087,N_23854,N_23894);
nand U24088 (N_24088,N_23938,N_23825);
or U24089 (N_24089,N_23925,N_23829);
nor U24090 (N_24090,N_23936,N_23836);
nor U24091 (N_24091,N_23856,N_23979);
or U24092 (N_24092,N_23924,N_23879);
nor U24093 (N_24093,N_23868,N_23817);
and U24094 (N_24094,N_23985,N_23961);
nor U24095 (N_24095,N_23906,N_23876);
and U24096 (N_24096,N_23912,N_23845);
xnor U24097 (N_24097,N_23904,N_23813);
nor U24098 (N_24098,N_23830,N_23970);
nor U24099 (N_24099,N_23910,N_23833);
nor U24100 (N_24100,N_23872,N_23854);
nor U24101 (N_24101,N_23894,N_23848);
nor U24102 (N_24102,N_23971,N_23993);
nor U24103 (N_24103,N_23861,N_23875);
nand U24104 (N_24104,N_23975,N_23828);
nor U24105 (N_24105,N_23966,N_23941);
or U24106 (N_24106,N_23958,N_23820);
or U24107 (N_24107,N_23998,N_23896);
or U24108 (N_24108,N_23959,N_23933);
xnor U24109 (N_24109,N_23951,N_23937);
or U24110 (N_24110,N_23985,N_23803);
nand U24111 (N_24111,N_23888,N_23969);
nor U24112 (N_24112,N_23903,N_23983);
nor U24113 (N_24113,N_23952,N_23880);
xor U24114 (N_24114,N_23835,N_23829);
and U24115 (N_24115,N_23874,N_23949);
or U24116 (N_24116,N_23829,N_23882);
or U24117 (N_24117,N_23871,N_23963);
xor U24118 (N_24118,N_23800,N_23837);
or U24119 (N_24119,N_23923,N_23906);
or U24120 (N_24120,N_23898,N_23845);
nor U24121 (N_24121,N_23887,N_23960);
xor U24122 (N_24122,N_23814,N_23985);
or U24123 (N_24123,N_23837,N_23950);
and U24124 (N_24124,N_23912,N_23859);
nor U24125 (N_24125,N_23953,N_23846);
xor U24126 (N_24126,N_23833,N_23986);
xnor U24127 (N_24127,N_23897,N_23947);
nand U24128 (N_24128,N_23909,N_23815);
nor U24129 (N_24129,N_23936,N_23993);
or U24130 (N_24130,N_23835,N_23888);
nor U24131 (N_24131,N_23894,N_23807);
nand U24132 (N_24132,N_23810,N_23854);
xnor U24133 (N_24133,N_23850,N_23979);
or U24134 (N_24134,N_23972,N_23911);
or U24135 (N_24135,N_23851,N_23896);
or U24136 (N_24136,N_23855,N_23802);
nor U24137 (N_24137,N_23868,N_23826);
xor U24138 (N_24138,N_23845,N_23951);
xnor U24139 (N_24139,N_23811,N_23964);
nor U24140 (N_24140,N_23873,N_23882);
nor U24141 (N_24141,N_23865,N_23843);
nand U24142 (N_24142,N_23893,N_23821);
and U24143 (N_24143,N_23830,N_23894);
or U24144 (N_24144,N_23807,N_23852);
or U24145 (N_24145,N_23819,N_23812);
or U24146 (N_24146,N_23803,N_23821);
and U24147 (N_24147,N_23964,N_23918);
and U24148 (N_24148,N_23986,N_23841);
nor U24149 (N_24149,N_23968,N_23999);
nand U24150 (N_24150,N_23963,N_23867);
nor U24151 (N_24151,N_23927,N_23810);
or U24152 (N_24152,N_23940,N_23941);
xor U24153 (N_24153,N_23859,N_23817);
or U24154 (N_24154,N_23954,N_23825);
and U24155 (N_24155,N_23961,N_23912);
and U24156 (N_24156,N_23986,N_23897);
and U24157 (N_24157,N_23996,N_23998);
nand U24158 (N_24158,N_23811,N_23923);
nand U24159 (N_24159,N_23975,N_23953);
nand U24160 (N_24160,N_23990,N_23891);
nand U24161 (N_24161,N_23915,N_23850);
nand U24162 (N_24162,N_23910,N_23869);
xnor U24163 (N_24163,N_23938,N_23967);
xor U24164 (N_24164,N_23815,N_23948);
nor U24165 (N_24165,N_23897,N_23917);
or U24166 (N_24166,N_23811,N_23966);
or U24167 (N_24167,N_23886,N_23817);
nand U24168 (N_24168,N_23850,N_23925);
or U24169 (N_24169,N_23988,N_23837);
nor U24170 (N_24170,N_23868,N_23871);
and U24171 (N_24171,N_23958,N_23872);
and U24172 (N_24172,N_23846,N_23918);
xor U24173 (N_24173,N_23981,N_23923);
and U24174 (N_24174,N_23999,N_23897);
nand U24175 (N_24175,N_23881,N_23847);
xnor U24176 (N_24176,N_23964,N_23884);
nor U24177 (N_24177,N_23832,N_23890);
nor U24178 (N_24178,N_23828,N_23874);
nand U24179 (N_24179,N_23936,N_23938);
nand U24180 (N_24180,N_23883,N_23886);
and U24181 (N_24181,N_23809,N_23853);
nor U24182 (N_24182,N_23924,N_23945);
xor U24183 (N_24183,N_23884,N_23905);
or U24184 (N_24184,N_23844,N_23929);
and U24185 (N_24185,N_23967,N_23896);
nor U24186 (N_24186,N_23951,N_23854);
and U24187 (N_24187,N_23990,N_23808);
xor U24188 (N_24188,N_23978,N_23833);
xor U24189 (N_24189,N_23998,N_23853);
nand U24190 (N_24190,N_23984,N_23909);
xnor U24191 (N_24191,N_23866,N_23816);
or U24192 (N_24192,N_23984,N_23892);
nand U24193 (N_24193,N_23836,N_23985);
nor U24194 (N_24194,N_23932,N_23800);
nor U24195 (N_24195,N_23835,N_23920);
and U24196 (N_24196,N_23923,N_23822);
xor U24197 (N_24197,N_23957,N_23836);
and U24198 (N_24198,N_23837,N_23859);
nand U24199 (N_24199,N_23868,N_23803);
xor U24200 (N_24200,N_24120,N_24198);
or U24201 (N_24201,N_24137,N_24105);
nor U24202 (N_24202,N_24014,N_24054);
or U24203 (N_24203,N_24085,N_24192);
or U24204 (N_24204,N_24111,N_24051);
nand U24205 (N_24205,N_24112,N_24182);
nand U24206 (N_24206,N_24037,N_24009);
nor U24207 (N_24207,N_24130,N_24074);
nor U24208 (N_24208,N_24007,N_24185);
and U24209 (N_24209,N_24033,N_24132);
nand U24210 (N_24210,N_24151,N_24189);
and U24211 (N_24211,N_24179,N_24031);
nor U24212 (N_24212,N_24155,N_24034);
nand U24213 (N_24213,N_24177,N_24024);
nor U24214 (N_24214,N_24138,N_24049);
xnor U24215 (N_24215,N_24047,N_24119);
nor U24216 (N_24216,N_24157,N_24025);
xor U24217 (N_24217,N_24013,N_24063);
or U24218 (N_24218,N_24030,N_24067);
xor U24219 (N_24219,N_24070,N_24069);
and U24220 (N_24220,N_24149,N_24032);
or U24221 (N_24221,N_24108,N_24133);
and U24222 (N_24222,N_24175,N_24090);
or U24223 (N_24223,N_24172,N_24023);
or U24224 (N_24224,N_24183,N_24164);
nand U24225 (N_24225,N_24064,N_24003);
and U24226 (N_24226,N_24059,N_24180);
xnor U24227 (N_24227,N_24015,N_24081);
or U24228 (N_24228,N_24102,N_24077);
or U24229 (N_24229,N_24147,N_24004);
xor U24230 (N_24230,N_24056,N_24026);
and U24231 (N_24231,N_24052,N_24163);
and U24232 (N_24232,N_24103,N_24018);
xnor U24233 (N_24233,N_24193,N_24017);
nor U24234 (N_24234,N_24199,N_24131);
and U24235 (N_24235,N_24098,N_24011);
nand U24236 (N_24236,N_24082,N_24053);
and U24237 (N_24237,N_24041,N_24065);
and U24238 (N_24238,N_24099,N_24076);
nor U24239 (N_24239,N_24171,N_24184);
and U24240 (N_24240,N_24190,N_24143);
xor U24241 (N_24241,N_24044,N_24062);
xor U24242 (N_24242,N_24122,N_24021);
and U24243 (N_24243,N_24170,N_24168);
xnor U24244 (N_24244,N_24161,N_24048);
nor U24245 (N_24245,N_24110,N_24087);
and U24246 (N_24246,N_24186,N_24006);
and U24247 (N_24247,N_24040,N_24142);
or U24248 (N_24248,N_24154,N_24084);
nand U24249 (N_24249,N_24022,N_24005);
and U24250 (N_24250,N_24117,N_24057);
and U24251 (N_24251,N_24101,N_24129);
and U24252 (N_24252,N_24043,N_24141);
nand U24253 (N_24253,N_24066,N_24036);
or U24254 (N_24254,N_24071,N_24008);
nand U24255 (N_24255,N_24197,N_24126);
xor U24256 (N_24256,N_24097,N_24121);
nand U24257 (N_24257,N_24079,N_24093);
and U24258 (N_24258,N_24114,N_24086);
xor U24259 (N_24259,N_24176,N_24152);
nor U24260 (N_24260,N_24109,N_24106);
and U24261 (N_24261,N_24083,N_24095);
nor U24262 (N_24262,N_24035,N_24160);
nor U24263 (N_24263,N_24038,N_24165);
or U24264 (N_24264,N_24148,N_24107);
nand U24265 (N_24265,N_24156,N_24089);
and U24266 (N_24266,N_24104,N_24055);
nor U24267 (N_24267,N_24140,N_24146);
and U24268 (N_24268,N_24159,N_24092);
nor U24269 (N_24269,N_24173,N_24058);
and U24270 (N_24270,N_24123,N_24128);
or U24271 (N_24271,N_24118,N_24050);
nor U24272 (N_24272,N_24150,N_24042);
and U24273 (N_24273,N_24196,N_24124);
or U24274 (N_24274,N_24039,N_24075);
and U24275 (N_24275,N_24169,N_24135);
and U24276 (N_24276,N_24045,N_24029);
nor U24277 (N_24277,N_24191,N_24012);
nand U24278 (N_24278,N_24115,N_24116);
nand U24279 (N_24279,N_24019,N_24073);
nor U24280 (N_24280,N_24127,N_24100);
nand U24281 (N_24281,N_24174,N_24078);
and U24282 (N_24282,N_24016,N_24027);
or U24283 (N_24283,N_24060,N_24088);
nor U24284 (N_24284,N_24144,N_24194);
nor U24285 (N_24285,N_24139,N_24153);
and U24286 (N_24286,N_24136,N_24188);
and U24287 (N_24287,N_24072,N_24167);
xor U24288 (N_24288,N_24162,N_24145);
nor U24289 (N_24289,N_24166,N_24061);
xnor U24290 (N_24290,N_24068,N_24125);
nand U24291 (N_24291,N_24080,N_24091);
nor U24292 (N_24292,N_24113,N_24096);
xor U24293 (N_24293,N_24195,N_24028);
nor U24294 (N_24294,N_24001,N_24094);
nor U24295 (N_24295,N_24187,N_24002);
nor U24296 (N_24296,N_24020,N_24010);
and U24297 (N_24297,N_24181,N_24158);
nand U24298 (N_24298,N_24046,N_24178);
nand U24299 (N_24299,N_24000,N_24134);
nand U24300 (N_24300,N_24169,N_24046);
xor U24301 (N_24301,N_24130,N_24129);
xor U24302 (N_24302,N_24023,N_24138);
or U24303 (N_24303,N_24109,N_24100);
and U24304 (N_24304,N_24100,N_24079);
xnor U24305 (N_24305,N_24057,N_24120);
xor U24306 (N_24306,N_24033,N_24119);
or U24307 (N_24307,N_24117,N_24032);
xnor U24308 (N_24308,N_24118,N_24120);
and U24309 (N_24309,N_24071,N_24153);
xor U24310 (N_24310,N_24061,N_24106);
nor U24311 (N_24311,N_24100,N_24034);
and U24312 (N_24312,N_24174,N_24037);
or U24313 (N_24313,N_24184,N_24150);
nand U24314 (N_24314,N_24050,N_24036);
nor U24315 (N_24315,N_24147,N_24140);
or U24316 (N_24316,N_24146,N_24086);
and U24317 (N_24317,N_24144,N_24164);
and U24318 (N_24318,N_24035,N_24106);
nand U24319 (N_24319,N_24085,N_24124);
and U24320 (N_24320,N_24019,N_24101);
or U24321 (N_24321,N_24193,N_24182);
and U24322 (N_24322,N_24192,N_24137);
or U24323 (N_24323,N_24107,N_24130);
or U24324 (N_24324,N_24017,N_24032);
nor U24325 (N_24325,N_24147,N_24110);
nor U24326 (N_24326,N_24141,N_24073);
and U24327 (N_24327,N_24122,N_24190);
or U24328 (N_24328,N_24186,N_24096);
nand U24329 (N_24329,N_24160,N_24146);
or U24330 (N_24330,N_24008,N_24158);
xor U24331 (N_24331,N_24105,N_24086);
or U24332 (N_24332,N_24069,N_24095);
nand U24333 (N_24333,N_24194,N_24147);
nor U24334 (N_24334,N_24042,N_24022);
xnor U24335 (N_24335,N_24023,N_24062);
nand U24336 (N_24336,N_24055,N_24120);
xnor U24337 (N_24337,N_24042,N_24188);
nor U24338 (N_24338,N_24179,N_24024);
nand U24339 (N_24339,N_24038,N_24155);
or U24340 (N_24340,N_24145,N_24179);
or U24341 (N_24341,N_24160,N_24062);
and U24342 (N_24342,N_24134,N_24180);
nor U24343 (N_24343,N_24033,N_24183);
nand U24344 (N_24344,N_24169,N_24002);
nand U24345 (N_24345,N_24119,N_24198);
or U24346 (N_24346,N_24111,N_24082);
nand U24347 (N_24347,N_24092,N_24052);
nand U24348 (N_24348,N_24148,N_24108);
nor U24349 (N_24349,N_24169,N_24110);
xnor U24350 (N_24350,N_24143,N_24048);
nand U24351 (N_24351,N_24112,N_24098);
and U24352 (N_24352,N_24044,N_24132);
or U24353 (N_24353,N_24015,N_24128);
and U24354 (N_24354,N_24151,N_24146);
nand U24355 (N_24355,N_24047,N_24165);
nor U24356 (N_24356,N_24077,N_24013);
or U24357 (N_24357,N_24129,N_24176);
xor U24358 (N_24358,N_24170,N_24175);
nor U24359 (N_24359,N_24095,N_24137);
and U24360 (N_24360,N_24098,N_24076);
and U24361 (N_24361,N_24146,N_24155);
or U24362 (N_24362,N_24039,N_24090);
or U24363 (N_24363,N_24092,N_24045);
xnor U24364 (N_24364,N_24122,N_24079);
nor U24365 (N_24365,N_24117,N_24171);
and U24366 (N_24366,N_24121,N_24100);
nand U24367 (N_24367,N_24013,N_24049);
and U24368 (N_24368,N_24009,N_24198);
xor U24369 (N_24369,N_24018,N_24127);
nor U24370 (N_24370,N_24104,N_24159);
nand U24371 (N_24371,N_24093,N_24037);
nor U24372 (N_24372,N_24063,N_24056);
nand U24373 (N_24373,N_24154,N_24003);
xor U24374 (N_24374,N_24065,N_24181);
or U24375 (N_24375,N_24137,N_24084);
xor U24376 (N_24376,N_24156,N_24158);
nor U24377 (N_24377,N_24032,N_24036);
nand U24378 (N_24378,N_24123,N_24014);
nor U24379 (N_24379,N_24040,N_24143);
or U24380 (N_24380,N_24028,N_24133);
or U24381 (N_24381,N_24042,N_24166);
and U24382 (N_24382,N_24067,N_24106);
and U24383 (N_24383,N_24183,N_24045);
nor U24384 (N_24384,N_24148,N_24041);
xnor U24385 (N_24385,N_24098,N_24006);
or U24386 (N_24386,N_24007,N_24083);
or U24387 (N_24387,N_24146,N_24144);
xnor U24388 (N_24388,N_24022,N_24142);
nor U24389 (N_24389,N_24031,N_24120);
xor U24390 (N_24390,N_24067,N_24078);
nor U24391 (N_24391,N_24090,N_24188);
or U24392 (N_24392,N_24123,N_24174);
nor U24393 (N_24393,N_24099,N_24056);
or U24394 (N_24394,N_24069,N_24068);
nand U24395 (N_24395,N_24197,N_24110);
nand U24396 (N_24396,N_24131,N_24108);
nor U24397 (N_24397,N_24050,N_24128);
or U24398 (N_24398,N_24156,N_24157);
xor U24399 (N_24399,N_24006,N_24165);
xor U24400 (N_24400,N_24229,N_24284);
and U24401 (N_24401,N_24207,N_24324);
nor U24402 (N_24402,N_24340,N_24396);
nand U24403 (N_24403,N_24275,N_24354);
or U24404 (N_24404,N_24247,N_24294);
xnor U24405 (N_24405,N_24338,N_24240);
and U24406 (N_24406,N_24225,N_24333);
xor U24407 (N_24407,N_24305,N_24383);
xnor U24408 (N_24408,N_24315,N_24318);
or U24409 (N_24409,N_24223,N_24379);
nand U24410 (N_24410,N_24287,N_24266);
and U24411 (N_24411,N_24334,N_24367);
and U24412 (N_24412,N_24355,N_24281);
xnor U24413 (N_24413,N_24264,N_24216);
and U24414 (N_24414,N_24361,N_24375);
nand U24415 (N_24415,N_24337,N_24364);
nor U24416 (N_24416,N_24389,N_24262);
nand U24417 (N_24417,N_24344,N_24370);
or U24418 (N_24418,N_24203,N_24283);
and U24419 (N_24419,N_24329,N_24306);
and U24420 (N_24420,N_24200,N_24269);
or U24421 (N_24421,N_24254,N_24292);
xnor U24422 (N_24422,N_24356,N_24279);
nor U24423 (N_24423,N_24213,N_24303);
nand U24424 (N_24424,N_24335,N_24362);
xor U24425 (N_24425,N_24282,N_24257);
xor U24426 (N_24426,N_24301,N_24388);
or U24427 (N_24427,N_24360,N_24273);
xor U24428 (N_24428,N_24321,N_24365);
nand U24429 (N_24429,N_24323,N_24206);
or U24430 (N_24430,N_24382,N_24304);
and U24431 (N_24431,N_24296,N_24252);
or U24432 (N_24432,N_24218,N_24395);
and U24433 (N_24433,N_24231,N_24378);
xor U24434 (N_24434,N_24313,N_24299);
nand U24435 (N_24435,N_24276,N_24278);
and U24436 (N_24436,N_24272,N_24298);
nand U24437 (N_24437,N_24236,N_24307);
and U24438 (N_24438,N_24285,N_24235);
and U24439 (N_24439,N_24258,N_24268);
and U24440 (N_24440,N_24267,N_24221);
and U24441 (N_24441,N_24316,N_24357);
nand U24442 (N_24442,N_24393,N_24255);
nor U24443 (N_24443,N_24397,N_24309);
nand U24444 (N_24444,N_24241,N_24342);
nand U24445 (N_24445,N_24398,N_24336);
xnor U24446 (N_24446,N_24244,N_24208);
nor U24447 (N_24447,N_24302,N_24261);
nor U24448 (N_24448,N_24217,N_24271);
or U24449 (N_24449,N_24234,N_24341);
nor U24450 (N_24450,N_24256,N_24385);
nor U24451 (N_24451,N_24343,N_24376);
and U24452 (N_24452,N_24295,N_24246);
nor U24453 (N_24453,N_24274,N_24384);
and U24454 (N_24454,N_24347,N_24214);
or U24455 (N_24455,N_24249,N_24238);
or U24456 (N_24456,N_24399,N_24326);
and U24457 (N_24457,N_24265,N_24352);
or U24458 (N_24458,N_24359,N_24270);
and U24459 (N_24459,N_24259,N_24394);
nand U24460 (N_24460,N_24286,N_24319);
nand U24461 (N_24461,N_24366,N_24260);
nand U24462 (N_24462,N_24381,N_24320);
xnor U24463 (N_24463,N_24392,N_24350);
nor U24464 (N_24464,N_24215,N_24205);
or U24465 (N_24465,N_24339,N_24368);
nor U24466 (N_24466,N_24293,N_24387);
nand U24467 (N_24467,N_24290,N_24325);
and U24468 (N_24468,N_24243,N_24377);
and U24469 (N_24469,N_24317,N_24351);
nor U24470 (N_24470,N_24369,N_24291);
nor U24471 (N_24471,N_24311,N_24239);
or U24472 (N_24472,N_24374,N_24288);
xor U24473 (N_24473,N_24328,N_24226);
or U24474 (N_24474,N_24330,N_24228);
or U24475 (N_24475,N_24363,N_24227);
nor U24476 (N_24476,N_24212,N_24220);
or U24477 (N_24477,N_24391,N_24353);
or U24478 (N_24478,N_24209,N_24358);
xor U24479 (N_24479,N_24245,N_24277);
nor U24480 (N_24480,N_24251,N_24250);
nor U24481 (N_24481,N_24230,N_24233);
and U24482 (N_24482,N_24308,N_24371);
and U24483 (N_24483,N_24248,N_24312);
nor U24484 (N_24484,N_24348,N_24300);
or U24485 (N_24485,N_24222,N_24310);
and U24486 (N_24486,N_24253,N_24332);
and U24487 (N_24487,N_24314,N_24280);
nor U24488 (N_24488,N_24390,N_24327);
nor U24489 (N_24489,N_24237,N_24204);
and U24490 (N_24490,N_24242,N_24232);
and U24491 (N_24491,N_24349,N_24202);
or U24492 (N_24492,N_24322,N_24373);
and U24493 (N_24493,N_24210,N_24219);
and U24494 (N_24494,N_24372,N_24297);
nand U24495 (N_24495,N_24263,N_24201);
nor U24496 (N_24496,N_24380,N_24211);
and U24497 (N_24497,N_24289,N_24346);
and U24498 (N_24498,N_24224,N_24331);
nand U24499 (N_24499,N_24345,N_24386);
nor U24500 (N_24500,N_24202,N_24264);
and U24501 (N_24501,N_24293,N_24290);
and U24502 (N_24502,N_24241,N_24294);
and U24503 (N_24503,N_24206,N_24302);
xnor U24504 (N_24504,N_24353,N_24226);
and U24505 (N_24505,N_24334,N_24278);
or U24506 (N_24506,N_24271,N_24365);
nand U24507 (N_24507,N_24265,N_24384);
xnor U24508 (N_24508,N_24396,N_24211);
nand U24509 (N_24509,N_24205,N_24338);
nor U24510 (N_24510,N_24288,N_24285);
or U24511 (N_24511,N_24355,N_24236);
nand U24512 (N_24512,N_24243,N_24351);
nand U24513 (N_24513,N_24397,N_24365);
xnor U24514 (N_24514,N_24228,N_24376);
nor U24515 (N_24515,N_24299,N_24391);
nand U24516 (N_24516,N_24239,N_24348);
and U24517 (N_24517,N_24285,N_24345);
or U24518 (N_24518,N_24350,N_24278);
xor U24519 (N_24519,N_24384,N_24373);
xnor U24520 (N_24520,N_24332,N_24387);
and U24521 (N_24521,N_24314,N_24358);
or U24522 (N_24522,N_24261,N_24363);
or U24523 (N_24523,N_24234,N_24397);
or U24524 (N_24524,N_24355,N_24232);
nor U24525 (N_24525,N_24332,N_24361);
and U24526 (N_24526,N_24356,N_24221);
nor U24527 (N_24527,N_24248,N_24339);
or U24528 (N_24528,N_24324,N_24253);
and U24529 (N_24529,N_24291,N_24318);
nand U24530 (N_24530,N_24304,N_24272);
or U24531 (N_24531,N_24345,N_24205);
nand U24532 (N_24532,N_24360,N_24291);
nand U24533 (N_24533,N_24307,N_24226);
nor U24534 (N_24534,N_24257,N_24299);
or U24535 (N_24535,N_24278,N_24205);
xor U24536 (N_24536,N_24227,N_24370);
xnor U24537 (N_24537,N_24382,N_24274);
xor U24538 (N_24538,N_24260,N_24343);
or U24539 (N_24539,N_24387,N_24241);
nor U24540 (N_24540,N_24245,N_24284);
and U24541 (N_24541,N_24348,N_24269);
and U24542 (N_24542,N_24383,N_24205);
xnor U24543 (N_24543,N_24221,N_24282);
or U24544 (N_24544,N_24266,N_24296);
nand U24545 (N_24545,N_24288,N_24383);
xnor U24546 (N_24546,N_24264,N_24242);
nand U24547 (N_24547,N_24329,N_24393);
nand U24548 (N_24548,N_24258,N_24348);
xor U24549 (N_24549,N_24398,N_24275);
nor U24550 (N_24550,N_24343,N_24307);
nand U24551 (N_24551,N_24321,N_24294);
nand U24552 (N_24552,N_24206,N_24238);
nor U24553 (N_24553,N_24297,N_24324);
or U24554 (N_24554,N_24345,N_24369);
nand U24555 (N_24555,N_24296,N_24328);
xor U24556 (N_24556,N_24390,N_24370);
xnor U24557 (N_24557,N_24224,N_24234);
xor U24558 (N_24558,N_24350,N_24273);
and U24559 (N_24559,N_24227,N_24381);
or U24560 (N_24560,N_24381,N_24318);
or U24561 (N_24561,N_24263,N_24307);
or U24562 (N_24562,N_24252,N_24352);
or U24563 (N_24563,N_24352,N_24277);
nand U24564 (N_24564,N_24395,N_24364);
xnor U24565 (N_24565,N_24350,N_24204);
nand U24566 (N_24566,N_24200,N_24386);
and U24567 (N_24567,N_24226,N_24383);
nand U24568 (N_24568,N_24275,N_24337);
nand U24569 (N_24569,N_24319,N_24367);
xor U24570 (N_24570,N_24382,N_24302);
nor U24571 (N_24571,N_24204,N_24366);
or U24572 (N_24572,N_24327,N_24352);
or U24573 (N_24573,N_24292,N_24268);
xor U24574 (N_24574,N_24374,N_24365);
and U24575 (N_24575,N_24338,N_24212);
or U24576 (N_24576,N_24201,N_24248);
or U24577 (N_24577,N_24206,N_24210);
or U24578 (N_24578,N_24326,N_24324);
and U24579 (N_24579,N_24330,N_24295);
xor U24580 (N_24580,N_24286,N_24242);
nand U24581 (N_24581,N_24265,N_24296);
nor U24582 (N_24582,N_24224,N_24217);
and U24583 (N_24583,N_24388,N_24307);
or U24584 (N_24584,N_24246,N_24201);
nor U24585 (N_24585,N_24339,N_24333);
or U24586 (N_24586,N_24324,N_24394);
xnor U24587 (N_24587,N_24258,N_24231);
nor U24588 (N_24588,N_24297,N_24234);
nor U24589 (N_24589,N_24386,N_24347);
and U24590 (N_24590,N_24322,N_24272);
and U24591 (N_24591,N_24300,N_24258);
nor U24592 (N_24592,N_24211,N_24303);
or U24593 (N_24593,N_24362,N_24338);
nand U24594 (N_24594,N_24283,N_24209);
nor U24595 (N_24595,N_24370,N_24268);
xor U24596 (N_24596,N_24236,N_24340);
nand U24597 (N_24597,N_24395,N_24205);
xnor U24598 (N_24598,N_24227,N_24220);
and U24599 (N_24599,N_24216,N_24282);
nor U24600 (N_24600,N_24512,N_24518);
nand U24601 (N_24601,N_24531,N_24419);
nand U24602 (N_24602,N_24492,N_24465);
xor U24603 (N_24603,N_24573,N_24427);
or U24604 (N_24604,N_24469,N_24549);
nor U24605 (N_24605,N_24446,N_24451);
and U24606 (N_24606,N_24428,N_24527);
nand U24607 (N_24607,N_24410,N_24405);
xnor U24608 (N_24608,N_24424,N_24448);
nor U24609 (N_24609,N_24436,N_24420);
nand U24610 (N_24610,N_24430,N_24473);
and U24611 (N_24611,N_24443,N_24460);
or U24612 (N_24612,N_24514,N_24407);
xor U24613 (N_24613,N_24484,N_24541);
or U24614 (N_24614,N_24454,N_24523);
and U24615 (N_24615,N_24526,N_24572);
or U24616 (N_24616,N_24571,N_24552);
nor U24617 (N_24617,N_24429,N_24455);
nand U24618 (N_24618,N_24506,N_24592);
xor U24619 (N_24619,N_24548,N_24519);
and U24620 (N_24620,N_24432,N_24445);
and U24621 (N_24621,N_24599,N_24452);
xor U24622 (N_24622,N_24555,N_24488);
xnor U24623 (N_24623,N_24578,N_24494);
nor U24624 (N_24624,N_24564,N_24476);
and U24625 (N_24625,N_24516,N_24467);
and U24626 (N_24626,N_24595,N_24550);
nor U24627 (N_24627,N_24579,N_24404);
or U24628 (N_24628,N_24418,N_24498);
and U24629 (N_24629,N_24584,N_24447);
nor U24630 (N_24630,N_24528,N_24577);
nor U24631 (N_24631,N_24534,N_24400);
nand U24632 (N_24632,N_24504,N_24496);
nand U24633 (N_24633,N_24450,N_24524);
and U24634 (N_24634,N_24435,N_24487);
nand U24635 (N_24635,N_24547,N_24583);
or U24636 (N_24636,N_24456,N_24569);
xnor U24637 (N_24637,N_24440,N_24585);
and U24638 (N_24638,N_24414,N_24511);
xnor U24639 (N_24639,N_24520,N_24507);
or U24640 (N_24640,N_24489,N_24480);
nand U24641 (N_24641,N_24542,N_24590);
nand U24642 (N_24642,N_24551,N_24500);
xor U24643 (N_24643,N_24425,N_24543);
nor U24644 (N_24644,N_24475,N_24403);
or U24645 (N_24645,N_24491,N_24597);
xor U24646 (N_24646,N_24482,N_24457);
and U24647 (N_24647,N_24545,N_24556);
xnor U24648 (N_24648,N_24536,N_24563);
or U24649 (N_24649,N_24412,N_24529);
nand U24650 (N_24650,N_24561,N_24477);
and U24651 (N_24651,N_24463,N_24509);
and U24652 (N_24652,N_24434,N_24576);
nand U24653 (N_24653,N_24401,N_24553);
nor U24654 (N_24654,N_24513,N_24416);
or U24655 (N_24655,N_24406,N_24437);
nor U24656 (N_24656,N_24530,N_24537);
nand U24657 (N_24657,N_24411,N_24433);
xnor U24658 (N_24658,N_24483,N_24468);
xnor U24659 (N_24659,N_24567,N_24581);
and U24660 (N_24660,N_24438,N_24517);
nor U24661 (N_24661,N_24464,N_24409);
xor U24662 (N_24662,N_24408,N_24495);
nand U24663 (N_24663,N_24574,N_24589);
nand U24664 (N_24664,N_24580,N_24402);
nand U24665 (N_24665,N_24540,N_24413);
or U24666 (N_24666,N_24490,N_24485);
and U24667 (N_24667,N_24538,N_24522);
and U24668 (N_24668,N_24486,N_24544);
nand U24669 (N_24669,N_24591,N_24535);
nand U24670 (N_24670,N_24557,N_24449);
or U24671 (N_24671,N_24417,N_24479);
xor U24672 (N_24672,N_24565,N_24558);
xnor U24673 (N_24673,N_24415,N_24532);
nand U24674 (N_24674,N_24466,N_24423);
nor U24675 (N_24675,N_24586,N_24470);
or U24676 (N_24676,N_24501,N_24525);
xnor U24677 (N_24677,N_24575,N_24499);
nor U24678 (N_24678,N_24588,N_24594);
or U24679 (N_24679,N_24503,N_24442);
nor U24680 (N_24680,N_24431,N_24497);
or U24681 (N_24681,N_24453,N_24539);
nand U24682 (N_24682,N_24439,N_24598);
nor U24683 (N_24683,N_24510,N_24461);
or U24684 (N_24684,N_24582,N_24508);
and U24685 (N_24685,N_24546,N_24587);
nand U24686 (N_24686,N_24441,N_24478);
nor U24687 (N_24687,N_24422,N_24481);
nand U24688 (N_24688,N_24459,N_24471);
nor U24689 (N_24689,N_24596,N_24502);
xnor U24690 (N_24690,N_24554,N_24515);
nor U24691 (N_24691,N_24474,N_24426);
nor U24692 (N_24692,N_24560,N_24521);
nor U24693 (N_24693,N_24444,N_24462);
and U24694 (N_24694,N_24559,N_24593);
nand U24695 (N_24695,N_24533,N_24505);
nand U24696 (N_24696,N_24562,N_24493);
nand U24697 (N_24697,N_24570,N_24458);
xnor U24698 (N_24698,N_24472,N_24421);
nand U24699 (N_24699,N_24568,N_24566);
xor U24700 (N_24700,N_24498,N_24425);
xor U24701 (N_24701,N_24413,N_24578);
xnor U24702 (N_24702,N_24566,N_24598);
or U24703 (N_24703,N_24533,N_24564);
nand U24704 (N_24704,N_24490,N_24579);
nand U24705 (N_24705,N_24555,N_24427);
nand U24706 (N_24706,N_24556,N_24415);
xnor U24707 (N_24707,N_24506,N_24570);
nand U24708 (N_24708,N_24497,N_24458);
nor U24709 (N_24709,N_24578,N_24597);
or U24710 (N_24710,N_24471,N_24566);
or U24711 (N_24711,N_24511,N_24577);
nand U24712 (N_24712,N_24478,N_24452);
nor U24713 (N_24713,N_24567,N_24445);
xor U24714 (N_24714,N_24476,N_24541);
nor U24715 (N_24715,N_24522,N_24407);
or U24716 (N_24716,N_24460,N_24426);
nor U24717 (N_24717,N_24572,N_24412);
nor U24718 (N_24718,N_24533,N_24577);
and U24719 (N_24719,N_24465,N_24464);
and U24720 (N_24720,N_24453,N_24543);
and U24721 (N_24721,N_24594,N_24465);
nand U24722 (N_24722,N_24424,N_24470);
and U24723 (N_24723,N_24443,N_24495);
and U24724 (N_24724,N_24476,N_24486);
or U24725 (N_24725,N_24480,N_24496);
nor U24726 (N_24726,N_24518,N_24483);
nor U24727 (N_24727,N_24422,N_24536);
nor U24728 (N_24728,N_24447,N_24500);
xnor U24729 (N_24729,N_24442,N_24437);
nor U24730 (N_24730,N_24424,N_24549);
and U24731 (N_24731,N_24480,N_24504);
nand U24732 (N_24732,N_24549,N_24407);
xnor U24733 (N_24733,N_24464,N_24439);
and U24734 (N_24734,N_24435,N_24518);
and U24735 (N_24735,N_24446,N_24518);
nand U24736 (N_24736,N_24508,N_24593);
and U24737 (N_24737,N_24513,N_24509);
and U24738 (N_24738,N_24430,N_24551);
or U24739 (N_24739,N_24478,N_24566);
and U24740 (N_24740,N_24436,N_24495);
xor U24741 (N_24741,N_24490,N_24460);
and U24742 (N_24742,N_24472,N_24423);
nor U24743 (N_24743,N_24532,N_24493);
and U24744 (N_24744,N_24534,N_24467);
or U24745 (N_24745,N_24407,N_24422);
or U24746 (N_24746,N_24593,N_24455);
xnor U24747 (N_24747,N_24542,N_24546);
or U24748 (N_24748,N_24552,N_24461);
nand U24749 (N_24749,N_24489,N_24497);
or U24750 (N_24750,N_24439,N_24470);
or U24751 (N_24751,N_24501,N_24537);
or U24752 (N_24752,N_24503,N_24402);
or U24753 (N_24753,N_24429,N_24569);
xor U24754 (N_24754,N_24450,N_24484);
and U24755 (N_24755,N_24598,N_24462);
nor U24756 (N_24756,N_24576,N_24487);
or U24757 (N_24757,N_24498,N_24507);
or U24758 (N_24758,N_24565,N_24570);
or U24759 (N_24759,N_24507,N_24405);
nor U24760 (N_24760,N_24569,N_24415);
nor U24761 (N_24761,N_24405,N_24429);
xor U24762 (N_24762,N_24522,N_24586);
nand U24763 (N_24763,N_24535,N_24433);
xnor U24764 (N_24764,N_24445,N_24435);
xor U24765 (N_24765,N_24484,N_24473);
or U24766 (N_24766,N_24493,N_24523);
nand U24767 (N_24767,N_24531,N_24548);
and U24768 (N_24768,N_24433,N_24473);
and U24769 (N_24769,N_24534,N_24524);
nand U24770 (N_24770,N_24570,N_24569);
nand U24771 (N_24771,N_24400,N_24439);
nor U24772 (N_24772,N_24525,N_24508);
nand U24773 (N_24773,N_24532,N_24498);
xor U24774 (N_24774,N_24415,N_24418);
xnor U24775 (N_24775,N_24508,N_24437);
and U24776 (N_24776,N_24570,N_24541);
or U24777 (N_24777,N_24498,N_24540);
nor U24778 (N_24778,N_24504,N_24495);
nand U24779 (N_24779,N_24489,N_24560);
xor U24780 (N_24780,N_24410,N_24431);
or U24781 (N_24781,N_24599,N_24416);
or U24782 (N_24782,N_24583,N_24573);
nor U24783 (N_24783,N_24437,N_24513);
nor U24784 (N_24784,N_24579,N_24452);
nor U24785 (N_24785,N_24566,N_24532);
nand U24786 (N_24786,N_24421,N_24504);
xor U24787 (N_24787,N_24555,N_24583);
xnor U24788 (N_24788,N_24480,N_24442);
or U24789 (N_24789,N_24599,N_24542);
nor U24790 (N_24790,N_24505,N_24591);
or U24791 (N_24791,N_24457,N_24418);
nand U24792 (N_24792,N_24513,N_24586);
xor U24793 (N_24793,N_24500,N_24591);
or U24794 (N_24794,N_24458,N_24517);
nand U24795 (N_24795,N_24519,N_24553);
xor U24796 (N_24796,N_24564,N_24408);
and U24797 (N_24797,N_24595,N_24567);
nand U24798 (N_24798,N_24500,N_24575);
xor U24799 (N_24799,N_24464,N_24567);
nand U24800 (N_24800,N_24702,N_24732);
nand U24801 (N_24801,N_24787,N_24601);
or U24802 (N_24802,N_24723,N_24794);
nor U24803 (N_24803,N_24775,N_24687);
nand U24804 (N_24804,N_24634,N_24665);
and U24805 (N_24805,N_24609,N_24683);
and U24806 (N_24806,N_24790,N_24606);
or U24807 (N_24807,N_24777,N_24776);
or U24808 (N_24808,N_24624,N_24604);
nor U24809 (N_24809,N_24742,N_24792);
or U24810 (N_24810,N_24641,N_24797);
nand U24811 (N_24811,N_24663,N_24664);
nor U24812 (N_24812,N_24607,N_24786);
nor U24813 (N_24813,N_24636,N_24671);
or U24814 (N_24814,N_24645,N_24713);
nor U24815 (N_24815,N_24795,N_24791);
nor U24816 (N_24816,N_24615,N_24623);
nand U24817 (N_24817,N_24639,N_24744);
nand U24818 (N_24818,N_24751,N_24774);
and U24819 (N_24819,N_24640,N_24709);
and U24820 (N_24820,N_24763,N_24772);
or U24821 (N_24821,N_24685,N_24686);
or U24822 (N_24822,N_24660,N_24614);
nor U24823 (N_24823,N_24613,N_24753);
and U24824 (N_24824,N_24661,N_24632);
and U24825 (N_24825,N_24612,N_24755);
nor U24826 (N_24826,N_24779,N_24629);
or U24827 (N_24827,N_24611,N_24712);
xor U24828 (N_24828,N_24616,N_24711);
or U24829 (N_24829,N_24635,N_24745);
nor U24830 (N_24830,N_24789,N_24602);
or U24831 (N_24831,N_24621,N_24691);
nor U24832 (N_24832,N_24720,N_24778);
xnor U24833 (N_24833,N_24741,N_24637);
or U24834 (N_24834,N_24669,N_24701);
or U24835 (N_24835,N_24750,N_24788);
xor U24836 (N_24836,N_24680,N_24708);
nor U24837 (N_24837,N_24650,N_24649);
and U24838 (N_24838,N_24655,N_24603);
and U24839 (N_24839,N_24688,N_24656);
or U24840 (N_24840,N_24674,N_24676);
nor U24841 (N_24841,N_24608,N_24785);
xor U24842 (N_24842,N_24622,N_24766);
xnor U24843 (N_24843,N_24796,N_24662);
nor U24844 (N_24844,N_24678,N_24717);
nor U24845 (N_24845,N_24705,N_24600);
or U24846 (N_24846,N_24798,N_24773);
nor U24847 (N_24847,N_24710,N_24667);
nand U24848 (N_24848,N_24625,N_24679);
nand U24849 (N_24849,N_24738,N_24716);
nand U24850 (N_24850,N_24781,N_24756);
nor U24851 (N_24851,N_24700,N_24689);
and U24852 (N_24852,N_24721,N_24644);
or U24853 (N_24853,N_24731,N_24771);
or U24854 (N_24854,N_24677,N_24758);
and U24855 (N_24855,N_24737,N_24743);
xor U24856 (N_24856,N_24715,N_24668);
nand U24857 (N_24857,N_24768,N_24722);
xnor U24858 (N_24858,N_24724,N_24695);
or U24859 (N_24859,N_24651,N_24770);
nand U24860 (N_24860,N_24648,N_24659);
or U24861 (N_24861,N_24675,N_24799);
nand U24862 (N_24862,N_24699,N_24767);
nor U24863 (N_24863,N_24620,N_24749);
or U24864 (N_24864,N_24682,N_24793);
or U24865 (N_24865,N_24706,N_24626);
or U24866 (N_24866,N_24681,N_24714);
or U24867 (N_24867,N_24617,N_24734);
nor U24868 (N_24868,N_24765,N_24754);
or U24869 (N_24869,N_24725,N_24666);
or U24870 (N_24870,N_24692,N_24654);
xnor U24871 (N_24871,N_24698,N_24752);
nand U24872 (N_24872,N_24704,N_24757);
nand U24873 (N_24873,N_24739,N_24647);
xor U24874 (N_24874,N_24761,N_24673);
nand U24875 (N_24875,N_24719,N_24782);
nor U24876 (N_24876,N_24670,N_24638);
xnor U24877 (N_24877,N_24653,N_24633);
nor U24878 (N_24878,N_24630,N_24759);
xnor U24879 (N_24879,N_24736,N_24627);
or U24880 (N_24880,N_24610,N_24733);
nor U24881 (N_24881,N_24652,N_24619);
nand U24882 (N_24882,N_24628,N_24740);
nor U24883 (N_24883,N_24728,N_24707);
and U24884 (N_24884,N_24642,N_24727);
or U24885 (N_24885,N_24703,N_24726);
and U24886 (N_24886,N_24784,N_24693);
xor U24887 (N_24887,N_24780,N_24746);
nor U24888 (N_24888,N_24657,N_24631);
nand U24889 (N_24889,N_24694,N_24760);
nor U24890 (N_24890,N_24684,N_24646);
nand U24891 (N_24891,N_24729,N_24769);
xor U24892 (N_24892,N_24697,N_24762);
nor U24893 (N_24893,N_24690,N_24748);
nand U24894 (N_24894,N_24696,N_24658);
xor U24895 (N_24895,N_24747,N_24730);
and U24896 (N_24896,N_24764,N_24605);
nand U24897 (N_24897,N_24672,N_24783);
nor U24898 (N_24898,N_24643,N_24718);
nand U24899 (N_24899,N_24618,N_24735);
xnor U24900 (N_24900,N_24775,N_24766);
and U24901 (N_24901,N_24639,N_24687);
or U24902 (N_24902,N_24749,N_24619);
xor U24903 (N_24903,N_24672,N_24615);
and U24904 (N_24904,N_24659,N_24628);
and U24905 (N_24905,N_24607,N_24614);
or U24906 (N_24906,N_24765,N_24743);
or U24907 (N_24907,N_24693,N_24772);
nand U24908 (N_24908,N_24774,N_24626);
xnor U24909 (N_24909,N_24782,N_24793);
nor U24910 (N_24910,N_24775,N_24790);
nand U24911 (N_24911,N_24702,N_24613);
and U24912 (N_24912,N_24783,N_24768);
xor U24913 (N_24913,N_24667,N_24624);
nor U24914 (N_24914,N_24690,N_24630);
or U24915 (N_24915,N_24613,N_24734);
and U24916 (N_24916,N_24687,N_24770);
nor U24917 (N_24917,N_24706,N_24649);
and U24918 (N_24918,N_24715,N_24797);
nor U24919 (N_24919,N_24795,N_24670);
nand U24920 (N_24920,N_24692,N_24764);
xor U24921 (N_24921,N_24623,N_24694);
xor U24922 (N_24922,N_24662,N_24654);
xor U24923 (N_24923,N_24721,N_24687);
nand U24924 (N_24924,N_24677,N_24674);
or U24925 (N_24925,N_24795,N_24749);
nor U24926 (N_24926,N_24753,N_24794);
or U24927 (N_24927,N_24690,N_24717);
and U24928 (N_24928,N_24782,N_24798);
xnor U24929 (N_24929,N_24766,N_24685);
nor U24930 (N_24930,N_24728,N_24787);
and U24931 (N_24931,N_24626,N_24759);
xor U24932 (N_24932,N_24722,N_24687);
xnor U24933 (N_24933,N_24603,N_24791);
or U24934 (N_24934,N_24672,N_24665);
and U24935 (N_24935,N_24783,N_24693);
nor U24936 (N_24936,N_24643,N_24784);
nor U24937 (N_24937,N_24734,N_24631);
nor U24938 (N_24938,N_24704,N_24614);
or U24939 (N_24939,N_24627,N_24733);
xnor U24940 (N_24940,N_24610,N_24692);
nor U24941 (N_24941,N_24762,N_24752);
or U24942 (N_24942,N_24667,N_24793);
nor U24943 (N_24943,N_24745,N_24731);
and U24944 (N_24944,N_24610,N_24708);
and U24945 (N_24945,N_24697,N_24702);
nor U24946 (N_24946,N_24613,N_24627);
nand U24947 (N_24947,N_24612,N_24739);
nor U24948 (N_24948,N_24711,N_24762);
nor U24949 (N_24949,N_24603,N_24619);
xor U24950 (N_24950,N_24648,N_24725);
and U24951 (N_24951,N_24798,N_24690);
or U24952 (N_24952,N_24782,N_24775);
xor U24953 (N_24953,N_24620,N_24653);
or U24954 (N_24954,N_24740,N_24625);
and U24955 (N_24955,N_24761,N_24709);
nand U24956 (N_24956,N_24777,N_24769);
nor U24957 (N_24957,N_24726,N_24759);
or U24958 (N_24958,N_24712,N_24681);
or U24959 (N_24959,N_24651,N_24641);
or U24960 (N_24960,N_24733,N_24668);
nand U24961 (N_24961,N_24642,N_24662);
nand U24962 (N_24962,N_24767,N_24790);
nand U24963 (N_24963,N_24749,N_24651);
nor U24964 (N_24964,N_24614,N_24604);
nor U24965 (N_24965,N_24626,N_24649);
and U24966 (N_24966,N_24762,N_24686);
nand U24967 (N_24967,N_24685,N_24742);
nand U24968 (N_24968,N_24717,N_24788);
nand U24969 (N_24969,N_24624,N_24766);
or U24970 (N_24970,N_24621,N_24721);
nor U24971 (N_24971,N_24668,N_24644);
or U24972 (N_24972,N_24611,N_24663);
nor U24973 (N_24973,N_24690,N_24781);
or U24974 (N_24974,N_24756,N_24648);
and U24975 (N_24975,N_24775,N_24740);
nand U24976 (N_24976,N_24712,N_24716);
or U24977 (N_24977,N_24672,N_24685);
and U24978 (N_24978,N_24733,N_24712);
or U24979 (N_24979,N_24649,N_24681);
xor U24980 (N_24980,N_24736,N_24728);
xnor U24981 (N_24981,N_24799,N_24720);
xor U24982 (N_24982,N_24655,N_24747);
nand U24983 (N_24983,N_24793,N_24758);
xnor U24984 (N_24984,N_24758,N_24689);
or U24985 (N_24985,N_24633,N_24738);
nand U24986 (N_24986,N_24765,N_24679);
and U24987 (N_24987,N_24714,N_24759);
and U24988 (N_24988,N_24737,N_24640);
nand U24989 (N_24989,N_24660,N_24758);
or U24990 (N_24990,N_24710,N_24642);
xor U24991 (N_24991,N_24657,N_24738);
nor U24992 (N_24992,N_24605,N_24666);
nor U24993 (N_24993,N_24732,N_24668);
nand U24994 (N_24994,N_24780,N_24683);
nand U24995 (N_24995,N_24618,N_24783);
and U24996 (N_24996,N_24664,N_24737);
nor U24997 (N_24997,N_24724,N_24699);
nand U24998 (N_24998,N_24756,N_24604);
nor U24999 (N_24999,N_24773,N_24766);
nor UO_0 (O_0,N_24856,N_24876);
xor UO_1 (O_1,N_24961,N_24878);
nand UO_2 (O_2,N_24820,N_24858);
nor UO_3 (O_3,N_24921,N_24995);
nand UO_4 (O_4,N_24854,N_24932);
or UO_5 (O_5,N_24885,N_24819);
and UO_6 (O_6,N_24974,N_24803);
and UO_7 (O_7,N_24825,N_24865);
or UO_8 (O_8,N_24866,N_24840);
and UO_9 (O_9,N_24928,N_24907);
xor UO_10 (O_10,N_24835,N_24807);
xor UO_11 (O_11,N_24908,N_24852);
or UO_12 (O_12,N_24801,N_24813);
or UO_13 (O_13,N_24849,N_24903);
and UO_14 (O_14,N_24844,N_24979);
nand UO_15 (O_15,N_24843,N_24897);
xor UO_16 (O_16,N_24947,N_24900);
nand UO_17 (O_17,N_24906,N_24926);
or UO_18 (O_18,N_24971,N_24923);
or UO_19 (O_19,N_24955,N_24954);
or UO_20 (O_20,N_24817,N_24957);
or UO_21 (O_21,N_24983,N_24806);
or UO_22 (O_22,N_24821,N_24829);
xnor UO_23 (O_23,N_24833,N_24892);
xor UO_24 (O_24,N_24952,N_24940);
nor UO_25 (O_25,N_24826,N_24924);
xnor UO_26 (O_26,N_24999,N_24818);
nand UO_27 (O_27,N_24816,N_24902);
nor UO_28 (O_28,N_24901,N_24815);
nand UO_29 (O_29,N_24977,N_24989);
nand UO_30 (O_30,N_24836,N_24981);
or UO_31 (O_31,N_24920,N_24934);
xor UO_32 (O_32,N_24860,N_24905);
nor UO_33 (O_33,N_24883,N_24972);
or UO_34 (O_34,N_24822,N_24808);
xnor UO_35 (O_35,N_24848,N_24839);
or UO_36 (O_36,N_24873,N_24916);
nand UO_37 (O_37,N_24964,N_24889);
or UO_38 (O_38,N_24863,N_24986);
or UO_39 (O_39,N_24811,N_24824);
or UO_40 (O_40,N_24967,N_24851);
nand UO_41 (O_41,N_24935,N_24992);
or UO_42 (O_42,N_24890,N_24944);
nand UO_43 (O_43,N_24917,N_24870);
nor UO_44 (O_44,N_24978,N_24948);
xnor UO_45 (O_45,N_24909,N_24953);
or UO_46 (O_46,N_24973,N_24842);
nor UO_47 (O_47,N_24894,N_24918);
or UO_48 (O_48,N_24927,N_24874);
and UO_49 (O_49,N_24800,N_24846);
nor UO_50 (O_50,N_24936,N_24888);
nor UO_51 (O_51,N_24975,N_24845);
xnor UO_52 (O_52,N_24879,N_24984);
nor UO_53 (O_53,N_24956,N_24832);
nand UO_54 (O_54,N_24875,N_24886);
nand UO_55 (O_55,N_24976,N_24834);
nand UO_56 (O_56,N_24862,N_24922);
xor UO_57 (O_57,N_24869,N_24855);
and UO_58 (O_58,N_24871,N_24881);
nand UO_59 (O_59,N_24904,N_24831);
and UO_60 (O_60,N_24830,N_24857);
or UO_61 (O_61,N_24861,N_24930);
nand UO_62 (O_62,N_24962,N_24910);
or UO_63 (O_63,N_24837,N_24912);
and UO_64 (O_64,N_24805,N_24893);
nor UO_65 (O_65,N_24877,N_24994);
nor UO_66 (O_66,N_24823,N_24958);
xor UO_67 (O_67,N_24943,N_24827);
or UO_68 (O_68,N_24991,N_24993);
or UO_69 (O_69,N_24949,N_24915);
or UO_70 (O_70,N_24996,N_24945);
xor UO_71 (O_71,N_24941,N_24828);
xor UO_72 (O_72,N_24887,N_24929);
nor UO_73 (O_73,N_24931,N_24859);
and UO_74 (O_74,N_24970,N_24997);
nand UO_75 (O_75,N_24937,N_24914);
and UO_76 (O_76,N_24899,N_24872);
and UO_77 (O_77,N_24853,N_24960);
xor UO_78 (O_78,N_24850,N_24802);
nor UO_79 (O_79,N_24847,N_24884);
nor UO_80 (O_80,N_24987,N_24867);
and UO_81 (O_81,N_24864,N_24950);
and UO_82 (O_82,N_24919,N_24809);
xnor UO_83 (O_83,N_24968,N_24939);
or UO_84 (O_84,N_24959,N_24988);
xnor UO_85 (O_85,N_24969,N_24804);
nor UO_86 (O_86,N_24810,N_24882);
xor UO_87 (O_87,N_24980,N_24998);
and UO_88 (O_88,N_24895,N_24946);
nor UO_89 (O_89,N_24868,N_24942);
nand UO_90 (O_90,N_24938,N_24990);
or UO_91 (O_91,N_24911,N_24965);
or UO_92 (O_92,N_24933,N_24812);
or UO_93 (O_93,N_24982,N_24814);
nor UO_94 (O_94,N_24891,N_24963);
nand UO_95 (O_95,N_24925,N_24966);
and UO_96 (O_96,N_24841,N_24985);
nor UO_97 (O_97,N_24913,N_24838);
and UO_98 (O_98,N_24898,N_24951);
nand UO_99 (O_99,N_24896,N_24880);
and UO_100 (O_100,N_24849,N_24927);
xnor UO_101 (O_101,N_24990,N_24853);
or UO_102 (O_102,N_24910,N_24879);
or UO_103 (O_103,N_24844,N_24988);
xnor UO_104 (O_104,N_24864,N_24841);
or UO_105 (O_105,N_24945,N_24826);
xor UO_106 (O_106,N_24878,N_24855);
nor UO_107 (O_107,N_24836,N_24868);
nand UO_108 (O_108,N_24893,N_24957);
nor UO_109 (O_109,N_24891,N_24995);
nor UO_110 (O_110,N_24933,N_24841);
nor UO_111 (O_111,N_24928,N_24911);
nand UO_112 (O_112,N_24913,N_24934);
nand UO_113 (O_113,N_24886,N_24980);
nor UO_114 (O_114,N_24909,N_24832);
xor UO_115 (O_115,N_24965,N_24994);
and UO_116 (O_116,N_24845,N_24822);
xnor UO_117 (O_117,N_24870,N_24974);
nand UO_118 (O_118,N_24819,N_24943);
xor UO_119 (O_119,N_24968,N_24870);
nand UO_120 (O_120,N_24859,N_24924);
nor UO_121 (O_121,N_24972,N_24800);
xor UO_122 (O_122,N_24950,N_24800);
xnor UO_123 (O_123,N_24908,N_24823);
nor UO_124 (O_124,N_24874,N_24992);
or UO_125 (O_125,N_24858,N_24826);
nand UO_126 (O_126,N_24857,N_24874);
nand UO_127 (O_127,N_24991,N_24960);
and UO_128 (O_128,N_24847,N_24905);
or UO_129 (O_129,N_24875,N_24919);
xnor UO_130 (O_130,N_24922,N_24964);
and UO_131 (O_131,N_24971,N_24916);
xor UO_132 (O_132,N_24974,N_24859);
xnor UO_133 (O_133,N_24822,N_24847);
nor UO_134 (O_134,N_24829,N_24899);
nand UO_135 (O_135,N_24849,N_24864);
or UO_136 (O_136,N_24820,N_24852);
xor UO_137 (O_137,N_24981,N_24951);
xnor UO_138 (O_138,N_24956,N_24803);
nor UO_139 (O_139,N_24975,N_24808);
or UO_140 (O_140,N_24823,N_24980);
and UO_141 (O_141,N_24864,N_24839);
nand UO_142 (O_142,N_24842,N_24862);
xor UO_143 (O_143,N_24888,N_24945);
and UO_144 (O_144,N_24957,N_24826);
nor UO_145 (O_145,N_24866,N_24935);
or UO_146 (O_146,N_24852,N_24835);
nand UO_147 (O_147,N_24822,N_24900);
nand UO_148 (O_148,N_24898,N_24939);
and UO_149 (O_149,N_24830,N_24854);
or UO_150 (O_150,N_24903,N_24830);
nor UO_151 (O_151,N_24914,N_24891);
and UO_152 (O_152,N_24901,N_24928);
nor UO_153 (O_153,N_24941,N_24892);
xnor UO_154 (O_154,N_24893,N_24969);
nand UO_155 (O_155,N_24932,N_24946);
or UO_156 (O_156,N_24971,N_24863);
xor UO_157 (O_157,N_24860,N_24995);
nor UO_158 (O_158,N_24982,N_24989);
xor UO_159 (O_159,N_24992,N_24997);
nor UO_160 (O_160,N_24968,N_24881);
or UO_161 (O_161,N_24924,N_24951);
and UO_162 (O_162,N_24827,N_24852);
and UO_163 (O_163,N_24941,N_24975);
nand UO_164 (O_164,N_24942,N_24858);
xor UO_165 (O_165,N_24960,N_24893);
and UO_166 (O_166,N_24901,N_24826);
xnor UO_167 (O_167,N_24858,N_24811);
or UO_168 (O_168,N_24883,N_24879);
and UO_169 (O_169,N_24893,N_24875);
nand UO_170 (O_170,N_24858,N_24860);
or UO_171 (O_171,N_24848,N_24825);
and UO_172 (O_172,N_24811,N_24902);
nand UO_173 (O_173,N_24810,N_24951);
nand UO_174 (O_174,N_24920,N_24849);
nand UO_175 (O_175,N_24903,N_24804);
or UO_176 (O_176,N_24912,N_24948);
xor UO_177 (O_177,N_24993,N_24963);
and UO_178 (O_178,N_24869,N_24868);
or UO_179 (O_179,N_24856,N_24888);
nor UO_180 (O_180,N_24960,N_24802);
and UO_181 (O_181,N_24838,N_24910);
and UO_182 (O_182,N_24876,N_24859);
xor UO_183 (O_183,N_24815,N_24966);
xnor UO_184 (O_184,N_24927,N_24859);
nand UO_185 (O_185,N_24889,N_24849);
or UO_186 (O_186,N_24985,N_24995);
nor UO_187 (O_187,N_24861,N_24896);
or UO_188 (O_188,N_24987,N_24850);
nor UO_189 (O_189,N_24851,N_24864);
nor UO_190 (O_190,N_24801,N_24805);
or UO_191 (O_191,N_24883,N_24982);
nor UO_192 (O_192,N_24839,N_24842);
nand UO_193 (O_193,N_24849,N_24916);
or UO_194 (O_194,N_24820,N_24928);
or UO_195 (O_195,N_24870,N_24929);
or UO_196 (O_196,N_24880,N_24953);
nor UO_197 (O_197,N_24969,N_24946);
and UO_198 (O_198,N_24877,N_24881);
or UO_199 (O_199,N_24856,N_24813);
nand UO_200 (O_200,N_24974,N_24928);
and UO_201 (O_201,N_24821,N_24897);
nand UO_202 (O_202,N_24995,N_24905);
and UO_203 (O_203,N_24955,N_24971);
xor UO_204 (O_204,N_24990,N_24996);
nor UO_205 (O_205,N_24901,N_24809);
xor UO_206 (O_206,N_24865,N_24967);
or UO_207 (O_207,N_24801,N_24899);
xnor UO_208 (O_208,N_24990,N_24988);
nand UO_209 (O_209,N_24996,N_24906);
xor UO_210 (O_210,N_24857,N_24901);
nand UO_211 (O_211,N_24915,N_24944);
and UO_212 (O_212,N_24926,N_24841);
nor UO_213 (O_213,N_24872,N_24957);
and UO_214 (O_214,N_24978,N_24864);
and UO_215 (O_215,N_24808,N_24820);
nand UO_216 (O_216,N_24902,N_24956);
or UO_217 (O_217,N_24862,N_24865);
or UO_218 (O_218,N_24982,N_24926);
and UO_219 (O_219,N_24863,N_24821);
or UO_220 (O_220,N_24812,N_24843);
nand UO_221 (O_221,N_24946,N_24862);
nor UO_222 (O_222,N_24824,N_24964);
or UO_223 (O_223,N_24810,N_24955);
nor UO_224 (O_224,N_24866,N_24805);
nor UO_225 (O_225,N_24946,N_24801);
xor UO_226 (O_226,N_24983,N_24829);
and UO_227 (O_227,N_24851,N_24858);
xnor UO_228 (O_228,N_24942,N_24885);
or UO_229 (O_229,N_24867,N_24836);
xor UO_230 (O_230,N_24929,N_24908);
xnor UO_231 (O_231,N_24884,N_24994);
and UO_232 (O_232,N_24938,N_24918);
xnor UO_233 (O_233,N_24804,N_24818);
nand UO_234 (O_234,N_24817,N_24811);
or UO_235 (O_235,N_24966,N_24986);
nor UO_236 (O_236,N_24801,N_24933);
or UO_237 (O_237,N_24942,N_24850);
nor UO_238 (O_238,N_24964,N_24987);
or UO_239 (O_239,N_24890,N_24984);
nand UO_240 (O_240,N_24861,N_24947);
xor UO_241 (O_241,N_24939,N_24992);
or UO_242 (O_242,N_24946,N_24829);
nor UO_243 (O_243,N_24966,N_24826);
or UO_244 (O_244,N_24881,N_24875);
or UO_245 (O_245,N_24888,N_24939);
nor UO_246 (O_246,N_24955,N_24909);
nor UO_247 (O_247,N_24910,N_24898);
nand UO_248 (O_248,N_24954,N_24812);
and UO_249 (O_249,N_24955,N_24960);
xor UO_250 (O_250,N_24808,N_24907);
nand UO_251 (O_251,N_24958,N_24884);
or UO_252 (O_252,N_24984,N_24908);
or UO_253 (O_253,N_24802,N_24832);
and UO_254 (O_254,N_24936,N_24926);
xor UO_255 (O_255,N_24887,N_24979);
nor UO_256 (O_256,N_24966,N_24850);
xnor UO_257 (O_257,N_24861,N_24853);
nor UO_258 (O_258,N_24943,N_24959);
and UO_259 (O_259,N_24819,N_24800);
and UO_260 (O_260,N_24968,N_24950);
or UO_261 (O_261,N_24804,N_24857);
or UO_262 (O_262,N_24860,N_24812);
nand UO_263 (O_263,N_24926,N_24820);
nand UO_264 (O_264,N_24829,N_24813);
or UO_265 (O_265,N_24965,N_24822);
xnor UO_266 (O_266,N_24919,N_24983);
nand UO_267 (O_267,N_24907,N_24823);
nor UO_268 (O_268,N_24886,N_24958);
nand UO_269 (O_269,N_24976,N_24871);
nand UO_270 (O_270,N_24936,N_24871);
and UO_271 (O_271,N_24973,N_24869);
nand UO_272 (O_272,N_24941,N_24980);
and UO_273 (O_273,N_24997,N_24899);
or UO_274 (O_274,N_24877,N_24870);
nor UO_275 (O_275,N_24957,N_24979);
and UO_276 (O_276,N_24947,N_24866);
nand UO_277 (O_277,N_24860,N_24935);
nor UO_278 (O_278,N_24946,N_24863);
nand UO_279 (O_279,N_24846,N_24925);
nand UO_280 (O_280,N_24872,N_24878);
or UO_281 (O_281,N_24901,N_24962);
nand UO_282 (O_282,N_24833,N_24834);
and UO_283 (O_283,N_24826,N_24946);
nand UO_284 (O_284,N_24907,N_24870);
nor UO_285 (O_285,N_24990,N_24830);
nand UO_286 (O_286,N_24942,N_24908);
and UO_287 (O_287,N_24828,N_24980);
and UO_288 (O_288,N_24866,N_24880);
and UO_289 (O_289,N_24818,N_24986);
or UO_290 (O_290,N_24846,N_24983);
xor UO_291 (O_291,N_24997,N_24826);
or UO_292 (O_292,N_24920,N_24900);
or UO_293 (O_293,N_24899,N_24851);
nand UO_294 (O_294,N_24820,N_24822);
or UO_295 (O_295,N_24884,N_24899);
nand UO_296 (O_296,N_24885,N_24822);
nor UO_297 (O_297,N_24889,N_24832);
or UO_298 (O_298,N_24825,N_24997);
xnor UO_299 (O_299,N_24963,N_24996);
or UO_300 (O_300,N_24991,N_24929);
nand UO_301 (O_301,N_24846,N_24902);
or UO_302 (O_302,N_24900,N_24825);
or UO_303 (O_303,N_24913,N_24920);
nor UO_304 (O_304,N_24951,N_24950);
or UO_305 (O_305,N_24857,N_24835);
and UO_306 (O_306,N_24986,N_24830);
and UO_307 (O_307,N_24855,N_24888);
xor UO_308 (O_308,N_24935,N_24955);
and UO_309 (O_309,N_24846,N_24945);
xnor UO_310 (O_310,N_24938,N_24944);
xnor UO_311 (O_311,N_24923,N_24862);
or UO_312 (O_312,N_24988,N_24826);
nor UO_313 (O_313,N_24989,N_24855);
nand UO_314 (O_314,N_24998,N_24897);
nor UO_315 (O_315,N_24938,N_24833);
nor UO_316 (O_316,N_24838,N_24934);
xor UO_317 (O_317,N_24949,N_24883);
nand UO_318 (O_318,N_24808,N_24961);
and UO_319 (O_319,N_24975,N_24997);
xnor UO_320 (O_320,N_24993,N_24962);
xnor UO_321 (O_321,N_24854,N_24983);
or UO_322 (O_322,N_24913,N_24967);
nor UO_323 (O_323,N_24932,N_24813);
or UO_324 (O_324,N_24899,N_24982);
nor UO_325 (O_325,N_24985,N_24971);
nor UO_326 (O_326,N_24891,N_24909);
and UO_327 (O_327,N_24908,N_24951);
nor UO_328 (O_328,N_24888,N_24827);
xnor UO_329 (O_329,N_24920,N_24889);
or UO_330 (O_330,N_24971,N_24865);
and UO_331 (O_331,N_24827,N_24871);
and UO_332 (O_332,N_24934,N_24965);
or UO_333 (O_333,N_24810,N_24823);
or UO_334 (O_334,N_24900,N_24999);
nand UO_335 (O_335,N_24820,N_24985);
nand UO_336 (O_336,N_24966,N_24914);
nand UO_337 (O_337,N_24858,N_24999);
or UO_338 (O_338,N_24861,N_24878);
nand UO_339 (O_339,N_24970,N_24931);
xnor UO_340 (O_340,N_24989,N_24824);
or UO_341 (O_341,N_24976,N_24865);
or UO_342 (O_342,N_24988,N_24811);
nor UO_343 (O_343,N_24984,N_24932);
and UO_344 (O_344,N_24807,N_24916);
nand UO_345 (O_345,N_24972,N_24859);
or UO_346 (O_346,N_24830,N_24901);
xor UO_347 (O_347,N_24809,N_24906);
or UO_348 (O_348,N_24814,N_24921);
or UO_349 (O_349,N_24999,N_24856);
xor UO_350 (O_350,N_24884,N_24865);
nor UO_351 (O_351,N_24945,N_24983);
nor UO_352 (O_352,N_24842,N_24970);
or UO_353 (O_353,N_24879,N_24954);
nand UO_354 (O_354,N_24803,N_24954);
and UO_355 (O_355,N_24970,N_24898);
nand UO_356 (O_356,N_24864,N_24867);
nor UO_357 (O_357,N_24825,N_24879);
nand UO_358 (O_358,N_24861,N_24846);
and UO_359 (O_359,N_24970,N_24979);
xor UO_360 (O_360,N_24931,N_24932);
xnor UO_361 (O_361,N_24813,N_24907);
or UO_362 (O_362,N_24818,N_24867);
and UO_363 (O_363,N_24861,N_24948);
and UO_364 (O_364,N_24937,N_24818);
nor UO_365 (O_365,N_24847,N_24886);
xor UO_366 (O_366,N_24956,N_24937);
xor UO_367 (O_367,N_24972,N_24860);
nand UO_368 (O_368,N_24917,N_24937);
nand UO_369 (O_369,N_24962,N_24809);
and UO_370 (O_370,N_24923,N_24941);
xor UO_371 (O_371,N_24891,N_24967);
nor UO_372 (O_372,N_24954,N_24875);
nor UO_373 (O_373,N_24873,N_24932);
and UO_374 (O_374,N_24885,N_24980);
and UO_375 (O_375,N_24977,N_24840);
xnor UO_376 (O_376,N_24873,N_24819);
nor UO_377 (O_377,N_24994,N_24915);
or UO_378 (O_378,N_24855,N_24942);
nor UO_379 (O_379,N_24997,N_24892);
nor UO_380 (O_380,N_24872,N_24809);
or UO_381 (O_381,N_24972,N_24823);
nor UO_382 (O_382,N_24845,N_24897);
nand UO_383 (O_383,N_24930,N_24866);
nand UO_384 (O_384,N_24927,N_24809);
nor UO_385 (O_385,N_24924,N_24948);
nand UO_386 (O_386,N_24900,N_24997);
xor UO_387 (O_387,N_24915,N_24956);
or UO_388 (O_388,N_24908,N_24898);
and UO_389 (O_389,N_24905,N_24866);
nor UO_390 (O_390,N_24872,N_24852);
nand UO_391 (O_391,N_24820,N_24816);
or UO_392 (O_392,N_24885,N_24835);
nand UO_393 (O_393,N_24894,N_24926);
nor UO_394 (O_394,N_24931,N_24927);
nand UO_395 (O_395,N_24805,N_24918);
xnor UO_396 (O_396,N_24854,N_24838);
nand UO_397 (O_397,N_24945,N_24978);
and UO_398 (O_398,N_24930,N_24813);
and UO_399 (O_399,N_24963,N_24972);
xnor UO_400 (O_400,N_24922,N_24934);
nand UO_401 (O_401,N_24969,N_24878);
or UO_402 (O_402,N_24931,N_24948);
xor UO_403 (O_403,N_24847,N_24867);
nand UO_404 (O_404,N_24907,N_24801);
nand UO_405 (O_405,N_24891,N_24911);
and UO_406 (O_406,N_24918,N_24848);
or UO_407 (O_407,N_24916,N_24801);
and UO_408 (O_408,N_24817,N_24887);
xnor UO_409 (O_409,N_24920,N_24998);
xor UO_410 (O_410,N_24968,N_24935);
nor UO_411 (O_411,N_24861,N_24941);
nor UO_412 (O_412,N_24988,N_24958);
nand UO_413 (O_413,N_24937,N_24987);
xnor UO_414 (O_414,N_24826,N_24875);
nor UO_415 (O_415,N_24816,N_24990);
xnor UO_416 (O_416,N_24932,N_24909);
nor UO_417 (O_417,N_24888,N_24966);
xnor UO_418 (O_418,N_24805,N_24980);
or UO_419 (O_419,N_24999,N_24935);
xnor UO_420 (O_420,N_24888,N_24879);
and UO_421 (O_421,N_24912,N_24865);
xnor UO_422 (O_422,N_24844,N_24912);
and UO_423 (O_423,N_24878,N_24874);
and UO_424 (O_424,N_24929,N_24821);
xor UO_425 (O_425,N_24910,N_24829);
and UO_426 (O_426,N_24864,N_24982);
or UO_427 (O_427,N_24871,N_24884);
or UO_428 (O_428,N_24938,N_24922);
nor UO_429 (O_429,N_24821,N_24958);
or UO_430 (O_430,N_24995,N_24914);
xnor UO_431 (O_431,N_24939,N_24981);
and UO_432 (O_432,N_24877,N_24983);
nand UO_433 (O_433,N_24968,N_24977);
nand UO_434 (O_434,N_24832,N_24803);
xor UO_435 (O_435,N_24984,N_24834);
and UO_436 (O_436,N_24890,N_24909);
or UO_437 (O_437,N_24800,N_24933);
nand UO_438 (O_438,N_24954,N_24948);
and UO_439 (O_439,N_24972,N_24845);
xnor UO_440 (O_440,N_24843,N_24967);
or UO_441 (O_441,N_24848,N_24819);
or UO_442 (O_442,N_24936,N_24915);
nand UO_443 (O_443,N_24805,N_24861);
and UO_444 (O_444,N_24899,N_24842);
xor UO_445 (O_445,N_24895,N_24856);
nand UO_446 (O_446,N_24889,N_24999);
or UO_447 (O_447,N_24831,N_24896);
nand UO_448 (O_448,N_24846,N_24911);
nor UO_449 (O_449,N_24892,N_24860);
nand UO_450 (O_450,N_24971,N_24903);
nand UO_451 (O_451,N_24972,N_24933);
xor UO_452 (O_452,N_24925,N_24996);
nor UO_453 (O_453,N_24872,N_24842);
nand UO_454 (O_454,N_24965,N_24979);
nand UO_455 (O_455,N_24800,N_24868);
nand UO_456 (O_456,N_24878,N_24956);
or UO_457 (O_457,N_24966,N_24913);
xnor UO_458 (O_458,N_24908,N_24944);
xnor UO_459 (O_459,N_24896,N_24846);
nor UO_460 (O_460,N_24980,N_24881);
nand UO_461 (O_461,N_24802,N_24929);
or UO_462 (O_462,N_24842,N_24845);
nor UO_463 (O_463,N_24888,N_24809);
xnor UO_464 (O_464,N_24912,N_24972);
and UO_465 (O_465,N_24881,N_24803);
or UO_466 (O_466,N_24821,N_24918);
xnor UO_467 (O_467,N_24852,N_24880);
xnor UO_468 (O_468,N_24967,N_24846);
and UO_469 (O_469,N_24967,N_24973);
nor UO_470 (O_470,N_24818,N_24840);
nand UO_471 (O_471,N_24994,N_24856);
and UO_472 (O_472,N_24875,N_24933);
or UO_473 (O_473,N_24935,N_24954);
and UO_474 (O_474,N_24803,N_24963);
or UO_475 (O_475,N_24896,N_24830);
or UO_476 (O_476,N_24966,N_24917);
nand UO_477 (O_477,N_24955,N_24835);
or UO_478 (O_478,N_24870,N_24815);
nor UO_479 (O_479,N_24876,N_24829);
xor UO_480 (O_480,N_24977,N_24812);
nand UO_481 (O_481,N_24819,N_24879);
xnor UO_482 (O_482,N_24815,N_24939);
nand UO_483 (O_483,N_24911,N_24881);
and UO_484 (O_484,N_24815,N_24918);
and UO_485 (O_485,N_24883,N_24990);
and UO_486 (O_486,N_24807,N_24878);
nand UO_487 (O_487,N_24993,N_24982);
or UO_488 (O_488,N_24904,N_24919);
and UO_489 (O_489,N_24982,N_24802);
and UO_490 (O_490,N_24913,N_24974);
xnor UO_491 (O_491,N_24830,N_24845);
or UO_492 (O_492,N_24953,N_24931);
nor UO_493 (O_493,N_24810,N_24933);
or UO_494 (O_494,N_24983,N_24865);
and UO_495 (O_495,N_24904,N_24808);
or UO_496 (O_496,N_24998,N_24999);
and UO_497 (O_497,N_24839,N_24818);
and UO_498 (O_498,N_24842,N_24938);
or UO_499 (O_499,N_24928,N_24997);
and UO_500 (O_500,N_24862,N_24819);
xnor UO_501 (O_501,N_24815,N_24830);
or UO_502 (O_502,N_24885,N_24987);
xor UO_503 (O_503,N_24873,N_24935);
nand UO_504 (O_504,N_24821,N_24896);
xnor UO_505 (O_505,N_24966,N_24877);
nand UO_506 (O_506,N_24939,N_24865);
or UO_507 (O_507,N_24936,N_24947);
xor UO_508 (O_508,N_24934,N_24874);
or UO_509 (O_509,N_24847,N_24934);
and UO_510 (O_510,N_24943,N_24872);
nor UO_511 (O_511,N_24888,N_24850);
or UO_512 (O_512,N_24814,N_24953);
nor UO_513 (O_513,N_24875,N_24890);
or UO_514 (O_514,N_24820,N_24917);
nor UO_515 (O_515,N_24941,N_24905);
nand UO_516 (O_516,N_24810,N_24927);
nand UO_517 (O_517,N_24801,N_24878);
or UO_518 (O_518,N_24935,N_24843);
and UO_519 (O_519,N_24951,N_24866);
or UO_520 (O_520,N_24977,N_24853);
and UO_521 (O_521,N_24931,N_24842);
nand UO_522 (O_522,N_24951,N_24855);
nor UO_523 (O_523,N_24822,N_24921);
and UO_524 (O_524,N_24969,N_24996);
and UO_525 (O_525,N_24866,N_24962);
or UO_526 (O_526,N_24975,N_24803);
and UO_527 (O_527,N_24908,N_24824);
nor UO_528 (O_528,N_24989,N_24861);
xor UO_529 (O_529,N_24986,N_24911);
xnor UO_530 (O_530,N_24821,N_24809);
nand UO_531 (O_531,N_24836,N_24948);
or UO_532 (O_532,N_24924,N_24983);
xnor UO_533 (O_533,N_24960,N_24870);
and UO_534 (O_534,N_24873,N_24843);
xnor UO_535 (O_535,N_24995,N_24928);
xor UO_536 (O_536,N_24874,N_24972);
nor UO_537 (O_537,N_24908,N_24953);
or UO_538 (O_538,N_24982,N_24845);
and UO_539 (O_539,N_24817,N_24944);
and UO_540 (O_540,N_24946,N_24903);
and UO_541 (O_541,N_24960,N_24978);
nor UO_542 (O_542,N_24807,N_24928);
nor UO_543 (O_543,N_24821,N_24931);
and UO_544 (O_544,N_24978,N_24956);
or UO_545 (O_545,N_24857,N_24960);
or UO_546 (O_546,N_24883,N_24963);
nor UO_547 (O_547,N_24868,N_24883);
or UO_548 (O_548,N_24829,N_24907);
or UO_549 (O_549,N_24824,N_24998);
xor UO_550 (O_550,N_24991,N_24831);
or UO_551 (O_551,N_24999,N_24876);
nor UO_552 (O_552,N_24913,N_24873);
nor UO_553 (O_553,N_24907,N_24844);
nor UO_554 (O_554,N_24826,N_24805);
and UO_555 (O_555,N_24811,N_24922);
nor UO_556 (O_556,N_24829,N_24901);
or UO_557 (O_557,N_24813,N_24911);
and UO_558 (O_558,N_24968,N_24946);
and UO_559 (O_559,N_24815,N_24945);
or UO_560 (O_560,N_24876,N_24962);
nand UO_561 (O_561,N_24876,N_24984);
or UO_562 (O_562,N_24935,N_24975);
xnor UO_563 (O_563,N_24969,N_24823);
xnor UO_564 (O_564,N_24918,N_24831);
or UO_565 (O_565,N_24928,N_24881);
xor UO_566 (O_566,N_24801,N_24840);
and UO_567 (O_567,N_24855,N_24920);
or UO_568 (O_568,N_24860,N_24910);
nor UO_569 (O_569,N_24994,N_24940);
xnor UO_570 (O_570,N_24835,N_24995);
and UO_571 (O_571,N_24985,N_24850);
nor UO_572 (O_572,N_24814,N_24927);
or UO_573 (O_573,N_24858,N_24901);
nor UO_574 (O_574,N_24960,N_24932);
xnor UO_575 (O_575,N_24920,N_24892);
nand UO_576 (O_576,N_24837,N_24863);
nor UO_577 (O_577,N_24940,N_24835);
or UO_578 (O_578,N_24832,N_24999);
or UO_579 (O_579,N_24820,N_24836);
and UO_580 (O_580,N_24826,N_24934);
nand UO_581 (O_581,N_24822,N_24974);
xor UO_582 (O_582,N_24869,N_24981);
nand UO_583 (O_583,N_24962,N_24977);
xor UO_584 (O_584,N_24886,N_24975);
nand UO_585 (O_585,N_24929,N_24901);
nand UO_586 (O_586,N_24863,N_24939);
or UO_587 (O_587,N_24872,N_24944);
nand UO_588 (O_588,N_24903,N_24846);
nand UO_589 (O_589,N_24930,N_24850);
nand UO_590 (O_590,N_24827,N_24979);
or UO_591 (O_591,N_24886,N_24879);
or UO_592 (O_592,N_24873,N_24884);
xor UO_593 (O_593,N_24941,N_24970);
or UO_594 (O_594,N_24979,N_24893);
xor UO_595 (O_595,N_24958,N_24955);
or UO_596 (O_596,N_24804,N_24801);
nand UO_597 (O_597,N_24998,N_24957);
xor UO_598 (O_598,N_24939,N_24834);
and UO_599 (O_599,N_24915,N_24997);
nand UO_600 (O_600,N_24846,N_24873);
nor UO_601 (O_601,N_24941,N_24800);
nor UO_602 (O_602,N_24980,N_24890);
or UO_603 (O_603,N_24985,N_24831);
xor UO_604 (O_604,N_24911,N_24900);
nand UO_605 (O_605,N_24909,N_24936);
nor UO_606 (O_606,N_24962,N_24908);
or UO_607 (O_607,N_24828,N_24865);
xnor UO_608 (O_608,N_24972,N_24967);
or UO_609 (O_609,N_24893,N_24860);
nor UO_610 (O_610,N_24858,N_24853);
xor UO_611 (O_611,N_24825,N_24881);
xnor UO_612 (O_612,N_24900,N_24866);
and UO_613 (O_613,N_24897,N_24828);
and UO_614 (O_614,N_24973,N_24815);
nor UO_615 (O_615,N_24870,N_24822);
or UO_616 (O_616,N_24906,N_24860);
or UO_617 (O_617,N_24866,N_24950);
or UO_618 (O_618,N_24868,N_24950);
nor UO_619 (O_619,N_24878,N_24928);
xnor UO_620 (O_620,N_24998,N_24831);
or UO_621 (O_621,N_24969,N_24954);
nand UO_622 (O_622,N_24872,N_24904);
and UO_623 (O_623,N_24823,N_24867);
nand UO_624 (O_624,N_24914,N_24980);
or UO_625 (O_625,N_24899,N_24839);
and UO_626 (O_626,N_24822,N_24826);
xnor UO_627 (O_627,N_24978,N_24867);
nand UO_628 (O_628,N_24803,N_24806);
and UO_629 (O_629,N_24834,N_24808);
xor UO_630 (O_630,N_24885,N_24831);
or UO_631 (O_631,N_24955,N_24963);
xnor UO_632 (O_632,N_24802,N_24837);
or UO_633 (O_633,N_24830,N_24859);
nand UO_634 (O_634,N_24999,N_24873);
xnor UO_635 (O_635,N_24874,N_24811);
and UO_636 (O_636,N_24836,N_24845);
or UO_637 (O_637,N_24844,N_24874);
and UO_638 (O_638,N_24937,N_24820);
nand UO_639 (O_639,N_24876,N_24937);
and UO_640 (O_640,N_24826,N_24844);
and UO_641 (O_641,N_24925,N_24831);
xor UO_642 (O_642,N_24852,N_24806);
nor UO_643 (O_643,N_24934,N_24807);
or UO_644 (O_644,N_24860,N_24865);
nor UO_645 (O_645,N_24803,N_24902);
xnor UO_646 (O_646,N_24981,N_24944);
nand UO_647 (O_647,N_24821,N_24978);
nand UO_648 (O_648,N_24824,N_24858);
nand UO_649 (O_649,N_24973,N_24936);
nor UO_650 (O_650,N_24901,N_24889);
xnor UO_651 (O_651,N_24978,N_24818);
and UO_652 (O_652,N_24980,N_24859);
xor UO_653 (O_653,N_24953,N_24980);
nor UO_654 (O_654,N_24856,N_24841);
xnor UO_655 (O_655,N_24924,N_24836);
xor UO_656 (O_656,N_24918,N_24872);
nand UO_657 (O_657,N_24809,N_24955);
or UO_658 (O_658,N_24890,N_24991);
and UO_659 (O_659,N_24915,N_24844);
nor UO_660 (O_660,N_24997,N_24930);
nor UO_661 (O_661,N_24814,N_24954);
and UO_662 (O_662,N_24996,N_24932);
or UO_663 (O_663,N_24812,N_24904);
and UO_664 (O_664,N_24818,N_24865);
or UO_665 (O_665,N_24954,N_24872);
xor UO_666 (O_666,N_24888,N_24886);
or UO_667 (O_667,N_24964,N_24810);
and UO_668 (O_668,N_24813,N_24927);
xor UO_669 (O_669,N_24817,N_24925);
and UO_670 (O_670,N_24887,N_24909);
or UO_671 (O_671,N_24800,N_24983);
and UO_672 (O_672,N_24913,N_24806);
or UO_673 (O_673,N_24919,N_24885);
nor UO_674 (O_674,N_24990,N_24889);
xnor UO_675 (O_675,N_24824,N_24902);
or UO_676 (O_676,N_24888,N_24910);
nor UO_677 (O_677,N_24978,N_24957);
and UO_678 (O_678,N_24848,N_24842);
nand UO_679 (O_679,N_24808,N_24864);
or UO_680 (O_680,N_24975,N_24971);
nand UO_681 (O_681,N_24835,N_24831);
nand UO_682 (O_682,N_24906,N_24821);
and UO_683 (O_683,N_24949,N_24964);
nor UO_684 (O_684,N_24890,N_24934);
and UO_685 (O_685,N_24867,N_24906);
nand UO_686 (O_686,N_24989,N_24841);
nand UO_687 (O_687,N_24951,N_24976);
or UO_688 (O_688,N_24853,N_24879);
and UO_689 (O_689,N_24982,N_24900);
or UO_690 (O_690,N_24974,N_24935);
nand UO_691 (O_691,N_24912,N_24888);
and UO_692 (O_692,N_24970,N_24843);
or UO_693 (O_693,N_24811,N_24999);
xor UO_694 (O_694,N_24943,N_24826);
xor UO_695 (O_695,N_24862,N_24835);
nor UO_696 (O_696,N_24912,N_24862);
nand UO_697 (O_697,N_24960,N_24966);
nor UO_698 (O_698,N_24839,N_24974);
nor UO_699 (O_699,N_24915,N_24924);
xor UO_700 (O_700,N_24902,N_24989);
and UO_701 (O_701,N_24975,N_24802);
nor UO_702 (O_702,N_24834,N_24940);
xor UO_703 (O_703,N_24989,N_24984);
and UO_704 (O_704,N_24871,N_24938);
or UO_705 (O_705,N_24890,N_24904);
nand UO_706 (O_706,N_24987,N_24853);
nor UO_707 (O_707,N_24859,N_24945);
nand UO_708 (O_708,N_24889,N_24899);
nand UO_709 (O_709,N_24984,N_24993);
and UO_710 (O_710,N_24916,N_24828);
and UO_711 (O_711,N_24972,N_24842);
or UO_712 (O_712,N_24896,N_24933);
or UO_713 (O_713,N_24865,N_24984);
or UO_714 (O_714,N_24820,N_24900);
xor UO_715 (O_715,N_24975,N_24879);
nand UO_716 (O_716,N_24982,N_24910);
or UO_717 (O_717,N_24884,N_24945);
and UO_718 (O_718,N_24825,N_24898);
nand UO_719 (O_719,N_24905,N_24933);
nor UO_720 (O_720,N_24812,N_24923);
nand UO_721 (O_721,N_24823,N_24962);
xor UO_722 (O_722,N_24882,N_24901);
nand UO_723 (O_723,N_24962,N_24934);
and UO_724 (O_724,N_24912,N_24914);
or UO_725 (O_725,N_24869,N_24893);
or UO_726 (O_726,N_24816,N_24974);
nor UO_727 (O_727,N_24972,N_24813);
nand UO_728 (O_728,N_24837,N_24896);
and UO_729 (O_729,N_24877,N_24845);
nor UO_730 (O_730,N_24973,N_24926);
nor UO_731 (O_731,N_24862,N_24803);
and UO_732 (O_732,N_24828,N_24885);
nor UO_733 (O_733,N_24939,N_24951);
xnor UO_734 (O_734,N_24998,N_24900);
nand UO_735 (O_735,N_24844,N_24882);
nor UO_736 (O_736,N_24937,N_24844);
or UO_737 (O_737,N_24950,N_24804);
and UO_738 (O_738,N_24865,N_24890);
and UO_739 (O_739,N_24828,N_24844);
or UO_740 (O_740,N_24990,N_24837);
or UO_741 (O_741,N_24879,N_24823);
xor UO_742 (O_742,N_24828,N_24843);
and UO_743 (O_743,N_24837,N_24801);
xnor UO_744 (O_744,N_24994,N_24926);
nand UO_745 (O_745,N_24802,N_24987);
xnor UO_746 (O_746,N_24848,N_24942);
nor UO_747 (O_747,N_24862,N_24911);
nor UO_748 (O_748,N_24900,N_24975);
nand UO_749 (O_749,N_24914,N_24821);
and UO_750 (O_750,N_24984,N_24948);
and UO_751 (O_751,N_24812,N_24979);
and UO_752 (O_752,N_24843,N_24846);
nand UO_753 (O_753,N_24893,N_24925);
nor UO_754 (O_754,N_24961,N_24896);
and UO_755 (O_755,N_24994,N_24872);
nor UO_756 (O_756,N_24824,N_24853);
nor UO_757 (O_757,N_24939,N_24853);
xor UO_758 (O_758,N_24934,N_24811);
and UO_759 (O_759,N_24883,N_24940);
nor UO_760 (O_760,N_24883,N_24855);
nand UO_761 (O_761,N_24907,N_24871);
and UO_762 (O_762,N_24928,N_24945);
nand UO_763 (O_763,N_24935,N_24921);
nand UO_764 (O_764,N_24997,N_24953);
and UO_765 (O_765,N_24879,N_24895);
xor UO_766 (O_766,N_24830,N_24996);
xor UO_767 (O_767,N_24931,N_24906);
xor UO_768 (O_768,N_24854,N_24853);
nand UO_769 (O_769,N_24904,N_24876);
nor UO_770 (O_770,N_24871,N_24917);
or UO_771 (O_771,N_24891,N_24875);
and UO_772 (O_772,N_24834,N_24997);
nor UO_773 (O_773,N_24850,N_24867);
or UO_774 (O_774,N_24878,N_24999);
and UO_775 (O_775,N_24900,N_24808);
nor UO_776 (O_776,N_24834,N_24970);
nand UO_777 (O_777,N_24849,N_24946);
and UO_778 (O_778,N_24902,N_24813);
and UO_779 (O_779,N_24820,N_24901);
and UO_780 (O_780,N_24840,N_24879);
or UO_781 (O_781,N_24972,N_24979);
or UO_782 (O_782,N_24882,N_24960);
nor UO_783 (O_783,N_24843,N_24936);
or UO_784 (O_784,N_24834,N_24853);
xor UO_785 (O_785,N_24931,N_24920);
nor UO_786 (O_786,N_24941,N_24997);
or UO_787 (O_787,N_24851,N_24994);
nor UO_788 (O_788,N_24967,N_24911);
xor UO_789 (O_789,N_24923,N_24886);
nor UO_790 (O_790,N_24804,N_24892);
nor UO_791 (O_791,N_24946,N_24951);
nand UO_792 (O_792,N_24803,N_24920);
xnor UO_793 (O_793,N_24951,N_24888);
and UO_794 (O_794,N_24914,N_24957);
or UO_795 (O_795,N_24865,N_24914);
nor UO_796 (O_796,N_24957,N_24949);
nor UO_797 (O_797,N_24871,N_24837);
or UO_798 (O_798,N_24840,N_24934);
nor UO_799 (O_799,N_24961,N_24850);
xor UO_800 (O_800,N_24956,N_24805);
or UO_801 (O_801,N_24980,N_24812);
or UO_802 (O_802,N_24928,N_24900);
nor UO_803 (O_803,N_24839,N_24964);
and UO_804 (O_804,N_24863,N_24951);
nor UO_805 (O_805,N_24808,N_24947);
nand UO_806 (O_806,N_24957,N_24834);
and UO_807 (O_807,N_24960,N_24850);
xor UO_808 (O_808,N_24981,N_24986);
nand UO_809 (O_809,N_24892,N_24998);
nor UO_810 (O_810,N_24877,N_24919);
and UO_811 (O_811,N_24978,N_24940);
and UO_812 (O_812,N_24998,N_24804);
and UO_813 (O_813,N_24810,N_24982);
and UO_814 (O_814,N_24813,N_24837);
xor UO_815 (O_815,N_24998,N_24928);
nor UO_816 (O_816,N_24891,N_24925);
nor UO_817 (O_817,N_24881,N_24920);
nor UO_818 (O_818,N_24913,N_24932);
nand UO_819 (O_819,N_24823,N_24911);
nor UO_820 (O_820,N_24970,N_24959);
and UO_821 (O_821,N_24946,N_24873);
or UO_822 (O_822,N_24805,N_24991);
and UO_823 (O_823,N_24961,N_24817);
and UO_824 (O_824,N_24845,N_24923);
xor UO_825 (O_825,N_24967,N_24933);
xor UO_826 (O_826,N_24882,N_24862);
nand UO_827 (O_827,N_24980,N_24928);
nand UO_828 (O_828,N_24852,N_24814);
nor UO_829 (O_829,N_24941,N_24904);
and UO_830 (O_830,N_24984,N_24874);
nand UO_831 (O_831,N_24853,N_24847);
or UO_832 (O_832,N_24835,N_24802);
and UO_833 (O_833,N_24836,N_24874);
and UO_834 (O_834,N_24960,N_24822);
xor UO_835 (O_835,N_24924,N_24975);
nand UO_836 (O_836,N_24880,N_24910);
and UO_837 (O_837,N_24835,N_24980);
nand UO_838 (O_838,N_24855,N_24881);
xor UO_839 (O_839,N_24907,N_24916);
and UO_840 (O_840,N_24803,N_24841);
or UO_841 (O_841,N_24890,N_24916);
and UO_842 (O_842,N_24806,N_24925);
or UO_843 (O_843,N_24978,N_24938);
xnor UO_844 (O_844,N_24803,N_24819);
xor UO_845 (O_845,N_24824,N_24969);
nor UO_846 (O_846,N_24844,N_24987);
nor UO_847 (O_847,N_24988,N_24918);
or UO_848 (O_848,N_24961,N_24950);
nand UO_849 (O_849,N_24858,N_24817);
xnor UO_850 (O_850,N_24892,N_24912);
or UO_851 (O_851,N_24918,N_24890);
nor UO_852 (O_852,N_24908,N_24868);
nor UO_853 (O_853,N_24924,N_24815);
nor UO_854 (O_854,N_24951,N_24853);
nand UO_855 (O_855,N_24901,N_24818);
nor UO_856 (O_856,N_24954,N_24836);
nor UO_857 (O_857,N_24937,N_24872);
xnor UO_858 (O_858,N_24849,N_24934);
nand UO_859 (O_859,N_24948,N_24980);
xor UO_860 (O_860,N_24881,N_24860);
nand UO_861 (O_861,N_24988,N_24925);
nand UO_862 (O_862,N_24888,N_24898);
nor UO_863 (O_863,N_24817,N_24946);
xor UO_864 (O_864,N_24839,N_24968);
nand UO_865 (O_865,N_24886,N_24902);
nor UO_866 (O_866,N_24907,N_24814);
and UO_867 (O_867,N_24949,N_24941);
nand UO_868 (O_868,N_24936,N_24824);
xnor UO_869 (O_869,N_24930,N_24833);
or UO_870 (O_870,N_24948,N_24842);
nand UO_871 (O_871,N_24976,N_24810);
xor UO_872 (O_872,N_24903,N_24934);
xnor UO_873 (O_873,N_24925,N_24876);
and UO_874 (O_874,N_24978,N_24930);
and UO_875 (O_875,N_24869,N_24885);
and UO_876 (O_876,N_24844,N_24823);
nand UO_877 (O_877,N_24878,N_24830);
nand UO_878 (O_878,N_24978,N_24926);
and UO_879 (O_879,N_24961,N_24988);
xnor UO_880 (O_880,N_24982,N_24867);
nand UO_881 (O_881,N_24901,N_24851);
nor UO_882 (O_882,N_24829,N_24939);
nor UO_883 (O_883,N_24942,N_24959);
nor UO_884 (O_884,N_24985,N_24941);
or UO_885 (O_885,N_24971,N_24997);
or UO_886 (O_886,N_24894,N_24885);
or UO_887 (O_887,N_24826,N_24900);
xnor UO_888 (O_888,N_24861,N_24893);
nor UO_889 (O_889,N_24857,N_24818);
and UO_890 (O_890,N_24942,N_24958);
or UO_891 (O_891,N_24812,N_24955);
nand UO_892 (O_892,N_24830,N_24886);
and UO_893 (O_893,N_24996,N_24855);
nor UO_894 (O_894,N_24969,N_24935);
nand UO_895 (O_895,N_24959,N_24882);
nor UO_896 (O_896,N_24956,N_24813);
nand UO_897 (O_897,N_24983,N_24802);
xnor UO_898 (O_898,N_24995,N_24919);
or UO_899 (O_899,N_24938,N_24975);
and UO_900 (O_900,N_24832,N_24920);
xor UO_901 (O_901,N_24832,N_24837);
nor UO_902 (O_902,N_24849,N_24815);
xor UO_903 (O_903,N_24807,N_24989);
nor UO_904 (O_904,N_24954,N_24898);
nor UO_905 (O_905,N_24863,N_24959);
nor UO_906 (O_906,N_24833,N_24822);
xnor UO_907 (O_907,N_24841,N_24850);
or UO_908 (O_908,N_24965,N_24902);
and UO_909 (O_909,N_24810,N_24986);
nor UO_910 (O_910,N_24946,N_24976);
and UO_911 (O_911,N_24938,N_24832);
or UO_912 (O_912,N_24846,N_24974);
nand UO_913 (O_913,N_24831,N_24859);
or UO_914 (O_914,N_24840,N_24834);
and UO_915 (O_915,N_24885,N_24830);
nand UO_916 (O_916,N_24856,N_24896);
nand UO_917 (O_917,N_24833,N_24978);
or UO_918 (O_918,N_24951,N_24948);
and UO_919 (O_919,N_24834,N_24832);
nor UO_920 (O_920,N_24976,N_24959);
or UO_921 (O_921,N_24952,N_24851);
xnor UO_922 (O_922,N_24973,N_24814);
and UO_923 (O_923,N_24826,N_24962);
and UO_924 (O_924,N_24877,N_24909);
nand UO_925 (O_925,N_24885,N_24979);
nor UO_926 (O_926,N_24973,N_24862);
nand UO_927 (O_927,N_24850,N_24903);
and UO_928 (O_928,N_24868,N_24842);
or UO_929 (O_929,N_24805,N_24984);
nor UO_930 (O_930,N_24969,N_24944);
xor UO_931 (O_931,N_24942,N_24953);
or UO_932 (O_932,N_24925,N_24956);
and UO_933 (O_933,N_24804,N_24806);
xnor UO_934 (O_934,N_24811,N_24807);
nand UO_935 (O_935,N_24908,N_24883);
nor UO_936 (O_936,N_24885,N_24876);
xnor UO_937 (O_937,N_24857,N_24862);
and UO_938 (O_938,N_24993,N_24860);
nor UO_939 (O_939,N_24818,N_24970);
nor UO_940 (O_940,N_24808,N_24895);
xnor UO_941 (O_941,N_24976,N_24852);
or UO_942 (O_942,N_24990,N_24818);
nand UO_943 (O_943,N_24900,N_24889);
xor UO_944 (O_944,N_24979,N_24930);
xor UO_945 (O_945,N_24953,N_24972);
nand UO_946 (O_946,N_24874,N_24917);
nor UO_947 (O_947,N_24858,N_24896);
xor UO_948 (O_948,N_24885,N_24982);
nand UO_949 (O_949,N_24828,N_24973);
xor UO_950 (O_950,N_24903,N_24969);
and UO_951 (O_951,N_24842,N_24813);
nand UO_952 (O_952,N_24971,N_24815);
nand UO_953 (O_953,N_24851,N_24953);
or UO_954 (O_954,N_24870,N_24844);
and UO_955 (O_955,N_24958,N_24994);
nand UO_956 (O_956,N_24904,N_24994);
xnor UO_957 (O_957,N_24813,N_24929);
xor UO_958 (O_958,N_24951,N_24875);
or UO_959 (O_959,N_24965,N_24973);
or UO_960 (O_960,N_24901,N_24977);
xor UO_961 (O_961,N_24884,N_24836);
nor UO_962 (O_962,N_24949,N_24950);
nand UO_963 (O_963,N_24961,N_24844);
nor UO_964 (O_964,N_24953,N_24867);
or UO_965 (O_965,N_24847,N_24802);
nand UO_966 (O_966,N_24967,N_24861);
nand UO_967 (O_967,N_24843,N_24852);
xnor UO_968 (O_968,N_24898,N_24807);
xor UO_969 (O_969,N_24923,N_24884);
nand UO_970 (O_970,N_24805,N_24855);
nand UO_971 (O_971,N_24942,N_24870);
nor UO_972 (O_972,N_24911,N_24913);
or UO_973 (O_973,N_24860,N_24840);
nand UO_974 (O_974,N_24942,N_24981);
nor UO_975 (O_975,N_24804,N_24929);
nor UO_976 (O_976,N_24821,N_24970);
nor UO_977 (O_977,N_24807,N_24965);
nor UO_978 (O_978,N_24908,N_24937);
nand UO_979 (O_979,N_24810,N_24889);
xnor UO_980 (O_980,N_24867,N_24809);
xor UO_981 (O_981,N_24997,N_24807);
nand UO_982 (O_982,N_24945,N_24935);
or UO_983 (O_983,N_24850,N_24983);
and UO_984 (O_984,N_24817,N_24964);
nand UO_985 (O_985,N_24824,N_24866);
or UO_986 (O_986,N_24894,N_24843);
and UO_987 (O_987,N_24844,N_24963);
xnor UO_988 (O_988,N_24989,N_24957);
xnor UO_989 (O_989,N_24950,N_24995);
nand UO_990 (O_990,N_24971,N_24960);
and UO_991 (O_991,N_24841,N_24919);
or UO_992 (O_992,N_24950,N_24875);
nor UO_993 (O_993,N_24811,N_24808);
xnor UO_994 (O_994,N_24972,N_24891);
nor UO_995 (O_995,N_24804,N_24863);
nor UO_996 (O_996,N_24978,N_24985);
xor UO_997 (O_997,N_24844,N_24958);
or UO_998 (O_998,N_24973,N_24924);
xnor UO_999 (O_999,N_24833,N_24937);
or UO_1000 (O_1000,N_24867,N_24828);
nand UO_1001 (O_1001,N_24823,N_24895);
nor UO_1002 (O_1002,N_24881,N_24954);
and UO_1003 (O_1003,N_24880,N_24993);
nor UO_1004 (O_1004,N_24834,N_24992);
nor UO_1005 (O_1005,N_24871,N_24971);
and UO_1006 (O_1006,N_24901,N_24853);
nor UO_1007 (O_1007,N_24800,N_24822);
nand UO_1008 (O_1008,N_24832,N_24828);
nor UO_1009 (O_1009,N_24854,N_24824);
nand UO_1010 (O_1010,N_24925,N_24992);
nor UO_1011 (O_1011,N_24980,N_24814);
nor UO_1012 (O_1012,N_24822,N_24823);
nand UO_1013 (O_1013,N_24817,N_24890);
and UO_1014 (O_1014,N_24836,N_24964);
and UO_1015 (O_1015,N_24906,N_24947);
or UO_1016 (O_1016,N_24969,N_24975);
or UO_1017 (O_1017,N_24961,N_24853);
xnor UO_1018 (O_1018,N_24880,N_24912);
or UO_1019 (O_1019,N_24815,N_24829);
and UO_1020 (O_1020,N_24991,N_24904);
nand UO_1021 (O_1021,N_24920,N_24853);
nor UO_1022 (O_1022,N_24973,N_24982);
nand UO_1023 (O_1023,N_24940,N_24967);
xnor UO_1024 (O_1024,N_24932,N_24933);
or UO_1025 (O_1025,N_24825,N_24833);
or UO_1026 (O_1026,N_24811,N_24859);
xor UO_1027 (O_1027,N_24996,N_24949);
or UO_1028 (O_1028,N_24955,N_24852);
and UO_1029 (O_1029,N_24810,N_24854);
nor UO_1030 (O_1030,N_24886,N_24929);
xnor UO_1031 (O_1031,N_24846,N_24927);
and UO_1032 (O_1032,N_24856,N_24924);
and UO_1033 (O_1033,N_24888,N_24978);
nand UO_1034 (O_1034,N_24847,N_24959);
and UO_1035 (O_1035,N_24815,N_24827);
or UO_1036 (O_1036,N_24948,N_24927);
and UO_1037 (O_1037,N_24977,N_24846);
xor UO_1038 (O_1038,N_24861,N_24976);
and UO_1039 (O_1039,N_24858,N_24955);
nor UO_1040 (O_1040,N_24810,N_24827);
nand UO_1041 (O_1041,N_24888,N_24847);
xnor UO_1042 (O_1042,N_24840,N_24911);
xor UO_1043 (O_1043,N_24940,N_24857);
nand UO_1044 (O_1044,N_24836,N_24949);
xor UO_1045 (O_1045,N_24879,N_24863);
nand UO_1046 (O_1046,N_24873,N_24800);
nor UO_1047 (O_1047,N_24985,N_24877);
xor UO_1048 (O_1048,N_24842,N_24811);
nand UO_1049 (O_1049,N_24914,N_24825);
xor UO_1050 (O_1050,N_24922,N_24900);
and UO_1051 (O_1051,N_24844,N_24803);
and UO_1052 (O_1052,N_24829,N_24999);
nand UO_1053 (O_1053,N_24832,N_24885);
nor UO_1054 (O_1054,N_24898,N_24815);
nor UO_1055 (O_1055,N_24932,N_24954);
xnor UO_1056 (O_1056,N_24866,N_24881);
or UO_1057 (O_1057,N_24911,N_24833);
or UO_1058 (O_1058,N_24901,N_24934);
or UO_1059 (O_1059,N_24906,N_24987);
or UO_1060 (O_1060,N_24841,N_24938);
xor UO_1061 (O_1061,N_24938,N_24819);
or UO_1062 (O_1062,N_24852,N_24999);
and UO_1063 (O_1063,N_24954,N_24910);
nor UO_1064 (O_1064,N_24801,N_24896);
and UO_1065 (O_1065,N_24905,N_24960);
nand UO_1066 (O_1066,N_24998,N_24985);
nand UO_1067 (O_1067,N_24920,N_24800);
nand UO_1068 (O_1068,N_24898,N_24839);
or UO_1069 (O_1069,N_24844,N_24921);
or UO_1070 (O_1070,N_24912,N_24964);
nand UO_1071 (O_1071,N_24947,N_24908);
xor UO_1072 (O_1072,N_24990,N_24827);
nor UO_1073 (O_1073,N_24868,N_24861);
nand UO_1074 (O_1074,N_24904,N_24845);
xnor UO_1075 (O_1075,N_24957,N_24813);
xnor UO_1076 (O_1076,N_24860,N_24925);
and UO_1077 (O_1077,N_24860,N_24859);
or UO_1078 (O_1078,N_24953,N_24845);
nand UO_1079 (O_1079,N_24870,N_24989);
nor UO_1080 (O_1080,N_24988,N_24808);
xnor UO_1081 (O_1081,N_24923,N_24983);
and UO_1082 (O_1082,N_24846,N_24965);
nand UO_1083 (O_1083,N_24965,N_24891);
and UO_1084 (O_1084,N_24977,N_24942);
nor UO_1085 (O_1085,N_24941,N_24807);
nand UO_1086 (O_1086,N_24953,N_24921);
nand UO_1087 (O_1087,N_24830,N_24898);
nand UO_1088 (O_1088,N_24925,N_24958);
nand UO_1089 (O_1089,N_24898,N_24865);
nand UO_1090 (O_1090,N_24874,N_24991);
nor UO_1091 (O_1091,N_24996,N_24818);
and UO_1092 (O_1092,N_24840,N_24903);
or UO_1093 (O_1093,N_24838,N_24876);
and UO_1094 (O_1094,N_24847,N_24958);
or UO_1095 (O_1095,N_24921,N_24949);
nand UO_1096 (O_1096,N_24918,N_24954);
or UO_1097 (O_1097,N_24860,N_24975);
nor UO_1098 (O_1098,N_24868,N_24867);
or UO_1099 (O_1099,N_24978,N_24877);
xor UO_1100 (O_1100,N_24999,N_24986);
nor UO_1101 (O_1101,N_24815,N_24822);
and UO_1102 (O_1102,N_24862,N_24957);
nor UO_1103 (O_1103,N_24831,N_24879);
or UO_1104 (O_1104,N_24834,N_24974);
and UO_1105 (O_1105,N_24920,N_24897);
nor UO_1106 (O_1106,N_24845,N_24876);
and UO_1107 (O_1107,N_24889,N_24993);
xor UO_1108 (O_1108,N_24839,N_24863);
nor UO_1109 (O_1109,N_24970,N_24867);
or UO_1110 (O_1110,N_24903,N_24853);
and UO_1111 (O_1111,N_24992,N_24887);
and UO_1112 (O_1112,N_24895,N_24861);
or UO_1113 (O_1113,N_24940,N_24820);
and UO_1114 (O_1114,N_24990,N_24873);
nand UO_1115 (O_1115,N_24828,N_24801);
nor UO_1116 (O_1116,N_24952,N_24875);
or UO_1117 (O_1117,N_24961,N_24970);
nor UO_1118 (O_1118,N_24977,N_24896);
nand UO_1119 (O_1119,N_24997,N_24833);
xnor UO_1120 (O_1120,N_24930,N_24802);
nor UO_1121 (O_1121,N_24878,N_24817);
or UO_1122 (O_1122,N_24860,N_24836);
or UO_1123 (O_1123,N_24883,N_24977);
nor UO_1124 (O_1124,N_24826,N_24804);
nand UO_1125 (O_1125,N_24929,N_24863);
or UO_1126 (O_1126,N_24958,N_24826);
and UO_1127 (O_1127,N_24811,N_24850);
and UO_1128 (O_1128,N_24921,N_24924);
or UO_1129 (O_1129,N_24804,N_24995);
and UO_1130 (O_1130,N_24946,N_24935);
and UO_1131 (O_1131,N_24887,N_24801);
and UO_1132 (O_1132,N_24898,N_24886);
or UO_1133 (O_1133,N_24943,N_24890);
or UO_1134 (O_1134,N_24944,N_24809);
or UO_1135 (O_1135,N_24873,N_24817);
xor UO_1136 (O_1136,N_24896,N_24915);
nand UO_1137 (O_1137,N_24900,N_24902);
xor UO_1138 (O_1138,N_24940,N_24984);
and UO_1139 (O_1139,N_24896,N_24995);
nand UO_1140 (O_1140,N_24815,N_24919);
or UO_1141 (O_1141,N_24847,N_24932);
and UO_1142 (O_1142,N_24877,N_24958);
or UO_1143 (O_1143,N_24924,N_24940);
nand UO_1144 (O_1144,N_24800,N_24825);
or UO_1145 (O_1145,N_24818,N_24983);
nand UO_1146 (O_1146,N_24917,N_24876);
nand UO_1147 (O_1147,N_24959,N_24930);
and UO_1148 (O_1148,N_24968,N_24982);
xnor UO_1149 (O_1149,N_24935,N_24965);
nand UO_1150 (O_1150,N_24852,N_24948);
or UO_1151 (O_1151,N_24893,N_24993);
nand UO_1152 (O_1152,N_24907,N_24974);
xnor UO_1153 (O_1153,N_24836,N_24985);
and UO_1154 (O_1154,N_24832,N_24998);
xor UO_1155 (O_1155,N_24816,N_24964);
nand UO_1156 (O_1156,N_24910,N_24871);
nor UO_1157 (O_1157,N_24912,N_24900);
or UO_1158 (O_1158,N_24861,N_24995);
nand UO_1159 (O_1159,N_24820,N_24891);
nand UO_1160 (O_1160,N_24894,N_24969);
and UO_1161 (O_1161,N_24929,N_24898);
and UO_1162 (O_1162,N_24878,N_24862);
nor UO_1163 (O_1163,N_24835,N_24926);
and UO_1164 (O_1164,N_24964,N_24960);
or UO_1165 (O_1165,N_24945,N_24977);
and UO_1166 (O_1166,N_24998,N_24877);
or UO_1167 (O_1167,N_24956,N_24973);
or UO_1168 (O_1168,N_24828,N_24929);
nor UO_1169 (O_1169,N_24998,N_24967);
or UO_1170 (O_1170,N_24866,N_24872);
xor UO_1171 (O_1171,N_24900,N_24800);
or UO_1172 (O_1172,N_24958,N_24841);
nand UO_1173 (O_1173,N_24867,N_24962);
xnor UO_1174 (O_1174,N_24902,N_24817);
or UO_1175 (O_1175,N_24824,N_24886);
nor UO_1176 (O_1176,N_24878,N_24932);
nand UO_1177 (O_1177,N_24861,N_24907);
xor UO_1178 (O_1178,N_24847,N_24876);
nor UO_1179 (O_1179,N_24990,N_24891);
nand UO_1180 (O_1180,N_24854,N_24852);
nor UO_1181 (O_1181,N_24940,N_24852);
xor UO_1182 (O_1182,N_24843,N_24978);
xor UO_1183 (O_1183,N_24877,N_24825);
xnor UO_1184 (O_1184,N_24885,N_24805);
and UO_1185 (O_1185,N_24825,N_24897);
or UO_1186 (O_1186,N_24853,N_24866);
xnor UO_1187 (O_1187,N_24827,N_24850);
nand UO_1188 (O_1188,N_24859,N_24884);
xor UO_1189 (O_1189,N_24935,N_24893);
and UO_1190 (O_1190,N_24877,N_24844);
xnor UO_1191 (O_1191,N_24851,N_24997);
or UO_1192 (O_1192,N_24980,N_24879);
xnor UO_1193 (O_1193,N_24866,N_24847);
or UO_1194 (O_1194,N_24801,N_24815);
and UO_1195 (O_1195,N_24943,N_24878);
xor UO_1196 (O_1196,N_24828,N_24861);
and UO_1197 (O_1197,N_24831,N_24970);
xnor UO_1198 (O_1198,N_24973,N_24802);
and UO_1199 (O_1199,N_24905,N_24914);
or UO_1200 (O_1200,N_24918,N_24818);
and UO_1201 (O_1201,N_24919,N_24883);
and UO_1202 (O_1202,N_24931,N_24837);
nor UO_1203 (O_1203,N_24863,N_24873);
and UO_1204 (O_1204,N_24922,N_24852);
and UO_1205 (O_1205,N_24906,N_24976);
and UO_1206 (O_1206,N_24986,N_24947);
xnor UO_1207 (O_1207,N_24884,N_24941);
and UO_1208 (O_1208,N_24908,N_24835);
nor UO_1209 (O_1209,N_24822,N_24871);
xor UO_1210 (O_1210,N_24821,N_24924);
nand UO_1211 (O_1211,N_24801,N_24855);
and UO_1212 (O_1212,N_24805,N_24838);
xnor UO_1213 (O_1213,N_24919,N_24804);
or UO_1214 (O_1214,N_24943,N_24865);
or UO_1215 (O_1215,N_24832,N_24824);
nand UO_1216 (O_1216,N_24997,N_24933);
nor UO_1217 (O_1217,N_24849,N_24900);
and UO_1218 (O_1218,N_24940,N_24855);
nor UO_1219 (O_1219,N_24877,N_24874);
xor UO_1220 (O_1220,N_24805,N_24807);
xor UO_1221 (O_1221,N_24865,N_24990);
nand UO_1222 (O_1222,N_24948,N_24907);
xor UO_1223 (O_1223,N_24913,N_24840);
or UO_1224 (O_1224,N_24813,N_24819);
or UO_1225 (O_1225,N_24848,N_24821);
xor UO_1226 (O_1226,N_24886,N_24992);
nand UO_1227 (O_1227,N_24924,N_24893);
or UO_1228 (O_1228,N_24906,N_24874);
and UO_1229 (O_1229,N_24874,N_24875);
nor UO_1230 (O_1230,N_24886,N_24908);
or UO_1231 (O_1231,N_24999,N_24954);
nor UO_1232 (O_1232,N_24885,N_24806);
or UO_1233 (O_1233,N_24821,N_24836);
or UO_1234 (O_1234,N_24985,N_24903);
and UO_1235 (O_1235,N_24805,N_24841);
nand UO_1236 (O_1236,N_24972,N_24843);
nand UO_1237 (O_1237,N_24929,N_24974);
or UO_1238 (O_1238,N_24817,N_24992);
or UO_1239 (O_1239,N_24837,N_24842);
xnor UO_1240 (O_1240,N_24939,N_24860);
xor UO_1241 (O_1241,N_24947,N_24909);
nor UO_1242 (O_1242,N_24993,N_24841);
and UO_1243 (O_1243,N_24897,N_24832);
nand UO_1244 (O_1244,N_24879,N_24900);
and UO_1245 (O_1245,N_24833,N_24817);
nor UO_1246 (O_1246,N_24975,N_24882);
and UO_1247 (O_1247,N_24928,N_24890);
nand UO_1248 (O_1248,N_24822,N_24936);
nor UO_1249 (O_1249,N_24928,N_24876);
nand UO_1250 (O_1250,N_24944,N_24986);
nor UO_1251 (O_1251,N_24954,N_24816);
nand UO_1252 (O_1252,N_24957,N_24951);
and UO_1253 (O_1253,N_24828,N_24970);
or UO_1254 (O_1254,N_24894,N_24808);
xnor UO_1255 (O_1255,N_24869,N_24970);
and UO_1256 (O_1256,N_24806,N_24961);
nand UO_1257 (O_1257,N_24895,N_24911);
nor UO_1258 (O_1258,N_24835,N_24968);
or UO_1259 (O_1259,N_24953,N_24933);
or UO_1260 (O_1260,N_24863,N_24915);
xnor UO_1261 (O_1261,N_24848,N_24887);
nor UO_1262 (O_1262,N_24983,N_24914);
or UO_1263 (O_1263,N_24966,N_24976);
nand UO_1264 (O_1264,N_24817,N_24828);
nand UO_1265 (O_1265,N_24950,N_24953);
nand UO_1266 (O_1266,N_24920,N_24939);
nor UO_1267 (O_1267,N_24817,N_24929);
and UO_1268 (O_1268,N_24959,N_24885);
or UO_1269 (O_1269,N_24987,N_24904);
nor UO_1270 (O_1270,N_24815,N_24840);
nand UO_1271 (O_1271,N_24956,N_24873);
xnor UO_1272 (O_1272,N_24914,N_24894);
or UO_1273 (O_1273,N_24917,N_24901);
nand UO_1274 (O_1274,N_24989,N_24809);
nor UO_1275 (O_1275,N_24863,N_24894);
xnor UO_1276 (O_1276,N_24910,N_24990);
and UO_1277 (O_1277,N_24936,N_24878);
xnor UO_1278 (O_1278,N_24895,N_24828);
xor UO_1279 (O_1279,N_24859,N_24923);
nor UO_1280 (O_1280,N_24858,N_24906);
and UO_1281 (O_1281,N_24919,N_24864);
xnor UO_1282 (O_1282,N_24872,N_24862);
nand UO_1283 (O_1283,N_24877,N_24995);
nor UO_1284 (O_1284,N_24960,N_24818);
nor UO_1285 (O_1285,N_24983,N_24874);
or UO_1286 (O_1286,N_24972,N_24998);
nor UO_1287 (O_1287,N_24970,N_24902);
nor UO_1288 (O_1288,N_24859,N_24845);
nand UO_1289 (O_1289,N_24857,N_24932);
xnor UO_1290 (O_1290,N_24828,N_24942);
or UO_1291 (O_1291,N_24815,N_24859);
xnor UO_1292 (O_1292,N_24927,N_24925);
nand UO_1293 (O_1293,N_24887,N_24873);
xnor UO_1294 (O_1294,N_24979,N_24817);
nand UO_1295 (O_1295,N_24979,N_24989);
or UO_1296 (O_1296,N_24899,N_24861);
xor UO_1297 (O_1297,N_24809,N_24889);
or UO_1298 (O_1298,N_24986,N_24819);
or UO_1299 (O_1299,N_24941,N_24955);
xor UO_1300 (O_1300,N_24928,N_24871);
and UO_1301 (O_1301,N_24978,N_24897);
and UO_1302 (O_1302,N_24872,N_24835);
and UO_1303 (O_1303,N_24816,N_24984);
nand UO_1304 (O_1304,N_24873,N_24896);
nor UO_1305 (O_1305,N_24839,N_24965);
nor UO_1306 (O_1306,N_24910,N_24856);
nor UO_1307 (O_1307,N_24959,N_24914);
and UO_1308 (O_1308,N_24949,N_24820);
nand UO_1309 (O_1309,N_24980,N_24860);
nand UO_1310 (O_1310,N_24939,N_24814);
xor UO_1311 (O_1311,N_24912,N_24899);
nor UO_1312 (O_1312,N_24831,N_24858);
nor UO_1313 (O_1313,N_24960,N_24827);
or UO_1314 (O_1314,N_24901,N_24913);
and UO_1315 (O_1315,N_24934,N_24825);
and UO_1316 (O_1316,N_24928,N_24804);
nor UO_1317 (O_1317,N_24878,N_24837);
or UO_1318 (O_1318,N_24985,N_24879);
xor UO_1319 (O_1319,N_24919,N_24891);
nand UO_1320 (O_1320,N_24814,N_24879);
nor UO_1321 (O_1321,N_24859,N_24989);
nand UO_1322 (O_1322,N_24952,N_24968);
nand UO_1323 (O_1323,N_24864,N_24995);
xnor UO_1324 (O_1324,N_24940,N_24912);
and UO_1325 (O_1325,N_24905,N_24875);
nand UO_1326 (O_1326,N_24850,N_24953);
nand UO_1327 (O_1327,N_24828,N_24912);
or UO_1328 (O_1328,N_24811,N_24998);
nor UO_1329 (O_1329,N_24880,N_24899);
nor UO_1330 (O_1330,N_24982,N_24917);
and UO_1331 (O_1331,N_24886,N_24890);
xor UO_1332 (O_1332,N_24950,N_24835);
nor UO_1333 (O_1333,N_24825,N_24986);
xor UO_1334 (O_1334,N_24843,N_24847);
xor UO_1335 (O_1335,N_24829,N_24891);
or UO_1336 (O_1336,N_24802,N_24986);
nand UO_1337 (O_1337,N_24945,N_24849);
nand UO_1338 (O_1338,N_24832,N_24841);
or UO_1339 (O_1339,N_24899,N_24965);
xnor UO_1340 (O_1340,N_24996,N_24930);
nand UO_1341 (O_1341,N_24853,N_24872);
and UO_1342 (O_1342,N_24990,N_24806);
and UO_1343 (O_1343,N_24987,N_24988);
or UO_1344 (O_1344,N_24925,N_24837);
or UO_1345 (O_1345,N_24832,N_24928);
and UO_1346 (O_1346,N_24890,N_24914);
or UO_1347 (O_1347,N_24833,N_24984);
nand UO_1348 (O_1348,N_24893,N_24838);
and UO_1349 (O_1349,N_24817,N_24864);
or UO_1350 (O_1350,N_24802,N_24880);
nand UO_1351 (O_1351,N_24850,N_24908);
nand UO_1352 (O_1352,N_24859,N_24951);
and UO_1353 (O_1353,N_24808,N_24827);
or UO_1354 (O_1354,N_24889,N_24927);
nand UO_1355 (O_1355,N_24906,N_24815);
or UO_1356 (O_1356,N_24975,N_24823);
nor UO_1357 (O_1357,N_24919,N_24895);
nand UO_1358 (O_1358,N_24969,N_24869);
xor UO_1359 (O_1359,N_24956,N_24817);
and UO_1360 (O_1360,N_24926,N_24911);
nand UO_1361 (O_1361,N_24838,N_24992);
and UO_1362 (O_1362,N_24956,N_24989);
nor UO_1363 (O_1363,N_24903,N_24878);
and UO_1364 (O_1364,N_24954,N_24959);
or UO_1365 (O_1365,N_24958,N_24898);
nand UO_1366 (O_1366,N_24946,N_24925);
nor UO_1367 (O_1367,N_24942,N_24876);
nor UO_1368 (O_1368,N_24976,N_24841);
and UO_1369 (O_1369,N_24877,N_24905);
or UO_1370 (O_1370,N_24922,N_24980);
nor UO_1371 (O_1371,N_24892,N_24966);
nor UO_1372 (O_1372,N_24850,N_24848);
nand UO_1373 (O_1373,N_24919,N_24986);
nand UO_1374 (O_1374,N_24977,N_24837);
nor UO_1375 (O_1375,N_24864,N_24934);
and UO_1376 (O_1376,N_24873,N_24833);
nand UO_1377 (O_1377,N_24971,N_24949);
and UO_1378 (O_1378,N_24897,N_24915);
xnor UO_1379 (O_1379,N_24883,N_24801);
xor UO_1380 (O_1380,N_24827,N_24921);
or UO_1381 (O_1381,N_24885,N_24810);
and UO_1382 (O_1382,N_24956,N_24952);
nor UO_1383 (O_1383,N_24853,N_24962);
nor UO_1384 (O_1384,N_24943,N_24982);
nor UO_1385 (O_1385,N_24810,N_24864);
nand UO_1386 (O_1386,N_24997,N_24875);
xnor UO_1387 (O_1387,N_24867,N_24883);
nor UO_1388 (O_1388,N_24900,N_24858);
xor UO_1389 (O_1389,N_24966,N_24900);
nor UO_1390 (O_1390,N_24828,N_24857);
xor UO_1391 (O_1391,N_24831,N_24806);
nor UO_1392 (O_1392,N_24823,N_24800);
nand UO_1393 (O_1393,N_24978,N_24973);
nand UO_1394 (O_1394,N_24858,N_24850);
nand UO_1395 (O_1395,N_24818,N_24977);
nand UO_1396 (O_1396,N_24826,N_24939);
and UO_1397 (O_1397,N_24863,N_24949);
and UO_1398 (O_1398,N_24887,N_24853);
nand UO_1399 (O_1399,N_24982,N_24969);
nor UO_1400 (O_1400,N_24804,N_24909);
and UO_1401 (O_1401,N_24829,N_24980);
nand UO_1402 (O_1402,N_24819,N_24966);
nor UO_1403 (O_1403,N_24871,N_24803);
xnor UO_1404 (O_1404,N_24903,N_24811);
xor UO_1405 (O_1405,N_24883,N_24857);
and UO_1406 (O_1406,N_24984,N_24873);
nor UO_1407 (O_1407,N_24974,N_24881);
xnor UO_1408 (O_1408,N_24862,N_24984);
or UO_1409 (O_1409,N_24943,N_24848);
and UO_1410 (O_1410,N_24865,N_24904);
and UO_1411 (O_1411,N_24915,N_24937);
or UO_1412 (O_1412,N_24842,N_24900);
nand UO_1413 (O_1413,N_24989,N_24888);
nor UO_1414 (O_1414,N_24831,N_24898);
and UO_1415 (O_1415,N_24971,N_24958);
nor UO_1416 (O_1416,N_24817,N_24842);
or UO_1417 (O_1417,N_24907,N_24913);
nor UO_1418 (O_1418,N_24846,N_24819);
xor UO_1419 (O_1419,N_24802,N_24990);
nor UO_1420 (O_1420,N_24832,N_24862);
nor UO_1421 (O_1421,N_24847,N_24900);
and UO_1422 (O_1422,N_24847,N_24883);
xor UO_1423 (O_1423,N_24912,N_24834);
xnor UO_1424 (O_1424,N_24911,N_24849);
nand UO_1425 (O_1425,N_24871,N_24924);
nand UO_1426 (O_1426,N_24997,N_24842);
and UO_1427 (O_1427,N_24813,N_24866);
and UO_1428 (O_1428,N_24816,N_24873);
nand UO_1429 (O_1429,N_24835,N_24943);
nand UO_1430 (O_1430,N_24915,N_24941);
or UO_1431 (O_1431,N_24967,N_24892);
nor UO_1432 (O_1432,N_24869,N_24968);
and UO_1433 (O_1433,N_24818,N_24855);
or UO_1434 (O_1434,N_24805,N_24955);
nor UO_1435 (O_1435,N_24854,N_24954);
nand UO_1436 (O_1436,N_24972,N_24877);
xnor UO_1437 (O_1437,N_24957,N_24959);
and UO_1438 (O_1438,N_24910,N_24837);
xnor UO_1439 (O_1439,N_24874,N_24858);
and UO_1440 (O_1440,N_24961,N_24956);
nand UO_1441 (O_1441,N_24827,N_24819);
nor UO_1442 (O_1442,N_24806,N_24855);
nand UO_1443 (O_1443,N_24866,N_24841);
nand UO_1444 (O_1444,N_24969,N_24814);
or UO_1445 (O_1445,N_24870,N_24826);
or UO_1446 (O_1446,N_24805,N_24949);
and UO_1447 (O_1447,N_24903,N_24858);
and UO_1448 (O_1448,N_24814,N_24985);
or UO_1449 (O_1449,N_24894,N_24903);
nor UO_1450 (O_1450,N_24960,N_24890);
nor UO_1451 (O_1451,N_24962,N_24869);
nor UO_1452 (O_1452,N_24879,N_24857);
xnor UO_1453 (O_1453,N_24861,N_24921);
nand UO_1454 (O_1454,N_24896,N_24951);
or UO_1455 (O_1455,N_24805,N_24946);
and UO_1456 (O_1456,N_24834,N_24961);
and UO_1457 (O_1457,N_24950,N_24813);
xnor UO_1458 (O_1458,N_24933,N_24824);
xor UO_1459 (O_1459,N_24935,N_24939);
or UO_1460 (O_1460,N_24965,N_24929);
nand UO_1461 (O_1461,N_24828,N_24928);
nand UO_1462 (O_1462,N_24889,N_24967);
and UO_1463 (O_1463,N_24984,N_24963);
nand UO_1464 (O_1464,N_24942,N_24983);
nand UO_1465 (O_1465,N_24951,N_24804);
nand UO_1466 (O_1466,N_24987,N_24804);
nand UO_1467 (O_1467,N_24822,N_24882);
and UO_1468 (O_1468,N_24816,N_24843);
or UO_1469 (O_1469,N_24946,N_24986);
nand UO_1470 (O_1470,N_24826,N_24940);
xor UO_1471 (O_1471,N_24981,N_24840);
or UO_1472 (O_1472,N_24828,N_24924);
or UO_1473 (O_1473,N_24816,N_24821);
xnor UO_1474 (O_1474,N_24838,N_24981);
and UO_1475 (O_1475,N_24976,N_24904);
nor UO_1476 (O_1476,N_24805,N_24977);
or UO_1477 (O_1477,N_24913,N_24987);
nor UO_1478 (O_1478,N_24915,N_24821);
xor UO_1479 (O_1479,N_24978,N_24850);
xnor UO_1480 (O_1480,N_24832,N_24852);
and UO_1481 (O_1481,N_24827,N_24880);
or UO_1482 (O_1482,N_24818,N_24854);
and UO_1483 (O_1483,N_24988,N_24882);
and UO_1484 (O_1484,N_24801,N_24875);
nor UO_1485 (O_1485,N_24839,N_24800);
nand UO_1486 (O_1486,N_24983,N_24852);
and UO_1487 (O_1487,N_24836,N_24876);
nor UO_1488 (O_1488,N_24984,N_24901);
nand UO_1489 (O_1489,N_24993,N_24950);
or UO_1490 (O_1490,N_24925,N_24897);
and UO_1491 (O_1491,N_24852,N_24937);
nand UO_1492 (O_1492,N_24961,N_24945);
nor UO_1493 (O_1493,N_24994,N_24989);
and UO_1494 (O_1494,N_24872,N_24807);
xnor UO_1495 (O_1495,N_24800,N_24964);
xnor UO_1496 (O_1496,N_24973,N_24993);
or UO_1497 (O_1497,N_24881,N_24942);
nor UO_1498 (O_1498,N_24916,N_24825);
or UO_1499 (O_1499,N_24846,N_24823);
xnor UO_1500 (O_1500,N_24898,N_24894);
nor UO_1501 (O_1501,N_24907,N_24972);
nand UO_1502 (O_1502,N_24896,N_24870);
xor UO_1503 (O_1503,N_24822,N_24878);
nor UO_1504 (O_1504,N_24935,N_24896);
xor UO_1505 (O_1505,N_24885,N_24901);
and UO_1506 (O_1506,N_24843,N_24811);
nand UO_1507 (O_1507,N_24992,N_24986);
or UO_1508 (O_1508,N_24976,N_24875);
xor UO_1509 (O_1509,N_24949,N_24965);
and UO_1510 (O_1510,N_24806,N_24875);
and UO_1511 (O_1511,N_24957,N_24997);
and UO_1512 (O_1512,N_24958,N_24987);
nor UO_1513 (O_1513,N_24984,N_24915);
or UO_1514 (O_1514,N_24868,N_24857);
and UO_1515 (O_1515,N_24986,N_24808);
nand UO_1516 (O_1516,N_24923,N_24842);
or UO_1517 (O_1517,N_24915,N_24940);
xnor UO_1518 (O_1518,N_24987,N_24914);
nand UO_1519 (O_1519,N_24941,N_24839);
and UO_1520 (O_1520,N_24835,N_24854);
and UO_1521 (O_1521,N_24982,N_24971);
nand UO_1522 (O_1522,N_24955,N_24988);
xor UO_1523 (O_1523,N_24884,N_24900);
and UO_1524 (O_1524,N_24969,N_24865);
xnor UO_1525 (O_1525,N_24855,N_24954);
nor UO_1526 (O_1526,N_24899,N_24875);
and UO_1527 (O_1527,N_24842,N_24846);
or UO_1528 (O_1528,N_24856,N_24902);
and UO_1529 (O_1529,N_24840,N_24898);
xor UO_1530 (O_1530,N_24800,N_24896);
nand UO_1531 (O_1531,N_24843,N_24963);
and UO_1532 (O_1532,N_24996,N_24892);
nor UO_1533 (O_1533,N_24956,N_24917);
and UO_1534 (O_1534,N_24848,N_24945);
xor UO_1535 (O_1535,N_24870,N_24802);
and UO_1536 (O_1536,N_24915,N_24993);
and UO_1537 (O_1537,N_24889,N_24860);
or UO_1538 (O_1538,N_24956,N_24971);
nor UO_1539 (O_1539,N_24804,N_24809);
nand UO_1540 (O_1540,N_24902,N_24858);
nor UO_1541 (O_1541,N_24998,N_24948);
and UO_1542 (O_1542,N_24824,N_24872);
nand UO_1543 (O_1543,N_24864,N_24968);
nand UO_1544 (O_1544,N_24901,N_24808);
xnor UO_1545 (O_1545,N_24903,N_24922);
and UO_1546 (O_1546,N_24886,N_24820);
and UO_1547 (O_1547,N_24901,N_24983);
nor UO_1548 (O_1548,N_24996,N_24942);
nor UO_1549 (O_1549,N_24916,N_24891);
nand UO_1550 (O_1550,N_24976,N_24847);
nand UO_1551 (O_1551,N_24866,N_24851);
or UO_1552 (O_1552,N_24823,N_24883);
xnor UO_1553 (O_1553,N_24992,N_24878);
nand UO_1554 (O_1554,N_24937,N_24859);
xor UO_1555 (O_1555,N_24821,N_24980);
nor UO_1556 (O_1556,N_24860,N_24801);
or UO_1557 (O_1557,N_24937,N_24838);
xnor UO_1558 (O_1558,N_24996,N_24983);
or UO_1559 (O_1559,N_24947,N_24825);
xor UO_1560 (O_1560,N_24908,N_24904);
xor UO_1561 (O_1561,N_24855,N_24917);
nand UO_1562 (O_1562,N_24931,N_24813);
or UO_1563 (O_1563,N_24828,N_24894);
nor UO_1564 (O_1564,N_24808,N_24889);
or UO_1565 (O_1565,N_24858,N_24882);
nand UO_1566 (O_1566,N_24958,N_24918);
xnor UO_1567 (O_1567,N_24996,N_24852);
xor UO_1568 (O_1568,N_24968,N_24956);
or UO_1569 (O_1569,N_24989,N_24960);
xor UO_1570 (O_1570,N_24912,N_24890);
or UO_1571 (O_1571,N_24950,N_24965);
and UO_1572 (O_1572,N_24955,N_24857);
xnor UO_1573 (O_1573,N_24937,N_24918);
nor UO_1574 (O_1574,N_24922,N_24928);
nand UO_1575 (O_1575,N_24904,N_24971);
xor UO_1576 (O_1576,N_24926,N_24977);
or UO_1577 (O_1577,N_24818,N_24873);
and UO_1578 (O_1578,N_24850,N_24849);
nand UO_1579 (O_1579,N_24926,N_24813);
or UO_1580 (O_1580,N_24878,N_24951);
nand UO_1581 (O_1581,N_24886,N_24901);
nor UO_1582 (O_1582,N_24836,N_24917);
or UO_1583 (O_1583,N_24822,N_24950);
nand UO_1584 (O_1584,N_24950,N_24888);
nand UO_1585 (O_1585,N_24889,N_24905);
nand UO_1586 (O_1586,N_24879,N_24921);
or UO_1587 (O_1587,N_24946,N_24992);
nand UO_1588 (O_1588,N_24952,N_24923);
xor UO_1589 (O_1589,N_24977,N_24981);
nor UO_1590 (O_1590,N_24810,N_24944);
or UO_1591 (O_1591,N_24814,N_24891);
or UO_1592 (O_1592,N_24933,N_24888);
xor UO_1593 (O_1593,N_24963,N_24946);
nand UO_1594 (O_1594,N_24893,N_24971);
or UO_1595 (O_1595,N_24810,N_24994);
nand UO_1596 (O_1596,N_24802,N_24997);
nor UO_1597 (O_1597,N_24889,N_24963);
xnor UO_1598 (O_1598,N_24896,N_24966);
xnor UO_1599 (O_1599,N_24840,N_24899);
nand UO_1600 (O_1600,N_24875,N_24958);
xnor UO_1601 (O_1601,N_24993,N_24876);
xor UO_1602 (O_1602,N_24976,N_24889);
nand UO_1603 (O_1603,N_24961,N_24901);
nand UO_1604 (O_1604,N_24821,N_24933);
nand UO_1605 (O_1605,N_24962,N_24912);
nor UO_1606 (O_1606,N_24981,N_24894);
nor UO_1607 (O_1607,N_24945,N_24821);
xnor UO_1608 (O_1608,N_24873,N_24944);
or UO_1609 (O_1609,N_24926,N_24963);
xor UO_1610 (O_1610,N_24968,N_24840);
nand UO_1611 (O_1611,N_24819,N_24924);
or UO_1612 (O_1612,N_24913,N_24972);
or UO_1613 (O_1613,N_24995,N_24888);
nor UO_1614 (O_1614,N_24970,N_24906);
and UO_1615 (O_1615,N_24819,N_24847);
xnor UO_1616 (O_1616,N_24814,N_24895);
nor UO_1617 (O_1617,N_24861,N_24952);
xor UO_1618 (O_1618,N_24928,N_24931);
nor UO_1619 (O_1619,N_24822,N_24930);
and UO_1620 (O_1620,N_24968,N_24976);
or UO_1621 (O_1621,N_24877,N_24863);
nand UO_1622 (O_1622,N_24806,N_24928);
nor UO_1623 (O_1623,N_24956,N_24947);
and UO_1624 (O_1624,N_24800,N_24859);
nand UO_1625 (O_1625,N_24915,N_24837);
or UO_1626 (O_1626,N_24976,N_24869);
and UO_1627 (O_1627,N_24844,N_24868);
or UO_1628 (O_1628,N_24966,N_24861);
nand UO_1629 (O_1629,N_24959,N_24924);
and UO_1630 (O_1630,N_24968,N_24879);
nor UO_1631 (O_1631,N_24992,N_24888);
xor UO_1632 (O_1632,N_24991,N_24998);
and UO_1633 (O_1633,N_24812,N_24978);
nor UO_1634 (O_1634,N_24905,N_24934);
or UO_1635 (O_1635,N_24956,N_24810);
or UO_1636 (O_1636,N_24900,N_24851);
nor UO_1637 (O_1637,N_24875,N_24996);
and UO_1638 (O_1638,N_24859,N_24953);
and UO_1639 (O_1639,N_24809,N_24814);
or UO_1640 (O_1640,N_24951,N_24996);
or UO_1641 (O_1641,N_24969,N_24928);
xnor UO_1642 (O_1642,N_24816,N_24952);
or UO_1643 (O_1643,N_24800,N_24911);
nor UO_1644 (O_1644,N_24998,N_24851);
and UO_1645 (O_1645,N_24948,N_24879);
xor UO_1646 (O_1646,N_24812,N_24937);
nor UO_1647 (O_1647,N_24800,N_24970);
or UO_1648 (O_1648,N_24852,N_24949);
nor UO_1649 (O_1649,N_24900,N_24951);
nor UO_1650 (O_1650,N_24856,N_24901);
xor UO_1651 (O_1651,N_24992,N_24905);
or UO_1652 (O_1652,N_24967,N_24870);
nand UO_1653 (O_1653,N_24924,N_24997);
and UO_1654 (O_1654,N_24862,N_24800);
xor UO_1655 (O_1655,N_24855,N_24808);
nand UO_1656 (O_1656,N_24808,N_24823);
nand UO_1657 (O_1657,N_24820,N_24954);
nand UO_1658 (O_1658,N_24840,N_24993);
or UO_1659 (O_1659,N_24921,N_24859);
nand UO_1660 (O_1660,N_24946,N_24893);
nand UO_1661 (O_1661,N_24929,N_24857);
nand UO_1662 (O_1662,N_24944,N_24961);
nand UO_1663 (O_1663,N_24805,N_24933);
xor UO_1664 (O_1664,N_24814,N_24820);
nor UO_1665 (O_1665,N_24949,N_24943);
nor UO_1666 (O_1666,N_24808,N_24875);
and UO_1667 (O_1667,N_24956,N_24839);
nor UO_1668 (O_1668,N_24902,N_24921);
nand UO_1669 (O_1669,N_24964,N_24838);
nand UO_1670 (O_1670,N_24865,N_24847);
or UO_1671 (O_1671,N_24806,N_24991);
or UO_1672 (O_1672,N_24998,N_24929);
and UO_1673 (O_1673,N_24903,N_24815);
and UO_1674 (O_1674,N_24955,N_24867);
and UO_1675 (O_1675,N_24892,N_24861);
nor UO_1676 (O_1676,N_24938,N_24844);
or UO_1677 (O_1677,N_24880,N_24971);
nand UO_1678 (O_1678,N_24876,N_24875);
and UO_1679 (O_1679,N_24929,N_24822);
nor UO_1680 (O_1680,N_24806,N_24878);
nor UO_1681 (O_1681,N_24964,N_24924);
nor UO_1682 (O_1682,N_24988,N_24970);
and UO_1683 (O_1683,N_24828,N_24971);
or UO_1684 (O_1684,N_24877,N_24886);
xnor UO_1685 (O_1685,N_24885,N_24909);
nand UO_1686 (O_1686,N_24944,N_24826);
xnor UO_1687 (O_1687,N_24883,N_24836);
or UO_1688 (O_1688,N_24843,N_24913);
xnor UO_1689 (O_1689,N_24832,N_24813);
xor UO_1690 (O_1690,N_24811,N_24871);
or UO_1691 (O_1691,N_24921,N_24998);
xor UO_1692 (O_1692,N_24891,N_24867);
or UO_1693 (O_1693,N_24813,N_24851);
and UO_1694 (O_1694,N_24965,N_24873);
or UO_1695 (O_1695,N_24838,N_24995);
or UO_1696 (O_1696,N_24845,N_24808);
xnor UO_1697 (O_1697,N_24841,N_24844);
nand UO_1698 (O_1698,N_24948,N_24841);
nand UO_1699 (O_1699,N_24815,N_24907);
nand UO_1700 (O_1700,N_24938,N_24882);
nor UO_1701 (O_1701,N_24858,N_24857);
nor UO_1702 (O_1702,N_24946,N_24815);
nand UO_1703 (O_1703,N_24889,N_24887);
and UO_1704 (O_1704,N_24945,N_24873);
and UO_1705 (O_1705,N_24863,N_24809);
xor UO_1706 (O_1706,N_24990,N_24902);
and UO_1707 (O_1707,N_24951,N_24949);
and UO_1708 (O_1708,N_24948,N_24811);
xnor UO_1709 (O_1709,N_24901,N_24969);
or UO_1710 (O_1710,N_24882,N_24921);
nor UO_1711 (O_1711,N_24955,N_24821);
or UO_1712 (O_1712,N_24860,N_24931);
nand UO_1713 (O_1713,N_24863,N_24844);
xnor UO_1714 (O_1714,N_24899,N_24854);
xnor UO_1715 (O_1715,N_24835,N_24982);
xor UO_1716 (O_1716,N_24961,N_24803);
or UO_1717 (O_1717,N_24886,N_24947);
nand UO_1718 (O_1718,N_24980,N_24903);
xnor UO_1719 (O_1719,N_24974,N_24912);
nor UO_1720 (O_1720,N_24894,N_24893);
xor UO_1721 (O_1721,N_24845,N_24881);
and UO_1722 (O_1722,N_24871,N_24848);
and UO_1723 (O_1723,N_24879,N_24800);
xnor UO_1724 (O_1724,N_24905,N_24958);
and UO_1725 (O_1725,N_24816,N_24912);
nand UO_1726 (O_1726,N_24903,N_24962);
xnor UO_1727 (O_1727,N_24981,N_24873);
nand UO_1728 (O_1728,N_24915,N_24849);
and UO_1729 (O_1729,N_24866,N_24831);
and UO_1730 (O_1730,N_24979,N_24834);
or UO_1731 (O_1731,N_24956,N_24864);
nand UO_1732 (O_1732,N_24911,N_24941);
or UO_1733 (O_1733,N_24931,N_24972);
xor UO_1734 (O_1734,N_24807,N_24981);
nor UO_1735 (O_1735,N_24926,N_24920);
xor UO_1736 (O_1736,N_24821,N_24954);
nor UO_1737 (O_1737,N_24984,N_24997);
and UO_1738 (O_1738,N_24949,N_24942);
nand UO_1739 (O_1739,N_24933,N_24978);
and UO_1740 (O_1740,N_24954,N_24971);
xnor UO_1741 (O_1741,N_24871,N_24991);
nand UO_1742 (O_1742,N_24817,N_24985);
xnor UO_1743 (O_1743,N_24905,N_24819);
nor UO_1744 (O_1744,N_24947,N_24810);
nor UO_1745 (O_1745,N_24877,N_24898);
nor UO_1746 (O_1746,N_24962,N_24897);
nand UO_1747 (O_1747,N_24848,N_24973);
nand UO_1748 (O_1748,N_24824,N_24972);
xnor UO_1749 (O_1749,N_24918,N_24813);
and UO_1750 (O_1750,N_24972,N_24996);
nor UO_1751 (O_1751,N_24947,N_24940);
nor UO_1752 (O_1752,N_24818,N_24843);
and UO_1753 (O_1753,N_24904,N_24948);
and UO_1754 (O_1754,N_24902,N_24810);
and UO_1755 (O_1755,N_24917,N_24935);
nor UO_1756 (O_1756,N_24984,N_24869);
nand UO_1757 (O_1757,N_24853,N_24967);
and UO_1758 (O_1758,N_24815,N_24841);
nor UO_1759 (O_1759,N_24831,N_24947);
or UO_1760 (O_1760,N_24992,N_24932);
or UO_1761 (O_1761,N_24866,N_24972);
or UO_1762 (O_1762,N_24818,N_24952);
nand UO_1763 (O_1763,N_24896,N_24950);
xnor UO_1764 (O_1764,N_24928,N_24803);
and UO_1765 (O_1765,N_24801,N_24994);
nand UO_1766 (O_1766,N_24938,N_24963);
nor UO_1767 (O_1767,N_24997,N_24849);
and UO_1768 (O_1768,N_24969,N_24904);
nor UO_1769 (O_1769,N_24833,N_24901);
nor UO_1770 (O_1770,N_24926,N_24918);
nor UO_1771 (O_1771,N_24856,N_24814);
xnor UO_1772 (O_1772,N_24992,N_24981);
nand UO_1773 (O_1773,N_24853,N_24952);
nand UO_1774 (O_1774,N_24810,N_24966);
and UO_1775 (O_1775,N_24912,N_24906);
and UO_1776 (O_1776,N_24810,N_24892);
nand UO_1777 (O_1777,N_24996,N_24954);
nand UO_1778 (O_1778,N_24806,N_24967);
xor UO_1779 (O_1779,N_24951,N_24963);
or UO_1780 (O_1780,N_24987,N_24929);
or UO_1781 (O_1781,N_24978,N_24979);
or UO_1782 (O_1782,N_24954,N_24847);
and UO_1783 (O_1783,N_24894,N_24886);
and UO_1784 (O_1784,N_24809,N_24977);
and UO_1785 (O_1785,N_24807,N_24867);
nand UO_1786 (O_1786,N_24849,N_24949);
or UO_1787 (O_1787,N_24895,N_24887);
and UO_1788 (O_1788,N_24973,N_24948);
or UO_1789 (O_1789,N_24997,N_24857);
nor UO_1790 (O_1790,N_24969,N_24887);
or UO_1791 (O_1791,N_24931,N_24912);
nand UO_1792 (O_1792,N_24870,N_24889);
or UO_1793 (O_1793,N_24864,N_24886);
or UO_1794 (O_1794,N_24825,N_24862);
nor UO_1795 (O_1795,N_24867,N_24855);
nand UO_1796 (O_1796,N_24961,N_24908);
nor UO_1797 (O_1797,N_24964,N_24929);
xor UO_1798 (O_1798,N_24985,N_24888);
or UO_1799 (O_1799,N_24824,N_24967);
nor UO_1800 (O_1800,N_24880,N_24838);
xnor UO_1801 (O_1801,N_24855,N_24903);
xor UO_1802 (O_1802,N_24934,N_24943);
xor UO_1803 (O_1803,N_24983,N_24893);
or UO_1804 (O_1804,N_24922,N_24991);
xnor UO_1805 (O_1805,N_24882,N_24840);
nand UO_1806 (O_1806,N_24834,N_24848);
or UO_1807 (O_1807,N_24929,N_24926);
or UO_1808 (O_1808,N_24998,N_24996);
and UO_1809 (O_1809,N_24912,N_24911);
nand UO_1810 (O_1810,N_24860,N_24963);
and UO_1811 (O_1811,N_24886,N_24979);
or UO_1812 (O_1812,N_24888,N_24926);
or UO_1813 (O_1813,N_24994,N_24864);
nor UO_1814 (O_1814,N_24983,N_24939);
nand UO_1815 (O_1815,N_24978,N_24900);
nand UO_1816 (O_1816,N_24831,N_24909);
nand UO_1817 (O_1817,N_24814,N_24964);
and UO_1818 (O_1818,N_24914,N_24856);
nand UO_1819 (O_1819,N_24998,N_24997);
nor UO_1820 (O_1820,N_24894,N_24850);
and UO_1821 (O_1821,N_24807,N_24999);
or UO_1822 (O_1822,N_24890,N_24978);
xnor UO_1823 (O_1823,N_24949,N_24844);
or UO_1824 (O_1824,N_24973,N_24856);
and UO_1825 (O_1825,N_24812,N_24833);
nor UO_1826 (O_1826,N_24969,N_24834);
xor UO_1827 (O_1827,N_24974,N_24848);
xor UO_1828 (O_1828,N_24901,N_24944);
nor UO_1829 (O_1829,N_24827,N_24942);
xnor UO_1830 (O_1830,N_24814,N_24941);
and UO_1831 (O_1831,N_24939,N_24841);
nor UO_1832 (O_1832,N_24968,N_24883);
and UO_1833 (O_1833,N_24988,N_24804);
nand UO_1834 (O_1834,N_24982,N_24841);
and UO_1835 (O_1835,N_24815,N_24997);
nor UO_1836 (O_1836,N_24946,N_24880);
or UO_1837 (O_1837,N_24871,N_24814);
and UO_1838 (O_1838,N_24838,N_24986);
nor UO_1839 (O_1839,N_24958,N_24982);
nor UO_1840 (O_1840,N_24851,N_24863);
nor UO_1841 (O_1841,N_24904,N_24950);
xnor UO_1842 (O_1842,N_24974,N_24989);
nand UO_1843 (O_1843,N_24952,N_24844);
nor UO_1844 (O_1844,N_24863,N_24937);
xor UO_1845 (O_1845,N_24824,N_24809);
nand UO_1846 (O_1846,N_24904,N_24888);
nand UO_1847 (O_1847,N_24899,N_24878);
xnor UO_1848 (O_1848,N_24959,N_24890);
xor UO_1849 (O_1849,N_24823,N_24976);
or UO_1850 (O_1850,N_24828,N_24875);
nor UO_1851 (O_1851,N_24902,N_24943);
and UO_1852 (O_1852,N_24936,N_24816);
nand UO_1853 (O_1853,N_24910,N_24892);
nand UO_1854 (O_1854,N_24825,N_24849);
nor UO_1855 (O_1855,N_24962,N_24862);
xor UO_1856 (O_1856,N_24995,N_24848);
xnor UO_1857 (O_1857,N_24977,N_24844);
nand UO_1858 (O_1858,N_24849,N_24989);
nor UO_1859 (O_1859,N_24921,N_24885);
nand UO_1860 (O_1860,N_24864,N_24907);
nand UO_1861 (O_1861,N_24835,N_24906);
or UO_1862 (O_1862,N_24904,N_24984);
and UO_1863 (O_1863,N_24939,N_24927);
nor UO_1864 (O_1864,N_24863,N_24896);
nand UO_1865 (O_1865,N_24966,N_24968);
nand UO_1866 (O_1866,N_24927,N_24999);
nor UO_1867 (O_1867,N_24986,N_24850);
xor UO_1868 (O_1868,N_24997,N_24968);
and UO_1869 (O_1869,N_24873,N_24928);
or UO_1870 (O_1870,N_24950,N_24873);
nor UO_1871 (O_1871,N_24820,N_24837);
xnor UO_1872 (O_1872,N_24952,N_24826);
nor UO_1873 (O_1873,N_24979,N_24862);
or UO_1874 (O_1874,N_24911,N_24959);
nand UO_1875 (O_1875,N_24850,N_24831);
xor UO_1876 (O_1876,N_24869,N_24920);
nand UO_1877 (O_1877,N_24942,N_24852);
and UO_1878 (O_1878,N_24834,N_24894);
or UO_1879 (O_1879,N_24859,N_24929);
nand UO_1880 (O_1880,N_24810,N_24918);
nor UO_1881 (O_1881,N_24937,N_24873);
and UO_1882 (O_1882,N_24812,N_24814);
or UO_1883 (O_1883,N_24843,N_24864);
nand UO_1884 (O_1884,N_24931,N_24886);
nand UO_1885 (O_1885,N_24965,N_24971);
and UO_1886 (O_1886,N_24956,N_24863);
xor UO_1887 (O_1887,N_24959,N_24921);
nand UO_1888 (O_1888,N_24935,N_24979);
xor UO_1889 (O_1889,N_24895,N_24892);
xor UO_1890 (O_1890,N_24844,N_24846);
nand UO_1891 (O_1891,N_24926,N_24989);
nor UO_1892 (O_1892,N_24936,N_24978);
nand UO_1893 (O_1893,N_24999,N_24847);
nor UO_1894 (O_1894,N_24915,N_24898);
or UO_1895 (O_1895,N_24986,N_24976);
nand UO_1896 (O_1896,N_24956,N_24859);
and UO_1897 (O_1897,N_24922,N_24926);
nand UO_1898 (O_1898,N_24938,N_24920);
nor UO_1899 (O_1899,N_24977,N_24824);
and UO_1900 (O_1900,N_24934,N_24865);
xnor UO_1901 (O_1901,N_24803,N_24808);
nor UO_1902 (O_1902,N_24848,N_24869);
nor UO_1903 (O_1903,N_24922,N_24896);
nor UO_1904 (O_1904,N_24838,N_24940);
or UO_1905 (O_1905,N_24988,N_24890);
xor UO_1906 (O_1906,N_24970,N_24841);
nand UO_1907 (O_1907,N_24866,N_24981);
nand UO_1908 (O_1908,N_24812,N_24887);
nor UO_1909 (O_1909,N_24984,N_24986);
and UO_1910 (O_1910,N_24899,N_24985);
and UO_1911 (O_1911,N_24941,N_24872);
nor UO_1912 (O_1912,N_24883,N_24928);
nand UO_1913 (O_1913,N_24913,N_24812);
and UO_1914 (O_1914,N_24871,N_24834);
nor UO_1915 (O_1915,N_24909,N_24881);
and UO_1916 (O_1916,N_24892,N_24928);
and UO_1917 (O_1917,N_24882,N_24879);
and UO_1918 (O_1918,N_24897,N_24810);
or UO_1919 (O_1919,N_24944,N_24843);
or UO_1920 (O_1920,N_24833,N_24962);
xor UO_1921 (O_1921,N_24949,N_24845);
nor UO_1922 (O_1922,N_24822,N_24911);
and UO_1923 (O_1923,N_24959,N_24833);
nand UO_1924 (O_1924,N_24820,N_24871);
nand UO_1925 (O_1925,N_24905,N_24926);
nand UO_1926 (O_1926,N_24962,N_24861);
or UO_1927 (O_1927,N_24827,N_24886);
and UO_1928 (O_1928,N_24838,N_24905);
xor UO_1929 (O_1929,N_24918,N_24930);
and UO_1930 (O_1930,N_24963,N_24835);
xor UO_1931 (O_1931,N_24929,N_24976);
nand UO_1932 (O_1932,N_24939,N_24873);
nand UO_1933 (O_1933,N_24823,N_24894);
or UO_1934 (O_1934,N_24948,N_24997);
or UO_1935 (O_1935,N_24824,N_24993);
nor UO_1936 (O_1936,N_24879,N_24997);
nand UO_1937 (O_1937,N_24804,N_24923);
nand UO_1938 (O_1938,N_24849,N_24812);
xor UO_1939 (O_1939,N_24864,N_24899);
nand UO_1940 (O_1940,N_24839,N_24926);
or UO_1941 (O_1941,N_24875,N_24959);
xnor UO_1942 (O_1942,N_24825,N_24895);
xor UO_1943 (O_1943,N_24865,N_24856);
xnor UO_1944 (O_1944,N_24947,N_24935);
nor UO_1945 (O_1945,N_24829,N_24993);
nor UO_1946 (O_1946,N_24820,N_24877);
nor UO_1947 (O_1947,N_24826,N_24971);
xor UO_1948 (O_1948,N_24838,N_24881);
xnor UO_1949 (O_1949,N_24974,N_24910);
nor UO_1950 (O_1950,N_24831,N_24938);
or UO_1951 (O_1951,N_24916,N_24954);
nor UO_1952 (O_1952,N_24988,N_24897);
nor UO_1953 (O_1953,N_24864,N_24917);
xor UO_1954 (O_1954,N_24845,N_24805);
xnor UO_1955 (O_1955,N_24985,N_24933);
xnor UO_1956 (O_1956,N_24840,N_24868);
nor UO_1957 (O_1957,N_24801,N_24959);
and UO_1958 (O_1958,N_24975,N_24875);
and UO_1959 (O_1959,N_24934,N_24921);
nor UO_1960 (O_1960,N_24973,N_24966);
nand UO_1961 (O_1961,N_24974,N_24997);
nand UO_1962 (O_1962,N_24930,N_24999);
nand UO_1963 (O_1963,N_24894,N_24984);
xnor UO_1964 (O_1964,N_24935,N_24959);
xor UO_1965 (O_1965,N_24812,N_24941);
or UO_1966 (O_1966,N_24948,N_24909);
and UO_1967 (O_1967,N_24966,N_24989);
nand UO_1968 (O_1968,N_24872,N_24820);
and UO_1969 (O_1969,N_24951,N_24990);
xor UO_1970 (O_1970,N_24891,N_24961);
nor UO_1971 (O_1971,N_24952,N_24993);
nand UO_1972 (O_1972,N_24813,N_24937);
or UO_1973 (O_1973,N_24881,N_24879);
or UO_1974 (O_1974,N_24993,N_24983);
nor UO_1975 (O_1975,N_24956,N_24890);
xnor UO_1976 (O_1976,N_24891,N_24817);
xnor UO_1977 (O_1977,N_24949,N_24902);
or UO_1978 (O_1978,N_24963,N_24949);
and UO_1979 (O_1979,N_24903,N_24921);
xnor UO_1980 (O_1980,N_24991,N_24899);
or UO_1981 (O_1981,N_24930,N_24949);
or UO_1982 (O_1982,N_24877,N_24923);
nand UO_1983 (O_1983,N_24935,N_24808);
nand UO_1984 (O_1984,N_24862,N_24843);
and UO_1985 (O_1985,N_24977,N_24933);
or UO_1986 (O_1986,N_24947,N_24959);
and UO_1987 (O_1987,N_24957,N_24828);
nor UO_1988 (O_1988,N_24926,N_24807);
or UO_1989 (O_1989,N_24881,N_24882);
and UO_1990 (O_1990,N_24954,N_24818);
and UO_1991 (O_1991,N_24909,N_24876);
and UO_1992 (O_1992,N_24817,N_24907);
xnor UO_1993 (O_1993,N_24956,N_24903);
nand UO_1994 (O_1994,N_24911,N_24982);
or UO_1995 (O_1995,N_24996,N_24863);
and UO_1996 (O_1996,N_24936,N_24873);
and UO_1997 (O_1997,N_24847,N_24896);
xor UO_1998 (O_1998,N_24815,N_24933);
xor UO_1999 (O_1999,N_24971,N_24804);
nor UO_2000 (O_2000,N_24943,N_24871);
or UO_2001 (O_2001,N_24927,N_24902);
nand UO_2002 (O_2002,N_24996,N_24823);
and UO_2003 (O_2003,N_24909,N_24996);
xor UO_2004 (O_2004,N_24913,N_24883);
nor UO_2005 (O_2005,N_24847,N_24945);
or UO_2006 (O_2006,N_24818,N_24841);
nand UO_2007 (O_2007,N_24893,N_24913);
xor UO_2008 (O_2008,N_24888,N_24938);
nor UO_2009 (O_2009,N_24999,N_24917);
nand UO_2010 (O_2010,N_24800,N_24875);
and UO_2011 (O_2011,N_24919,N_24806);
nor UO_2012 (O_2012,N_24969,N_24801);
or UO_2013 (O_2013,N_24937,N_24802);
or UO_2014 (O_2014,N_24978,N_24881);
and UO_2015 (O_2015,N_24983,N_24863);
nor UO_2016 (O_2016,N_24892,N_24813);
xor UO_2017 (O_2017,N_24815,N_24867);
xor UO_2018 (O_2018,N_24875,N_24930);
nor UO_2019 (O_2019,N_24946,N_24875);
xnor UO_2020 (O_2020,N_24949,N_24961);
nor UO_2021 (O_2021,N_24966,N_24820);
nand UO_2022 (O_2022,N_24943,N_24897);
and UO_2023 (O_2023,N_24972,N_24934);
and UO_2024 (O_2024,N_24806,N_24975);
and UO_2025 (O_2025,N_24820,N_24874);
nor UO_2026 (O_2026,N_24932,N_24814);
or UO_2027 (O_2027,N_24907,N_24956);
nor UO_2028 (O_2028,N_24926,N_24917);
nor UO_2029 (O_2029,N_24923,N_24932);
and UO_2030 (O_2030,N_24974,N_24815);
and UO_2031 (O_2031,N_24806,N_24811);
nand UO_2032 (O_2032,N_24815,N_24916);
or UO_2033 (O_2033,N_24973,N_24878);
nor UO_2034 (O_2034,N_24808,N_24902);
and UO_2035 (O_2035,N_24833,N_24995);
or UO_2036 (O_2036,N_24976,N_24997);
and UO_2037 (O_2037,N_24986,N_24967);
xnor UO_2038 (O_2038,N_24829,N_24808);
nand UO_2039 (O_2039,N_24936,N_24900);
xor UO_2040 (O_2040,N_24979,N_24852);
nor UO_2041 (O_2041,N_24832,N_24983);
xnor UO_2042 (O_2042,N_24912,N_24920);
and UO_2043 (O_2043,N_24850,N_24898);
and UO_2044 (O_2044,N_24814,N_24961);
or UO_2045 (O_2045,N_24912,N_24864);
and UO_2046 (O_2046,N_24983,N_24884);
and UO_2047 (O_2047,N_24801,N_24982);
and UO_2048 (O_2048,N_24821,N_24833);
or UO_2049 (O_2049,N_24904,N_24927);
and UO_2050 (O_2050,N_24986,N_24813);
xnor UO_2051 (O_2051,N_24992,N_24990);
nand UO_2052 (O_2052,N_24926,N_24878);
nor UO_2053 (O_2053,N_24832,N_24906);
nand UO_2054 (O_2054,N_24814,N_24951);
nor UO_2055 (O_2055,N_24811,N_24927);
and UO_2056 (O_2056,N_24815,N_24832);
nand UO_2057 (O_2057,N_24845,N_24803);
nor UO_2058 (O_2058,N_24942,N_24967);
nand UO_2059 (O_2059,N_24889,N_24852);
xor UO_2060 (O_2060,N_24967,N_24879);
and UO_2061 (O_2061,N_24948,N_24876);
or UO_2062 (O_2062,N_24853,N_24818);
and UO_2063 (O_2063,N_24983,N_24876);
and UO_2064 (O_2064,N_24852,N_24804);
nand UO_2065 (O_2065,N_24955,N_24952);
or UO_2066 (O_2066,N_24992,N_24822);
nand UO_2067 (O_2067,N_24967,N_24817);
and UO_2068 (O_2068,N_24994,N_24993);
and UO_2069 (O_2069,N_24896,N_24991);
or UO_2070 (O_2070,N_24996,N_24913);
xor UO_2071 (O_2071,N_24936,N_24846);
nand UO_2072 (O_2072,N_24851,N_24809);
or UO_2073 (O_2073,N_24995,N_24912);
or UO_2074 (O_2074,N_24945,N_24809);
and UO_2075 (O_2075,N_24924,N_24829);
xor UO_2076 (O_2076,N_24953,N_24966);
nor UO_2077 (O_2077,N_24860,N_24822);
nand UO_2078 (O_2078,N_24880,N_24814);
nand UO_2079 (O_2079,N_24876,N_24837);
or UO_2080 (O_2080,N_24872,N_24942);
or UO_2081 (O_2081,N_24949,N_24806);
nand UO_2082 (O_2082,N_24832,N_24943);
nand UO_2083 (O_2083,N_24977,N_24813);
nor UO_2084 (O_2084,N_24928,N_24970);
or UO_2085 (O_2085,N_24888,N_24873);
nand UO_2086 (O_2086,N_24979,N_24955);
nand UO_2087 (O_2087,N_24913,N_24870);
nor UO_2088 (O_2088,N_24981,N_24850);
nor UO_2089 (O_2089,N_24895,N_24893);
xnor UO_2090 (O_2090,N_24976,N_24925);
xor UO_2091 (O_2091,N_24867,N_24988);
or UO_2092 (O_2092,N_24993,N_24914);
or UO_2093 (O_2093,N_24886,N_24996);
and UO_2094 (O_2094,N_24950,N_24849);
and UO_2095 (O_2095,N_24890,N_24888);
nand UO_2096 (O_2096,N_24941,N_24882);
and UO_2097 (O_2097,N_24957,N_24904);
nor UO_2098 (O_2098,N_24925,N_24816);
or UO_2099 (O_2099,N_24868,N_24826);
nand UO_2100 (O_2100,N_24841,N_24923);
nor UO_2101 (O_2101,N_24943,N_24956);
and UO_2102 (O_2102,N_24964,N_24908);
and UO_2103 (O_2103,N_24950,N_24940);
xnor UO_2104 (O_2104,N_24816,N_24916);
xor UO_2105 (O_2105,N_24901,N_24935);
xor UO_2106 (O_2106,N_24851,N_24889);
nor UO_2107 (O_2107,N_24956,N_24822);
xor UO_2108 (O_2108,N_24850,N_24902);
nand UO_2109 (O_2109,N_24983,N_24864);
or UO_2110 (O_2110,N_24966,N_24979);
or UO_2111 (O_2111,N_24990,N_24914);
nand UO_2112 (O_2112,N_24979,N_24953);
xor UO_2113 (O_2113,N_24941,N_24852);
nand UO_2114 (O_2114,N_24852,N_24825);
nor UO_2115 (O_2115,N_24953,N_24812);
xnor UO_2116 (O_2116,N_24810,N_24858);
nor UO_2117 (O_2117,N_24904,N_24940);
xnor UO_2118 (O_2118,N_24903,N_24957);
nor UO_2119 (O_2119,N_24962,N_24835);
or UO_2120 (O_2120,N_24860,N_24918);
or UO_2121 (O_2121,N_24935,N_24863);
xor UO_2122 (O_2122,N_24988,N_24895);
nor UO_2123 (O_2123,N_24894,N_24869);
and UO_2124 (O_2124,N_24961,N_24858);
or UO_2125 (O_2125,N_24893,N_24809);
nor UO_2126 (O_2126,N_24965,N_24925);
or UO_2127 (O_2127,N_24952,N_24873);
and UO_2128 (O_2128,N_24860,N_24943);
or UO_2129 (O_2129,N_24887,N_24880);
xor UO_2130 (O_2130,N_24849,N_24902);
xor UO_2131 (O_2131,N_24847,N_24916);
and UO_2132 (O_2132,N_24958,N_24804);
or UO_2133 (O_2133,N_24930,N_24904);
and UO_2134 (O_2134,N_24820,N_24856);
or UO_2135 (O_2135,N_24857,N_24950);
and UO_2136 (O_2136,N_24881,N_24898);
xnor UO_2137 (O_2137,N_24947,N_24957);
or UO_2138 (O_2138,N_24808,N_24814);
nand UO_2139 (O_2139,N_24952,N_24860);
xor UO_2140 (O_2140,N_24832,N_24848);
nand UO_2141 (O_2141,N_24829,N_24834);
xnor UO_2142 (O_2142,N_24812,N_24965);
nor UO_2143 (O_2143,N_24962,N_24920);
xor UO_2144 (O_2144,N_24952,N_24920);
nand UO_2145 (O_2145,N_24818,N_24876);
xor UO_2146 (O_2146,N_24865,N_24814);
xor UO_2147 (O_2147,N_24922,N_24824);
and UO_2148 (O_2148,N_24976,N_24883);
nand UO_2149 (O_2149,N_24912,N_24886);
nor UO_2150 (O_2150,N_24802,N_24968);
nor UO_2151 (O_2151,N_24830,N_24809);
nor UO_2152 (O_2152,N_24985,N_24950);
nand UO_2153 (O_2153,N_24839,N_24891);
and UO_2154 (O_2154,N_24989,N_24992);
nand UO_2155 (O_2155,N_24983,N_24808);
and UO_2156 (O_2156,N_24872,N_24839);
nand UO_2157 (O_2157,N_24855,N_24829);
nor UO_2158 (O_2158,N_24857,N_24992);
xnor UO_2159 (O_2159,N_24848,N_24854);
or UO_2160 (O_2160,N_24904,N_24968);
and UO_2161 (O_2161,N_24916,N_24913);
and UO_2162 (O_2162,N_24837,N_24978);
or UO_2163 (O_2163,N_24801,N_24908);
or UO_2164 (O_2164,N_24965,N_24904);
or UO_2165 (O_2165,N_24801,N_24856);
and UO_2166 (O_2166,N_24950,N_24915);
or UO_2167 (O_2167,N_24846,N_24930);
nand UO_2168 (O_2168,N_24871,N_24841);
nor UO_2169 (O_2169,N_24815,N_24819);
nand UO_2170 (O_2170,N_24804,N_24821);
xnor UO_2171 (O_2171,N_24896,N_24895);
nand UO_2172 (O_2172,N_24829,N_24863);
nand UO_2173 (O_2173,N_24825,N_24954);
and UO_2174 (O_2174,N_24816,N_24836);
xnor UO_2175 (O_2175,N_24872,N_24831);
and UO_2176 (O_2176,N_24800,N_24915);
or UO_2177 (O_2177,N_24910,N_24845);
or UO_2178 (O_2178,N_24963,N_24991);
nor UO_2179 (O_2179,N_24893,N_24837);
and UO_2180 (O_2180,N_24850,N_24890);
nor UO_2181 (O_2181,N_24890,N_24827);
xor UO_2182 (O_2182,N_24916,N_24951);
nand UO_2183 (O_2183,N_24832,N_24812);
and UO_2184 (O_2184,N_24934,N_24904);
nor UO_2185 (O_2185,N_24860,N_24816);
nand UO_2186 (O_2186,N_24841,N_24895);
and UO_2187 (O_2187,N_24906,N_24875);
nand UO_2188 (O_2188,N_24824,N_24876);
or UO_2189 (O_2189,N_24855,N_24998);
and UO_2190 (O_2190,N_24855,N_24839);
and UO_2191 (O_2191,N_24922,N_24883);
xor UO_2192 (O_2192,N_24840,N_24833);
and UO_2193 (O_2193,N_24825,N_24974);
xnor UO_2194 (O_2194,N_24914,N_24974);
nand UO_2195 (O_2195,N_24996,N_24922);
nand UO_2196 (O_2196,N_24863,N_24940);
nand UO_2197 (O_2197,N_24845,N_24821);
xor UO_2198 (O_2198,N_24902,N_24861);
xnor UO_2199 (O_2199,N_24830,N_24995);
or UO_2200 (O_2200,N_24921,N_24971);
nor UO_2201 (O_2201,N_24845,N_24958);
nor UO_2202 (O_2202,N_24920,N_24864);
and UO_2203 (O_2203,N_24941,N_24930);
or UO_2204 (O_2204,N_24964,N_24883);
nor UO_2205 (O_2205,N_24836,N_24923);
or UO_2206 (O_2206,N_24988,N_24848);
or UO_2207 (O_2207,N_24880,N_24817);
nand UO_2208 (O_2208,N_24954,N_24958);
nor UO_2209 (O_2209,N_24975,N_24930);
or UO_2210 (O_2210,N_24833,N_24944);
nand UO_2211 (O_2211,N_24909,N_24862);
nor UO_2212 (O_2212,N_24918,N_24914);
xnor UO_2213 (O_2213,N_24894,N_24819);
nor UO_2214 (O_2214,N_24887,N_24908);
and UO_2215 (O_2215,N_24828,N_24887);
nand UO_2216 (O_2216,N_24960,N_24831);
xor UO_2217 (O_2217,N_24858,N_24895);
or UO_2218 (O_2218,N_24985,N_24905);
and UO_2219 (O_2219,N_24982,N_24970);
and UO_2220 (O_2220,N_24914,N_24926);
nor UO_2221 (O_2221,N_24855,N_24846);
xnor UO_2222 (O_2222,N_24922,N_24863);
or UO_2223 (O_2223,N_24929,N_24949);
nor UO_2224 (O_2224,N_24979,N_24986);
nor UO_2225 (O_2225,N_24863,N_24801);
xor UO_2226 (O_2226,N_24842,N_24984);
nor UO_2227 (O_2227,N_24955,N_24989);
and UO_2228 (O_2228,N_24904,N_24928);
nand UO_2229 (O_2229,N_24991,N_24892);
nand UO_2230 (O_2230,N_24984,N_24832);
and UO_2231 (O_2231,N_24951,N_24912);
nor UO_2232 (O_2232,N_24959,N_24949);
xor UO_2233 (O_2233,N_24975,N_24990);
xor UO_2234 (O_2234,N_24993,N_24838);
nor UO_2235 (O_2235,N_24855,N_24971);
nand UO_2236 (O_2236,N_24826,N_24803);
xnor UO_2237 (O_2237,N_24872,N_24854);
and UO_2238 (O_2238,N_24842,N_24957);
and UO_2239 (O_2239,N_24973,N_24881);
or UO_2240 (O_2240,N_24897,N_24853);
nand UO_2241 (O_2241,N_24822,N_24903);
xnor UO_2242 (O_2242,N_24834,N_24946);
nand UO_2243 (O_2243,N_24887,N_24857);
nand UO_2244 (O_2244,N_24856,N_24823);
nor UO_2245 (O_2245,N_24941,N_24968);
nand UO_2246 (O_2246,N_24917,N_24893);
and UO_2247 (O_2247,N_24967,N_24983);
nor UO_2248 (O_2248,N_24907,N_24811);
xnor UO_2249 (O_2249,N_24939,N_24857);
or UO_2250 (O_2250,N_24888,N_24919);
or UO_2251 (O_2251,N_24962,N_24917);
and UO_2252 (O_2252,N_24857,N_24899);
and UO_2253 (O_2253,N_24823,N_24829);
nand UO_2254 (O_2254,N_24904,N_24870);
xor UO_2255 (O_2255,N_24927,N_24879);
nand UO_2256 (O_2256,N_24963,N_24846);
or UO_2257 (O_2257,N_24867,N_24882);
xnor UO_2258 (O_2258,N_24917,N_24878);
and UO_2259 (O_2259,N_24979,N_24976);
nor UO_2260 (O_2260,N_24969,N_24977);
nor UO_2261 (O_2261,N_24820,N_24804);
nor UO_2262 (O_2262,N_24927,N_24972);
nor UO_2263 (O_2263,N_24884,N_24955);
nand UO_2264 (O_2264,N_24909,N_24801);
nand UO_2265 (O_2265,N_24803,N_24838);
nand UO_2266 (O_2266,N_24962,N_24838);
and UO_2267 (O_2267,N_24820,N_24880);
nor UO_2268 (O_2268,N_24961,N_24855);
nand UO_2269 (O_2269,N_24823,N_24841);
or UO_2270 (O_2270,N_24975,N_24856);
nand UO_2271 (O_2271,N_24934,N_24848);
xor UO_2272 (O_2272,N_24856,N_24897);
nand UO_2273 (O_2273,N_24879,N_24940);
and UO_2274 (O_2274,N_24939,N_24938);
nand UO_2275 (O_2275,N_24896,N_24936);
xor UO_2276 (O_2276,N_24932,N_24958);
nand UO_2277 (O_2277,N_24996,N_24890);
or UO_2278 (O_2278,N_24851,N_24977);
xnor UO_2279 (O_2279,N_24854,N_24804);
nand UO_2280 (O_2280,N_24867,N_24972);
and UO_2281 (O_2281,N_24924,N_24841);
and UO_2282 (O_2282,N_24936,N_24807);
nor UO_2283 (O_2283,N_24851,N_24831);
nand UO_2284 (O_2284,N_24978,N_24829);
and UO_2285 (O_2285,N_24858,N_24936);
xnor UO_2286 (O_2286,N_24887,N_24903);
xnor UO_2287 (O_2287,N_24997,N_24855);
or UO_2288 (O_2288,N_24883,N_24805);
xnor UO_2289 (O_2289,N_24936,N_24844);
or UO_2290 (O_2290,N_24868,N_24941);
nand UO_2291 (O_2291,N_24816,N_24961);
nor UO_2292 (O_2292,N_24814,N_24919);
nor UO_2293 (O_2293,N_24987,N_24967);
or UO_2294 (O_2294,N_24918,N_24917);
nand UO_2295 (O_2295,N_24970,N_24855);
and UO_2296 (O_2296,N_24852,N_24856);
xor UO_2297 (O_2297,N_24944,N_24889);
and UO_2298 (O_2298,N_24970,N_24915);
nand UO_2299 (O_2299,N_24900,N_24980);
and UO_2300 (O_2300,N_24862,N_24864);
xor UO_2301 (O_2301,N_24957,N_24871);
xor UO_2302 (O_2302,N_24844,N_24944);
or UO_2303 (O_2303,N_24825,N_24969);
or UO_2304 (O_2304,N_24994,N_24814);
nand UO_2305 (O_2305,N_24863,N_24912);
or UO_2306 (O_2306,N_24807,N_24890);
and UO_2307 (O_2307,N_24817,N_24854);
or UO_2308 (O_2308,N_24804,N_24849);
nand UO_2309 (O_2309,N_24878,N_24857);
and UO_2310 (O_2310,N_24831,N_24867);
or UO_2311 (O_2311,N_24893,N_24936);
nor UO_2312 (O_2312,N_24889,N_24878);
nand UO_2313 (O_2313,N_24915,N_24980);
nor UO_2314 (O_2314,N_24838,N_24927);
nor UO_2315 (O_2315,N_24961,N_24862);
or UO_2316 (O_2316,N_24857,N_24988);
and UO_2317 (O_2317,N_24955,N_24864);
or UO_2318 (O_2318,N_24865,N_24889);
or UO_2319 (O_2319,N_24957,N_24863);
nand UO_2320 (O_2320,N_24952,N_24883);
and UO_2321 (O_2321,N_24928,N_24956);
nand UO_2322 (O_2322,N_24843,N_24925);
xor UO_2323 (O_2323,N_24936,N_24959);
xor UO_2324 (O_2324,N_24806,N_24942);
nand UO_2325 (O_2325,N_24868,N_24846);
xnor UO_2326 (O_2326,N_24993,N_24927);
and UO_2327 (O_2327,N_24966,N_24996);
and UO_2328 (O_2328,N_24809,N_24827);
or UO_2329 (O_2329,N_24807,N_24879);
xor UO_2330 (O_2330,N_24907,N_24977);
or UO_2331 (O_2331,N_24933,N_24858);
nand UO_2332 (O_2332,N_24847,N_24968);
xor UO_2333 (O_2333,N_24925,N_24856);
nor UO_2334 (O_2334,N_24920,N_24973);
or UO_2335 (O_2335,N_24812,N_24905);
nor UO_2336 (O_2336,N_24870,N_24964);
xor UO_2337 (O_2337,N_24890,N_24929);
xnor UO_2338 (O_2338,N_24840,N_24973);
nand UO_2339 (O_2339,N_24845,N_24889);
nand UO_2340 (O_2340,N_24847,N_24972);
and UO_2341 (O_2341,N_24857,N_24889);
or UO_2342 (O_2342,N_24833,N_24860);
xor UO_2343 (O_2343,N_24804,N_24975);
nor UO_2344 (O_2344,N_24958,N_24808);
nor UO_2345 (O_2345,N_24974,N_24878);
and UO_2346 (O_2346,N_24939,N_24910);
xor UO_2347 (O_2347,N_24841,N_24966);
xnor UO_2348 (O_2348,N_24898,N_24977);
xnor UO_2349 (O_2349,N_24860,N_24839);
xor UO_2350 (O_2350,N_24824,N_24983);
or UO_2351 (O_2351,N_24888,N_24803);
nand UO_2352 (O_2352,N_24927,N_24924);
or UO_2353 (O_2353,N_24903,N_24984);
and UO_2354 (O_2354,N_24934,N_24800);
or UO_2355 (O_2355,N_24845,N_24852);
nor UO_2356 (O_2356,N_24877,N_24915);
xnor UO_2357 (O_2357,N_24941,N_24924);
or UO_2358 (O_2358,N_24996,N_24927);
and UO_2359 (O_2359,N_24945,N_24923);
or UO_2360 (O_2360,N_24906,N_24890);
xnor UO_2361 (O_2361,N_24817,N_24806);
nand UO_2362 (O_2362,N_24842,N_24886);
nor UO_2363 (O_2363,N_24846,N_24841);
and UO_2364 (O_2364,N_24893,N_24911);
xnor UO_2365 (O_2365,N_24829,N_24860);
xnor UO_2366 (O_2366,N_24930,N_24916);
nand UO_2367 (O_2367,N_24980,N_24808);
xor UO_2368 (O_2368,N_24980,N_24963);
xor UO_2369 (O_2369,N_24840,N_24867);
and UO_2370 (O_2370,N_24989,N_24968);
and UO_2371 (O_2371,N_24915,N_24945);
and UO_2372 (O_2372,N_24838,N_24875);
nand UO_2373 (O_2373,N_24823,N_24835);
nor UO_2374 (O_2374,N_24988,N_24951);
or UO_2375 (O_2375,N_24815,N_24992);
or UO_2376 (O_2376,N_24853,N_24935);
xor UO_2377 (O_2377,N_24886,N_24941);
and UO_2378 (O_2378,N_24960,N_24951);
nand UO_2379 (O_2379,N_24836,N_24890);
and UO_2380 (O_2380,N_24934,N_24952);
nor UO_2381 (O_2381,N_24866,N_24884);
or UO_2382 (O_2382,N_24969,N_24877);
or UO_2383 (O_2383,N_24800,N_24802);
nand UO_2384 (O_2384,N_24846,N_24905);
xor UO_2385 (O_2385,N_24869,N_24847);
and UO_2386 (O_2386,N_24830,N_24856);
xnor UO_2387 (O_2387,N_24916,N_24928);
or UO_2388 (O_2388,N_24831,N_24964);
nor UO_2389 (O_2389,N_24881,N_24902);
or UO_2390 (O_2390,N_24944,N_24900);
nand UO_2391 (O_2391,N_24840,N_24896);
nand UO_2392 (O_2392,N_24875,N_24889);
nor UO_2393 (O_2393,N_24946,N_24802);
xor UO_2394 (O_2394,N_24958,N_24890);
or UO_2395 (O_2395,N_24829,N_24953);
nor UO_2396 (O_2396,N_24939,N_24866);
nand UO_2397 (O_2397,N_24942,N_24936);
nand UO_2398 (O_2398,N_24973,N_24882);
or UO_2399 (O_2399,N_24882,N_24861);
nor UO_2400 (O_2400,N_24891,N_24804);
xor UO_2401 (O_2401,N_24908,N_24889);
nor UO_2402 (O_2402,N_24990,N_24847);
or UO_2403 (O_2403,N_24861,N_24862);
xnor UO_2404 (O_2404,N_24863,N_24854);
xor UO_2405 (O_2405,N_24895,N_24890);
nor UO_2406 (O_2406,N_24936,N_24953);
nor UO_2407 (O_2407,N_24867,N_24800);
xnor UO_2408 (O_2408,N_24855,N_24834);
xnor UO_2409 (O_2409,N_24881,N_24822);
xor UO_2410 (O_2410,N_24884,N_24823);
xor UO_2411 (O_2411,N_24935,N_24854);
or UO_2412 (O_2412,N_24810,N_24828);
xnor UO_2413 (O_2413,N_24942,N_24971);
nor UO_2414 (O_2414,N_24978,N_24977);
or UO_2415 (O_2415,N_24842,N_24807);
xor UO_2416 (O_2416,N_24819,N_24929);
or UO_2417 (O_2417,N_24810,N_24905);
or UO_2418 (O_2418,N_24815,N_24952);
nand UO_2419 (O_2419,N_24921,N_24976);
nand UO_2420 (O_2420,N_24881,N_24897);
nand UO_2421 (O_2421,N_24958,N_24816);
or UO_2422 (O_2422,N_24976,N_24927);
or UO_2423 (O_2423,N_24946,N_24847);
nor UO_2424 (O_2424,N_24972,N_24918);
or UO_2425 (O_2425,N_24908,N_24916);
nand UO_2426 (O_2426,N_24968,N_24973);
and UO_2427 (O_2427,N_24839,N_24816);
or UO_2428 (O_2428,N_24829,N_24968);
and UO_2429 (O_2429,N_24917,N_24932);
and UO_2430 (O_2430,N_24827,N_24953);
or UO_2431 (O_2431,N_24934,N_24912);
nand UO_2432 (O_2432,N_24837,N_24926);
and UO_2433 (O_2433,N_24913,N_24830);
xnor UO_2434 (O_2434,N_24876,N_24881);
nor UO_2435 (O_2435,N_24953,N_24985);
xnor UO_2436 (O_2436,N_24813,N_24881);
nand UO_2437 (O_2437,N_24906,N_24896);
and UO_2438 (O_2438,N_24821,N_24806);
and UO_2439 (O_2439,N_24986,N_24913);
xor UO_2440 (O_2440,N_24943,N_24940);
nand UO_2441 (O_2441,N_24999,N_24801);
nand UO_2442 (O_2442,N_24883,N_24953);
nor UO_2443 (O_2443,N_24811,N_24930);
nand UO_2444 (O_2444,N_24943,N_24914);
or UO_2445 (O_2445,N_24867,N_24854);
nand UO_2446 (O_2446,N_24964,N_24954);
and UO_2447 (O_2447,N_24897,N_24918);
and UO_2448 (O_2448,N_24926,N_24949);
nor UO_2449 (O_2449,N_24861,N_24950);
or UO_2450 (O_2450,N_24812,N_24824);
xor UO_2451 (O_2451,N_24930,N_24907);
xor UO_2452 (O_2452,N_24906,N_24807);
xnor UO_2453 (O_2453,N_24811,N_24923);
nor UO_2454 (O_2454,N_24950,N_24903);
and UO_2455 (O_2455,N_24808,N_24937);
xnor UO_2456 (O_2456,N_24920,N_24946);
nor UO_2457 (O_2457,N_24978,N_24819);
and UO_2458 (O_2458,N_24948,N_24856);
nor UO_2459 (O_2459,N_24867,N_24844);
or UO_2460 (O_2460,N_24892,N_24831);
nand UO_2461 (O_2461,N_24816,N_24859);
or UO_2462 (O_2462,N_24834,N_24856);
nand UO_2463 (O_2463,N_24952,N_24880);
xor UO_2464 (O_2464,N_24866,N_24908);
xor UO_2465 (O_2465,N_24886,N_24808);
nand UO_2466 (O_2466,N_24837,N_24916);
and UO_2467 (O_2467,N_24882,N_24978);
xnor UO_2468 (O_2468,N_24965,N_24982);
or UO_2469 (O_2469,N_24947,N_24834);
nand UO_2470 (O_2470,N_24861,N_24991);
nor UO_2471 (O_2471,N_24939,N_24858);
nand UO_2472 (O_2472,N_24851,N_24978);
or UO_2473 (O_2473,N_24939,N_24990);
xor UO_2474 (O_2474,N_24835,N_24840);
xnor UO_2475 (O_2475,N_24846,N_24932);
nor UO_2476 (O_2476,N_24977,N_24975);
xnor UO_2477 (O_2477,N_24977,N_24850);
nand UO_2478 (O_2478,N_24862,N_24953);
and UO_2479 (O_2479,N_24821,N_24895);
nand UO_2480 (O_2480,N_24978,N_24878);
nand UO_2481 (O_2481,N_24854,N_24909);
xnor UO_2482 (O_2482,N_24943,N_24803);
and UO_2483 (O_2483,N_24870,N_24915);
nor UO_2484 (O_2484,N_24818,N_24885);
nor UO_2485 (O_2485,N_24958,N_24814);
nand UO_2486 (O_2486,N_24915,N_24866);
and UO_2487 (O_2487,N_24861,N_24956);
nor UO_2488 (O_2488,N_24890,N_24924);
or UO_2489 (O_2489,N_24887,N_24940);
nor UO_2490 (O_2490,N_24927,N_24864);
or UO_2491 (O_2491,N_24923,N_24947);
xor UO_2492 (O_2492,N_24883,N_24915);
xnor UO_2493 (O_2493,N_24866,N_24822);
nand UO_2494 (O_2494,N_24943,N_24813);
nor UO_2495 (O_2495,N_24975,N_24864);
or UO_2496 (O_2496,N_24863,N_24917);
nor UO_2497 (O_2497,N_24823,N_24842);
and UO_2498 (O_2498,N_24874,N_24939);
or UO_2499 (O_2499,N_24934,N_24963);
nand UO_2500 (O_2500,N_24845,N_24838);
nand UO_2501 (O_2501,N_24814,N_24877);
and UO_2502 (O_2502,N_24826,N_24816);
or UO_2503 (O_2503,N_24842,N_24909);
and UO_2504 (O_2504,N_24945,N_24972);
nor UO_2505 (O_2505,N_24891,N_24950);
xor UO_2506 (O_2506,N_24916,N_24987);
xnor UO_2507 (O_2507,N_24807,N_24853);
or UO_2508 (O_2508,N_24893,N_24828);
or UO_2509 (O_2509,N_24814,N_24893);
and UO_2510 (O_2510,N_24898,N_24855);
nor UO_2511 (O_2511,N_24997,N_24903);
nand UO_2512 (O_2512,N_24934,N_24968);
xor UO_2513 (O_2513,N_24812,N_24922);
and UO_2514 (O_2514,N_24975,N_24878);
or UO_2515 (O_2515,N_24978,N_24992);
or UO_2516 (O_2516,N_24968,N_24800);
xor UO_2517 (O_2517,N_24895,N_24927);
nand UO_2518 (O_2518,N_24852,N_24956);
and UO_2519 (O_2519,N_24916,N_24909);
nand UO_2520 (O_2520,N_24903,N_24941);
and UO_2521 (O_2521,N_24825,N_24832);
and UO_2522 (O_2522,N_24813,N_24996);
nand UO_2523 (O_2523,N_24986,N_24912);
and UO_2524 (O_2524,N_24993,N_24820);
and UO_2525 (O_2525,N_24835,N_24939);
nor UO_2526 (O_2526,N_24958,N_24850);
and UO_2527 (O_2527,N_24992,N_24965);
nor UO_2528 (O_2528,N_24967,N_24925);
and UO_2529 (O_2529,N_24947,N_24918);
xnor UO_2530 (O_2530,N_24911,N_24998);
nor UO_2531 (O_2531,N_24844,N_24861);
and UO_2532 (O_2532,N_24951,N_24975);
xnor UO_2533 (O_2533,N_24985,N_24909);
nand UO_2534 (O_2534,N_24831,N_24861);
xor UO_2535 (O_2535,N_24849,N_24983);
nor UO_2536 (O_2536,N_24948,N_24850);
and UO_2537 (O_2537,N_24841,N_24972);
xor UO_2538 (O_2538,N_24931,N_24930);
and UO_2539 (O_2539,N_24916,N_24999);
or UO_2540 (O_2540,N_24910,N_24809);
nor UO_2541 (O_2541,N_24992,N_24848);
nor UO_2542 (O_2542,N_24838,N_24897);
xnor UO_2543 (O_2543,N_24912,N_24873);
nor UO_2544 (O_2544,N_24994,N_24802);
nor UO_2545 (O_2545,N_24832,N_24959);
xnor UO_2546 (O_2546,N_24991,N_24976);
nor UO_2547 (O_2547,N_24821,N_24923);
or UO_2548 (O_2548,N_24895,N_24906);
or UO_2549 (O_2549,N_24987,N_24826);
nand UO_2550 (O_2550,N_24891,N_24855);
or UO_2551 (O_2551,N_24983,N_24803);
nand UO_2552 (O_2552,N_24863,N_24954);
and UO_2553 (O_2553,N_24830,N_24914);
or UO_2554 (O_2554,N_24993,N_24845);
and UO_2555 (O_2555,N_24855,N_24859);
or UO_2556 (O_2556,N_24875,N_24847);
xor UO_2557 (O_2557,N_24891,N_24837);
nand UO_2558 (O_2558,N_24963,N_24836);
xnor UO_2559 (O_2559,N_24985,N_24894);
xor UO_2560 (O_2560,N_24909,N_24904);
nor UO_2561 (O_2561,N_24981,N_24845);
nor UO_2562 (O_2562,N_24996,N_24806);
xnor UO_2563 (O_2563,N_24802,N_24909);
or UO_2564 (O_2564,N_24929,N_24885);
nor UO_2565 (O_2565,N_24887,N_24910);
nand UO_2566 (O_2566,N_24999,N_24891);
and UO_2567 (O_2567,N_24834,N_24835);
xnor UO_2568 (O_2568,N_24995,N_24941);
and UO_2569 (O_2569,N_24977,N_24836);
nor UO_2570 (O_2570,N_24832,N_24905);
nor UO_2571 (O_2571,N_24821,N_24993);
nor UO_2572 (O_2572,N_24878,N_24962);
and UO_2573 (O_2573,N_24929,N_24905);
or UO_2574 (O_2574,N_24988,N_24968);
and UO_2575 (O_2575,N_24987,N_24991);
nand UO_2576 (O_2576,N_24833,N_24987);
nor UO_2577 (O_2577,N_24965,N_24975);
or UO_2578 (O_2578,N_24936,N_24982);
nand UO_2579 (O_2579,N_24843,N_24836);
xor UO_2580 (O_2580,N_24945,N_24900);
xnor UO_2581 (O_2581,N_24877,N_24861);
or UO_2582 (O_2582,N_24999,N_24938);
and UO_2583 (O_2583,N_24844,N_24926);
nor UO_2584 (O_2584,N_24938,N_24942);
nand UO_2585 (O_2585,N_24898,N_24897);
nor UO_2586 (O_2586,N_24947,N_24905);
or UO_2587 (O_2587,N_24825,N_24887);
and UO_2588 (O_2588,N_24935,N_24870);
nand UO_2589 (O_2589,N_24997,N_24869);
nand UO_2590 (O_2590,N_24870,N_24976);
nor UO_2591 (O_2591,N_24868,N_24820);
nor UO_2592 (O_2592,N_24922,N_24869);
or UO_2593 (O_2593,N_24838,N_24909);
xor UO_2594 (O_2594,N_24938,N_24967);
nor UO_2595 (O_2595,N_24805,N_24911);
xnor UO_2596 (O_2596,N_24930,N_24982);
or UO_2597 (O_2597,N_24941,N_24958);
and UO_2598 (O_2598,N_24869,N_24930);
or UO_2599 (O_2599,N_24887,N_24935);
and UO_2600 (O_2600,N_24878,N_24803);
xnor UO_2601 (O_2601,N_24813,N_24806);
xor UO_2602 (O_2602,N_24947,N_24864);
xnor UO_2603 (O_2603,N_24921,N_24919);
nor UO_2604 (O_2604,N_24901,N_24813);
nor UO_2605 (O_2605,N_24917,N_24952);
or UO_2606 (O_2606,N_24816,N_24834);
nor UO_2607 (O_2607,N_24839,N_24904);
xnor UO_2608 (O_2608,N_24854,N_24813);
nor UO_2609 (O_2609,N_24983,N_24960);
or UO_2610 (O_2610,N_24813,N_24839);
nand UO_2611 (O_2611,N_24840,N_24967);
and UO_2612 (O_2612,N_24830,N_24924);
or UO_2613 (O_2613,N_24991,N_24939);
nand UO_2614 (O_2614,N_24948,N_24999);
nor UO_2615 (O_2615,N_24858,N_24909);
or UO_2616 (O_2616,N_24937,N_24827);
xor UO_2617 (O_2617,N_24880,N_24871);
or UO_2618 (O_2618,N_24842,N_24891);
and UO_2619 (O_2619,N_24973,N_24979);
xor UO_2620 (O_2620,N_24876,N_24865);
nand UO_2621 (O_2621,N_24969,N_24884);
xor UO_2622 (O_2622,N_24913,N_24803);
and UO_2623 (O_2623,N_24893,N_24891);
nand UO_2624 (O_2624,N_24981,N_24997);
nand UO_2625 (O_2625,N_24883,N_24865);
and UO_2626 (O_2626,N_24979,N_24849);
nor UO_2627 (O_2627,N_24847,N_24828);
and UO_2628 (O_2628,N_24919,N_24935);
nor UO_2629 (O_2629,N_24900,N_24802);
nor UO_2630 (O_2630,N_24810,N_24815);
xnor UO_2631 (O_2631,N_24802,N_24822);
nand UO_2632 (O_2632,N_24923,N_24905);
and UO_2633 (O_2633,N_24941,N_24961);
and UO_2634 (O_2634,N_24940,N_24955);
nor UO_2635 (O_2635,N_24819,N_24809);
and UO_2636 (O_2636,N_24887,N_24912);
xor UO_2637 (O_2637,N_24846,N_24858);
and UO_2638 (O_2638,N_24841,N_24804);
xnor UO_2639 (O_2639,N_24891,N_24996);
xor UO_2640 (O_2640,N_24834,N_24954);
nor UO_2641 (O_2641,N_24999,N_24871);
or UO_2642 (O_2642,N_24907,N_24955);
xor UO_2643 (O_2643,N_24873,N_24827);
nor UO_2644 (O_2644,N_24999,N_24843);
nand UO_2645 (O_2645,N_24940,N_24982);
or UO_2646 (O_2646,N_24972,N_24938);
nand UO_2647 (O_2647,N_24872,N_24888);
or UO_2648 (O_2648,N_24862,N_24887);
xnor UO_2649 (O_2649,N_24981,N_24890);
xnor UO_2650 (O_2650,N_24887,N_24882);
and UO_2651 (O_2651,N_24940,N_24854);
nor UO_2652 (O_2652,N_24918,N_24903);
xnor UO_2653 (O_2653,N_24957,N_24911);
xor UO_2654 (O_2654,N_24944,N_24913);
xor UO_2655 (O_2655,N_24804,N_24972);
and UO_2656 (O_2656,N_24800,N_24987);
xnor UO_2657 (O_2657,N_24838,N_24974);
or UO_2658 (O_2658,N_24876,N_24968);
nor UO_2659 (O_2659,N_24905,N_24880);
or UO_2660 (O_2660,N_24811,N_24816);
nand UO_2661 (O_2661,N_24996,N_24871);
xnor UO_2662 (O_2662,N_24996,N_24856);
and UO_2663 (O_2663,N_24869,N_24801);
nor UO_2664 (O_2664,N_24852,N_24830);
or UO_2665 (O_2665,N_24899,N_24841);
and UO_2666 (O_2666,N_24963,N_24994);
or UO_2667 (O_2667,N_24872,N_24889);
and UO_2668 (O_2668,N_24846,N_24845);
or UO_2669 (O_2669,N_24888,N_24947);
and UO_2670 (O_2670,N_24983,N_24892);
nand UO_2671 (O_2671,N_24802,N_24851);
nand UO_2672 (O_2672,N_24972,N_24948);
xor UO_2673 (O_2673,N_24908,N_24993);
or UO_2674 (O_2674,N_24811,N_24997);
xor UO_2675 (O_2675,N_24953,N_24879);
xnor UO_2676 (O_2676,N_24966,N_24883);
and UO_2677 (O_2677,N_24823,N_24836);
and UO_2678 (O_2678,N_24812,N_24851);
nand UO_2679 (O_2679,N_24898,N_24980);
nor UO_2680 (O_2680,N_24861,N_24802);
nor UO_2681 (O_2681,N_24839,N_24890);
or UO_2682 (O_2682,N_24980,N_24950);
nand UO_2683 (O_2683,N_24802,N_24866);
or UO_2684 (O_2684,N_24977,N_24841);
nand UO_2685 (O_2685,N_24862,N_24987);
nor UO_2686 (O_2686,N_24867,N_24826);
nor UO_2687 (O_2687,N_24824,N_24884);
or UO_2688 (O_2688,N_24833,N_24904);
and UO_2689 (O_2689,N_24979,N_24811);
xor UO_2690 (O_2690,N_24946,N_24813);
or UO_2691 (O_2691,N_24992,N_24913);
or UO_2692 (O_2692,N_24847,N_24834);
or UO_2693 (O_2693,N_24862,N_24994);
xor UO_2694 (O_2694,N_24883,N_24974);
nor UO_2695 (O_2695,N_24862,N_24817);
xnor UO_2696 (O_2696,N_24911,N_24944);
nand UO_2697 (O_2697,N_24814,N_24991);
or UO_2698 (O_2698,N_24885,N_24844);
nand UO_2699 (O_2699,N_24824,N_24856);
nor UO_2700 (O_2700,N_24965,N_24826);
and UO_2701 (O_2701,N_24871,N_24995);
nand UO_2702 (O_2702,N_24971,N_24917);
and UO_2703 (O_2703,N_24805,N_24998);
nor UO_2704 (O_2704,N_24876,N_24964);
nand UO_2705 (O_2705,N_24817,N_24973);
and UO_2706 (O_2706,N_24930,N_24969);
and UO_2707 (O_2707,N_24985,N_24815);
nand UO_2708 (O_2708,N_24924,N_24803);
xnor UO_2709 (O_2709,N_24825,N_24831);
and UO_2710 (O_2710,N_24955,N_24836);
and UO_2711 (O_2711,N_24843,N_24903);
and UO_2712 (O_2712,N_24894,N_24978);
or UO_2713 (O_2713,N_24925,N_24904);
and UO_2714 (O_2714,N_24935,N_24862);
nor UO_2715 (O_2715,N_24996,N_24917);
nand UO_2716 (O_2716,N_24866,N_24929);
nor UO_2717 (O_2717,N_24896,N_24955);
or UO_2718 (O_2718,N_24849,N_24835);
or UO_2719 (O_2719,N_24921,N_24826);
or UO_2720 (O_2720,N_24909,N_24941);
and UO_2721 (O_2721,N_24969,N_24938);
nor UO_2722 (O_2722,N_24811,N_24951);
nor UO_2723 (O_2723,N_24937,N_24816);
nor UO_2724 (O_2724,N_24893,N_24826);
xnor UO_2725 (O_2725,N_24974,N_24889);
and UO_2726 (O_2726,N_24812,N_24820);
xnor UO_2727 (O_2727,N_24810,N_24850);
nor UO_2728 (O_2728,N_24843,N_24996);
nor UO_2729 (O_2729,N_24945,N_24912);
xor UO_2730 (O_2730,N_24831,N_24833);
nand UO_2731 (O_2731,N_24955,N_24949);
or UO_2732 (O_2732,N_24933,N_24995);
nor UO_2733 (O_2733,N_24884,N_24930);
and UO_2734 (O_2734,N_24852,N_24846);
nor UO_2735 (O_2735,N_24802,N_24801);
nand UO_2736 (O_2736,N_24854,N_24843);
nand UO_2737 (O_2737,N_24815,N_24855);
and UO_2738 (O_2738,N_24844,N_24804);
xor UO_2739 (O_2739,N_24883,N_24997);
and UO_2740 (O_2740,N_24895,N_24851);
nand UO_2741 (O_2741,N_24929,N_24940);
or UO_2742 (O_2742,N_24815,N_24957);
and UO_2743 (O_2743,N_24954,N_24888);
nor UO_2744 (O_2744,N_24802,N_24922);
and UO_2745 (O_2745,N_24907,N_24802);
nand UO_2746 (O_2746,N_24909,N_24926);
or UO_2747 (O_2747,N_24898,N_24955);
nor UO_2748 (O_2748,N_24905,N_24855);
nor UO_2749 (O_2749,N_24941,N_24829);
xnor UO_2750 (O_2750,N_24813,N_24811);
nor UO_2751 (O_2751,N_24933,N_24956);
nand UO_2752 (O_2752,N_24850,N_24962);
nor UO_2753 (O_2753,N_24935,N_24849);
or UO_2754 (O_2754,N_24996,N_24956);
xor UO_2755 (O_2755,N_24811,N_24981);
and UO_2756 (O_2756,N_24931,N_24969);
nor UO_2757 (O_2757,N_24978,N_24887);
xnor UO_2758 (O_2758,N_24916,N_24811);
nor UO_2759 (O_2759,N_24800,N_24948);
or UO_2760 (O_2760,N_24981,N_24975);
xnor UO_2761 (O_2761,N_24820,N_24973);
and UO_2762 (O_2762,N_24921,N_24926);
xor UO_2763 (O_2763,N_24968,N_24930);
or UO_2764 (O_2764,N_24824,N_24917);
nand UO_2765 (O_2765,N_24863,N_24919);
nand UO_2766 (O_2766,N_24838,N_24885);
nor UO_2767 (O_2767,N_24945,N_24863);
or UO_2768 (O_2768,N_24816,N_24832);
or UO_2769 (O_2769,N_24904,N_24851);
nand UO_2770 (O_2770,N_24937,N_24904);
nand UO_2771 (O_2771,N_24835,N_24816);
nor UO_2772 (O_2772,N_24817,N_24822);
nand UO_2773 (O_2773,N_24941,N_24937);
nor UO_2774 (O_2774,N_24991,N_24836);
and UO_2775 (O_2775,N_24936,N_24825);
nor UO_2776 (O_2776,N_24817,N_24876);
or UO_2777 (O_2777,N_24898,N_24938);
nor UO_2778 (O_2778,N_24939,N_24958);
nand UO_2779 (O_2779,N_24991,N_24944);
and UO_2780 (O_2780,N_24972,N_24958);
and UO_2781 (O_2781,N_24907,N_24837);
nor UO_2782 (O_2782,N_24978,N_24976);
and UO_2783 (O_2783,N_24983,N_24830);
nor UO_2784 (O_2784,N_24855,N_24851);
nand UO_2785 (O_2785,N_24834,N_24879);
nor UO_2786 (O_2786,N_24845,N_24939);
nand UO_2787 (O_2787,N_24853,N_24801);
xnor UO_2788 (O_2788,N_24891,N_24803);
or UO_2789 (O_2789,N_24986,N_24905);
xnor UO_2790 (O_2790,N_24937,N_24964);
nor UO_2791 (O_2791,N_24960,N_24896);
nand UO_2792 (O_2792,N_24984,N_24875);
xnor UO_2793 (O_2793,N_24982,N_24987);
nor UO_2794 (O_2794,N_24970,N_24949);
xor UO_2795 (O_2795,N_24960,N_24957);
nor UO_2796 (O_2796,N_24863,N_24834);
or UO_2797 (O_2797,N_24900,N_24968);
or UO_2798 (O_2798,N_24941,N_24893);
xnor UO_2799 (O_2799,N_24981,N_24854);
nand UO_2800 (O_2800,N_24832,N_24915);
or UO_2801 (O_2801,N_24992,N_24916);
nand UO_2802 (O_2802,N_24843,N_24814);
nand UO_2803 (O_2803,N_24875,N_24988);
nor UO_2804 (O_2804,N_24892,N_24962);
and UO_2805 (O_2805,N_24918,N_24846);
xnor UO_2806 (O_2806,N_24978,N_24847);
nand UO_2807 (O_2807,N_24903,N_24998);
nand UO_2808 (O_2808,N_24877,N_24902);
nor UO_2809 (O_2809,N_24810,N_24941);
or UO_2810 (O_2810,N_24900,N_24964);
and UO_2811 (O_2811,N_24989,N_24921);
or UO_2812 (O_2812,N_24967,N_24993);
and UO_2813 (O_2813,N_24835,N_24846);
xnor UO_2814 (O_2814,N_24837,N_24847);
or UO_2815 (O_2815,N_24853,N_24905);
or UO_2816 (O_2816,N_24959,N_24952);
xnor UO_2817 (O_2817,N_24913,N_24879);
or UO_2818 (O_2818,N_24921,N_24930);
or UO_2819 (O_2819,N_24912,N_24859);
nor UO_2820 (O_2820,N_24854,N_24949);
nand UO_2821 (O_2821,N_24914,N_24906);
nand UO_2822 (O_2822,N_24970,N_24980);
and UO_2823 (O_2823,N_24897,N_24823);
and UO_2824 (O_2824,N_24881,N_24989);
nor UO_2825 (O_2825,N_24948,N_24906);
and UO_2826 (O_2826,N_24919,N_24817);
or UO_2827 (O_2827,N_24934,N_24929);
nand UO_2828 (O_2828,N_24837,N_24860);
and UO_2829 (O_2829,N_24812,N_24864);
nor UO_2830 (O_2830,N_24982,N_24995);
and UO_2831 (O_2831,N_24890,N_24896);
nand UO_2832 (O_2832,N_24946,N_24882);
xor UO_2833 (O_2833,N_24836,N_24979);
nand UO_2834 (O_2834,N_24845,N_24833);
xnor UO_2835 (O_2835,N_24893,N_24866);
nand UO_2836 (O_2836,N_24938,N_24977);
and UO_2837 (O_2837,N_24854,N_24938);
nand UO_2838 (O_2838,N_24894,N_24837);
nor UO_2839 (O_2839,N_24931,N_24936);
and UO_2840 (O_2840,N_24957,N_24996);
and UO_2841 (O_2841,N_24932,N_24851);
or UO_2842 (O_2842,N_24827,N_24999);
nor UO_2843 (O_2843,N_24917,N_24848);
xnor UO_2844 (O_2844,N_24956,N_24897);
or UO_2845 (O_2845,N_24904,N_24889);
nand UO_2846 (O_2846,N_24886,N_24916);
and UO_2847 (O_2847,N_24987,N_24889);
xor UO_2848 (O_2848,N_24832,N_24967);
or UO_2849 (O_2849,N_24955,N_24847);
nand UO_2850 (O_2850,N_24825,N_24906);
and UO_2851 (O_2851,N_24845,N_24858);
or UO_2852 (O_2852,N_24824,N_24962);
xnor UO_2853 (O_2853,N_24985,N_24865);
xor UO_2854 (O_2854,N_24896,N_24884);
and UO_2855 (O_2855,N_24922,N_24989);
nand UO_2856 (O_2856,N_24913,N_24968);
and UO_2857 (O_2857,N_24992,N_24911);
nand UO_2858 (O_2858,N_24961,N_24899);
and UO_2859 (O_2859,N_24963,N_24979);
nor UO_2860 (O_2860,N_24964,N_24884);
and UO_2861 (O_2861,N_24888,N_24964);
nor UO_2862 (O_2862,N_24862,N_24950);
xor UO_2863 (O_2863,N_24886,N_24806);
or UO_2864 (O_2864,N_24931,N_24916);
or UO_2865 (O_2865,N_24857,N_24935);
and UO_2866 (O_2866,N_24932,N_24809);
or UO_2867 (O_2867,N_24896,N_24815);
and UO_2868 (O_2868,N_24969,N_24883);
nor UO_2869 (O_2869,N_24882,N_24996);
nand UO_2870 (O_2870,N_24964,N_24873);
and UO_2871 (O_2871,N_24880,N_24895);
and UO_2872 (O_2872,N_24914,N_24899);
nand UO_2873 (O_2873,N_24927,N_24910);
nor UO_2874 (O_2874,N_24843,N_24880);
or UO_2875 (O_2875,N_24984,N_24980);
nor UO_2876 (O_2876,N_24840,N_24856);
or UO_2877 (O_2877,N_24824,N_24851);
xor UO_2878 (O_2878,N_24873,N_24914);
nand UO_2879 (O_2879,N_24827,N_24900);
or UO_2880 (O_2880,N_24896,N_24954);
and UO_2881 (O_2881,N_24892,N_24866);
nor UO_2882 (O_2882,N_24808,N_24859);
xor UO_2883 (O_2883,N_24939,N_24901);
or UO_2884 (O_2884,N_24977,N_24979);
or UO_2885 (O_2885,N_24824,N_24991);
nor UO_2886 (O_2886,N_24817,N_24884);
nor UO_2887 (O_2887,N_24972,N_24978);
xnor UO_2888 (O_2888,N_24891,N_24802);
nor UO_2889 (O_2889,N_24990,N_24801);
or UO_2890 (O_2890,N_24865,N_24880);
nor UO_2891 (O_2891,N_24854,N_24921);
nor UO_2892 (O_2892,N_24850,N_24873);
or UO_2893 (O_2893,N_24864,N_24845);
xnor UO_2894 (O_2894,N_24987,N_24808);
nand UO_2895 (O_2895,N_24949,N_24919);
and UO_2896 (O_2896,N_24844,N_24941);
or UO_2897 (O_2897,N_24945,N_24917);
nand UO_2898 (O_2898,N_24965,N_24951);
nand UO_2899 (O_2899,N_24814,N_24828);
and UO_2900 (O_2900,N_24937,N_24916);
and UO_2901 (O_2901,N_24962,N_24998);
or UO_2902 (O_2902,N_24889,N_24929);
nor UO_2903 (O_2903,N_24864,N_24963);
nor UO_2904 (O_2904,N_24993,N_24856);
nor UO_2905 (O_2905,N_24855,N_24895);
nand UO_2906 (O_2906,N_24905,N_24977);
nand UO_2907 (O_2907,N_24875,N_24898);
nand UO_2908 (O_2908,N_24868,N_24928);
nor UO_2909 (O_2909,N_24950,N_24819);
and UO_2910 (O_2910,N_24925,N_24894);
xnor UO_2911 (O_2911,N_24961,N_24960);
and UO_2912 (O_2912,N_24923,N_24834);
nor UO_2913 (O_2913,N_24835,N_24833);
and UO_2914 (O_2914,N_24934,N_24845);
nor UO_2915 (O_2915,N_24945,N_24894);
nand UO_2916 (O_2916,N_24808,N_24848);
or UO_2917 (O_2917,N_24991,N_24978);
xnor UO_2918 (O_2918,N_24886,N_24837);
nand UO_2919 (O_2919,N_24980,N_24877);
or UO_2920 (O_2920,N_24893,N_24973);
nor UO_2921 (O_2921,N_24885,N_24845);
nor UO_2922 (O_2922,N_24929,N_24874);
xor UO_2923 (O_2923,N_24913,N_24877);
or UO_2924 (O_2924,N_24904,N_24945);
xor UO_2925 (O_2925,N_24801,N_24874);
and UO_2926 (O_2926,N_24932,N_24927);
xor UO_2927 (O_2927,N_24831,N_24986);
nand UO_2928 (O_2928,N_24888,N_24810);
nand UO_2929 (O_2929,N_24816,N_24930);
nand UO_2930 (O_2930,N_24867,N_24802);
and UO_2931 (O_2931,N_24981,N_24979);
or UO_2932 (O_2932,N_24949,N_24889);
nor UO_2933 (O_2933,N_24805,N_24904);
xnor UO_2934 (O_2934,N_24827,N_24927);
or UO_2935 (O_2935,N_24964,N_24829);
nand UO_2936 (O_2936,N_24867,N_24926);
xnor UO_2937 (O_2937,N_24934,N_24961);
xnor UO_2938 (O_2938,N_24820,N_24944);
and UO_2939 (O_2939,N_24988,N_24976);
nand UO_2940 (O_2940,N_24960,N_24921);
nor UO_2941 (O_2941,N_24917,N_24809);
nand UO_2942 (O_2942,N_24978,N_24811);
or UO_2943 (O_2943,N_24982,N_24997);
nor UO_2944 (O_2944,N_24803,N_24863);
or UO_2945 (O_2945,N_24900,N_24959);
xnor UO_2946 (O_2946,N_24948,N_24853);
nand UO_2947 (O_2947,N_24885,N_24891);
xor UO_2948 (O_2948,N_24812,N_24848);
or UO_2949 (O_2949,N_24880,N_24837);
nor UO_2950 (O_2950,N_24806,N_24953);
and UO_2951 (O_2951,N_24962,N_24942);
xnor UO_2952 (O_2952,N_24911,N_24827);
nor UO_2953 (O_2953,N_24802,N_24827);
xor UO_2954 (O_2954,N_24879,N_24899);
xnor UO_2955 (O_2955,N_24974,N_24851);
and UO_2956 (O_2956,N_24886,N_24802);
xnor UO_2957 (O_2957,N_24973,N_24868);
nand UO_2958 (O_2958,N_24837,N_24855);
xor UO_2959 (O_2959,N_24875,N_24839);
xnor UO_2960 (O_2960,N_24858,N_24924);
and UO_2961 (O_2961,N_24866,N_24992);
xnor UO_2962 (O_2962,N_24924,N_24918);
or UO_2963 (O_2963,N_24989,N_24834);
nand UO_2964 (O_2964,N_24810,N_24876);
and UO_2965 (O_2965,N_24917,N_24927);
nor UO_2966 (O_2966,N_24815,N_24853);
and UO_2967 (O_2967,N_24881,N_24946);
xor UO_2968 (O_2968,N_24980,N_24837);
and UO_2969 (O_2969,N_24924,N_24894);
xor UO_2970 (O_2970,N_24892,N_24842);
or UO_2971 (O_2971,N_24998,N_24803);
nand UO_2972 (O_2972,N_24808,N_24861);
xor UO_2973 (O_2973,N_24915,N_24923);
or UO_2974 (O_2974,N_24946,N_24999);
nand UO_2975 (O_2975,N_24920,N_24949);
xnor UO_2976 (O_2976,N_24967,N_24805);
and UO_2977 (O_2977,N_24907,N_24950);
or UO_2978 (O_2978,N_24980,N_24883);
and UO_2979 (O_2979,N_24889,N_24829);
or UO_2980 (O_2980,N_24869,N_24945);
or UO_2981 (O_2981,N_24815,N_24883);
xor UO_2982 (O_2982,N_24930,N_24977);
nand UO_2983 (O_2983,N_24966,N_24958);
or UO_2984 (O_2984,N_24983,N_24862);
and UO_2985 (O_2985,N_24812,N_24825);
nor UO_2986 (O_2986,N_24815,N_24812);
and UO_2987 (O_2987,N_24899,N_24800);
xor UO_2988 (O_2988,N_24949,N_24858);
or UO_2989 (O_2989,N_24877,N_24920);
or UO_2990 (O_2990,N_24993,N_24886);
xor UO_2991 (O_2991,N_24818,N_24826);
nand UO_2992 (O_2992,N_24985,N_24984);
or UO_2993 (O_2993,N_24935,N_24932);
and UO_2994 (O_2994,N_24860,N_24932);
nand UO_2995 (O_2995,N_24950,N_24954);
xor UO_2996 (O_2996,N_24988,N_24862);
and UO_2997 (O_2997,N_24989,N_24980);
nand UO_2998 (O_2998,N_24940,N_24814);
nand UO_2999 (O_2999,N_24901,N_24945);
endmodule