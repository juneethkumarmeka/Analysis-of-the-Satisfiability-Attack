module basic_1000_10000_1500_4_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_934,In_437);
xor U1 (N_1,In_570,In_92);
or U2 (N_2,In_891,In_396);
nor U3 (N_3,In_988,In_864);
xor U4 (N_4,In_556,In_498);
nand U5 (N_5,In_381,In_832);
or U6 (N_6,In_523,In_945);
nand U7 (N_7,In_179,In_0);
and U8 (N_8,In_554,In_350);
and U9 (N_9,In_526,In_339);
and U10 (N_10,In_737,In_641);
and U11 (N_11,In_302,In_297);
nor U12 (N_12,In_427,In_163);
and U13 (N_13,In_95,In_728);
or U14 (N_14,In_568,In_135);
xnor U15 (N_15,In_458,In_720);
nor U16 (N_16,In_606,In_488);
or U17 (N_17,In_117,In_979);
xnor U18 (N_18,In_764,In_436);
nor U19 (N_19,In_848,In_112);
nor U20 (N_20,In_463,In_462);
xor U21 (N_21,In_304,In_83);
xnor U22 (N_22,In_331,In_303);
or U23 (N_23,In_477,In_226);
nand U24 (N_24,In_445,In_403);
xor U25 (N_25,In_310,In_134);
and U26 (N_26,In_991,In_999);
nand U27 (N_27,In_371,In_993);
nor U28 (N_28,In_459,In_334);
nor U29 (N_29,In_697,In_305);
xnor U30 (N_30,In_485,In_46);
xnor U31 (N_31,In_825,In_851);
and U32 (N_32,In_673,In_104);
nor U33 (N_33,In_642,In_274);
nor U34 (N_34,In_600,In_654);
xor U35 (N_35,In_343,In_312);
nor U36 (N_36,In_480,In_726);
or U37 (N_37,In_996,In_174);
nor U38 (N_38,In_421,In_52);
xnor U39 (N_39,In_60,In_633);
xor U40 (N_40,In_789,In_820);
or U41 (N_41,In_625,In_430);
and U42 (N_42,In_181,In_894);
or U43 (N_43,In_35,In_301);
and U44 (N_44,In_861,In_186);
nand U45 (N_45,In_797,In_839);
or U46 (N_46,In_845,In_241);
and U47 (N_47,In_583,In_729);
nand U48 (N_48,In_951,In_218);
nand U49 (N_49,In_145,In_318);
and U50 (N_50,In_139,In_317);
and U51 (N_51,In_6,In_567);
and U52 (N_52,In_147,In_746);
or U53 (N_53,In_569,In_667);
xnor U54 (N_54,In_860,In_285);
xnor U55 (N_55,In_683,In_877);
or U56 (N_56,In_206,In_224);
nand U57 (N_57,In_661,In_249);
and U58 (N_58,In_389,In_363);
or U59 (N_59,In_639,In_479);
or U60 (N_60,In_131,In_70);
nand U61 (N_61,In_233,In_31);
nor U62 (N_62,In_596,In_98);
nor U63 (N_63,In_250,In_33);
nor U64 (N_64,In_399,In_743);
nor U65 (N_65,In_816,In_874);
or U66 (N_66,In_702,In_539);
nor U67 (N_67,In_838,In_947);
nand U68 (N_68,In_45,In_414);
or U69 (N_69,In_366,In_563);
and U70 (N_70,In_785,In_169);
nor U71 (N_71,In_308,In_342);
and U72 (N_72,In_916,In_635);
xor U73 (N_73,In_184,In_928);
xor U74 (N_74,In_122,In_679);
xnor U75 (N_75,In_209,In_895);
nor U76 (N_76,In_686,In_741);
and U77 (N_77,In_230,In_292);
xnor U78 (N_78,In_144,In_976);
xnor U79 (N_79,In_193,In_791);
or U80 (N_80,In_82,In_689);
nand U81 (N_81,In_751,In_504);
nand U82 (N_82,In_202,In_532);
xor U83 (N_83,In_938,In_182);
or U84 (N_84,In_101,In_244);
xor U85 (N_85,In_293,In_943);
nor U86 (N_86,In_843,In_971);
xnor U87 (N_87,In_452,In_377);
or U88 (N_88,In_829,In_752);
nor U89 (N_89,In_196,In_234);
xor U90 (N_90,In_946,In_63);
nor U91 (N_91,In_256,In_869);
or U92 (N_92,In_964,In_676);
and U93 (N_93,In_713,In_10);
xor U94 (N_94,In_309,In_509);
nand U95 (N_95,In_681,In_191);
nor U96 (N_96,In_219,In_836);
xnor U97 (N_97,In_529,In_538);
nand U98 (N_98,In_264,In_662);
or U99 (N_99,In_253,In_392);
nor U100 (N_100,In_141,In_517);
and U101 (N_101,In_175,In_906);
and U102 (N_102,In_688,In_449);
xnor U103 (N_103,In_631,In_800);
nand U104 (N_104,In_878,In_914);
and U105 (N_105,In_856,In_168);
nand U106 (N_106,In_613,In_283);
or U107 (N_107,In_893,In_769);
and U108 (N_108,In_59,In_411);
nor U109 (N_109,In_106,In_8);
or U110 (N_110,In_963,In_486);
or U111 (N_111,In_849,In_133);
nor U112 (N_112,In_275,In_448);
xnor U113 (N_113,In_37,In_99);
nor U114 (N_114,In_56,In_794);
and U115 (N_115,In_513,In_238);
or U116 (N_116,In_502,In_936);
nor U117 (N_117,In_278,In_602);
or U118 (N_118,In_624,In_398);
or U119 (N_119,In_153,In_261);
or U120 (N_120,In_346,In_390);
xor U121 (N_121,In_775,In_332);
nand U122 (N_122,In_232,In_587);
nand U123 (N_123,In_680,In_972);
and U124 (N_124,In_454,In_973);
nand U125 (N_125,In_551,In_723);
nand U126 (N_126,In_722,In_997);
nor U127 (N_127,In_508,In_5);
and U128 (N_128,In_362,In_432);
or U129 (N_129,In_798,In_473);
nand U130 (N_130,In_79,In_647);
nor U131 (N_131,In_322,In_474);
xor U132 (N_132,In_176,In_614);
nor U133 (N_133,In_585,In_691);
xor U134 (N_134,In_985,In_211);
xor U135 (N_135,In_354,In_382);
or U136 (N_136,In_656,In_792);
nand U137 (N_137,In_657,In_749);
and U138 (N_138,In_648,In_300);
nand U139 (N_139,In_113,In_81);
nor U140 (N_140,In_565,In_566);
xor U141 (N_141,In_511,In_588);
nand U142 (N_142,In_388,In_665);
xnor U143 (N_143,In_26,In_571);
and U144 (N_144,In_365,In_802);
nand U145 (N_145,In_137,In_690);
and U146 (N_146,In_368,In_968);
xor U147 (N_147,In_952,In_151);
nand U148 (N_148,In_840,In_937);
nor U149 (N_149,In_594,In_97);
xnor U150 (N_150,In_160,In_774);
nor U151 (N_151,In_361,In_505);
xor U152 (N_152,In_883,In_919);
and U153 (N_153,In_959,In_240);
xor U154 (N_154,In_801,In_889);
and U155 (N_155,In_197,In_172);
xnor U156 (N_156,In_49,In_767);
and U157 (N_157,In_482,In_68);
nor U158 (N_158,In_91,In_61);
nand U159 (N_159,In_161,In_955);
or U160 (N_160,In_875,In_140);
or U161 (N_161,In_696,In_188);
xor U162 (N_162,In_214,In_57);
nand U163 (N_163,In_653,In_666);
xnor U164 (N_164,In_216,In_143);
xor U165 (N_165,In_675,In_74);
nor U166 (N_166,In_48,In_649);
nand U167 (N_167,In_251,In_965);
nor U168 (N_168,In_779,In_616);
nand U169 (N_169,In_351,In_902);
nand U170 (N_170,In_948,In_898);
or U171 (N_171,In_822,In_194);
nor U172 (N_172,In_407,In_730);
nand U173 (N_173,In_886,In_13);
or U174 (N_174,In_373,In_263);
nand U175 (N_175,In_525,In_711);
and U176 (N_176,In_533,In_17);
and U177 (N_177,In_467,In_913);
or U178 (N_178,In_531,In_977);
nand U179 (N_179,In_475,In_917);
xnor U180 (N_180,In_761,In_957);
and U181 (N_181,In_591,In_827);
nand U182 (N_182,In_423,In_198);
nor U183 (N_183,In_327,In_205);
or U184 (N_184,In_821,In_367);
nand U185 (N_185,In_41,In_557);
and U186 (N_186,In_506,In_772);
nor U187 (N_187,In_88,In_21);
nand U188 (N_188,In_280,In_180);
and U189 (N_189,In_541,In_905);
or U190 (N_190,In_215,In_788);
and U191 (N_191,In_73,In_727);
nor U192 (N_192,In_950,In_818);
or U193 (N_193,In_86,In_805);
or U194 (N_194,In_469,In_124);
and U195 (N_195,In_259,In_966);
nand U196 (N_196,In_989,In_406);
and U197 (N_197,In_518,In_72);
and U198 (N_198,In_384,In_415);
or U199 (N_199,In_337,In_933);
xor U200 (N_200,In_111,In_806);
nor U201 (N_201,In_830,In_495);
xor U202 (N_202,In_926,In_987);
and U203 (N_203,In_441,In_753);
or U204 (N_204,In_353,In_273);
or U205 (N_205,In_745,In_929);
nand U206 (N_206,In_659,In_413);
xnor U207 (N_207,In_815,In_246);
xnor U208 (N_208,In_148,In_739);
xor U209 (N_209,In_235,In_416);
and U210 (N_210,In_760,In_412);
or U211 (N_211,In_766,In_961);
or U212 (N_212,In_858,In_763);
and U213 (N_213,In_289,In_636);
nand U214 (N_214,In_582,In_885);
nor U215 (N_215,In_4,In_655);
xnor U216 (N_216,In_786,In_379);
and U217 (N_217,In_975,In_721);
xnor U218 (N_218,In_494,In_632);
nor U219 (N_219,In_155,In_530);
and U220 (N_220,In_408,In_378);
nor U221 (N_221,In_790,In_684);
xor U222 (N_222,In_804,In_547);
and U223 (N_223,In_94,In_510);
xor U224 (N_224,In_440,In_497);
xor U225 (N_225,In_619,In_370);
nor U226 (N_226,In_247,In_484);
or U227 (N_227,In_626,In_281);
xor U228 (N_228,In_707,In_778);
xnor U229 (N_229,In_941,In_225);
xor U230 (N_230,In_62,In_734);
nand U231 (N_231,In_844,In_55);
and U232 (N_232,In_694,In_863);
nor U233 (N_233,In_114,In_67);
or U234 (N_234,In_853,In_574);
and U235 (N_235,In_515,In_284);
xnor U236 (N_236,In_740,In_121);
xnor U237 (N_237,In_426,In_699);
or U238 (N_238,In_835,In_693);
nor U239 (N_239,In_277,In_341);
xor U240 (N_240,In_298,In_444);
or U241 (N_241,In_23,In_76);
and U242 (N_242,In_781,In_190);
nor U243 (N_243,In_931,In_347);
xnor U244 (N_244,In_357,In_773);
and U245 (N_245,In_149,In_622);
xnor U246 (N_246,In_220,In_3);
and U247 (N_247,In_254,In_607);
and U248 (N_248,In_324,In_50);
nor U249 (N_249,In_876,In_66);
or U250 (N_250,In_813,In_704);
nor U251 (N_251,In_80,In_643);
nand U252 (N_252,In_335,In_663);
nor U253 (N_253,In_701,In_425);
xor U254 (N_254,In_2,In_672);
and U255 (N_255,In_669,In_383);
and U256 (N_256,In_524,In_290);
xor U257 (N_257,In_754,In_901);
nand U258 (N_258,In_712,In_276);
nand U259 (N_259,In_265,In_204);
and U260 (N_260,In_439,In_500);
and U261 (N_261,In_345,In_34);
and U262 (N_262,In_603,In_958);
or U263 (N_263,In_719,In_930);
xor U264 (N_264,In_271,In_550);
nor U265 (N_265,In_455,In_824);
xnor U266 (N_266,In_269,In_18);
nand U267 (N_267,In_814,In_595);
xnor U268 (N_268,In_579,In_857);
nand U269 (N_269,In_323,In_200);
or U270 (N_270,In_629,In_572);
nand U271 (N_271,In_146,In_252);
or U272 (N_272,In_167,In_674);
or U273 (N_273,In_255,In_904);
nand U274 (N_274,In_282,In_921);
nor U275 (N_275,In_879,In_733);
xor U276 (N_276,In_534,In_442);
nand U277 (N_277,In_640,In_808);
xnor U278 (N_278,In_450,In_553);
or U279 (N_279,In_39,In_424);
or U280 (N_280,In_810,In_356);
nand U281 (N_281,In_294,In_288);
and U282 (N_282,In_385,In_328);
xnor U283 (N_283,In_248,In_36);
and U284 (N_284,In_725,In_29);
nor U285 (N_285,In_490,In_742);
or U286 (N_286,In_142,In_77);
nor U287 (N_287,In_872,In_942);
xnor U288 (N_288,In_521,In_223);
nand U289 (N_289,In_42,In_333);
xor U290 (N_290,In_978,In_478);
or U291 (N_291,In_84,In_201);
or U292 (N_292,In_664,In_589);
and U293 (N_293,In_854,In_833);
and U294 (N_294,In_710,In_27);
xnor U295 (N_295,In_897,In_545);
or U296 (N_296,In_164,In_492);
xor U297 (N_297,In_446,In_803);
nand U298 (N_298,In_157,In_910);
xor U299 (N_299,In_750,In_239);
xnor U300 (N_300,In_108,In_562);
or U301 (N_301,In_771,In_348);
xnor U302 (N_302,In_586,In_758);
xnor U303 (N_303,In_336,In_981);
xnor U304 (N_304,In_796,In_575);
nand U305 (N_305,In_115,In_837);
nand U306 (N_306,In_394,In_892);
xnor U307 (N_307,In_28,In_391);
nand U308 (N_308,In_687,In_866);
nor U309 (N_309,In_708,In_460);
nor U310 (N_310,In_850,In_811);
xor U311 (N_311,In_862,In_173);
nand U312 (N_312,In_355,In_868);
xnor U313 (N_313,In_576,In_842);
nor U314 (N_314,In_888,In_192);
xnor U315 (N_315,In_116,In_907);
and U316 (N_316,In_402,In_501);
xor U317 (N_317,In_590,In_735);
nand U318 (N_318,In_162,In_852);
or U319 (N_319,In_349,In_100);
xnor U320 (N_320,In_682,In_266);
and U321 (N_321,In_471,In_499);
and U322 (N_322,In_468,In_11);
nand U323 (N_323,In_387,In_599);
and U324 (N_324,In_890,In_306);
nor U325 (N_325,In_243,In_685);
nor U326 (N_326,In_185,In_608);
or U327 (N_327,In_522,In_369);
or U328 (N_328,In_560,In_299);
or U329 (N_329,In_549,In_177);
or U330 (N_330,In_552,In_130);
nand U331 (N_331,In_321,In_109);
xor U332 (N_332,In_364,In_660);
nand U333 (N_333,In_834,In_823);
and U334 (N_334,In_717,In_986);
xor U335 (N_335,In_592,In_736);
and U336 (N_336,In_940,In_970);
or U337 (N_337,In_85,In_405);
nor U338 (N_338,In_698,In_507);
nand U339 (N_339,In_123,In_212);
xnor U340 (N_340,In_410,In_69);
and U341 (N_341,In_136,In_543);
or U342 (N_342,In_765,In_924);
and U343 (N_343,In_677,In_604);
or U344 (N_344,In_555,In_998);
nand U345 (N_345,In_923,In_418);
or U346 (N_346,In_903,In_24);
xor U347 (N_347,In_447,In_873);
nand U348 (N_348,In_757,In_841);
nor U349 (N_349,In_314,In_340);
nand U350 (N_350,In_623,In_171);
nor U351 (N_351,In_967,In_210);
nand U352 (N_352,In_953,In_434);
and U353 (N_353,In_644,In_195);
nor U354 (N_354,In_496,In_828);
nand U355 (N_355,In_457,In_561);
and U356 (N_356,In_465,In_296);
or U357 (N_357,In_609,In_325);
xnor U358 (N_358,In_150,In_612);
xor U359 (N_359,In_756,In_922);
and U360 (N_360,In_896,In_199);
and U361 (N_361,In_96,In_311);
or U362 (N_362,In_78,In_925);
xor U363 (N_363,In_213,In_537);
nor U364 (N_364,In_127,In_295);
nor U365 (N_365,In_528,In_19);
and U366 (N_366,In_634,In_705);
nand U367 (N_367,In_714,In_451);
nor U368 (N_368,In_983,In_154);
or U369 (N_369,In_481,In_208);
nand U370 (N_370,In_16,In_32);
nor U371 (N_371,In_287,In_747);
nor U372 (N_372,In_880,In_927);
or U373 (N_373,In_152,In_9);
and U374 (N_374,In_584,In_787);
and U375 (N_375,In_386,In_939);
and U376 (N_376,In_315,In_268);
nor U377 (N_377,In_102,In_187);
nor U378 (N_378,In_170,In_65);
or U379 (N_379,In_435,In_540);
nor U380 (N_380,In_548,In_491);
or U381 (N_381,In_25,In_75);
xor U382 (N_382,In_38,In_64);
and U383 (N_383,In_90,In_670);
nand U384 (N_384,In_846,In_47);
and U385 (N_385,In_260,In_912);
xor U386 (N_386,In_703,In_718);
xor U387 (N_387,In_443,In_519);
xor U388 (N_388,In_855,In_692);
and U389 (N_389,In_453,In_493);
xnor U390 (N_390,In_770,In_706);
or U391 (N_391,In_994,In_165);
or U392 (N_392,In_417,In_795);
nand U393 (N_393,In_716,In_126);
or U394 (N_394,In_630,In_159);
nor U395 (N_395,In_558,In_954);
and U396 (N_396,In_372,In_125);
and U397 (N_397,In_884,In_270);
and U398 (N_398,In_593,In_807);
or U399 (N_399,In_578,In_87);
or U400 (N_400,In_542,In_628);
xnor U401 (N_401,In_782,In_470);
xnor U402 (N_402,In_918,In_573);
or U403 (N_403,In_819,In_227);
nor U404 (N_404,In_535,In_646);
nand U405 (N_405,In_419,In_44);
xor U406 (N_406,In_944,In_668);
nand U407 (N_407,In_605,In_228);
and U408 (N_408,In_236,In_960);
or U409 (N_409,In_611,In_54);
and U410 (N_410,In_71,In_974);
xor U411 (N_411,In_330,In_272);
and U412 (N_412,In_621,In_615);
or U413 (N_413,In_598,In_380);
or U414 (N_414,In_637,In_119);
xnor U415 (N_415,In_620,In_516);
and U416 (N_416,In_128,In_645);
and U417 (N_417,In_783,In_617);
or U418 (N_418,In_438,In_319);
nand U419 (N_419,In_344,In_103);
nand U420 (N_420,In_709,In_110);
xnor U421 (N_421,In_536,In_279);
nand U422 (N_422,In_658,In_237);
or U423 (N_423,In_732,In_51);
xor U424 (N_424,In_222,In_360);
and U425 (N_425,In_326,In_376);
or U426 (N_426,In_487,In_118);
nand U427 (N_427,In_678,In_132);
xor U428 (N_428,In_105,In_597);
nor U429 (N_429,In_738,In_920);
xnor U430 (N_430,In_428,In_397);
and U431 (N_431,In_867,In_881);
nor U432 (N_432,In_258,In_14);
nand U433 (N_433,In_338,In_564);
and U434 (N_434,In_207,In_984);
nand U435 (N_435,In_242,In_93);
nand U436 (N_436,In_776,In_189);
nor U437 (N_437,In_178,In_433);
nand U438 (N_438,In_514,In_650);
nor U439 (N_439,In_431,In_217);
or U440 (N_440,In_724,In_871);
xor U441 (N_441,In_887,In_262);
nand U442 (N_442,In_581,In_393);
or U443 (N_443,In_908,In_826);
nand U444 (N_444,In_882,In_358);
and U445 (N_445,In_329,In_30);
nand U446 (N_446,In_731,In_320);
xnor U447 (N_447,In_992,In_183);
nand U448 (N_448,In_969,In_291);
nand U449 (N_449,In_456,In_400);
or U450 (N_450,In_245,In_464);
and U451 (N_451,In_831,In_762);
or U452 (N_452,In_809,In_638);
xor U453 (N_453,In_847,In_58);
and U454 (N_454,In_651,In_12);
or U455 (N_455,In_352,In_267);
nor U456 (N_456,In_375,In_374);
xnor U457 (N_457,In_286,In_627);
nor U458 (N_458,In_20,In_817);
xor U459 (N_459,In_40,In_715);
and U460 (N_460,In_221,In_949);
and U461 (N_461,In_53,In_755);
nor U462 (N_462,In_422,In_409);
or U463 (N_463,In_956,In_671);
xor U464 (N_464,In_229,In_489);
nand U465 (N_465,In_935,In_777);
xnor U466 (N_466,In_527,In_618);
xor U467 (N_467,In_695,In_503);
xnor U468 (N_468,In_784,In_476);
nor U469 (N_469,In_395,In_793);
xnor U470 (N_470,In_932,In_483);
or U471 (N_471,In_865,In_138);
and U472 (N_472,In_420,In_129);
nand U473 (N_473,In_859,In_401);
or U474 (N_474,In_15,In_915);
and U475 (N_475,In_980,In_472);
and U476 (N_476,In_544,In_107);
nand U477 (N_477,In_359,In_156);
nand U478 (N_478,In_799,In_744);
and U479 (N_479,In_120,In_461);
or U480 (N_480,In_466,In_158);
and U481 (N_481,In_909,In_759);
xor U482 (N_482,In_900,In_911);
or U483 (N_483,In_870,In_512);
xor U484 (N_484,In_780,In_1);
nor U485 (N_485,In_313,In_982);
or U486 (N_486,In_899,In_577);
nand U487 (N_487,In_580,In_610);
xor U488 (N_488,In_546,In_962);
and U489 (N_489,In_404,In_43);
and U490 (N_490,In_748,In_990);
or U491 (N_491,In_166,In_995);
xor U492 (N_492,In_316,In_22);
nand U493 (N_493,In_700,In_231);
xnor U494 (N_494,In_812,In_307);
and U495 (N_495,In_520,In_89);
nand U496 (N_496,In_601,In_652);
xor U497 (N_497,In_203,In_7);
xor U498 (N_498,In_257,In_559);
nor U499 (N_499,In_429,In_768);
nand U500 (N_500,In_717,In_80);
or U501 (N_501,In_974,In_932);
xor U502 (N_502,In_337,In_988);
and U503 (N_503,In_983,In_649);
xnor U504 (N_504,In_718,In_164);
and U505 (N_505,In_117,In_573);
xnor U506 (N_506,In_270,In_710);
xor U507 (N_507,In_197,In_122);
nor U508 (N_508,In_48,In_370);
or U509 (N_509,In_170,In_917);
xnor U510 (N_510,In_785,In_448);
or U511 (N_511,In_365,In_492);
xor U512 (N_512,In_989,In_232);
or U513 (N_513,In_180,In_434);
or U514 (N_514,In_698,In_170);
nand U515 (N_515,In_557,In_747);
and U516 (N_516,In_792,In_452);
nor U517 (N_517,In_31,In_77);
and U518 (N_518,In_825,In_662);
nand U519 (N_519,In_573,In_690);
xor U520 (N_520,In_528,In_837);
nand U521 (N_521,In_560,In_873);
xnor U522 (N_522,In_77,In_546);
nand U523 (N_523,In_641,In_395);
nor U524 (N_524,In_556,In_451);
nor U525 (N_525,In_995,In_705);
and U526 (N_526,In_69,In_663);
or U527 (N_527,In_897,In_981);
xor U528 (N_528,In_542,In_721);
nand U529 (N_529,In_897,In_975);
or U530 (N_530,In_575,In_543);
nand U531 (N_531,In_832,In_962);
xor U532 (N_532,In_102,In_360);
and U533 (N_533,In_656,In_467);
xor U534 (N_534,In_709,In_789);
and U535 (N_535,In_194,In_247);
nor U536 (N_536,In_958,In_777);
nand U537 (N_537,In_626,In_304);
nand U538 (N_538,In_71,In_955);
xnor U539 (N_539,In_76,In_482);
nor U540 (N_540,In_567,In_775);
xor U541 (N_541,In_85,In_59);
nor U542 (N_542,In_38,In_993);
xnor U543 (N_543,In_289,In_15);
or U544 (N_544,In_221,In_303);
nand U545 (N_545,In_912,In_730);
nor U546 (N_546,In_58,In_659);
and U547 (N_547,In_887,In_94);
or U548 (N_548,In_251,In_64);
nor U549 (N_549,In_728,In_213);
and U550 (N_550,In_100,In_124);
nand U551 (N_551,In_290,In_702);
and U552 (N_552,In_574,In_610);
or U553 (N_553,In_50,In_427);
nand U554 (N_554,In_48,In_490);
nor U555 (N_555,In_43,In_109);
and U556 (N_556,In_779,In_803);
or U557 (N_557,In_459,In_834);
nand U558 (N_558,In_310,In_79);
nand U559 (N_559,In_752,In_563);
and U560 (N_560,In_757,In_883);
or U561 (N_561,In_280,In_622);
xor U562 (N_562,In_51,In_419);
nand U563 (N_563,In_45,In_265);
and U564 (N_564,In_728,In_83);
xnor U565 (N_565,In_948,In_828);
and U566 (N_566,In_472,In_753);
and U567 (N_567,In_674,In_467);
nor U568 (N_568,In_708,In_347);
nor U569 (N_569,In_819,In_621);
and U570 (N_570,In_459,In_663);
nor U571 (N_571,In_851,In_347);
nor U572 (N_572,In_282,In_589);
nand U573 (N_573,In_474,In_550);
or U574 (N_574,In_824,In_980);
xor U575 (N_575,In_742,In_250);
and U576 (N_576,In_77,In_971);
xor U577 (N_577,In_826,In_348);
nor U578 (N_578,In_703,In_391);
and U579 (N_579,In_902,In_490);
or U580 (N_580,In_164,In_350);
nor U581 (N_581,In_835,In_198);
or U582 (N_582,In_728,In_387);
and U583 (N_583,In_974,In_965);
xnor U584 (N_584,In_785,In_956);
nor U585 (N_585,In_19,In_652);
xor U586 (N_586,In_385,In_960);
and U587 (N_587,In_476,In_361);
or U588 (N_588,In_318,In_949);
nor U589 (N_589,In_286,In_765);
xor U590 (N_590,In_818,In_56);
and U591 (N_591,In_456,In_803);
or U592 (N_592,In_710,In_811);
xor U593 (N_593,In_394,In_708);
nor U594 (N_594,In_765,In_757);
or U595 (N_595,In_201,In_289);
or U596 (N_596,In_417,In_857);
nor U597 (N_597,In_752,In_706);
xor U598 (N_598,In_196,In_335);
nor U599 (N_599,In_88,In_120);
and U600 (N_600,In_311,In_606);
or U601 (N_601,In_256,In_329);
nor U602 (N_602,In_570,In_128);
and U603 (N_603,In_954,In_308);
nor U604 (N_604,In_842,In_315);
or U605 (N_605,In_940,In_5);
and U606 (N_606,In_426,In_403);
or U607 (N_607,In_153,In_416);
xor U608 (N_608,In_247,In_649);
and U609 (N_609,In_741,In_226);
and U610 (N_610,In_192,In_452);
and U611 (N_611,In_753,In_688);
or U612 (N_612,In_518,In_697);
and U613 (N_613,In_702,In_277);
nand U614 (N_614,In_530,In_745);
nand U615 (N_615,In_878,In_606);
xor U616 (N_616,In_585,In_617);
or U617 (N_617,In_768,In_834);
xnor U618 (N_618,In_159,In_201);
or U619 (N_619,In_994,In_304);
nor U620 (N_620,In_485,In_496);
nor U621 (N_621,In_225,In_350);
nor U622 (N_622,In_875,In_656);
and U623 (N_623,In_694,In_795);
nand U624 (N_624,In_590,In_258);
nand U625 (N_625,In_2,In_932);
nand U626 (N_626,In_424,In_104);
xor U627 (N_627,In_456,In_582);
or U628 (N_628,In_330,In_382);
xnor U629 (N_629,In_395,In_995);
nor U630 (N_630,In_533,In_31);
xor U631 (N_631,In_981,In_296);
and U632 (N_632,In_544,In_261);
nand U633 (N_633,In_894,In_657);
xnor U634 (N_634,In_741,In_582);
or U635 (N_635,In_294,In_525);
or U636 (N_636,In_962,In_269);
xor U637 (N_637,In_943,In_806);
nand U638 (N_638,In_452,In_45);
xor U639 (N_639,In_807,In_60);
nor U640 (N_640,In_889,In_681);
nand U641 (N_641,In_829,In_849);
nor U642 (N_642,In_855,In_766);
nand U643 (N_643,In_808,In_44);
nand U644 (N_644,In_256,In_483);
xnor U645 (N_645,In_260,In_721);
nand U646 (N_646,In_825,In_856);
or U647 (N_647,In_662,In_462);
nand U648 (N_648,In_241,In_429);
nand U649 (N_649,In_749,In_679);
or U650 (N_650,In_683,In_593);
and U651 (N_651,In_110,In_856);
xor U652 (N_652,In_203,In_166);
and U653 (N_653,In_692,In_380);
xnor U654 (N_654,In_693,In_574);
nor U655 (N_655,In_411,In_816);
or U656 (N_656,In_855,In_307);
nand U657 (N_657,In_870,In_529);
nand U658 (N_658,In_778,In_376);
nand U659 (N_659,In_774,In_918);
or U660 (N_660,In_966,In_34);
nor U661 (N_661,In_905,In_122);
xor U662 (N_662,In_293,In_54);
and U663 (N_663,In_31,In_865);
or U664 (N_664,In_117,In_262);
nor U665 (N_665,In_957,In_176);
xnor U666 (N_666,In_827,In_686);
and U667 (N_667,In_222,In_607);
and U668 (N_668,In_755,In_914);
nor U669 (N_669,In_98,In_622);
nor U670 (N_670,In_304,In_521);
and U671 (N_671,In_238,In_521);
or U672 (N_672,In_642,In_80);
nor U673 (N_673,In_593,In_293);
nand U674 (N_674,In_592,In_255);
nand U675 (N_675,In_918,In_416);
nand U676 (N_676,In_15,In_360);
nor U677 (N_677,In_646,In_903);
and U678 (N_678,In_490,In_712);
or U679 (N_679,In_550,In_872);
xor U680 (N_680,In_644,In_403);
xor U681 (N_681,In_574,In_933);
or U682 (N_682,In_986,In_16);
nand U683 (N_683,In_317,In_363);
and U684 (N_684,In_365,In_433);
and U685 (N_685,In_245,In_814);
nand U686 (N_686,In_373,In_783);
and U687 (N_687,In_982,In_228);
or U688 (N_688,In_362,In_760);
nand U689 (N_689,In_811,In_427);
or U690 (N_690,In_653,In_171);
nor U691 (N_691,In_361,In_480);
nor U692 (N_692,In_720,In_555);
nand U693 (N_693,In_448,In_433);
nand U694 (N_694,In_869,In_606);
or U695 (N_695,In_792,In_910);
nand U696 (N_696,In_618,In_130);
nor U697 (N_697,In_219,In_463);
nor U698 (N_698,In_194,In_288);
or U699 (N_699,In_183,In_333);
nand U700 (N_700,In_489,In_936);
or U701 (N_701,In_336,In_730);
or U702 (N_702,In_725,In_663);
or U703 (N_703,In_955,In_860);
nand U704 (N_704,In_92,In_522);
and U705 (N_705,In_102,In_870);
nand U706 (N_706,In_361,In_390);
nand U707 (N_707,In_957,In_131);
nand U708 (N_708,In_557,In_441);
and U709 (N_709,In_294,In_542);
xor U710 (N_710,In_252,In_491);
and U711 (N_711,In_120,In_82);
and U712 (N_712,In_838,In_210);
xnor U713 (N_713,In_16,In_541);
and U714 (N_714,In_928,In_766);
nor U715 (N_715,In_516,In_62);
nand U716 (N_716,In_492,In_915);
and U717 (N_717,In_853,In_946);
nor U718 (N_718,In_87,In_909);
nand U719 (N_719,In_126,In_243);
or U720 (N_720,In_787,In_168);
xnor U721 (N_721,In_231,In_338);
nor U722 (N_722,In_566,In_836);
and U723 (N_723,In_298,In_485);
or U724 (N_724,In_850,In_603);
xnor U725 (N_725,In_341,In_182);
xnor U726 (N_726,In_577,In_683);
nor U727 (N_727,In_741,In_966);
and U728 (N_728,In_202,In_763);
nor U729 (N_729,In_409,In_311);
or U730 (N_730,In_46,In_126);
xnor U731 (N_731,In_340,In_473);
nor U732 (N_732,In_381,In_431);
or U733 (N_733,In_691,In_30);
and U734 (N_734,In_249,In_96);
and U735 (N_735,In_768,In_928);
nand U736 (N_736,In_846,In_745);
or U737 (N_737,In_621,In_343);
nand U738 (N_738,In_293,In_448);
and U739 (N_739,In_214,In_925);
and U740 (N_740,In_826,In_992);
nand U741 (N_741,In_719,In_169);
nor U742 (N_742,In_101,In_79);
nand U743 (N_743,In_142,In_129);
or U744 (N_744,In_18,In_909);
nor U745 (N_745,In_739,In_400);
nor U746 (N_746,In_860,In_779);
xnor U747 (N_747,In_681,In_922);
nand U748 (N_748,In_11,In_190);
or U749 (N_749,In_556,In_676);
xor U750 (N_750,In_302,In_598);
nor U751 (N_751,In_945,In_41);
xor U752 (N_752,In_881,In_783);
nand U753 (N_753,In_114,In_987);
and U754 (N_754,In_948,In_224);
nand U755 (N_755,In_325,In_882);
or U756 (N_756,In_610,In_620);
xor U757 (N_757,In_849,In_571);
and U758 (N_758,In_467,In_163);
and U759 (N_759,In_393,In_807);
or U760 (N_760,In_974,In_363);
xor U761 (N_761,In_58,In_585);
and U762 (N_762,In_1,In_201);
nand U763 (N_763,In_375,In_394);
nand U764 (N_764,In_474,In_144);
or U765 (N_765,In_641,In_638);
nand U766 (N_766,In_776,In_716);
and U767 (N_767,In_766,In_919);
nor U768 (N_768,In_788,In_417);
xor U769 (N_769,In_429,In_611);
nand U770 (N_770,In_892,In_284);
or U771 (N_771,In_398,In_701);
or U772 (N_772,In_212,In_341);
nor U773 (N_773,In_158,In_111);
or U774 (N_774,In_472,In_283);
nand U775 (N_775,In_307,In_241);
xor U776 (N_776,In_397,In_661);
or U777 (N_777,In_263,In_80);
and U778 (N_778,In_5,In_878);
nor U779 (N_779,In_376,In_296);
and U780 (N_780,In_980,In_501);
xnor U781 (N_781,In_272,In_332);
or U782 (N_782,In_397,In_570);
xor U783 (N_783,In_650,In_110);
nor U784 (N_784,In_763,In_767);
nand U785 (N_785,In_542,In_817);
xor U786 (N_786,In_761,In_833);
nor U787 (N_787,In_691,In_66);
xor U788 (N_788,In_379,In_812);
nor U789 (N_789,In_501,In_394);
xor U790 (N_790,In_548,In_789);
nor U791 (N_791,In_489,In_993);
nand U792 (N_792,In_861,In_579);
and U793 (N_793,In_206,In_655);
nor U794 (N_794,In_964,In_435);
nand U795 (N_795,In_721,In_871);
nand U796 (N_796,In_50,In_787);
nor U797 (N_797,In_436,In_198);
nand U798 (N_798,In_413,In_985);
nor U799 (N_799,In_969,In_811);
or U800 (N_800,In_242,In_178);
nor U801 (N_801,In_894,In_425);
xor U802 (N_802,In_650,In_510);
and U803 (N_803,In_222,In_267);
and U804 (N_804,In_9,In_565);
xnor U805 (N_805,In_677,In_494);
xnor U806 (N_806,In_956,In_966);
and U807 (N_807,In_68,In_417);
and U808 (N_808,In_848,In_425);
and U809 (N_809,In_523,In_540);
xor U810 (N_810,In_662,In_388);
nor U811 (N_811,In_748,In_913);
nand U812 (N_812,In_17,In_739);
nand U813 (N_813,In_382,In_620);
nor U814 (N_814,In_386,In_670);
and U815 (N_815,In_753,In_57);
nor U816 (N_816,In_876,In_738);
nand U817 (N_817,In_821,In_629);
nor U818 (N_818,In_205,In_110);
or U819 (N_819,In_655,In_74);
or U820 (N_820,In_512,In_899);
nand U821 (N_821,In_951,In_94);
xnor U822 (N_822,In_719,In_824);
xor U823 (N_823,In_315,In_560);
nand U824 (N_824,In_840,In_738);
nor U825 (N_825,In_233,In_590);
or U826 (N_826,In_412,In_85);
nor U827 (N_827,In_472,In_625);
and U828 (N_828,In_241,In_626);
nand U829 (N_829,In_997,In_327);
or U830 (N_830,In_908,In_627);
xnor U831 (N_831,In_982,In_349);
or U832 (N_832,In_727,In_752);
xor U833 (N_833,In_500,In_956);
and U834 (N_834,In_333,In_691);
or U835 (N_835,In_742,In_747);
and U836 (N_836,In_629,In_117);
and U837 (N_837,In_495,In_512);
and U838 (N_838,In_300,In_461);
xor U839 (N_839,In_837,In_685);
or U840 (N_840,In_62,In_66);
and U841 (N_841,In_549,In_419);
nor U842 (N_842,In_734,In_497);
nor U843 (N_843,In_47,In_385);
xnor U844 (N_844,In_825,In_205);
xor U845 (N_845,In_184,In_561);
and U846 (N_846,In_913,In_487);
nor U847 (N_847,In_173,In_302);
xor U848 (N_848,In_73,In_553);
nor U849 (N_849,In_831,In_32);
or U850 (N_850,In_613,In_190);
and U851 (N_851,In_601,In_413);
xor U852 (N_852,In_181,In_665);
nor U853 (N_853,In_733,In_174);
xnor U854 (N_854,In_98,In_705);
nand U855 (N_855,In_613,In_264);
and U856 (N_856,In_877,In_495);
xor U857 (N_857,In_261,In_191);
and U858 (N_858,In_488,In_957);
xor U859 (N_859,In_222,In_929);
and U860 (N_860,In_831,In_209);
and U861 (N_861,In_56,In_184);
and U862 (N_862,In_340,In_94);
or U863 (N_863,In_669,In_209);
nor U864 (N_864,In_395,In_91);
and U865 (N_865,In_843,In_477);
and U866 (N_866,In_347,In_896);
or U867 (N_867,In_653,In_486);
nor U868 (N_868,In_292,In_139);
nor U869 (N_869,In_967,In_485);
xor U870 (N_870,In_99,In_488);
and U871 (N_871,In_882,In_261);
nor U872 (N_872,In_377,In_209);
and U873 (N_873,In_72,In_776);
xor U874 (N_874,In_761,In_169);
and U875 (N_875,In_40,In_991);
and U876 (N_876,In_733,In_865);
or U877 (N_877,In_515,In_413);
or U878 (N_878,In_452,In_766);
or U879 (N_879,In_257,In_511);
and U880 (N_880,In_45,In_757);
or U881 (N_881,In_890,In_784);
nor U882 (N_882,In_105,In_127);
nand U883 (N_883,In_975,In_793);
nand U884 (N_884,In_858,In_27);
nand U885 (N_885,In_81,In_641);
xnor U886 (N_886,In_683,In_504);
and U887 (N_887,In_945,In_151);
nor U888 (N_888,In_703,In_443);
nor U889 (N_889,In_410,In_790);
nor U890 (N_890,In_30,In_973);
and U891 (N_891,In_201,In_898);
and U892 (N_892,In_851,In_325);
xor U893 (N_893,In_312,In_323);
xor U894 (N_894,In_17,In_956);
and U895 (N_895,In_410,In_557);
nand U896 (N_896,In_446,In_132);
nor U897 (N_897,In_85,In_874);
xnor U898 (N_898,In_502,In_602);
nor U899 (N_899,In_559,In_669);
xnor U900 (N_900,In_879,In_773);
and U901 (N_901,In_332,In_95);
nor U902 (N_902,In_145,In_311);
and U903 (N_903,In_258,In_969);
nand U904 (N_904,In_34,In_414);
xnor U905 (N_905,In_808,In_908);
or U906 (N_906,In_67,In_782);
xor U907 (N_907,In_138,In_433);
xor U908 (N_908,In_745,In_124);
nand U909 (N_909,In_704,In_962);
or U910 (N_910,In_783,In_792);
nor U911 (N_911,In_88,In_130);
and U912 (N_912,In_657,In_116);
xnor U913 (N_913,In_66,In_560);
or U914 (N_914,In_963,In_184);
and U915 (N_915,In_522,In_12);
xor U916 (N_916,In_948,In_291);
or U917 (N_917,In_774,In_335);
xor U918 (N_918,In_500,In_670);
and U919 (N_919,In_607,In_605);
xnor U920 (N_920,In_775,In_688);
or U921 (N_921,In_773,In_398);
nor U922 (N_922,In_604,In_196);
and U923 (N_923,In_56,In_301);
xor U924 (N_924,In_118,In_867);
nand U925 (N_925,In_224,In_347);
and U926 (N_926,In_537,In_616);
nor U927 (N_927,In_487,In_907);
nand U928 (N_928,In_161,In_147);
nor U929 (N_929,In_185,In_243);
or U930 (N_930,In_57,In_866);
nor U931 (N_931,In_498,In_667);
nor U932 (N_932,In_69,In_327);
and U933 (N_933,In_849,In_568);
nor U934 (N_934,In_872,In_625);
or U935 (N_935,In_654,In_248);
xnor U936 (N_936,In_627,In_173);
and U937 (N_937,In_651,In_882);
nand U938 (N_938,In_230,In_673);
nor U939 (N_939,In_377,In_248);
xor U940 (N_940,In_846,In_860);
and U941 (N_941,In_270,In_945);
nand U942 (N_942,In_63,In_464);
or U943 (N_943,In_427,In_324);
xnor U944 (N_944,In_818,In_357);
and U945 (N_945,In_102,In_624);
and U946 (N_946,In_932,In_192);
xnor U947 (N_947,In_338,In_333);
and U948 (N_948,In_140,In_194);
nand U949 (N_949,In_889,In_551);
and U950 (N_950,In_533,In_30);
or U951 (N_951,In_518,In_937);
nor U952 (N_952,In_247,In_433);
or U953 (N_953,In_78,In_957);
nand U954 (N_954,In_988,In_198);
xnor U955 (N_955,In_245,In_252);
xnor U956 (N_956,In_29,In_178);
and U957 (N_957,In_45,In_525);
and U958 (N_958,In_569,In_458);
or U959 (N_959,In_338,In_387);
xor U960 (N_960,In_297,In_858);
or U961 (N_961,In_736,In_808);
and U962 (N_962,In_669,In_879);
and U963 (N_963,In_666,In_255);
and U964 (N_964,In_29,In_51);
nor U965 (N_965,In_762,In_671);
nand U966 (N_966,In_972,In_877);
xor U967 (N_967,In_84,In_510);
nand U968 (N_968,In_802,In_598);
nor U969 (N_969,In_679,In_978);
and U970 (N_970,In_189,In_448);
xnor U971 (N_971,In_217,In_808);
or U972 (N_972,In_558,In_990);
and U973 (N_973,In_522,In_234);
and U974 (N_974,In_118,In_526);
and U975 (N_975,In_868,In_314);
and U976 (N_976,In_677,In_209);
nor U977 (N_977,In_819,In_865);
or U978 (N_978,In_185,In_991);
nor U979 (N_979,In_192,In_672);
and U980 (N_980,In_514,In_258);
nand U981 (N_981,In_7,In_378);
nand U982 (N_982,In_709,In_204);
xnor U983 (N_983,In_319,In_135);
or U984 (N_984,In_457,In_780);
or U985 (N_985,In_590,In_268);
and U986 (N_986,In_791,In_682);
nor U987 (N_987,In_174,In_391);
nor U988 (N_988,In_952,In_917);
or U989 (N_989,In_468,In_643);
or U990 (N_990,In_693,In_679);
xor U991 (N_991,In_515,In_614);
xnor U992 (N_992,In_255,In_268);
xnor U993 (N_993,In_724,In_190);
xor U994 (N_994,In_598,In_989);
and U995 (N_995,In_505,In_333);
and U996 (N_996,In_937,In_82);
and U997 (N_997,In_277,In_591);
and U998 (N_998,In_335,In_694);
or U999 (N_999,In_964,In_333);
and U1000 (N_1000,In_735,In_670);
and U1001 (N_1001,In_143,In_81);
or U1002 (N_1002,In_679,In_358);
nand U1003 (N_1003,In_341,In_720);
xor U1004 (N_1004,In_42,In_840);
nand U1005 (N_1005,In_655,In_963);
or U1006 (N_1006,In_621,In_201);
nor U1007 (N_1007,In_512,In_485);
nor U1008 (N_1008,In_630,In_373);
and U1009 (N_1009,In_284,In_722);
and U1010 (N_1010,In_341,In_854);
or U1011 (N_1011,In_981,In_237);
and U1012 (N_1012,In_859,In_709);
and U1013 (N_1013,In_581,In_333);
and U1014 (N_1014,In_909,In_97);
xor U1015 (N_1015,In_627,In_300);
and U1016 (N_1016,In_11,In_845);
and U1017 (N_1017,In_745,In_220);
xor U1018 (N_1018,In_418,In_371);
nand U1019 (N_1019,In_421,In_1);
xor U1020 (N_1020,In_59,In_452);
or U1021 (N_1021,In_592,In_39);
or U1022 (N_1022,In_269,In_980);
nand U1023 (N_1023,In_298,In_267);
and U1024 (N_1024,In_981,In_47);
and U1025 (N_1025,In_660,In_875);
nand U1026 (N_1026,In_638,In_578);
xor U1027 (N_1027,In_570,In_447);
xor U1028 (N_1028,In_1,In_793);
xor U1029 (N_1029,In_436,In_985);
or U1030 (N_1030,In_638,In_576);
nor U1031 (N_1031,In_232,In_384);
xnor U1032 (N_1032,In_482,In_133);
and U1033 (N_1033,In_596,In_42);
xor U1034 (N_1034,In_172,In_345);
nor U1035 (N_1035,In_583,In_77);
or U1036 (N_1036,In_78,In_369);
or U1037 (N_1037,In_759,In_796);
xnor U1038 (N_1038,In_763,In_263);
nand U1039 (N_1039,In_834,In_234);
nor U1040 (N_1040,In_877,In_643);
nand U1041 (N_1041,In_847,In_718);
nor U1042 (N_1042,In_459,In_108);
nand U1043 (N_1043,In_54,In_918);
xor U1044 (N_1044,In_459,In_354);
or U1045 (N_1045,In_972,In_299);
xnor U1046 (N_1046,In_228,In_857);
and U1047 (N_1047,In_942,In_102);
xor U1048 (N_1048,In_544,In_601);
xor U1049 (N_1049,In_212,In_909);
xor U1050 (N_1050,In_11,In_272);
and U1051 (N_1051,In_675,In_248);
or U1052 (N_1052,In_99,In_649);
xor U1053 (N_1053,In_307,In_270);
xor U1054 (N_1054,In_682,In_958);
nor U1055 (N_1055,In_898,In_769);
nor U1056 (N_1056,In_178,In_658);
and U1057 (N_1057,In_548,In_48);
nor U1058 (N_1058,In_865,In_949);
xor U1059 (N_1059,In_821,In_381);
nand U1060 (N_1060,In_658,In_770);
xnor U1061 (N_1061,In_576,In_468);
nor U1062 (N_1062,In_397,In_245);
or U1063 (N_1063,In_392,In_870);
or U1064 (N_1064,In_59,In_555);
nor U1065 (N_1065,In_646,In_604);
or U1066 (N_1066,In_813,In_605);
or U1067 (N_1067,In_105,In_451);
nor U1068 (N_1068,In_591,In_549);
nor U1069 (N_1069,In_410,In_934);
or U1070 (N_1070,In_438,In_467);
nand U1071 (N_1071,In_497,In_623);
xor U1072 (N_1072,In_438,In_24);
and U1073 (N_1073,In_903,In_334);
nand U1074 (N_1074,In_137,In_372);
xor U1075 (N_1075,In_792,In_618);
and U1076 (N_1076,In_238,In_556);
nand U1077 (N_1077,In_799,In_85);
or U1078 (N_1078,In_664,In_442);
xnor U1079 (N_1079,In_94,In_39);
nor U1080 (N_1080,In_18,In_519);
xor U1081 (N_1081,In_768,In_342);
and U1082 (N_1082,In_17,In_820);
xor U1083 (N_1083,In_32,In_417);
nand U1084 (N_1084,In_282,In_826);
and U1085 (N_1085,In_908,In_153);
xnor U1086 (N_1086,In_150,In_624);
xor U1087 (N_1087,In_238,In_224);
and U1088 (N_1088,In_5,In_516);
or U1089 (N_1089,In_289,In_341);
nor U1090 (N_1090,In_995,In_865);
nand U1091 (N_1091,In_42,In_586);
and U1092 (N_1092,In_568,In_664);
nor U1093 (N_1093,In_749,In_831);
nand U1094 (N_1094,In_218,In_10);
nor U1095 (N_1095,In_907,In_212);
xnor U1096 (N_1096,In_124,In_825);
or U1097 (N_1097,In_461,In_783);
or U1098 (N_1098,In_724,In_163);
and U1099 (N_1099,In_406,In_507);
nand U1100 (N_1100,In_134,In_560);
nand U1101 (N_1101,In_470,In_737);
nand U1102 (N_1102,In_288,In_138);
or U1103 (N_1103,In_890,In_163);
nand U1104 (N_1104,In_799,In_443);
nand U1105 (N_1105,In_696,In_506);
and U1106 (N_1106,In_322,In_642);
xnor U1107 (N_1107,In_58,In_892);
nand U1108 (N_1108,In_856,In_77);
or U1109 (N_1109,In_225,In_398);
nor U1110 (N_1110,In_748,In_267);
or U1111 (N_1111,In_810,In_51);
nor U1112 (N_1112,In_962,In_203);
or U1113 (N_1113,In_198,In_492);
nor U1114 (N_1114,In_317,In_499);
or U1115 (N_1115,In_822,In_847);
and U1116 (N_1116,In_151,In_536);
xor U1117 (N_1117,In_214,In_555);
and U1118 (N_1118,In_331,In_386);
nor U1119 (N_1119,In_149,In_230);
and U1120 (N_1120,In_87,In_137);
and U1121 (N_1121,In_698,In_977);
nand U1122 (N_1122,In_369,In_576);
xor U1123 (N_1123,In_568,In_515);
nor U1124 (N_1124,In_484,In_199);
xor U1125 (N_1125,In_465,In_551);
or U1126 (N_1126,In_983,In_931);
and U1127 (N_1127,In_928,In_701);
nand U1128 (N_1128,In_739,In_963);
and U1129 (N_1129,In_588,In_77);
nand U1130 (N_1130,In_420,In_68);
xor U1131 (N_1131,In_422,In_310);
xor U1132 (N_1132,In_402,In_55);
nor U1133 (N_1133,In_26,In_921);
nor U1134 (N_1134,In_384,In_33);
nand U1135 (N_1135,In_724,In_759);
xor U1136 (N_1136,In_60,In_977);
nor U1137 (N_1137,In_451,In_317);
and U1138 (N_1138,In_100,In_351);
and U1139 (N_1139,In_463,In_445);
and U1140 (N_1140,In_498,In_662);
nor U1141 (N_1141,In_5,In_413);
and U1142 (N_1142,In_920,In_866);
nor U1143 (N_1143,In_948,In_583);
or U1144 (N_1144,In_206,In_987);
nor U1145 (N_1145,In_512,In_364);
nand U1146 (N_1146,In_121,In_779);
xnor U1147 (N_1147,In_838,In_614);
and U1148 (N_1148,In_630,In_323);
xnor U1149 (N_1149,In_302,In_555);
and U1150 (N_1150,In_150,In_188);
nand U1151 (N_1151,In_563,In_692);
or U1152 (N_1152,In_432,In_13);
xnor U1153 (N_1153,In_316,In_275);
or U1154 (N_1154,In_842,In_5);
and U1155 (N_1155,In_20,In_870);
or U1156 (N_1156,In_411,In_577);
nand U1157 (N_1157,In_443,In_127);
nand U1158 (N_1158,In_216,In_658);
or U1159 (N_1159,In_168,In_560);
nand U1160 (N_1160,In_398,In_61);
nand U1161 (N_1161,In_51,In_877);
and U1162 (N_1162,In_935,In_954);
and U1163 (N_1163,In_479,In_711);
xnor U1164 (N_1164,In_347,In_466);
nand U1165 (N_1165,In_45,In_195);
and U1166 (N_1166,In_150,In_254);
and U1167 (N_1167,In_271,In_732);
or U1168 (N_1168,In_828,In_641);
nand U1169 (N_1169,In_683,In_729);
xor U1170 (N_1170,In_828,In_296);
or U1171 (N_1171,In_721,In_256);
xnor U1172 (N_1172,In_921,In_328);
xnor U1173 (N_1173,In_149,In_601);
nor U1174 (N_1174,In_349,In_608);
nand U1175 (N_1175,In_356,In_426);
nand U1176 (N_1176,In_153,In_505);
and U1177 (N_1177,In_451,In_837);
nor U1178 (N_1178,In_994,In_95);
or U1179 (N_1179,In_910,In_190);
or U1180 (N_1180,In_831,In_373);
nand U1181 (N_1181,In_442,In_610);
and U1182 (N_1182,In_546,In_634);
or U1183 (N_1183,In_348,In_834);
nand U1184 (N_1184,In_269,In_285);
xnor U1185 (N_1185,In_961,In_505);
or U1186 (N_1186,In_116,In_534);
xnor U1187 (N_1187,In_265,In_936);
nor U1188 (N_1188,In_648,In_436);
nand U1189 (N_1189,In_49,In_709);
and U1190 (N_1190,In_838,In_434);
xnor U1191 (N_1191,In_922,In_426);
xor U1192 (N_1192,In_562,In_294);
xor U1193 (N_1193,In_142,In_543);
or U1194 (N_1194,In_374,In_833);
and U1195 (N_1195,In_980,In_364);
and U1196 (N_1196,In_428,In_188);
nand U1197 (N_1197,In_707,In_365);
xnor U1198 (N_1198,In_504,In_891);
nor U1199 (N_1199,In_276,In_360);
nand U1200 (N_1200,In_15,In_94);
nor U1201 (N_1201,In_463,In_13);
nor U1202 (N_1202,In_106,In_132);
and U1203 (N_1203,In_508,In_197);
and U1204 (N_1204,In_327,In_118);
xor U1205 (N_1205,In_424,In_902);
and U1206 (N_1206,In_961,In_657);
xor U1207 (N_1207,In_458,In_746);
nor U1208 (N_1208,In_433,In_493);
nor U1209 (N_1209,In_781,In_645);
xor U1210 (N_1210,In_41,In_32);
nand U1211 (N_1211,In_799,In_867);
nor U1212 (N_1212,In_809,In_281);
nor U1213 (N_1213,In_599,In_551);
nand U1214 (N_1214,In_193,In_260);
or U1215 (N_1215,In_248,In_287);
nand U1216 (N_1216,In_403,In_387);
and U1217 (N_1217,In_849,In_900);
and U1218 (N_1218,In_895,In_972);
nand U1219 (N_1219,In_283,In_649);
xor U1220 (N_1220,In_117,In_628);
xnor U1221 (N_1221,In_939,In_638);
or U1222 (N_1222,In_784,In_453);
nand U1223 (N_1223,In_549,In_211);
nand U1224 (N_1224,In_463,In_725);
and U1225 (N_1225,In_412,In_618);
nand U1226 (N_1226,In_272,In_129);
nand U1227 (N_1227,In_445,In_267);
and U1228 (N_1228,In_872,In_476);
nand U1229 (N_1229,In_366,In_247);
nor U1230 (N_1230,In_562,In_370);
nor U1231 (N_1231,In_384,In_375);
and U1232 (N_1232,In_633,In_866);
nor U1233 (N_1233,In_704,In_58);
nor U1234 (N_1234,In_667,In_687);
nor U1235 (N_1235,In_733,In_338);
or U1236 (N_1236,In_343,In_728);
or U1237 (N_1237,In_545,In_136);
nand U1238 (N_1238,In_11,In_301);
nor U1239 (N_1239,In_193,In_225);
xnor U1240 (N_1240,In_389,In_611);
xnor U1241 (N_1241,In_966,In_379);
xnor U1242 (N_1242,In_233,In_896);
or U1243 (N_1243,In_945,In_805);
xnor U1244 (N_1244,In_98,In_7);
xnor U1245 (N_1245,In_958,In_419);
nand U1246 (N_1246,In_79,In_995);
or U1247 (N_1247,In_341,In_514);
xnor U1248 (N_1248,In_444,In_772);
nor U1249 (N_1249,In_998,In_1);
and U1250 (N_1250,In_847,In_608);
xnor U1251 (N_1251,In_420,In_897);
and U1252 (N_1252,In_890,In_682);
xor U1253 (N_1253,In_360,In_346);
nand U1254 (N_1254,In_292,In_465);
and U1255 (N_1255,In_166,In_84);
xnor U1256 (N_1256,In_559,In_68);
xnor U1257 (N_1257,In_507,In_227);
and U1258 (N_1258,In_79,In_786);
nand U1259 (N_1259,In_136,In_827);
nand U1260 (N_1260,In_241,In_445);
and U1261 (N_1261,In_445,In_865);
or U1262 (N_1262,In_55,In_613);
nor U1263 (N_1263,In_152,In_797);
and U1264 (N_1264,In_517,In_664);
nor U1265 (N_1265,In_15,In_265);
and U1266 (N_1266,In_182,In_657);
or U1267 (N_1267,In_636,In_665);
or U1268 (N_1268,In_737,In_999);
xnor U1269 (N_1269,In_988,In_886);
or U1270 (N_1270,In_658,In_884);
or U1271 (N_1271,In_558,In_298);
nor U1272 (N_1272,In_183,In_89);
and U1273 (N_1273,In_336,In_916);
nand U1274 (N_1274,In_781,In_640);
xnor U1275 (N_1275,In_277,In_926);
nor U1276 (N_1276,In_659,In_113);
xnor U1277 (N_1277,In_457,In_249);
nand U1278 (N_1278,In_631,In_441);
xnor U1279 (N_1279,In_923,In_663);
xor U1280 (N_1280,In_847,In_763);
and U1281 (N_1281,In_700,In_295);
xnor U1282 (N_1282,In_41,In_163);
or U1283 (N_1283,In_672,In_54);
nor U1284 (N_1284,In_765,In_635);
or U1285 (N_1285,In_735,In_472);
and U1286 (N_1286,In_106,In_46);
or U1287 (N_1287,In_460,In_468);
nor U1288 (N_1288,In_67,In_169);
nor U1289 (N_1289,In_69,In_474);
nor U1290 (N_1290,In_632,In_566);
nor U1291 (N_1291,In_813,In_22);
nand U1292 (N_1292,In_114,In_113);
nor U1293 (N_1293,In_641,In_416);
nand U1294 (N_1294,In_953,In_580);
and U1295 (N_1295,In_393,In_281);
or U1296 (N_1296,In_248,In_682);
xor U1297 (N_1297,In_866,In_754);
nand U1298 (N_1298,In_945,In_654);
nand U1299 (N_1299,In_686,In_464);
nor U1300 (N_1300,In_32,In_604);
or U1301 (N_1301,In_602,In_636);
and U1302 (N_1302,In_332,In_96);
nand U1303 (N_1303,In_951,In_824);
or U1304 (N_1304,In_705,In_732);
nand U1305 (N_1305,In_502,In_457);
nand U1306 (N_1306,In_750,In_259);
nor U1307 (N_1307,In_850,In_109);
and U1308 (N_1308,In_810,In_299);
or U1309 (N_1309,In_93,In_466);
xnor U1310 (N_1310,In_375,In_425);
xnor U1311 (N_1311,In_801,In_264);
xnor U1312 (N_1312,In_239,In_201);
xnor U1313 (N_1313,In_37,In_887);
xnor U1314 (N_1314,In_610,In_20);
nand U1315 (N_1315,In_99,In_117);
nand U1316 (N_1316,In_988,In_250);
and U1317 (N_1317,In_671,In_785);
xnor U1318 (N_1318,In_594,In_389);
nand U1319 (N_1319,In_325,In_474);
nand U1320 (N_1320,In_821,In_225);
xnor U1321 (N_1321,In_870,In_619);
and U1322 (N_1322,In_366,In_997);
xnor U1323 (N_1323,In_734,In_43);
xor U1324 (N_1324,In_963,In_718);
nor U1325 (N_1325,In_379,In_755);
or U1326 (N_1326,In_415,In_66);
xor U1327 (N_1327,In_617,In_591);
or U1328 (N_1328,In_173,In_691);
or U1329 (N_1329,In_795,In_225);
xor U1330 (N_1330,In_205,In_7);
nor U1331 (N_1331,In_235,In_312);
and U1332 (N_1332,In_485,In_772);
and U1333 (N_1333,In_364,In_434);
and U1334 (N_1334,In_435,In_382);
and U1335 (N_1335,In_128,In_603);
or U1336 (N_1336,In_600,In_353);
or U1337 (N_1337,In_111,In_711);
nand U1338 (N_1338,In_216,In_585);
and U1339 (N_1339,In_593,In_411);
and U1340 (N_1340,In_896,In_964);
or U1341 (N_1341,In_365,In_567);
and U1342 (N_1342,In_721,In_973);
nand U1343 (N_1343,In_638,In_444);
nor U1344 (N_1344,In_825,In_601);
and U1345 (N_1345,In_12,In_600);
and U1346 (N_1346,In_993,In_815);
or U1347 (N_1347,In_319,In_228);
nand U1348 (N_1348,In_490,In_358);
and U1349 (N_1349,In_415,In_745);
or U1350 (N_1350,In_791,In_838);
nor U1351 (N_1351,In_182,In_200);
xor U1352 (N_1352,In_70,In_274);
nor U1353 (N_1353,In_630,In_409);
or U1354 (N_1354,In_995,In_616);
or U1355 (N_1355,In_54,In_17);
nand U1356 (N_1356,In_794,In_20);
xnor U1357 (N_1357,In_41,In_427);
nand U1358 (N_1358,In_487,In_636);
and U1359 (N_1359,In_75,In_431);
nor U1360 (N_1360,In_52,In_566);
and U1361 (N_1361,In_860,In_787);
xor U1362 (N_1362,In_423,In_883);
xnor U1363 (N_1363,In_758,In_763);
nand U1364 (N_1364,In_620,In_493);
nand U1365 (N_1365,In_917,In_787);
xnor U1366 (N_1366,In_321,In_87);
nand U1367 (N_1367,In_192,In_221);
nand U1368 (N_1368,In_458,In_225);
nor U1369 (N_1369,In_385,In_241);
nand U1370 (N_1370,In_635,In_805);
xnor U1371 (N_1371,In_481,In_626);
or U1372 (N_1372,In_169,In_870);
nand U1373 (N_1373,In_447,In_775);
and U1374 (N_1374,In_42,In_756);
nor U1375 (N_1375,In_267,In_2);
and U1376 (N_1376,In_295,In_306);
nand U1377 (N_1377,In_233,In_174);
nand U1378 (N_1378,In_886,In_144);
nand U1379 (N_1379,In_106,In_988);
nand U1380 (N_1380,In_877,In_779);
nor U1381 (N_1381,In_551,In_782);
nand U1382 (N_1382,In_822,In_323);
or U1383 (N_1383,In_601,In_659);
and U1384 (N_1384,In_155,In_59);
xnor U1385 (N_1385,In_917,In_797);
and U1386 (N_1386,In_216,In_877);
nor U1387 (N_1387,In_650,In_511);
nor U1388 (N_1388,In_397,In_148);
or U1389 (N_1389,In_124,In_839);
nor U1390 (N_1390,In_152,In_409);
and U1391 (N_1391,In_187,In_473);
nand U1392 (N_1392,In_907,In_343);
xor U1393 (N_1393,In_376,In_719);
xnor U1394 (N_1394,In_941,In_820);
or U1395 (N_1395,In_681,In_139);
nand U1396 (N_1396,In_175,In_542);
nor U1397 (N_1397,In_603,In_421);
nand U1398 (N_1398,In_618,In_888);
xor U1399 (N_1399,In_763,In_273);
nor U1400 (N_1400,In_391,In_756);
nand U1401 (N_1401,In_144,In_880);
nand U1402 (N_1402,In_178,In_22);
or U1403 (N_1403,In_69,In_426);
nand U1404 (N_1404,In_498,In_93);
and U1405 (N_1405,In_105,In_389);
nand U1406 (N_1406,In_174,In_563);
xnor U1407 (N_1407,In_912,In_708);
and U1408 (N_1408,In_392,In_492);
nand U1409 (N_1409,In_225,In_445);
xnor U1410 (N_1410,In_391,In_218);
nand U1411 (N_1411,In_152,In_407);
xor U1412 (N_1412,In_738,In_215);
nor U1413 (N_1413,In_47,In_911);
or U1414 (N_1414,In_375,In_100);
nand U1415 (N_1415,In_250,In_101);
xnor U1416 (N_1416,In_798,In_644);
or U1417 (N_1417,In_986,In_903);
nand U1418 (N_1418,In_763,In_617);
nor U1419 (N_1419,In_843,In_717);
nand U1420 (N_1420,In_44,In_441);
and U1421 (N_1421,In_697,In_889);
or U1422 (N_1422,In_442,In_236);
and U1423 (N_1423,In_886,In_154);
xnor U1424 (N_1424,In_798,In_741);
and U1425 (N_1425,In_387,In_519);
or U1426 (N_1426,In_353,In_722);
or U1427 (N_1427,In_871,In_78);
nor U1428 (N_1428,In_177,In_510);
and U1429 (N_1429,In_610,In_327);
nand U1430 (N_1430,In_47,In_927);
nand U1431 (N_1431,In_703,In_824);
or U1432 (N_1432,In_786,In_53);
nand U1433 (N_1433,In_905,In_401);
nor U1434 (N_1434,In_287,In_950);
xnor U1435 (N_1435,In_423,In_324);
nor U1436 (N_1436,In_480,In_325);
and U1437 (N_1437,In_857,In_732);
nand U1438 (N_1438,In_725,In_51);
xnor U1439 (N_1439,In_622,In_396);
nand U1440 (N_1440,In_615,In_201);
nand U1441 (N_1441,In_635,In_875);
nand U1442 (N_1442,In_609,In_119);
nor U1443 (N_1443,In_793,In_891);
and U1444 (N_1444,In_81,In_846);
xor U1445 (N_1445,In_696,In_947);
nand U1446 (N_1446,In_359,In_744);
nor U1447 (N_1447,In_667,In_134);
xnor U1448 (N_1448,In_45,In_78);
nand U1449 (N_1449,In_764,In_524);
and U1450 (N_1450,In_327,In_681);
and U1451 (N_1451,In_340,In_41);
and U1452 (N_1452,In_828,In_731);
xor U1453 (N_1453,In_524,In_283);
xnor U1454 (N_1454,In_662,In_798);
nor U1455 (N_1455,In_266,In_865);
or U1456 (N_1456,In_669,In_339);
xor U1457 (N_1457,In_76,In_122);
or U1458 (N_1458,In_866,In_489);
nor U1459 (N_1459,In_745,In_874);
nor U1460 (N_1460,In_199,In_531);
or U1461 (N_1461,In_603,In_736);
and U1462 (N_1462,In_329,In_381);
xor U1463 (N_1463,In_702,In_135);
xnor U1464 (N_1464,In_172,In_119);
or U1465 (N_1465,In_539,In_930);
and U1466 (N_1466,In_970,In_775);
nand U1467 (N_1467,In_803,In_815);
or U1468 (N_1468,In_353,In_450);
and U1469 (N_1469,In_112,In_705);
xor U1470 (N_1470,In_222,In_2);
and U1471 (N_1471,In_117,In_921);
nor U1472 (N_1472,In_761,In_181);
nor U1473 (N_1473,In_382,In_733);
xor U1474 (N_1474,In_965,In_601);
xor U1475 (N_1475,In_429,In_866);
nand U1476 (N_1476,In_2,In_6);
xor U1477 (N_1477,In_592,In_78);
and U1478 (N_1478,In_139,In_658);
or U1479 (N_1479,In_745,In_524);
nand U1480 (N_1480,In_582,In_917);
or U1481 (N_1481,In_687,In_717);
and U1482 (N_1482,In_976,In_923);
and U1483 (N_1483,In_169,In_141);
or U1484 (N_1484,In_78,In_830);
xnor U1485 (N_1485,In_533,In_91);
xor U1486 (N_1486,In_260,In_611);
nand U1487 (N_1487,In_657,In_460);
xnor U1488 (N_1488,In_303,In_8);
and U1489 (N_1489,In_697,In_257);
nand U1490 (N_1490,In_744,In_692);
and U1491 (N_1491,In_27,In_453);
nand U1492 (N_1492,In_286,In_557);
nand U1493 (N_1493,In_867,In_44);
nand U1494 (N_1494,In_970,In_212);
nand U1495 (N_1495,In_759,In_417);
or U1496 (N_1496,In_141,In_625);
nor U1497 (N_1497,In_366,In_936);
nand U1498 (N_1498,In_511,In_101);
and U1499 (N_1499,In_424,In_804);
or U1500 (N_1500,In_227,In_579);
nand U1501 (N_1501,In_417,In_99);
xnor U1502 (N_1502,In_133,In_937);
xor U1503 (N_1503,In_423,In_451);
xnor U1504 (N_1504,In_399,In_403);
or U1505 (N_1505,In_578,In_710);
and U1506 (N_1506,In_693,In_101);
and U1507 (N_1507,In_757,In_289);
nor U1508 (N_1508,In_299,In_711);
xnor U1509 (N_1509,In_414,In_39);
xor U1510 (N_1510,In_434,In_776);
nand U1511 (N_1511,In_540,In_967);
xor U1512 (N_1512,In_468,In_991);
and U1513 (N_1513,In_554,In_815);
or U1514 (N_1514,In_750,In_495);
and U1515 (N_1515,In_62,In_969);
nand U1516 (N_1516,In_206,In_462);
and U1517 (N_1517,In_52,In_140);
nor U1518 (N_1518,In_949,In_729);
and U1519 (N_1519,In_728,In_592);
xnor U1520 (N_1520,In_349,In_558);
or U1521 (N_1521,In_837,In_981);
xnor U1522 (N_1522,In_521,In_534);
nor U1523 (N_1523,In_137,In_752);
or U1524 (N_1524,In_868,In_491);
or U1525 (N_1525,In_812,In_791);
xor U1526 (N_1526,In_442,In_48);
xor U1527 (N_1527,In_603,In_255);
and U1528 (N_1528,In_62,In_455);
or U1529 (N_1529,In_643,In_110);
or U1530 (N_1530,In_512,In_353);
xor U1531 (N_1531,In_252,In_919);
xor U1532 (N_1532,In_906,In_512);
nor U1533 (N_1533,In_433,In_929);
or U1534 (N_1534,In_161,In_132);
xnor U1535 (N_1535,In_442,In_75);
nor U1536 (N_1536,In_329,In_194);
xor U1537 (N_1537,In_282,In_480);
and U1538 (N_1538,In_791,In_256);
or U1539 (N_1539,In_247,In_210);
nand U1540 (N_1540,In_598,In_44);
nand U1541 (N_1541,In_849,In_953);
nand U1542 (N_1542,In_162,In_850);
nand U1543 (N_1543,In_672,In_523);
and U1544 (N_1544,In_297,In_528);
and U1545 (N_1545,In_573,In_287);
xnor U1546 (N_1546,In_764,In_302);
xor U1547 (N_1547,In_618,In_368);
xor U1548 (N_1548,In_584,In_520);
nand U1549 (N_1549,In_263,In_768);
nand U1550 (N_1550,In_566,In_961);
xnor U1551 (N_1551,In_477,In_413);
and U1552 (N_1552,In_353,In_565);
nor U1553 (N_1553,In_761,In_865);
nor U1554 (N_1554,In_491,In_938);
nor U1555 (N_1555,In_595,In_524);
nand U1556 (N_1556,In_596,In_259);
nor U1557 (N_1557,In_69,In_239);
nand U1558 (N_1558,In_217,In_239);
nand U1559 (N_1559,In_469,In_130);
or U1560 (N_1560,In_364,In_853);
nor U1561 (N_1561,In_326,In_539);
xor U1562 (N_1562,In_886,In_710);
nand U1563 (N_1563,In_268,In_42);
and U1564 (N_1564,In_128,In_681);
or U1565 (N_1565,In_985,In_122);
nand U1566 (N_1566,In_308,In_852);
nand U1567 (N_1567,In_438,In_372);
nand U1568 (N_1568,In_874,In_977);
nand U1569 (N_1569,In_428,In_333);
or U1570 (N_1570,In_864,In_276);
xor U1571 (N_1571,In_804,In_130);
nor U1572 (N_1572,In_577,In_75);
nor U1573 (N_1573,In_546,In_173);
and U1574 (N_1574,In_796,In_605);
xor U1575 (N_1575,In_587,In_551);
or U1576 (N_1576,In_823,In_937);
xor U1577 (N_1577,In_516,In_84);
xor U1578 (N_1578,In_605,In_570);
nand U1579 (N_1579,In_726,In_618);
nand U1580 (N_1580,In_153,In_272);
or U1581 (N_1581,In_934,In_221);
nor U1582 (N_1582,In_729,In_901);
and U1583 (N_1583,In_568,In_595);
nor U1584 (N_1584,In_309,In_730);
and U1585 (N_1585,In_740,In_985);
xor U1586 (N_1586,In_769,In_767);
nand U1587 (N_1587,In_291,In_227);
nor U1588 (N_1588,In_790,In_461);
nor U1589 (N_1589,In_36,In_922);
nor U1590 (N_1590,In_499,In_398);
nor U1591 (N_1591,In_82,In_809);
or U1592 (N_1592,In_891,In_355);
nor U1593 (N_1593,In_187,In_808);
xor U1594 (N_1594,In_868,In_554);
xor U1595 (N_1595,In_299,In_378);
and U1596 (N_1596,In_310,In_402);
nor U1597 (N_1597,In_725,In_352);
or U1598 (N_1598,In_768,In_227);
or U1599 (N_1599,In_547,In_275);
xnor U1600 (N_1600,In_193,In_974);
and U1601 (N_1601,In_281,In_782);
nand U1602 (N_1602,In_608,In_476);
nand U1603 (N_1603,In_140,In_325);
or U1604 (N_1604,In_435,In_530);
or U1605 (N_1605,In_716,In_28);
or U1606 (N_1606,In_181,In_270);
nand U1607 (N_1607,In_995,In_615);
xor U1608 (N_1608,In_348,In_195);
and U1609 (N_1609,In_526,In_290);
nor U1610 (N_1610,In_139,In_765);
or U1611 (N_1611,In_121,In_921);
xor U1612 (N_1612,In_638,In_82);
xor U1613 (N_1613,In_615,In_217);
xnor U1614 (N_1614,In_659,In_245);
nor U1615 (N_1615,In_975,In_427);
xnor U1616 (N_1616,In_226,In_917);
nand U1617 (N_1617,In_32,In_563);
xnor U1618 (N_1618,In_511,In_941);
and U1619 (N_1619,In_804,In_761);
nand U1620 (N_1620,In_312,In_87);
nor U1621 (N_1621,In_141,In_1);
xnor U1622 (N_1622,In_549,In_983);
xor U1623 (N_1623,In_349,In_900);
and U1624 (N_1624,In_499,In_620);
nor U1625 (N_1625,In_162,In_297);
and U1626 (N_1626,In_465,In_451);
or U1627 (N_1627,In_353,In_465);
and U1628 (N_1628,In_996,In_601);
xor U1629 (N_1629,In_598,In_401);
nand U1630 (N_1630,In_74,In_822);
or U1631 (N_1631,In_602,In_114);
xnor U1632 (N_1632,In_907,In_673);
xor U1633 (N_1633,In_972,In_297);
nand U1634 (N_1634,In_905,In_847);
or U1635 (N_1635,In_331,In_898);
xnor U1636 (N_1636,In_537,In_602);
xnor U1637 (N_1637,In_167,In_83);
and U1638 (N_1638,In_580,In_659);
nand U1639 (N_1639,In_425,In_734);
xnor U1640 (N_1640,In_211,In_865);
and U1641 (N_1641,In_543,In_755);
xnor U1642 (N_1642,In_322,In_946);
or U1643 (N_1643,In_851,In_245);
or U1644 (N_1644,In_765,In_279);
nand U1645 (N_1645,In_166,In_382);
or U1646 (N_1646,In_827,In_344);
and U1647 (N_1647,In_580,In_203);
or U1648 (N_1648,In_208,In_854);
or U1649 (N_1649,In_264,In_599);
nand U1650 (N_1650,In_967,In_528);
nor U1651 (N_1651,In_446,In_245);
or U1652 (N_1652,In_251,In_867);
xor U1653 (N_1653,In_674,In_350);
or U1654 (N_1654,In_10,In_426);
or U1655 (N_1655,In_767,In_836);
or U1656 (N_1656,In_915,In_722);
xnor U1657 (N_1657,In_159,In_266);
or U1658 (N_1658,In_299,In_79);
nor U1659 (N_1659,In_311,In_822);
nor U1660 (N_1660,In_259,In_874);
and U1661 (N_1661,In_978,In_8);
xor U1662 (N_1662,In_959,In_441);
or U1663 (N_1663,In_392,In_473);
nand U1664 (N_1664,In_242,In_290);
nand U1665 (N_1665,In_395,In_170);
xor U1666 (N_1666,In_851,In_901);
nor U1667 (N_1667,In_903,In_442);
or U1668 (N_1668,In_726,In_643);
nor U1669 (N_1669,In_61,In_223);
nor U1670 (N_1670,In_423,In_409);
nand U1671 (N_1671,In_757,In_8);
nor U1672 (N_1672,In_873,In_344);
xnor U1673 (N_1673,In_337,In_738);
or U1674 (N_1674,In_148,In_204);
nor U1675 (N_1675,In_720,In_943);
and U1676 (N_1676,In_642,In_132);
nor U1677 (N_1677,In_755,In_539);
or U1678 (N_1678,In_273,In_127);
or U1679 (N_1679,In_618,In_801);
nor U1680 (N_1680,In_894,In_854);
nor U1681 (N_1681,In_162,In_101);
or U1682 (N_1682,In_453,In_972);
xnor U1683 (N_1683,In_549,In_146);
nand U1684 (N_1684,In_817,In_413);
xor U1685 (N_1685,In_128,In_731);
nand U1686 (N_1686,In_895,In_485);
xor U1687 (N_1687,In_476,In_743);
or U1688 (N_1688,In_645,In_295);
xnor U1689 (N_1689,In_572,In_52);
nand U1690 (N_1690,In_825,In_838);
nand U1691 (N_1691,In_508,In_569);
nor U1692 (N_1692,In_31,In_297);
and U1693 (N_1693,In_271,In_529);
or U1694 (N_1694,In_129,In_285);
and U1695 (N_1695,In_793,In_826);
xnor U1696 (N_1696,In_544,In_85);
and U1697 (N_1697,In_813,In_953);
xor U1698 (N_1698,In_130,In_742);
or U1699 (N_1699,In_369,In_363);
and U1700 (N_1700,In_156,In_966);
nand U1701 (N_1701,In_608,In_590);
xor U1702 (N_1702,In_313,In_491);
and U1703 (N_1703,In_349,In_134);
nor U1704 (N_1704,In_183,In_392);
or U1705 (N_1705,In_968,In_544);
nor U1706 (N_1706,In_870,In_427);
nand U1707 (N_1707,In_105,In_79);
and U1708 (N_1708,In_706,In_301);
or U1709 (N_1709,In_198,In_452);
nor U1710 (N_1710,In_413,In_516);
xor U1711 (N_1711,In_903,In_392);
or U1712 (N_1712,In_477,In_205);
xor U1713 (N_1713,In_857,In_253);
or U1714 (N_1714,In_414,In_134);
nor U1715 (N_1715,In_548,In_593);
xor U1716 (N_1716,In_954,In_786);
and U1717 (N_1717,In_649,In_943);
nand U1718 (N_1718,In_948,In_84);
nand U1719 (N_1719,In_429,In_333);
nor U1720 (N_1720,In_779,In_412);
nand U1721 (N_1721,In_45,In_36);
and U1722 (N_1722,In_593,In_684);
nor U1723 (N_1723,In_933,In_212);
nor U1724 (N_1724,In_907,In_601);
xnor U1725 (N_1725,In_948,In_218);
xor U1726 (N_1726,In_582,In_699);
and U1727 (N_1727,In_92,In_753);
nand U1728 (N_1728,In_895,In_417);
and U1729 (N_1729,In_580,In_126);
and U1730 (N_1730,In_458,In_349);
and U1731 (N_1731,In_565,In_384);
or U1732 (N_1732,In_37,In_728);
and U1733 (N_1733,In_310,In_132);
xnor U1734 (N_1734,In_537,In_187);
and U1735 (N_1735,In_820,In_760);
xnor U1736 (N_1736,In_377,In_216);
and U1737 (N_1737,In_855,In_874);
nand U1738 (N_1738,In_496,In_494);
or U1739 (N_1739,In_106,In_246);
nor U1740 (N_1740,In_682,In_914);
or U1741 (N_1741,In_317,In_698);
or U1742 (N_1742,In_566,In_591);
nand U1743 (N_1743,In_365,In_293);
nor U1744 (N_1744,In_732,In_21);
and U1745 (N_1745,In_459,In_675);
nor U1746 (N_1746,In_216,In_596);
xor U1747 (N_1747,In_934,In_198);
or U1748 (N_1748,In_61,In_879);
or U1749 (N_1749,In_25,In_239);
nand U1750 (N_1750,In_918,In_146);
nor U1751 (N_1751,In_602,In_233);
or U1752 (N_1752,In_778,In_774);
xnor U1753 (N_1753,In_764,In_229);
or U1754 (N_1754,In_939,In_961);
nor U1755 (N_1755,In_779,In_631);
and U1756 (N_1756,In_943,In_506);
nand U1757 (N_1757,In_206,In_954);
or U1758 (N_1758,In_482,In_371);
nand U1759 (N_1759,In_497,In_128);
and U1760 (N_1760,In_749,In_77);
or U1761 (N_1761,In_152,In_185);
and U1762 (N_1762,In_345,In_439);
nand U1763 (N_1763,In_325,In_331);
and U1764 (N_1764,In_440,In_836);
xnor U1765 (N_1765,In_398,In_514);
nand U1766 (N_1766,In_53,In_821);
or U1767 (N_1767,In_85,In_145);
and U1768 (N_1768,In_237,In_772);
xor U1769 (N_1769,In_965,In_827);
or U1770 (N_1770,In_12,In_26);
and U1771 (N_1771,In_106,In_12);
xor U1772 (N_1772,In_969,In_67);
or U1773 (N_1773,In_855,In_450);
nand U1774 (N_1774,In_508,In_732);
xor U1775 (N_1775,In_50,In_400);
nand U1776 (N_1776,In_773,In_637);
and U1777 (N_1777,In_995,In_729);
nand U1778 (N_1778,In_679,In_54);
or U1779 (N_1779,In_527,In_177);
xor U1780 (N_1780,In_875,In_237);
and U1781 (N_1781,In_380,In_337);
nor U1782 (N_1782,In_524,In_243);
and U1783 (N_1783,In_775,In_368);
or U1784 (N_1784,In_196,In_882);
xnor U1785 (N_1785,In_542,In_771);
nand U1786 (N_1786,In_34,In_599);
or U1787 (N_1787,In_835,In_876);
nor U1788 (N_1788,In_641,In_776);
and U1789 (N_1789,In_714,In_745);
xnor U1790 (N_1790,In_776,In_740);
nor U1791 (N_1791,In_955,In_523);
or U1792 (N_1792,In_535,In_139);
nand U1793 (N_1793,In_467,In_584);
nor U1794 (N_1794,In_388,In_805);
or U1795 (N_1795,In_358,In_29);
nand U1796 (N_1796,In_337,In_185);
nor U1797 (N_1797,In_514,In_110);
nand U1798 (N_1798,In_718,In_584);
nand U1799 (N_1799,In_177,In_388);
and U1800 (N_1800,In_557,In_278);
xor U1801 (N_1801,In_149,In_382);
and U1802 (N_1802,In_154,In_934);
and U1803 (N_1803,In_686,In_684);
and U1804 (N_1804,In_921,In_586);
or U1805 (N_1805,In_422,In_721);
nor U1806 (N_1806,In_495,In_147);
or U1807 (N_1807,In_869,In_602);
xnor U1808 (N_1808,In_455,In_125);
and U1809 (N_1809,In_923,In_234);
nand U1810 (N_1810,In_825,In_913);
nand U1811 (N_1811,In_631,In_193);
and U1812 (N_1812,In_65,In_325);
and U1813 (N_1813,In_486,In_388);
xor U1814 (N_1814,In_967,In_513);
xor U1815 (N_1815,In_401,In_701);
nand U1816 (N_1816,In_426,In_373);
nand U1817 (N_1817,In_647,In_883);
nor U1818 (N_1818,In_698,In_560);
nand U1819 (N_1819,In_632,In_909);
and U1820 (N_1820,In_446,In_702);
and U1821 (N_1821,In_846,In_793);
or U1822 (N_1822,In_114,In_832);
or U1823 (N_1823,In_563,In_661);
and U1824 (N_1824,In_728,In_700);
nand U1825 (N_1825,In_717,In_810);
and U1826 (N_1826,In_419,In_98);
and U1827 (N_1827,In_656,In_733);
xnor U1828 (N_1828,In_77,In_851);
xnor U1829 (N_1829,In_591,In_595);
and U1830 (N_1830,In_271,In_651);
nand U1831 (N_1831,In_567,In_700);
xnor U1832 (N_1832,In_840,In_140);
and U1833 (N_1833,In_883,In_728);
nor U1834 (N_1834,In_660,In_269);
nand U1835 (N_1835,In_661,In_102);
xor U1836 (N_1836,In_512,In_18);
or U1837 (N_1837,In_519,In_306);
xor U1838 (N_1838,In_89,In_153);
xor U1839 (N_1839,In_21,In_127);
xor U1840 (N_1840,In_493,In_763);
xor U1841 (N_1841,In_554,In_386);
nand U1842 (N_1842,In_95,In_901);
xor U1843 (N_1843,In_577,In_944);
and U1844 (N_1844,In_521,In_433);
xor U1845 (N_1845,In_770,In_287);
xnor U1846 (N_1846,In_336,In_211);
and U1847 (N_1847,In_198,In_356);
and U1848 (N_1848,In_693,In_956);
and U1849 (N_1849,In_384,In_329);
or U1850 (N_1850,In_402,In_155);
and U1851 (N_1851,In_277,In_71);
and U1852 (N_1852,In_164,In_805);
or U1853 (N_1853,In_3,In_503);
nand U1854 (N_1854,In_595,In_657);
and U1855 (N_1855,In_369,In_127);
or U1856 (N_1856,In_702,In_937);
and U1857 (N_1857,In_706,In_376);
or U1858 (N_1858,In_279,In_349);
nor U1859 (N_1859,In_688,In_29);
xnor U1860 (N_1860,In_457,In_533);
nand U1861 (N_1861,In_74,In_476);
xor U1862 (N_1862,In_241,In_706);
nand U1863 (N_1863,In_485,In_197);
xnor U1864 (N_1864,In_775,In_892);
nor U1865 (N_1865,In_986,In_553);
xor U1866 (N_1866,In_16,In_100);
nor U1867 (N_1867,In_802,In_974);
nand U1868 (N_1868,In_306,In_896);
nand U1869 (N_1869,In_387,In_132);
or U1870 (N_1870,In_169,In_518);
xnor U1871 (N_1871,In_478,In_143);
or U1872 (N_1872,In_746,In_138);
and U1873 (N_1873,In_99,In_342);
and U1874 (N_1874,In_919,In_945);
nor U1875 (N_1875,In_401,In_120);
and U1876 (N_1876,In_758,In_402);
nand U1877 (N_1877,In_458,In_512);
or U1878 (N_1878,In_166,In_539);
nor U1879 (N_1879,In_349,In_123);
and U1880 (N_1880,In_961,In_338);
and U1881 (N_1881,In_391,In_523);
nand U1882 (N_1882,In_441,In_455);
nand U1883 (N_1883,In_868,In_546);
or U1884 (N_1884,In_436,In_782);
and U1885 (N_1885,In_923,In_822);
and U1886 (N_1886,In_174,In_934);
or U1887 (N_1887,In_836,In_843);
xor U1888 (N_1888,In_416,In_289);
nand U1889 (N_1889,In_936,In_279);
and U1890 (N_1890,In_144,In_772);
nor U1891 (N_1891,In_835,In_129);
nand U1892 (N_1892,In_277,In_813);
or U1893 (N_1893,In_828,In_972);
xnor U1894 (N_1894,In_167,In_531);
and U1895 (N_1895,In_793,In_367);
or U1896 (N_1896,In_895,In_41);
or U1897 (N_1897,In_345,In_491);
or U1898 (N_1898,In_482,In_881);
or U1899 (N_1899,In_706,In_817);
nor U1900 (N_1900,In_523,In_977);
or U1901 (N_1901,In_365,In_39);
nand U1902 (N_1902,In_566,In_70);
or U1903 (N_1903,In_256,In_979);
or U1904 (N_1904,In_356,In_238);
or U1905 (N_1905,In_102,In_532);
or U1906 (N_1906,In_600,In_37);
xor U1907 (N_1907,In_204,In_744);
and U1908 (N_1908,In_306,In_390);
nand U1909 (N_1909,In_665,In_989);
or U1910 (N_1910,In_546,In_313);
and U1911 (N_1911,In_567,In_98);
nor U1912 (N_1912,In_247,In_232);
and U1913 (N_1913,In_105,In_49);
nand U1914 (N_1914,In_896,In_823);
and U1915 (N_1915,In_678,In_415);
xor U1916 (N_1916,In_98,In_924);
or U1917 (N_1917,In_511,In_574);
nor U1918 (N_1918,In_662,In_630);
or U1919 (N_1919,In_60,In_812);
and U1920 (N_1920,In_7,In_183);
nor U1921 (N_1921,In_316,In_486);
xnor U1922 (N_1922,In_826,In_665);
xor U1923 (N_1923,In_537,In_225);
and U1924 (N_1924,In_440,In_286);
and U1925 (N_1925,In_688,In_504);
nand U1926 (N_1926,In_801,In_415);
and U1927 (N_1927,In_746,In_489);
xor U1928 (N_1928,In_109,In_385);
and U1929 (N_1929,In_231,In_604);
xor U1930 (N_1930,In_558,In_65);
nand U1931 (N_1931,In_723,In_84);
or U1932 (N_1932,In_521,In_730);
nand U1933 (N_1933,In_354,In_288);
nor U1934 (N_1934,In_655,In_688);
xnor U1935 (N_1935,In_159,In_755);
and U1936 (N_1936,In_333,In_57);
xor U1937 (N_1937,In_121,In_368);
xnor U1938 (N_1938,In_657,In_849);
nor U1939 (N_1939,In_624,In_458);
and U1940 (N_1940,In_558,In_727);
nor U1941 (N_1941,In_702,In_16);
xor U1942 (N_1942,In_506,In_870);
xor U1943 (N_1943,In_126,In_103);
and U1944 (N_1944,In_775,In_382);
or U1945 (N_1945,In_22,In_638);
and U1946 (N_1946,In_834,In_284);
nand U1947 (N_1947,In_517,In_58);
nand U1948 (N_1948,In_330,In_97);
nand U1949 (N_1949,In_719,In_573);
nand U1950 (N_1950,In_216,In_83);
or U1951 (N_1951,In_374,In_116);
nor U1952 (N_1952,In_269,In_72);
and U1953 (N_1953,In_864,In_116);
or U1954 (N_1954,In_974,In_51);
xor U1955 (N_1955,In_135,In_407);
xor U1956 (N_1956,In_536,In_285);
nor U1957 (N_1957,In_339,In_100);
and U1958 (N_1958,In_176,In_817);
nor U1959 (N_1959,In_574,In_29);
or U1960 (N_1960,In_13,In_931);
xnor U1961 (N_1961,In_647,In_294);
and U1962 (N_1962,In_14,In_586);
and U1963 (N_1963,In_640,In_467);
nor U1964 (N_1964,In_747,In_353);
nor U1965 (N_1965,In_632,In_781);
xor U1966 (N_1966,In_762,In_746);
xnor U1967 (N_1967,In_898,In_68);
and U1968 (N_1968,In_277,In_914);
nor U1969 (N_1969,In_737,In_980);
and U1970 (N_1970,In_175,In_615);
nor U1971 (N_1971,In_928,In_85);
xor U1972 (N_1972,In_413,In_10);
nor U1973 (N_1973,In_117,In_291);
nand U1974 (N_1974,In_183,In_990);
nand U1975 (N_1975,In_490,In_718);
nor U1976 (N_1976,In_71,In_967);
nand U1977 (N_1977,In_493,In_226);
nand U1978 (N_1978,In_680,In_777);
or U1979 (N_1979,In_445,In_878);
nor U1980 (N_1980,In_329,In_404);
xnor U1981 (N_1981,In_876,In_160);
xnor U1982 (N_1982,In_899,In_256);
nor U1983 (N_1983,In_951,In_500);
and U1984 (N_1984,In_645,In_993);
or U1985 (N_1985,In_956,In_816);
and U1986 (N_1986,In_780,In_544);
or U1987 (N_1987,In_337,In_541);
nor U1988 (N_1988,In_292,In_443);
and U1989 (N_1989,In_927,In_637);
nand U1990 (N_1990,In_911,In_16);
nor U1991 (N_1991,In_868,In_664);
nand U1992 (N_1992,In_35,In_348);
nor U1993 (N_1993,In_653,In_133);
nor U1994 (N_1994,In_817,In_322);
and U1995 (N_1995,In_84,In_80);
xor U1996 (N_1996,In_477,In_95);
and U1997 (N_1997,In_951,In_568);
and U1998 (N_1998,In_103,In_381);
and U1999 (N_1999,In_840,In_478);
nand U2000 (N_2000,In_431,In_520);
or U2001 (N_2001,In_477,In_216);
nor U2002 (N_2002,In_793,In_94);
xor U2003 (N_2003,In_187,In_921);
nor U2004 (N_2004,In_538,In_380);
nor U2005 (N_2005,In_649,In_106);
nor U2006 (N_2006,In_867,In_806);
nor U2007 (N_2007,In_393,In_6);
or U2008 (N_2008,In_82,In_18);
nor U2009 (N_2009,In_41,In_827);
or U2010 (N_2010,In_658,In_609);
xnor U2011 (N_2011,In_278,In_420);
nor U2012 (N_2012,In_740,In_533);
nand U2013 (N_2013,In_694,In_590);
or U2014 (N_2014,In_653,In_589);
nor U2015 (N_2015,In_958,In_363);
xnor U2016 (N_2016,In_219,In_637);
or U2017 (N_2017,In_709,In_960);
nor U2018 (N_2018,In_295,In_979);
nor U2019 (N_2019,In_732,In_55);
nor U2020 (N_2020,In_147,In_583);
nand U2021 (N_2021,In_888,In_196);
and U2022 (N_2022,In_484,In_578);
nor U2023 (N_2023,In_413,In_900);
xnor U2024 (N_2024,In_856,In_101);
or U2025 (N_2025,In_394,In_65);
xnor U2026 (N_2026,In_720,In_80);
or U2027 (N_2027,In_279,In_477);
and U2028 (N_2028,In_749,In_501);
nand U2029 (N_2029,In_146,In_552);
nor U2030 (N_2030,In_633,In_64);
or U2031 (N_2031,In_703,In_575);
xnor U2032 (N_2032,In_433,In_887);
nand U2033 (N_2033,In_119,In_939);
or U2034 (N_2034,In_255,In_764);
xor U2035 (N_2035,In_938,In_894);
nor U2036 (N_2036,In_321,In_682);
or U2037 (N_2037,In_702,In_982);
nand U2038 (N_2038,In_236,In_842);
xor U2039 (N_2039,In_212,In_915);
or U2040 (N_2040,In_607,In_189);
nand U2041 (N_2041,In_914,In_209);
or U2042 (N_2042,In_746,In_636);
and U2043 (N_2043,In_532,In_409);
and U2044 (N_2044,In_442,In_766);
and U2045 (N_2045,In_171,In_410);
nand U2046 (N_2046,In_113,In_425);
or U2047 (N_2047,In_699,In_163);
nor U2048 (N_2048,In_254,In_335);
xor U2049 (N_2049,In_167,In_723);
nand U2050 (N_2050,In_301,In_594);
nor U2051 (N_2051,In_268,In_668);
nor U2052 (N_2052,In_463,In_315);
and U2053 (N_2053,In_563,In_51);
or U2054 (N_2054,In_631,In_121);
nand U2055 (N_2055,In_845,In_792);
and U2056 (N_2056,In_429,In_950);
and U2057 (N_2057,In_998,In_552);
xor U2058 (N_2058,In_65,In_68);
nand U2059 (N_2059,In_50,In_220);
nand U2060 (N_2060,In_500,In_331);
and U2061 (N_2061,In_564,In_710);
xnor U2062 (N_2062,In_301,In_307);
xnor U2063 (N_2063,In_751,In_122);
nand U2064 (N_2064,In_253,In_153);
and U2065 (N_2065,In_352,In_718);
nor U2066 (N_2066,In_257,In_399);
or U2067 (N_2067,In_53,In_16);
nand U2068 (N_2068,In_707,In_227);
xnor U2069 (N_2069,In_583,In_885);
and U2070 (N_2070,In_677,In_115);
and U2071 (N_2071,In_111,In_604);
and U2072 (N_2072,In_294,In_709);
nor U2073 (N_2073,In_323,In_265);
nand U2074 (N_2074,In_369,In_114);
nor U2075 (N_2075,In_789,In_961);
or U2076 (N_2076,In_374,In_993);
xor U2077 (N_2077,In_760,In_187);
nor U2078 (N_2078,In_477,In_2);
xnor U2079 (N_2079,In_875,In_730);
xnor U2080 (N_2080,In_851,In_144);
nand U2081 (N_2081,In_49,In_210);
nand U2082 (N_2082,In_313,In_459);
nand U2083 (N_2083,In_917,In_368);
nand U2084 (N_2084,In_564,In_840);
or U2085 (N_2085,In_115,In_158);
and U2086 (N_2086,In_665,In_269);
or U2087 (N_2087,In_86,In_641);
xor U2088 (N_2088,In_740,In_118);
xor U2089 (N_2089,In_588,In_861);
xor U2090 (N_2090,In_940,In_576);
nor U2091 (N_2091,In_564,In_997);
and U2092 (N_2092,In_904,In_146);
nor U2093 (N_2093,In_571,In_61);
xor U2094 (N_2094,In_409,In_468);
or U2095 (N_2095,In_712,In_293);
or U2096 (N_2096,In_373,In_264);
or U2097 (N_2097,In_738,In_844);
xnor U2098 (N_2098,In_6,In_3);
nand U2099 (N_2099,In_803,In_784);
and U2100 (N_2100,In_739,In_614);
or U2101 (N_2101,In_730,In_175);
xor U2102 (N_2102,In_675,In_627);
and U2103 (N_2103,In_396,In_934);
or U2104 (N_2104,In_946,In_407);
xnor U2105 (N_2105,In_389,In_572);
xnor U2106 (N_2106,In_904,In_806);
xor U2107 (N_2107,In_868,In_852);
or U2108 (N_2108,In_6,In_260);
xor U2109 (N_2109,In_133,In_442);
or U2110 (N_2110,In_783,In_46);
xnor U2111 (N_2111,In_293,In_952);
xnor U2112 (N_2112,In_165,In_528);
nor U2113 (N_2113,In_900,In_419);
and U2114 (N_2114,In_516,In_499);
xor U2115 (N_2115,In_269,In_937);
and U2116 (N_2116,In_997,In_737);
xor U2117 (N_2117,In_759,In_897);
nor U2118 (N_2118,In_358,In_288);
xnor U2119 (N_2119,In_429,In_731);
nor U2120 (N_2120,In_422,In_446);
xnor U2121 (N_2121,In_436,In_290);
xnor U2122 (N_2122,In_593,In_581);
or U2123 (N_2123,In_789,In_942);
or U2124 (N_2124,In_135,In_80);
nor U2125 (N_2125,In_530,In_230);
and U2126 (N_2126,In_529,In_506);
or U2127 (N_2127,In_159,In_300);
or U2128 (N_2128,In_688,In_25);
and U2129 (N_2129,In_989,In_904);
xnor U2130 (N_2130,In_329,In_264);
and U2131 (N_2131,In_744,In_806);
xor U2132 (N_2132,In_637,In_321);
nor U2133 (N_2133,In_621,In_707);
nand U2134 (N_2134,In_551,In_969);
xnor U2135 (N_2135,In_764,In_237);
or U2136 (N_2136,In_815,In_421);
nand U2137 (N_2137,In_697,In_781);
and U2138 (N_2138,In_1,In_78);
xor U2139 (N_2139,In_842,In_175);
nand U2140 (N_2140,In_572,In_150);
and U2141 (N_2141,In_981,In_151);
nand U2142 (N_2142,In_889,In_385);
or U2143 (N_2143,In_379,In_461);
nor U2144 (N_2144,In_842,In_198);
nand U2145 (N_2145,In_704,In_349);
or U2146 (N_2146,In_963,In_917);
or U2147 (N_2147,In_545,In_729);
and U2148 (N_2148,In_817,In_964);
nand U2149 (N_2149,In_758,In_345);
or U2150 (N_2150,In_15,In_88);
nand U2151 (N_2151,In_993,In_187);
or U2152 (N_2152,In_971,In_977);
nand U2153 (N_2153,In_466,In_797);
nor U2154 (N_2154,In_560,In_225);
nand U2155 (N_2155,In_935,In_270);
or U2156 (N_2156,In_326,In_41);
and U2157 (N_2157,In_953,In_900);
nand U2158 (N_2158,In_735,In_713);
xor U2159 (N_2159,In_934,In_153);
and U2160 (N_2160,In_205,In_977);
and U2161 (N_2161,In_676,In_683);
xnor U2162 (N_2162,In_428,In_931);
nor U2163 (N_2163,In_654,In_154);
and U2164 (N_2164,In_185,In_585);
or U2165 (N_2165,In_65,In_748);
xor U2166 (N_2166,In_746,In_156);
and U2167 (N_2167,In_721,In_128);
nand U2168 (N_2168,In_351,In_28);
or U2169 (N_2169,In_470,In_728);
nand U2170 (N_2170,In_536,In_801);
and U2171 (N_2171,In_466,In_109);
and U2172 (N_2172,In_953,In_219);
xor U2173 (N_2173,In_516,In_547);
nor U2174 (N_2174,In_949,In_736);
nor U2175 (N_2175,In_276,In_53);
or U2176 (N_2176,In_201,In_981);
or U2177 (N_2177,In_942,In_493);
nand U2178 (N_2178,In_354,In_151);
and U2179 (N_2179,In_558,In_472);
and U2180 (N_2180,In_925,In_923);
and U2181 (N_2181,In_912,In_539);
nand U2182 (N_2182,In_272,In_393);
nor U2183 (N_2183,In_920,In_609);
nor U2184 (N_2184,In_971,In_767);
nor U2185 (N_2185,In_996,In_949);
nand U2186 (N_2186,In_938,In_536);
xnor U2187 (N_2187,In_692,In_239);
xnor U2188 (N_2188,In_457,In_50);
nand U2189 (N_2189,In_195,In_47);
nor U2190 (N_2190,In_852,In_492);
or U2191 (N_2191,In_252,In_346);
or U2192 (N_2192,In_609,In_42);
or U2193 (N_2193,In_284,In_489);
xor U2194 (N_2194,In_800,In_44);
nor U2195 (N_2195,In_289,In_241);
nand U2196 (N_2196,In_355,In_414);
or U2197 (N_2197,In_642,In_122);
nor U2198 (N_2198,In_435,In_32);
xnor U2199 (N_2199,In_981,In_639);
nand U2200 (N_2200,In_944,In_280);
nor U2201 (N_2201,In_618,In_796);
and U2202 (N_2202,In_369,In_15);
nor U2203 (N_2203,In_242,In_521);
and U2204 (N_2204,In_339,In_928);
nand U2205 (N_2205,In_602,In_743);
xnor U2206 (N_2206,In_958,In_495);
or U2207 (N_2207,In_640,In_534);
or U2208 (N_2208,In_977,In_800);
nor U2209 (N_2209,In_23,In_390);
xnor U2210 (N_2210,In_848,In_546);
xnor U2211 (N_2211,In_589,In_367);
or U2212 (N_2212,In_253,In_381);
nand U2213 (N_2213,In_492,In_171);
nor U2214 (N_2214,In_304,In_736);
and U2215 (N_2215,In_6,In_597);
nor U2216 (N_2216,In_997,In_13);
or U2217 (N_2217,In_450,In_612);
nand U2218 (N_2218,In_333,In_99);
nand U2219 (N_2219,In_796,In_958);
xor U2220 (N_2220,In_842,In_978);
nor U2221 (N_2221,In_548,In_312);
or U2222 (N_2222,In_178,In_725);
and U2223 (N_2223,In_349,In_845);
nand U2224 (N_2224,In_537,In_638);
xor U2225 (N_2225,In_560,In_242);
nor U2226 (N_2226,In_677,In_980);
nor U2227 (N_2227,In_957,In_576);
xnor U2228 (N_2228,In_272,In_518);
xnor U2229 (N_2229,In_698,In_253);
and U2230 (N_2230,In_802,In_777);
nand U2231 (N_2231,In_420,In_337);
and U2232 (N_2232,In_362,In_733);
and U2233 (N_2233,In_795,In_720);
or U2234 (N_2234,In_706,In_815);
or U2235 (N_2235,In_703,In_589);
or U2236 (N_2236,In_745,In_122);
and U2237 (N_2237,In_458,In_851);
nor U2238 (N_2238,In_19,In_101);
or U2239 (N_2239,In_236,In_824);
xnor U2240 (N_2240,In_377,In_217);
xor U2241 (N_2241,In_481,In_435);
nand U2242 (N_2242,In_6,In_335);
nand U2243 (N_2243,In_376,In_672);
and U2244 (N_2244,In_227,In_288);
xnor U2245 (N_2245,In_624,In_126);
nand U2246 (N_2246,In_453,In_778);
nand U2247 (N_2247,In_406,In_590);
nand U2248 (N_2248,In_684,In_467);
nand U2249 (N_2249,In_157,In_97);
nor U2250 (N_2250,In_206,In_692);
nand U2251 (N_2251,In_938,In_461);
or U2252 (N_2252,In_973,In_576);
nand U2253 (N_2253,In_271,In_760);
and U2254 (N_2254,In_318,In_918);
and U2255 (N_2255,In_38,In_909);
xnor U2256 (N_2256,In_655,In_905);
nand U2257 (N_2257,In_717,In_214);
or U2258 (N_2258,In_421,In_401);
xor U2259 (N_2259,In_591,In_792);
xor U2260 (N_2260,In_364,In_441);
nor U2261 (N_2261,In_277,In_185);
nand U2262 (N_2262,In_666,In_774);
nand U2263 (N_2263,In_868,In_571);
and U2264 (N_2264,In_59,In_944);
xor U2265 (N_2265,In_939,In_183);
and U2266 (N_2266,In_829,In_290);
and U2267 (N_2267,In_357,In_837);
nand U2268 (N_2268,In_462,In_389);
and U2269 (N_2269,In_839,In_363);
or U2270 (N_2270,In_338,In_784);
nand U2271 (N_2271,In_393,In_283);
or U2272 (N_2272,In_124,In_743);
nor U2273 (N_2273,In_211,In_338);
or U2274 (N_2274,In_897,In_183);
nor U2275 (N_2275,In_424,In_743);
or U2276 (N_2276,In_973,In_645);
xnor U2277 (N_2277,In_537,In_965);
nor U2278 (N_2278,In_242,In_892);
nor U2279 (N_2279,In_14,In_914);
and U2280 (N_2280,In_515,In_734);
nor U2281 (N_2281,In_213,In_732);
or U2282 (N_2282,In_971,In_216);
nand U2283 (N_2283,In_925,In_441);
xnor U2284 (N_2284,In_248,In_609);
and U2285 (N_2285,In_143,In_383);
xor U2286 (N_2286,In_834,In_55);
xnor U2287 (N_2287,In_952,In_931);
or U2288 (N_2288,In_874,In_827);
or U2289 (N_2289,In_754,In_725);
xor U2290 (N_2290,In_318,In_196);
nand U2291 (N_2291,In_603,In_47);
or U2292 (N_2292,In_331,In_76);
nor U2293 (N_2293,In_785,In_981);
xnor U2294 (N_2294,In_438,In_330);
and U2295 (N_2295,In_916,In_794);
nor U2296 (N_2296,In_326,In_504);
nor U2297 (N_2297,In_158,In_544);
xor U2298 (N_2298,In_756,In_802);
nor U2299 (N_2299,In_587,In_511);
xor U2300 (N_2300,In_364,In_589);
nand U2301 (N_2301,In_85,In_951);
nand U2302 (N_2302,In_767,In_642);
nand U2303 (N_2303,In_570,In_863);
or U2304 (N_2304,In_241,In_685);
xor U2305 (N_2305,In_964,In_556);
and U2306 (N_2306,In_424,In_526);
and U2307 (N_2307,In_883,In_556);
or U2308 (N_2308,In_660,In_873);
nand U2309 (N_2309,In_820,In_164);
nand U2310 (N_2310,In_325,In_953);
and U2311 (N_2311,In_282,In_679);
nand U2312 (N_2312,In_665,In_956);
nor U2313 (N_2313,In_84,In_564);
nand U2314 (N_2314,In_84,In_734);
nand U2315 (N_2315,In_700,In_568);
nor U2316 (N_2316,In_620,In_730);
or U2317 (N_2317,In_423,In_190);
nor U2318 (N_2318,In_650,In_851);
xor U2319 (N_2319,In_903,In_418);
or U2320 (N_2320,In_258,In_383);
or U2321 (N_2321,In_281,In_369);
xnor U2322 (N_2322,In_317,In_717);
and U2323 (N_2323,In_955,In_262);
nor U2324 (N_2324,In_448,In_854);
nand U2325 (N_2325,In_395,In_690);
xor U2326 (N_2326,In_392,In_32);
xnor U2327 (N_2327,In_356,In_740);
nor U2328 (N_2328,In_234,In_314);
nor U2329 (N_2329,In_851,In_47);
nor U2330 (N_2330,In_174,In_922);
nand U2331 (N_2331,In_566,In_190);
or U2332 (N_2332,In_847,In_308);
and U2333 (N_2333,In_150,In_971);
nor U2334 (N_2334,In_145,In_763);
xor U2335 (N_2335,In_894,In_317);
or U2336 (N_2336,In_631,In_840);
or U2337 (N_2337,In_55,In_795);
nor U2338 (N_2338,In_333,In_364);
and U2339 (N_2339,In_631,In_273);
nand U2340 (N_2340,In_396,In_441);
or U2341 (N_2341,In_118,In_162);
nand U2342 (N_2342,In_322,In_194);
nand U2343 (N_2343,In_625,In_324);
xor U2344 (N_2344,In_641,In_581);
nand U2345 (N_2345,In_8,In_191);
nor U2346 (N_2346,In_504,In_185);
nand U2347 (N_2347,In_739,In_451);
nand U2348 (N_2348,In_340,In_80);
xnor U2349 (N_2349,In_639,In_731);
nor U2350 (N_2350,In_604,In_7);
nor U2351 (N_2351,In_479,In_394);
nor U2352 (N_2352,In_452,In_20);
xnor U2353 (N_2353,In_461,In_188);
xnor U2354 (N_2354,In_835,In_626);
or U2355 (N_2355,In_542,In_830);
and U2356 (N_2356,In_784,In_459);
nor U2357 (N_2357,In_556,In_289);
and U2358 (N_2358,In_734,In_217);
and U2359 (N_2359,In_296,In_234);
nand U2360 (N_2360,In_147,In_507);
xnor U2361 (N_2361,In_353,In_161);
or U2362 (N_2362,In_810,In_880);
and U2363 (N_2363,In_24,In_342);
or U2364 (N_2364,In_688,In_825);
or U2365 (N_2365,In_49,In_918);
xnor U2366 (N_2366,In_956,In_59);
or U2367 (N_2367,In_560,In_777);
nand U2368 (N_2368,In_942,In_603);
xnor U2369 (N_2369,In_210,In_725);
nor U2370 (N_2370,In_531,In_447);
xor U2371 (N_2371,In_75,In_564);
or U2372 (N_2372,In_930,In_899);
xnor U2373 (N_2373,In_760,In_609);
xnor U2374 (N_2374,In_559,In_335);
or U2375 (N_2375,In_327,In_449);
nand U2376 (N_2376,In_315,In_619);
xnor U2377 (N_2377,In_377,In_252);
or U2378 (N_2378,In_614,In_878);
nand U2379 (N_2379,In_997,In_141);
and U2380 (N_2380,In_288,In_948);
nor U2381 (N_2381,In_714,In_428);
and U2382 (N_2382,In_712,In_854);
or U2383 (N_2383,In_594,In_473);
and U2384 (N_2384,In_884,In_52);
and U2385 (N_2385,In_405,In_769);
nor U2386 (N_2386,In_349,In_711);
nand U2387 (N_2387,In_442,In_105);
nand U2388 (N_2388,In_892,In_783);
nand U2389 (N_2389,In_446,In_23);
nor U2390 (N_2390,In_328,In_602);
xor U2391 (N_2391,In_13,In_562);
nand U2392 (N_2392,In_930,In_168);
or U2393 (N_2393,In_49,In_196);
xor U2394 (N_2394,In_556,In_363);
nand U2395 (N_2395,In_758,In_465);
or U2396 (N_2396,In_455,In_236);
and U2397 (N_2397,In_7,In_864);
nor U2398 (N_2398,In_469,In_273);
nand U2399 (N_2399,In_455,In_422);
nand U2400 (N_2400,In_194,In_833);
and U2401 (N_2401,In_561,In_980);
nand U2402 (N_2402,In_689,In_545);
or U2403 (N_2403,In_125,In_866);
xor U2404 (N_2404,In_970,In_677);
nand U2405 (N_2405,In_566,In_838);
nor U2406 (N_2406,In_838,In_507);
nand U2407 (N_2407,In_141,In_2);
nor U2408 (N_2408,In_891,In_992);
or U2409 (N_2409,In_361,In_508);
or U2410 (N_2410,In_498,In_0);
xnor U2411 (N_2411,In_91,In_983);
nor U2412 (N_2412,In_823,In_153);
and U2413 (N_2413,In_383,In_872);
nor U2414 (N_2414,In_545,In_769);
and U2415 (N_2415,In_763,In_813);
and U2416 (N_2416,In_43,In_871);
nor U2417 (N_2417,In_232,In_357);
nor U2418 (N_2418,In_491,In_310);
xnor U2419 (N_2419,In_399,In_150);
and U2420 (N_2420,In_780,In_734);
nor U2421 (N_2421,In_333,In_975);
nor U2422 (N_2422,In_164,In_545);
nor U2423 (N_2423,In_504,In_888);
or U2424 (N_2424,In_943,In_919);
nor U2425 (N_2425,In_240,In_528);
xnor U2426 (N_2426,In_257,In_91);
nand U2427 (N_2427,In_381,In_896);
nand U2428 (N_2428,In_942,In_762);
nand U2429 (N_2429,In_669,In_906);
and U2430 (N_2430,In_139,In_721);
nand U2431 (N_2431,In_445,In_221);
or U2432 (N_2432,In_971,In_799);
xor U2433 (N_2433,In_4,In_929);
nor U2434 (N_2434,In_304,In_337);
or U2435 (N_2435,In_374,In_39);
or U2436 (N_2436,In_951,In_328);
or U2437 (N_2437,In_763,In_897);
and U2438 (N_2438,In_886,In_777);
nor U2439 (N_2439,In_292,In_177);
nand U2440 (N_2440,In_725,In_956);
xor U2441 (N_2441,In_372,In_54);
nor U2442 (N_2442,In_817,In_944);
nor U2443 (N_2443,In_818,In_241);
nor U2444 (N_2444,In_132,In_43);
xor U2445 (N_2445,In_409,In_104);
xnor U2446 (N_2446,In_938,In_8);
and U2447 (N_2447,In_520,In_617);
or U2448 (N_2448,In_195,In_905);
and U2449 (N_2449,In_782,In_826);
or U2450 (N_2450,In_748,In_335);
nand U2451 (N_2451,In_29,In_9);
nor U2452 (N_2452,In_116,In_190);
nor U2453 (N_2453,In_730,In_908);
xor U2454 (N_2454,In_355,In_693);
nand U2455 (N_2455,In_659,In_391);
xor U2456 (N_2456,In_142,In_505);
xnor U2457 (N_2457,In_258,In_369);
and U2458 (N_2458,In_477,In_831);
xnor U2459 (N_2459,In_910,In_892);
and U2460 (N_2460,In_264,In_619);
nand U2461 (N_2461,In_20,In_454);
or U2462 (N_2462,In_198,In_245);
and U2463 (N_2463,In_688,In_892);
nand U2464 (N_2464,In_833,In_464);
nand U2465 (N_2465,In_130,In_338);
and U2466 (N_2466,In_995,In_349);
or U2467 (N_2467,In_374,In_88);
and U2468 (N_2468,In_84,In_436);
or U2469 (N_2469,In_83,In_649);
and U2470 (N_2470,In_257,In_211);
and U2471 (N_2471,In_292,In_207);
xnor U2472 (N_2472,In_423,In_508);
xnor U2473 (N_2473,In_191,In_724);
nand U2474 (N_2474,In_543,In_56);
xor U2475 (N_2475,In_789,In_667);
nor U2476 (N_2476,In_519,In_227);
nor U2477 (N_2477,In_681,In_147);
nand U2478 (N_2478,In_725,In_300);
xor U2479 (N_2479,In_178,In_38);
or U2480 (N_2480,In_167,In_902);
xor U2481 (N_2481,In_900,In_590);
or U2482 (N_2482,In_896,In_486);
and U2483 (N_2483,In_130,In_980);
xnor U2484 (N_2484,In_624,In_8);
xnor U2485 (N_2485,In_225,In_394);
and U2486 (N_2486,In_295,In_950);
or U2487 (N_2487,In_262,In_378);
xor U2488 (N_2488,In_541,In_976);
nor U2489 (N_2489,In_314,In_546);
nand U2490 (N_2490,In_130,In_747);
xnor U2491 (N_2491,In_36,In_674);
nor U2492 (N_2492,In_632,In_550);
and U2493 (N_2493,In_272,In_71);
or U2494 (N_2494,In_63,In_860);
nor U2495 (N_2495,In_643,In_758);
nand U2496 (N_2496,In_967,In_679);
or U2497 (N_2497,In_818,In_347);
and U2498 (N_2498,In_851,In_890);
and U2499 (N_2499,In_406,In_34);
nor U2500 (N_2500,N_1693,N_932);
xor U2501 (N_2501,N_2008,N_1811);
nor U2502 (N_2502,N_695,N_1454);
nand U2503 (N_2503,N_502,N_1252);
and U2504 (N_2504,N_1527,N_1232);
and U2505 (N_2505,N_1519,N_2258);
and U2506 (N_2506,N_568,N_1215);
xor U2507 (N_2507,N_1395,N_1917);
xnor U2508 (N_2508,N_1826,N_750);
and U2509 (N_2509,N_538,N_896);
xnor U2510 (N_2510,N_897,N_1868);
or U2511 (N_2511,N_1406,N_638);
nand U2512 (N_2512,N_1067,N_636);
xor U2513 (N_2513,N_1746,N_88);
xor U2514 (N_2514,N_167,N_529);
xor U2515 (N_2515,N_1686,N_1995);
nor U2516 (N_2516,N_86,N_32);
or U2517 (N_2517,N_309,N_609);
xnor U2518 (N_2518,N_1038,N_2127);
xor U2519 (N_2519,N_849,N_2225);
and U2520 (N_2520,N_377,N_49);
and U2521 (N_2521,N_516,N_517);
and U2522 (N_2522,N_2015,N_1564);
nor U2523 (N_2523,N_295,N_105);
or U2524 (N_2524,N_1310,N_919);
nand U2525 (N_2525,N_890,N_1155);
or U2526 (N_2526,N_308,N_1325);
xor U2527 (N_2527,N_2484,N_1723);
and U2528 (N_2528,N_2451,N_1249);
nor U2529 (N_2529,N_2226,N_1034);
nand U2530 (N_2530,N_214,N_7);
and U2531 (N_2531,N_84,N_1084);
nand U2532 (N_2532,N_1961,N_1261);
and U2533 (N_2533,N_1577,N_1465);
nor U2534 (N_2534,N_725,N_2163);
or U2535 (N_2535,N_981,N_2269);
and U2536 (N_2536,N_1503,N_1547);
nand U2537 (N_2537,N_1624,N_465);
or U2538 (N_2538,N_1654,N_704);
and U2539 (N_2539,N_410,N_1182);
nand U2540 (N_2540,N_1389,N_2120);
and U2541 (N_2541,N_1025,N_1306);
or U2542 (N_2542,N_1890,N_2423);
or U2543 (N_2543,N_1715,N_2230);
and U2544 (N_2544,N_2236,N_1688);
nand U2545 (N_2545,N_1258,N_628);
nand U2546 (N_2546,N_576,N_1659);
or U2547 (N_2547,N_1081,N_408);
xor U2548 (N_2548,N_1426,N_531);
nand U2549 (N_2549,N_1922,N_795);
xnor U2550 (N_2550,N_2132,N_1728);
nand U2551 (N_2551,N_2465,N_539);
nor U2552 (N_2552,N_294,N_367);
nand U2553 (N_2553,N_2246,N_1499);
or U2554 (N_2554,N_2342,N_709);
and U2555 (N_2555,N_2149,N_1187);
nor U2556 (N_2556,N_33,N_671);
or U2557 (N_2557,N_255,N_2084);
xnor U2558 (N_2558,N_1488,N_1885);
xor U2559 (N_2559,N_1030,N_1866);
nor U2560 (N_2560,N_2444,N_1703);
and U2561 (N_2561,N_1440,N_2217);
nor U2562 (N_2562,N_2042,N_268);
nor U2563 (N_2563,N_1735,N_315);
or U2564 (N_2564,N_317,N_2142);
xnor U2565 (N_2565,N_1364,N_506);
xnor U2566 (N_2566,N_1991,N_943);
nor U2567 (N_2567,N_2277,N_1360);
nand U2568 (N_2568,N_37,N_1997);
nand U2569 (N_2569,N_2313,N_1611);
nor U2570 (N_2570,N_1640,N_1322);
and U2571 (N_2571,N_1127,N_11);
or U2572 (N_2572,N_555,N_690);
and U2573 (N_2573,N_349,N_2201);
or U2574 (N_2574,N_1248,N_1820);
or U2575 (N_2575,N_1619,N_1166);
nand U2576 (N_2576,N_549,N_1721);
and U2577 (N_2577,N_483,N_736);
nand U2578 (N_2578,N_2453,N_310);
nor U2579 (N_2579,N_2141,N_256);
or U2580 (N_2580,N_1633,N_1586);
nand U2581 (N_2581,N_976,N_420);
xor U2582 (N_2582,N_1348,N_754);
nor U2583 (N_2583,N_36,N_1705);
or U2584 (N_2584,N_683,N_888);
or U2585 (N_2585,N_1342,N_742);
or U2586 (N_2586,N_835,N_964);
nand U2587 (N_2587,N_1445,N_1904);
nor U2588 (N_2588,N_661,N_2394);
or U2589 (N_2589,N_2154,N_1908);
xnor U2590 (N_2590,N_1867,N_1637);
and U2591 (N_2591,N_14,N_1321);
or U2592 (N_2592,N_643,N_118);
and U2593 (N_2593,N_1651,N_1699);
nor U2594 (N_2594,N_1168,N_1761);
and U2595 (N_2595,N_8,N_2460);
nor U2596 (N_2596,N_867,N_448);
xnor U2597 (N_2597,N_594,N_724);
and U2598 (N_2598,N_1662,N_2454);
nor U2599 (N_2599,N_802,N_278);
nor U2600 (N_2600,N_148,N_1185);
and U2601 (N_2601,N_1143,N_1971);
xor U2602 (N_2602,N_1815,N_855);
or U2603 (N_2603,N_200,N_2382);
xor U2604 (N_2604,N_2026,N_1441);
nor U2605 (N_2605,N_2368,N_935);
and U2606 (N_2606,N_2208,N_1539);
and U2607 (N_2607,N_829,N_64);
and U2608 (N_2608,N_1158,N_519);
xor U2609 (N_2609,N_34,N_1119);
or U2610 (N_2610,N_1593,N_1114);
nand U2611 (N_2611,N_78,N_2206);
and U2612 (N_2612,N_1351,N_1159);
nor U2613 (N_2613,N_2278,N_891);
nor U2614 (N_2614,N_817,N_2261);
nand U2615 (N_2615,N_287,N_2346);
nor U2616 (N_2616,N_863,N_2104);
xor U2617 (N_2617,N_2310,N_391);
or U2618 (N_2618,N_1381,N_1457);
xor U2619 (N_2619,N_326,N_2094);
and U2620 (N_2620,N_2403,N_1965);
nand U2621 (N_2621,N_1007,N_955);
nand U2622 (N_2622,N_893,N_460);
nor U2623 (N_2623,N_1666,N_411);
nor U2624 (N_2624,N_1399,N_737);
nand U2625 (N_2625,N_1046,N_1966);
and U2626 (N_2626,N_2321,N_1006);
xor U2627 (N_2627,N_173,N_422);
nand U2628 (N_2628,N_1392,N_881);
and U2629 (N_2629,N_2404,N_137);
and U2630 (N_2630,N_1600,N_313);
or U2631 (N_2631,N_1111,N_1572);
or U2632 (N_2632,N_250,N_1663);
xnor U2633 (N_2633,N_670,N_899);
nand U2634 (N_2634,N_511,N_2020);
xor U2635 (N_2635,N_42,N_475);
nand U2636 (N_2636,N_366,N_1368);
or U2637 (N_2637,N_1412,N_2216);
xnor U2638 (N_2638,N_2352,N_1580);
or U2639 (N_2639,N_731,N_1959);
nand U2640 (N_2640,N_1596,N_1425);
xor U2641 (N_2641,N_1530,N_265);
nor U2642 (N_2642,N_1109,N_165);
xor U2643 (N_2643,N_844,N_2000);
nand U2644 (N_2644,N_325,N_1538);
or U2645 (N_2645,N_967,N_1635);
nor U2646 (N_2646,N_1860,N_1801);
and U2647 (N_2647,N_2472,N_106);
nor U2648 (N_2648,N_1671,N_330);
xor U2649 (N_2649,N_1018,N_53);
or U2650 (N_2650,N_542,N_1729);
nor U2651 (N_2651,N_755,N_895);
nor U2652 (N_2652,N_1759,N_1225);
nand U2653 (N_2653,N_2434,N_2390);
nand U2654 (N_2654,N_1978,N_2438);
nand U2655 (N_2655,N_3,N_1694);
xor U2656 (N_2656,N_633,N_1313);
nand U2657 (N_2657,N_1268,N_716);
nor U2658 (N_2658,N_1035,N_1308);
xnor U2659 (N_2659,N_253,N_1548);
xor U2660 (N_2660,N_1865,N_2088);
or U2661 (N_2661,N_1052,N_550);
xnor U2662 (N_2662,N_1123,N_2260);
xor U2663 (N_2663,N_455,N_2369);
and U2664 (N_2664,N_1171,N_757);
and U2665 (N_2665,N_699,N_320);
or U2666 (N_2666,N_288,N_807);
and U2667 (N_2667,N_462,N_1305);
nor U2668 (N_2668,N_231,N_1498);
nor U2669 (N_2669,N_299,N_756);
or U2670 (N_2670,N_306,N_2459);
xnor U2671 (N_2671,N_916,N_2044);
and U2672 (N_2672,N_814,N_177);
xor U2673 (N_2673,N_1089,N_908);
or U2674 (N_2674,N_1193,N_484);
nand U2675 (N_2675,N_1823,N_2265);
xor U2676 (N_2676,N_2147,N_813);
xnor U2677 (N_2677,N_1272,N_1743);
nor U2678 (N_2678,N_1575,N_124);
nand U2679 (N_2679,N_2467,N_449);
xor U2680 (N_2680,N_1960,N_1112);
nand U2681 (N_2681,N_642,N_67);
and U2682 (N_2682,N_438,N_780);
or U2683 (N_2683,N_2073,N_263);
and U2684 (N_2684,N_386,N_164);
xor U2685 (N_2685,N_2348,N_557);
and U2686 (N_2686,N_2435,N_1338);
nor U2687 (N_2687,N_1246,N_56);
and U2688 (N_2688,N_1757,N_2294);
nor U2689 (N_2689,N_676,N_1205);
or U2690 (N_2690,N_640,N_906);
nor U2691 (N_2691,N_1106,N_1181);
xnor U2692 (N_2692,N_1140,N_2340);
nor U2693 (N_2693,N_237,N_2220);
nor U2694 (N_2694,N_392,N_47);
nand U2695 (N_2695,N_645,N_1652);
nand U2696 (N_2696,N_1452,N_954);
nor U2697 (N_2697,N_902,N_1370);
nor U2698 (N_2698,N_1645,N_1667);
xor U2699 (N_2699,N_1913,N_1359);
nor U2700 (N_2700,N_2383,N_2327);
nor U2701 (N_2701,N_2036,N_564);
and U2702 (N_2702,N_2161,N_1022);
and U2703 (N_2703,N_1145,N_2419);
or U2704 (N_2704,N_436,N_280);
or U2705 (N_2705,N_1196,N_2136);
or U2706 (N_2706,N_903,N_433);
nand U2707 (N_2707,N_769,N_144);
nor U2708 (N_2708,N_1169,N_1615);
or U2709 (N_2709,N_2098,N_2409);
or U2710 (N_2710,N_806,N_646);
or U2711 (N_2711,N_247,N_1150);
nand U2712 (N_2712,N_454,N_2115);
xnor U2713 (N_2713,N_521,N_980);
xnor U2714 (N_2714,N_476,N_72);
nor U2715 (N_2715,N_752,N_602);
or U2716 (N_2716,N_857,N_1949);
nor U2717 (N_2717,N_533,N_1365);
nand U2718 (N_2718,N_27,N_1930);
or U2719 (N_2719,N_2179,N_1269);
nor U2720 (N_2720,N_2183,N_1554);
xnor U2721 (N_2721,N_712,N_2055);
nand U2722 (N_2722,N_1608,N_759);
or U2723 (N_2723,N_1096,N_1763);
and U2724 (N_2724,N_275,N_590);
or U2725 (N_2725,N_2481,N_641);
xnor U2726 (N_2726,N_1638,N_1891);
or U2727 (N_2727,N_1676,N_525);
and U2728 (N_2728,N_721,N_1576);
and U2729 (N_2729,N_809,N_1509);
and U2730 (N_2730,N_187,N_1481);
nand U2731 (N_2731,N_2070,N_1683);
and U2732 (N_2732,N_1453,N_477);
and U2733 (N_2733,N_1097,N_1798);
xor U2734 (N_2734,N_1433,N_1724);
or U2735 (N_2735,N_262,N_2167);
and U2736 (N_2736,N_421,N_1056);
nor U2737 (N_2737,N_1849,N_1354);
or U2738 (N_2738,N_1881,N_1814);
xnor U2739 (N_2739,N_73,N_1203);
xor U2740 (N_2740,N_223,N_2239);
nand U2741 (N_2741,N_761,N_149);
or U2742 (N_2742,N_2080,N_405);
nor U2743 (N_2743,N_946,N_672);
nor U2744 (N_2744,N_1386,N_1108);
nand U2745 (N_2745,N_1099,N_304);
and U2746 (N_2746,N_328,N_2013);
or U2747 (N_2747,N_1559,N_989);
and U2748 (N_2748,N_1719,N_1969);
nor U2749 (N_2749,N_584,N_1075);
or U2750 (N_2750,N_336,N_1905);
and U2751 (N_2751,N_950,N_2191);
xor U2752 (N_2752,N_493,N_1847);
xnor U2753 (N_2753,N_1256,N_782);
or U2754 (N_2754,N_1076,N_681);
nand U2755 (N_2755,N_2307,N_1679);
or U2756 (N_2756,N_2172,N_2218);
nand U2757 (N_2757,N_2338,N_2344);
and U2758 (N_2758,N_2447,N_1393);
nor U2759 (N_2759,N_1753,N_949);
xnor U2760 (N_2760,N_1648,N_1054);
nand U2761 (N_2761,N_2461,N_2181);
and U2762 (N_2762,N_738,N_378);
and U2763 (N_2763,N_456,N_2229);
xor U2764 (N_2764,N_2323,N_2030);
xnor U2765 (N_2765,N_928,N_577);
nand U2766 (N_2766,N_694,N_1449);
or U2767 (N_2767,N_1942,N_2466);
nor U2768 (N_2768,N_1478,N_234);
nand U2769 (N_2769,N_1768,N_1045);
nand U2770 (N_2770,N_1324,N_2114);
nand U2771 (N_2771,N_1574,N_1956);
nand U2772 (N_2772,N_2328,N_2279);
nor U2773 (N_2773,N_1973,N_730);
xnor U2774 (N_2774,N_122,N_1455);
nand U2775 (N_2775,N_504,N_1356);
xor U2776 (N_2776,N_1188,N_400);
nor U2777 (N_2777,N_1627,N_2072);
and U2778 (N_2778,N_717,N_1583);
nor U2779 (N_2779,N_70,N_2486);
and U2780 (N_2780,N_443,N_2306);
nor U2781 (N_2781,N_2199,N_1191);
or U2782 (N_2782,N_401,N_233);
xnor U2783 (N_2783,N_1825,N_398);
nor U2784 (N_2784,N_512,N_513);
and U2785 (N_2785,N_1431,N_2488);
nor U2786 (N_2786,N_2119,N_2109);
or U2787 (N_2787,N_350,N_1817);
xor U2788 (N_2788,N_1843,N_2405);
and U2789 (N_2789,N_1556,N_2320);
nor U2790 (N_2790,N_1220,N_1350);
nand U2791 (N_2791,N_2052,N_986);
and U2792 (N_2792,N_2384,N_936);
nand U2793 (N_2793,N_1852,N_1286);
or U2794 (N_2794,N_1216,N_457);
nand U2795 (N_2795,N_1563,N_771);
nor U2796 (N_2796,N_1420,N_792);
or U2797 (N_2797,N_1070,N_581);
nor U2798 (N_2798,N_79,N_657);
nor U2799 (N_2799,N_705,N_1599);
nand U2800 (N_2800,N_2339,N_1988);
or U2801 (N_2801,N_2326,N_693);
nor U2802 (N_2802,N_239,N_23);
xnor U2803 (N_2803,N_1788,N_103);
xor U2804 (N_2804,N_1065,N_1626);
and U2805 (N_2805,N_558,N_1019);
xnor U2806 (N_2806,N_828,N_1484);
nand U2807 (N_2807,N_1524,N_1260);
or U2808 (N_2808,N_1660,N_485);
and U2809 (N_2809,N_1585,N_1396);
and U2810 (N_2810,N_248,N_1689);
xnor U2811 (N_2811,N_2424,N_193);
or U2812 (N_2812,N_1806,N_1813);
nor U2813 (N_2813,N_1709,N_1295);
and U2814 (N_2814,N_1312,N_1841);
nor U2815 (N_2815,N_1601,N_1783);
xnor U2816 (N_2816,N_403,N_680);
and U2817 (N_2817,N_1243,N_2041);
xor U2818 (N_2818,N_251,N_1078);
xor U2819 (N_2819,N_2315,N_701);
nand U2820 (N_2820,N_2219,N_973);
nand U2821 (N_2821,N_60,N_2134);
and U2822 (N_2822,N_1644,N_138);
xnor U2823 (N_2823,N_1562,N_1299);
or U2824 (N_2824,N_885,N_1794);
or U2825 (N_2825,N_1511,N_473);
or U2826 (N_2826,N_940,N_1032);
nor U2827 (N_2827,N_2375,N_706);
xnor U2828 (N_2828,N_1733,N_861);
or U2829 (N_2829,N_686,N_1080);
and U2830 (N_2830,N_2268,N_1749);
nor U2831 (N_2831,N_191,N_2449);
and U2832 (N_2832,N_612,N_2416);
nor U2833 (N_2833,N_1598,N_1621);
xor U2834 (N_2834,N_2176,N_877);
and U2835 (N_2835,N_1818,N_2397);
nor U2836 (N_2836,N_2249,N_944);
nand U2837 (N_2837,N_2241,N_997);
and U2838 (N_2838,N_2097,N_1491);
or U2839 (N_2839,N_2064,N_242);
nor U2840 (N_2840,N_664,N_1822);
or U2841 (N_2841,N_162,N_1464);
xor U2842 (N_2842,N_2391,N_1702);
or U2843 (N_2843,N_2202,N_1409);
or U2844 (N_2844,N_2399,N_1394);
nor U2845 (N_2845,N_1289,N_1192);
nand U2846 (N_2846,N_1931,N_588);
and U2847 (N_2847,N_2290,N_823);
nor U2848 (N_2848,N_1899,N_824);
and U2849 (N_2849,N_2076,N_659);
xor U2850 (N_2850,N_1777,N_1320);
xnor U2851 (N_2851,N_1967,N_2221);
and U2852 (N_2852,N_2250,N_1963);
nand U2853 (N_2853,N_1643,N_348);
or U2854 (N_2854,N_1919,N_962);
xor U2855 (N_2855,N_62,N_1830);
xor U2856 (N_2856,N_161,N_1876);
xnor U2857 (N_2857,N_171,N_2464);
xnor U2858 (N_2858,N_930,N_1687);
and U2859 (N_2859,N_2113,N_563);
nor U2860 (N_2860,N_1871,N_218);
and U2861 (N_2861,N_1490,N_2002);
nor U2862 (N_2862,N_2308,N_1367);
nor U2863 (N_2863,N_2285,N_1769);
nand U2864 (N_2864,N_1063,N_1979);
and U2865 (N_2865,N_1578,N_2003);
or U2866 (N_2866,N_2446,N_2406);
or U2867 (N_2867,N_678,N_1254);
nor U2868 (N_2868,N_1456,N_48);
nand U2869 (N_2869,N_1026,N_2215);
nand U2870 (N_2870,N_2032,N_1234);
or U2871 (N_2871,N_1267,N_175);
and U2872 (N_2872,N_2180,N_1226);
and U2873 (N_2873,N_2355,N_1945);
nand U2874 (N_2874,N_562,N_69);
and U2875 (N_2875,N_963,N_1157);
or U2876 (N_2876,N_472,N_1402);
nor U2877 (N_2877,N_1906,N_1941);
xor U2878 (N_2878,N_1828,N_1873);
nand U2879 (N_2879,N_1069,N_1658);
or U2880 (N_2880,N_482,N_674);
nor U2881 (N_2881,N_254,N_1280);
or U2882 (N_2882,N_719,N_2425);
nand U2883 (N_2883,N_1008,N_1397);
and U2884 (N_2884,N_1605,N_673);
nor U2885 (N_2885,N_1824,N_1856);
nand U2886 (N_2886,N_763,N_1928);
nand U2887 (N_2887,N_1879,N_58);
nor U2888 (N_2888,N_1845,N_1537);
nor U2889 (N_2889,N_684,N_2233);
or U2890 (N_2890,N_2050,N_883);
nor U2891 (N_2891,N_1921,N_1408);
or U2892 (N_2892,N_1877,N_598);
xor U2893 (N_2893,N_580,N_338);
nand U2894 (N_2894,N_1533,N_1040);
and U2895 (N_2895,N_2232,N_876);
and U2896 (N_2896,N_266,N_221);
xnor U2897 (N_2897,N_2337,N_1482);
nand U2898 (N_2898,N_307,N_1137);
nor U2899 (N_2899,N_613,N_2116);
nor U2900 (N_2900,N_343,N_2146);
or U2901 (N_2901,N_1964,N_227);
and U2902 (N_2902,N_414,N_929);
or U2903 (N_2903,N_1668,N_1208);
nand U2904 (N_2904,N_1033,N_2187);
nand U2905 (N_2905,N_556,N_1403);
xor U2906 (N_2906,N_648,N_1095);
or U2907 (N_2907,N_1421,N_1303);
nand U2908 (N_2908,N_1,N_2238);
nand U2909 (N_2909,N_1128,N_2427);
or U2910 (N_2910,N_822,N_481);
xor U2911 (N_2911,N_318,N_1677);
xnor U2912 (N_2912,N_63,N_623);
nand U2913 (N_2913,N_1373,N_1602);
nor U2914 (N_2914,N_82,N_1469);
and U2915 (N_2915,N_1629,N_966);
nor U2916 (N_2916,N_2252,N_1450);
xnor U2917 (N_2917,N_1784,N_697);
or U2918 (N_2918,N_2398,N_1218);
nand U2919 (N_2919,N_195,N_2165);
or U2920 (N_2920,N_2392,N_492);
nor U2921 (N_2921,N_159,N_2031);
nand U2922 (N_2922,N_1855,N_958);
and U2923 (N_2923,N_2157,N_1976);
or U2924 (N_2924,N_1692,N_133);
and U2925 (N_2925,N_2067,N_2089);
xor U2926 (N_2926,N_241,N_1361);
nand U2927 (N_2927,N_184,N_2096);
and U2928 (N_2928,N_258,N_2156);
or U2929 (N_2929,N_2305,N_1907);
nand U2930 (N_2930,N_1549,N_1304);
xnor U2931 (N_2931,N_1797,N_707);
nand U2932 (N_2932,N_735,N_974);
xnor U2933 (N_2933,N_1088,N_87);
or U2934 (N_2934,N_2063,N_1641);
or U2935 (N_2935,N_1031,N_753);
xnor U2936 (N_2936,N_922,N_2062);
nand U2937 (N_2937,N_1521,N_746);
and U2938 (N_2938,N_2300,N_1613);
xnor U2939 (N_2939,N_1739,N_205);
and U2940 (N_2940,N_1786,N_495);
or U2941 (N_2941,N_1141,N_1766);
nor U2942 (N_2942,N_1116,N_1178);
nand U2943 (N_2943,N_751,N_1447);
nor U2944 (N_2944,N_249,N_571);
nor U2945 (N_2945,N_415,N_332);
xnor U2946 (N_2946,N_839,N_1102);
and U2947 (N_2947,N_2228,N_501);
and U2948 (N_2948,N_1413,N_119);
and U2949 (N_2949,N_1259,N_1147);
nand U2950 (N_2950,N_1535,N_1079);
or U2951 (N_2951,N_2168,N_991);
nand U2952 (N_2952,N_314,N_419);
nor U2953 (N_2953,N_154,N_1459);
or U2954 (N_2954,N_2235,N_2441);
nand U2955 (N_2955,N_146,N_2492);
nor U2956 (N_2956,N_601,N_1754);
nand U2957 (N_2957,N_1170,N_783);
and U2958 (N_2958,N_1020,N_188);
nor U2959 (N_2959,N_573,N_51);
and U2960 (N_2960,N_180,N_2332);
or U2961 (N_2961,N_2264,N_434);
nor U2962 (N_2962,N_1331,N_211);
nand U2963 (N_2963,N_351,N_2039);
and U2964 (N_2964,N_1916,N_1625);
xnor U2965 (N_2965,N_566,N_1347);
nand U2966 (N_2966,N_1091,N_2443);
or U2967 (N_2967,N_2359,N_125);
nor U2968 (N_2968,N_848,N_297);
and U2969 (N_2969,N_323,N_765);
nor U2970 (N_2970,N_786,N_904);
xnor U2971 (N_2971,N_800,N_1863);
and U2972 (N_2972,N_2038,N_1374);
xnor U2973 (N_2973,N_2011,N_1282);
nor U2974 (N_2974,N_1221,N_1180);
nand U2975 (N_2975,N_1557,N_1307);
nor U2976 (N_2976,N_727,N_2297);
or U2977 (N_2977,N_92,N_1179);
and U2978 (N_2978,N_1494,N_1840);
xor U2979 (N_2979,N_2282,N_1201);
nor U2980 (N_2980,N_820,N_489);
nor U2981 (N_2981,N_1567,N_772);
or U2982 (N_2982,N_101,N_459);
nor U2983 (N_2983,N_1257,N_1121);
xnor U2984 (N_2984,N_1051,N_1124);
nor U2985 (N_2985,N_1909,N_2366);
nor U2986 (N_2986,N_1375,N_1023);
and U2987 (N_2987,N_463,N_1691);
xnor U2988 (N_2988,N_559,N_1189);
and U2989 (N_2989,N_630,N_859);
nor U2990 (N_2990,N_113,N_1048);
or U2991 (N_2991,N_1785,N_261);
nand U2992 (N_2992,N_990,N_1834);
nor U2993 (N_2993,N_2099,N_2376);
and U2994 (N_2994,N_1592,N_959);
nor U2995 (N_2995,N_1740,N_808);
xor U2996 (N_2996,N_2170,N_2266);
and U2997 (N_2997,N_1085,N_1461);
xnor U2998 (N_2998,N_347,N_197);
or U2999 (N_2999,N_213,N_1398);
or U3000 (N_3000,N_740,N_1990);
nand U3001 (N_3001,N_2057,N_1750);
xor U3002 (N_3002,N_2267,N_9);
or U3003 (N_3003,N_1113,N_12);
nand U3004 (N_3004,N_1337,N_2445);
nor U3005 (N_3005,N_1987,N_1416);
xor U3006 (N_3006,N_2029,N_57);
or U3007 (N_3007,N_1198,N_189);
or U3008 (N_3008,N_6,N_131);
or U3009 (N_3009,N_91,N_353);
or U3010 (N_3010,N_781,N_284);
and U3011 (N_3011,N_76,N_1311);
xnor U3012 (N_3012,N_2001,N_634);
and U3013 (N_3013,N_953,N_1773);
nor U3014 (N_3014,N_2194,N_447);
or U3015 (N_3015,N_2009,N_865);
and U3016 (N_3016,N_799,N_1732);
or U3017 (N_3017,N_836,N_937);
or U3018 (N_3018,N_2185,N_2121);
and U3019 (N_3019,N_1297,N_2110);
or U3020 (N_3020,N_834,N_1776);
and U3021 (N_3021,N_2111,N_2259);
xnor U3022 (N_3022,N_2442,N_346);
nand U3023 (N_3023,N_1770,N_1912);
xnor U3024 (N_3024,N_1911,N_126);
nor U3025 (N_3025,N_1850,N_1133);
xnor U3026 (N_3026,N_1343,N_1875);
or U3027 (N_3027,N_1551,N_210);
xor U3028 (N_3028,N_948,N_1428);
nor U3029 (N_3029,N_651,N_198);
nand U3030 (N_3030,N_2408,N_1233);
or U3031 (N_3031,N_1632,N_153);
nand U3032 (N_3032,N_1086,N_2131);
nand U3033 (N_3033,N_1796,N_2177);
and U3034 (N_3034,N_669,N_530);
xnor U3035 (N_3035,N_208,N_873);
nand U3036 (N_3036,N_710,N_1027);
nand U3037 (N_3037,N_1836,N_2373);
nor U3038 (N_3038,N_743,N_845);
nor U3039 (N_3039,N_1595,N_388);
xnor U3040 (N_3040,N_675,N_2287);
nor U3041 (N_3041,N_300,N_203);
xnor U3042 (N_3042,N_246,N_1704);
and U3043 (N_3043,N_2496,N_979);
and U3044 (N_3044,N_933,N_383);
nor U3045 (N_3045,N_758,N_2137);
nor U3046 (N_3046,N_1832,N_352);
nor U3047 (N_3047,N_2389,N_1357);
or U3048 (N_3048,N_1610,N_1462);
xor U3049 (N_3049,N_1105,N_2316);
and U3050 (N_3050,N_2018,N_1223);
xor U3051 (N_3051,N_1385,N_851);
and U3052 (N_3052,N_1004,N_1029);
or U3053 (N_3053,N_1339,N_655);
nor U3054 (N_3054,N_281,N_1407);
nor U3055 (N_3055,N_114,N_1279);
nand U3056 (N_3056,N_259,N_647);
nand U3057 (N_3057,N_579,N_868);
xnor U3058 (N_3058,N_1742,N_541);
xnor U3059 (N_3059,N_2356,N_319);
and U3060 (N_3060,N_442,N_94);
or U3061 (N_3061,N_2203,N_1948);
and U3062 (N_3062,N_2049,N_965);
nor U3063 (N_3063,N_2289,N_1800);
or U3064 (N_3064,N_1090,N_961);
and U3065 (N_3065,N_2407,N_301);
and U3066 (N_3066,N_2489,N_837);
xnor U3067 (N_3067,N_2033,N_535);
nor U3068 (N_3068,N_1765,N_479);
and U3069 (N_3069,N_1092,N_1884);
xnor U3070 (N_3070,N_340,N_2410);
xor U3071 (N_3071,N_668,N_1036);
and U3072 (N_3072,N_1588,N_333);
nand U3073 (N_3073,N_217,N_2462);
nor U3074 (N_3074,N_1424,N_689);
nor U3075 (N_3075,N_30,N_1401);
xor U3076 (N_3076,N_748,N_1609);
xor U3077 (N_3077,N_894,N_708);
nand U3078 (N_3078,N_2173,N_24);
and U3079 (N_3079,N_1017,N_532);
nor U3080 (N_3080,N_1298,N_912);
and U3081 (N_3081,N_1842,N_993);
nor U3082 (N_3082,N_779,N_850);
and U3083 (N_3083,N_1047,N_1829);
and U3084 (N_3084,N_784,N_1504);
and U3085 (N_3085,N_158,N_335);
and U3086 (N_3086,N_703,N_487);
nor U3087 (N_3087,N_2335,N_745);
and U3088 (N_3088,N_1939,N_399);
xnor U3089 (N_3089,N_1589,N_616);
and U3090 (N_3090,N_413,N_1043);
xor U3091 (N_3091,N_526,N_1098);
nor U3092 (N_3092,N_626,N_1328);
nand U3093 (N_3093,N_244,N_975);
and U3094 (N_3094,N_1001,N_988);
xor U3095 (N_3095,N_130,N_1543);
nand U3096 (N_3096,N_1713,N_1423);
xnor U3097 (N_3097,N_1670,N_387);
xor U3098 (N_3098,N_1934,N_1411);
and U3099 (N_3099,N_1100,N_1838);
or U3100 (N_3100,N_1476,N_2336);
nand U3101 (N_3101,N_311,N_1695);
and U3102 (N_3102,N_2387,N_1958);
nand U3103 (N_3103,N_1992,N_572);
nand U3104 (N_3104,N_374,N_1898);
xnor U3105 (N_3105,N_1380,N_2061);
or U3106 (N_3106,N_151,N_1066);
nor U3107 (N_3107,N_2107,N_1244);
xnor U3108 (N_3108,N_1994,N_497);
xnor U3109 (N_3109,N_220,N_128);
and U3110 (N_3110,N_801,N_2411);
xor U3111 (N_3111,N_2248,N_2318);
xor U3112 (N_3112,N_446,N_1631);
nor U3113 (N_3113,N_662,N_1779);
or U3114 (N_3114,N_570,N_644);
nor U3115 (N_3115,N_1219,N_1214);
or U3116 (N_3116,N_1493,N_917);
and U3117 (N_3117,N_624,N_140);
nor U3118 (N_3118,N_774,N_589);
nand U3119 (N_3119,N_312,N_2106);
or U3120 (N_3120,N_1117,N_635);
xnor U3121 (N_3121,N_1540,N_423);
nor U3122 (N_3122,N_1405,N_787);
nand U3123 (N_3123,N_1782,N_1726);
nand U3124 (N_3124,N_2092,N_1467);
or U3125 (N_3125,N_1940,N_2130);
or U3126 (N_3126,N_1932,N_2074);
xnor U3127 (N_3127,N_1058,N_179);
or U3128 (N_3128,N_700,N_596);
nand U3129 (N_3129,N_915,N_1390);
nand U3130 (N_3130,N_1213,N_2412);
nand U3131 (N_3131,N_2380,N_826);
nand U3132 (N_3132,N_474,N_2023);
xnor U3133 (N_3133,N_44,N_1864);
or U3134 (N_3134,N_2448,N_1781);
nor U3135 (N_3135,N_2058,N_432);
nand U3136 (N_3136,N_1281,N_1851);
xnor U3137 (N_3137,N_1690,N_305);
or U3138 (N_3138,N_2028,N_264);
nor U3139 (N_3139,N_2331,N_1358);
nor U3140 (N_3140,N_1993,N_2498);
and U3141 (N_3141,N_649,N_1808);
or U3142 (N_3142,N_603,N_458);
or U3143 (N_3143,N_567,N_597);
xnor U3144 (N_3144,N_1448,N_2415);
xnor U3145 (N_3145,N_599,N_322);
nor U3146 (N_3146,N_1164,N_1273);
xnor U3147 (N_3147,N_2160,N_2150);
and U3148 (N_3148,N_1028,N_1384);
and U3149 (N_3149,N_1107,N_582);
nor U3150 (N_3150,N_1326,N_931);
or U3151 (N_3151,N_1064,N_1153);
xnor U3152 (N_3152,N_219,N_1486);
nor U3153 (N_3153,N_437,N_2100);
nand U3154 (N_3154,N_760,N_1622);
or U3155 (N_3155,N_886,N_870);
xor U3156 (N_3156,N_821,N_1315);
or U3157 (N_3157,N_2047,N_2334);
or U3158 (N_3158,N_605,N_1892);
nor U3159 (N_3159,N_277,N_2276);
xnor U3160 (N_3160,N_1861,N_1752);
and U3161 (N_3161,N_2086,N_394);
nand U3162 (N_3162,N_2400,N_2200);
nor U3163 (N_3163,N_0,N_80);
nor U3164 (N_3164,N_2463,N_1804);
and U3165 (N_3165,N_1327,N_1716);
nor U3166 (N_3166,N_1429,N_663);
and U3167 (N_3167,N_587,N_272);
xnor U3168 (N_3168,N_1377,N_1162);
and U3169 (N_3169,N_1333,N_1936);
nor U3170 (N_3170,N_1446,N_1334);
and U3171 (N_3171,N_794,N_134);
or U3172 (N_3172,N_552,N_1681);
or U3173 (N_3173,N_342,N_2480);
nand U3174 (N_3174,N_871,N_2299);
xnor U3175 (N_3175,N_274,N_380);
nand U3176 (N_3176,N_467,N_2417);
or U3177 (N_3177,N_1061,N_2312);
or U3178 (N_3178,N_1962,N_1487);
or U3179 (N_3179,N_1245,N_1561);
or U3180 (N_3180,N_376,N_412);
or U3181 (N_3181,N_2059,N_1953);
or U3182 (N_3182,N_2128,N_2066);
xor U3183 (N_3183,N_2253,N_1460);
or U3184 (N_3184,N_913,N_1947);
xnor U3185 (N_3185,N_337,N_494);
and U3186 (N_3186,N_1271,N_1073);
xnor U3187 (N_3187,N_911,N_55);
and U3188 (N_3188,N_147,N_1471);
or U3189 (N_3189,N_321,N_143);
nor U3190 (N_3190,N_155,N_1330);
or U3191 (N_3191,N_1522,N_2284);
or U3192 (N_3192,N_866,N_995);
nand U3193 (N_3193,N_1302,N_1546);
xor U3194 (N_3194,N_395,N_2014);
xnor U3195 (N_3195,N_172,N_2343);
or U3196 (N_3196,N_2019,N_574);
nor U3197 (N_3197,N_1565,N_341);
or U3198 (N_3198,N_406,N_2470);
or U3199 (N_3199,N_854,N_524);
nor U3200 (N_3200,N_790,N_1387);
and U3201 (N_3201,N_1523,N_653);
and U3202 (N_3202,N_289,N_1787);
and U3203 (N_3203,N_1810,N_1570);
and U3204 (N_3204,N_1514,N_2122);
nor U3205 (N_3205,N_1309,N_994);
or U3206 (N_3206,N_2071,N_98);
nor U3207 (N_3207,N_2469,N_951);
nand U3208 (N_3208,N_1039,N_1569);
and U3209 (N_3209,N_947,N_2010);
or U3210 (N_3210,N_1237,N_373);
or U3211 (N_3211,N_1736,N_1110);
nor U3212 (N_3212,N_586,N_1489);
and U3213 (N_3213,N_718,N_1597);
nand U3214 (N_3214,N_615,N_971);
xnor U3215 (N_3215,N_1854,N_520);
nand U3216 (N_3216,N_1050,N_920);
xnor U3217 (N_3217,N_2166,N_569);
nor U3218 (N_3218,N_747,N_480);
and U3219 (N_3219,N_81,N_1896);
nand U3220 (N_3220,N_2450,N_1870);
nor U3221 (N_3221,N_2124,N_770);
xor U3222 (N_3222,N_1914,N_293);
xnor U3223 (N_3223,N_331,N_1902);
and U3224 (N_3224,N_426,N_575);
or U3225 (N_3225,N_409,N_1792);
or U3226 (N_3226,N_825,N_1344);
nor U3227 (N_3227,N_1620,N_1925);
xor U3228 (N_3228,N_1647,N_1673);
nor U3229 (N_3229,N_1053,N_739);
xnor U3230 (N_3230,N_2090,N_1566);
xnor U3231 (N_3231,N_2118,N_2255);
xnor U3232 (N_3232,N_1607,N_593);
or U3233 (N_3233,N_2302,N_345);
nand U3234 (N_3234,N_238,N_121);
nand U3235 (N_3235,N_1714,N_54);
and U3236 (N_3236,N_658,N_921);
xnor U3237 (N_3237,N_500,N_1636);
or U3238 (N_3238,N_68,N_2197);
and U3239 (N_3239,N_1707,N_1165);
and U3240 (N_3240,N_749,N_245);
xor U3241 (N_3241,N_543,N_1661);
nand U3242 (N_3242,N_2169,N_2153);
and U3243 (N_3243,N_344,N_157);
nand U3244 (N_3244,N_2037,N_117);
and U3245 (N_3245,N_972,N_1266);
and U3246 (N_3246,N_1184,N_2237);
or U3247 (N_3247,N_1646,N_2175);
nand U3248 (N_3248,N_1163,N_16);
and U3249 (N_3249,N_548,N_1319);
nor U3250 (N_3250,N_206,N_561);
nand U3251 (N_3251,N_2087,N_1419);
and U3252 (N_3252,N_267,N_1270);
nand U3253 (N_3253,N_1346,N_1937);
xor U3254 (N_3254,N_793,N_923);
nand U3255 (N_3255,N_1122,N_2271);
and U3256 (N_3256,N_26,N_296);
xnor U3257 (N_3257,N_1174,N_430);
xnor U3258 (N_3258,N_1710,N_181);
xnor U3259 (N_3259,N_1087,N_29);
nor U3260 (N_3260,N_1650,N_2190);
xnor U3261 (N_3261,N_1748,N_1839);
nand U3262 (N_3262,N_1442,N_402);
nor U3263 (N_3263,N_141,N_987);
nor U3264 (N_3264,N_1410,N_1265);
nand U3265 (N_3265,N_1341,N_1483);
xor U3266 (N_3266,N_1685,N_762);
nor U3267 (N_3267,N_1731,N_1857);
or U3268 (N_3268,N_667,N_1217);
and U3269 (N_3269,N_970,N_595);
nor U3270 (N_3270,N_2151,N_243);
or U3271 (N_3271,N_2025,N_2351);
xnor U3272 (N_3272,N_1148,N_2456);
or U3273 (N_3273,N_853,N_677);
and U3274 (N_3274,N_1968,N_2440);
xnor U3275 (N_3275,N_327,N_1722);
xor U3276 (N_3276,N_2198,N_163);
xnor U3277 (N_3277,N_942,N_2487);
and U3278 (N_3278,N_2283,N_722);
nand U3279 (N_3279,N_1897,N_2140);
nor U3280 (N_3280,N_235,N_2251);
nand U3281 (N_3281,N_5,N_2035);
and U3282 (N_3282,N_1933,N_65);
nand U3283 (N_3283,N_889,N_229);
xnor U3284 (N_3284,N_1951,N_1427);
nor U3285 (N_3285,N_1176,N_1340);
or U3286 (N_3286,N_1649,N_1872);
xor U3287 (N_3287,N_190,N_1880);
and U3288 (N_3288,N_363,N_518);
xor U3289 (N_3289,N_1970,N_1718);
xor U3290 (N_3290,N_1552,N_2082);
and U3291 (N_3291,N_1131,N_240);
or U3292 (N_3292,N_1238,N_1915);
nor U3293 (N_3293,N_1526,N_1037);
or U3294 (N_3294,N_2189,N_1439);
nor U3295 (N_3295,N_687,N_831);
or U3296 (N_3296,N_1986,N_2256);
nand U3297 (N_3297,N_1138,N_1473);
and U3298 (N_3298,N_1981,N_618);
and U3299 (N_3299,N_1678,N_619);
and U3300 (N_3300,N_444,N_1156);
nor U3301 (N_3301,N_1977,N_1345);
nor U3302 (N_3302,N_1512,N_1093);
or U3303 (N_3303,N_2314,N_71);
nor U3304 (N_3304,N_2006,N_938);
nor U3305 (N_3305,N_1104,N_1846);
nand U3306 (N_3306,N_1206,N_2126);
and U3307 (N_3307,N_2139,N_1573);
xnor U3308 (N_3308,N_2045,N_1264);
and U3309 (N_3309,N_939,N_4);
xor U3310 (N_3310,N_2192,N_445);
and U3311 (N_3311,N_875,N_1404);
nand U3312 (N_3312,N_2457,N_1926);
and U3313 (N_3313,N_59,N_2354);
nor U3314 (N_3314,N_1837,N_2125);
xor U3315 (N_3315,N_1136,N_2048);
nor U3316 (N_3316,N_2091,N_232);
nand U3317 (N_3317,N_324,N_1443);
xor U3318 (N_3318,N_2304,N_1697);
xor U3319 (N_3319,N_1720,N_215);
or U3320 (N_3320,N_798,N_2105);
and U3321 (N_3321,N_1518,N_1130);
xnor U3322 (N_3322,N_186,N_1015);
nand U3323 (N_3323,N_2345,N_1082);
nand U3324 (N_3324,N_2288,N_1161);
nand U3325 (N_3325,N_282,N_2471);
or U3326 (N_3326,N_21,N_291);
xor U3327 (N_3327,N_1571,N_1011);
and U3328 (N_3328,N_390,N_1502);
or U3329 (N_3329,N_720,N_1332);
nor U3330 (N_3330,N_1468,N_2413);
and U3331 (N_3331,N_583,N_1183);
nor U3332 (N_3332,N_2273,N_1013);
and U3333 (N_3333,N_404,N_1400);
nor U3334 (N_3334,N_1591,N_1492);
nor U3335 (N_3335,N_882,N_418);
or U3336 (N_3336,N_2381,N_1186);
or U3337 (N_3337,N_368,N_832);
nand U3338 (N_3338,N_1528,N_713);
nor U3339 (N_3339,N_1895,N_1532);
and U3340 (N_3340,N_361,N_1653);
nor U3341 (N_3341,N_1698,N_874);
or U3342 (N_3342,N_2363,N_372);
nand U3343 (N_3343,N_732,N_1195);
or U3344 (N_3344,N_1950,N_1758);
xnor U3345 (N_3345,N_407,N_2231);
nor U3346 (N_3346,N_1239,N_2083);
and U3347 (N_3347,N_2458,N_2330);
nor U3348 (N_3348,N_339,N_109);
nand U3349 (N_3349,N_142,N_2436);
nor U3350 (N_3350,N_996,N_1444);
or U3351 (N_3351,N_1944,N_2081);
xor U3352 (N_3352,N_2291,N_1791);
xnor U3353 (N_3353,N_375,N_2499);
and U3354 (N_3354,N_1929,N_1594);
and U3355 (N_3355,N_804,N_1998);
nor U3356 (N_3356,N_688,N_356);
and U3357 (N_3357,N_1495,N_1438);
nor U3358 (N_3358,N_1154,N_1616);
or U3359 (N_3359,N_1207,N_1789);
xor U3360 (N_3360,N_610,N_290);
nand U3361 (N_3361,N_1294,N_1675);
xor U3362 (N_3362,N_608,N_2102);
nor U3363 (N_3363,N_1366,N_878);
nor U3364 (N_3364,N_1751,N_1231);
and U3365 (N_3365,N_1003,N_385);
nand U3366 (N_3366,N_2311,N_271);
nand U3367 (N_3367,N_1355,N_1508);
nor U3368 (N_3368,N_998,N_714);
nor U3369 (N_3369,N_427,N_478);
or U3370 (N_3370,N_650,N_1844);
nand U3371 (N_3371,N_2112,N_441);
nor U3372 (N_3372,N_1955,N_1199);
or U3373 (N_3373,N_1869,N_169);
xor U3374 (N_3374,N_471,N_2319);
and U3375 (N_3375,N_216,N_728);
xor U3376 (N_3376,N_2079,N_978);
nor U3377 (N_3377,N_1738,N_1149);
or U3378 (N_3378,N_1317,N_1276);
nand U3379 (N_3379,N_209,N_632);
nand U3380 (N_3380,N_1664,N_2429);
or U3381 (N_3381,N_1253,N_578);
or U3382 (N_3382,N_2362,N_1809);
nand U3383 (N_3383,N_120,N_1352);
nor U3384 (N_3384,N_166,N_2043);
and U3385 (N_3385,N_2468,N_2272);
nand U3386 (N_3386,N_515,N_2065);
nor U3387 (N_3387,N_1349,N_45);
nand U3388 (N_3388,N_316,N_499);
xor U3389 (N_3389,N_778,N_1263);
xnor U3390 (N_3390,N_329,N_1775);
nand U3391 (N_3391,N_2263,N_1525);
xor U3392 (N_3392,N_1886,N_1756);
and U3393 (N_3393,N_52,N_1236);
and U3394 (N_3394,N_1283,N_112);
or U3395 (N_3395,N_1744,N_1656);
nor U3396 (N_3396,N_2303,N_999);
or U3397 (N_3397,N_1505,N_2333);
nor U3398 (N_3398,N_1230,N_292);
and U3399 (N_3399,N_2123,N_2053);
or U3400 (N_3400,N_2196,N_1210);
nand U3401 (N_3401,N_1606,N_334);
nand U3402 (N_3402,N_1515,N_1466);
and U3403 (N_3403,N_2254,N_1432);
nand U3404 (N_3404,N_429,N_1318);
and U3405 (N_3405,N_815,N_490);
xnor U3406 (N_3406,N_2155,N_38);
nor U3407 (N_3407,N_840,N_1292);
xnor U3408 (N_3408,N_384,N_1684);
nand U3409 (N_3409,N_90,N_741);
or U3410 (N_3410,N_61,N_2);
or U3411 (N_3411,N_1727,N_2159);
and U3412 (N_3412,N_1274,N_1173);
or U3413 (N_3413,N_2034,N_696);
or U3414 (N_3414,N_910,N_371);
nor U3415 (N_3415,N_453,N_679);
xor U3416 (N_3416,N_461,N_303);
xnor U3417 (N_3417,N_1989,N_611);
nor U3418 (N_3418,N_614,N_2210);
and U3419 (N_3419,N_901,N_96);
xnor U3420 (N_3420,N_225,N_1024);
and U3421 (N_3421,N_968,N_1900);
xor U3422 (N_3422,N_629,N_2364);
or U3423 (N_3423,N_810,N_1202);
nand U3424 (N_3424,N_1858,N_1200);
nor U3425 (N_3425,N_360,N_1848);
or U3426 (N_3426,N_1553,N_302);
nor U3427 (N_3427,N_1010,N_156);
or U3428 (N_3428,N_498,N_960);
or U3429 (N_3429,N_1485,N_842);
xor U3430 (N_3430,N_1529,N_1655);
xor U3431 (N_3431,N_381,N_637);
and U3432 (N_3432,N_1391,N_2433);
or U3433 (N_3433,N_431,N_1760);
xor U3434 (N_3434,N_1544,N_1062);
nand U3435 (N_3435,N_1579,N_514);
and U3436 (N_3436,N_1434,N_1745);
xor U3437 (N_3437,N_439,N_393);
nand U3438 (N_3438,N_435,N_2222);
and U3439 (N_3439,N_1799,N_1451);
or U3440 (N_3440,N_362,N_2395);
or U3441 (N_3441,N_2093,N_2431);
nor U3442 (N_3442,N_2455,N_136);
xor U3443 (N_3443,N_617,N_2046);
nand U3444 (N_3444,N_2152,N_1151);
nand U3445 (N_3445,N_983,N_2075);
and U3446 (N_3446,N_660,N_838);
and U3447 (N_3447,N_508,N_192);
xor U3448 (N_3448,N_2372,N_766);
nor U3449 (N_3449,N_1680,N_1972);
xor U3450 (N_3450,N_1741,N_625);
nor U3451 (N_3451,N_2361,N_1383);
nand U3452 (N_3452,N_1167,N_2133);
nor U3453 (N_3453,N_665,N_2485);
or U3454 (N_3454,N_1550,N_2060);
xnor U3455 (N_3455,N_1329,N_123);
nand U3456 (N_3456,N_224,N_2432);
xor U3457 (N_3457,N_2275,N_2016);
or U3458 (N_3458,N_1336,N_1582);
nor U3459 (N_3459,N_469,N_791);
nand U3460 (N_3460,N_1827,N_785);
and U3461 (N_3461,N_1614,N_547);
nand U3462 (N_3462,N_486,N_726);
or U3463 (N_3463,N_507,N_1935);
nand U3464 (N_3464,N_2101,N_2021);
and U3465 (N_3465,N_1068,N_357);
xnor U3466 (N_3466,N_607,N_15);
or U3467 (N_3467,N_1819,N_715);
and U3468 (N_3468,N_1558,N_2262);
nand U3469 (N_3469,N_10,N_2365);
nand U3470 (N_3470,N_1755,N_1175);
nand U3471 (N_3471,N_1603,N_682);
nor U3472 (N_3472,N_2242,N_358);
xor U3473 (N_3473,N_1795,N_621);
and U3474 (N_3474,N_600,N_1975);
nand U3475 (N_3475,N_864,N_1816);
and U3476 (N_3476,N_2056,N_1772);
nand U3477 (N_3477,N_1889,N_41);
and U3478 (N_3478,N_226,N_818);
xnor U3479 (N_3479,N_1152,N_1984);
or U3480 (N_3480,N_816,N_2040);
nand U3481 (N_3481,N_1211,N_100);
xor U3482 (N_3482,N_1241,N_2209);
xnor U3483 (N_3483,N_666,N_370);
nand U3484 (N_3484,N_509,N_1144);
or U3485 (N_3485,N_2138,N_2295);
and U3486 (N_3486,N_279,N_1414);
xnor U3487 (N_3487,N_152,N_2012);
or U3488 (N_3488,N_20,N_178);
or U3489 (N_3489,N_50,N_622);
nand U3490 (N_3490,N_466,N_74);
nand U3491 (N_3491,N_2479,N_236);
or U3492 (N_3492,N_132,N_887);
or U3493 (N_3493,N_2247,N_631);
nor U3494 (N_3494,N_1835,N_116);
nand U3495 (N_3495,N_2193,N_2475);
xor U3496 (N_3496,N_1250,N_2207);
nand U3497 (N_3497,N_1125,N_982);
nor U3498 (N_3498,N_2135,N_1617);
nand U3499 (N_3499,N_428,N_2027);
nor U3500 (N_3500,N_160,N_1044);
nor U3501 (N_3501,N_269,N_1278);
or U3502 (N_3502,N_2494,N_639);
xor U3503 (N_3503,N_1132,N_2022);
nor U3504 (N_3504,N_2178,N_1172);
xnor U3505 (N_3505,N_528,N_1807);
xor U3506 (N_3506,N_1463,N_1229);
nand U3507 (N_3507,N_858,N_2005);
or U3508 (N_3508,N_2280,N_2418);
and U3509 (N_3509,N_1542,N_25);
xnor U3510 (N_3510,N_1500,N_95);
and U3511 (N_3511,N_451,N_1496);
and U3512 (N_3512,N_510,N_416);
and U3513 (N_3513,N_2349,N_396);
nor U3514 (N_3514,N_918,N_46);
xor U3515 (N_3515,N_627,N_1938);
nor U3516 (N_3516,N_2371,N_464);
nand U3517 (N_3517,N_424,N_764);
nand U3518 (N_3518,N_1118,N_2144);
and U3519 (N_3519,N_2085,N_1190);
nand U3520 (N_3520,N_1764,N_1296);
and U3521 (N_3521,N_606,N_1101);
and U3522 (N_3522,N_174,N_1251);
xnor U3523 (N_3523,N_2491,N_2357);
or U3524 (N_3524,N_812,N_1115);
and U3525 (N_3525,N_1730,N_2227);
nor U3526 (N_3526,N_2162,N_1639);
xnor U3527 (N_3527,N_1074,N_2428);
or U3528 (N_3528,N_1793,N_2421);
nor U3529 (N_3529,N_2414,N_230);
or U3530 (N_3530,N_734,N_1146);
or U3531 (N_3531,N_397,N_252);
nor U3532 (N_3532,N_2069,N_2377);
and U3533 (N_3533,N_491,N_591);
and U3534 (N_3534,N_1568,N_2309);
nor U3535 (N_3535,N_2426,N_534);
nor U3536 (N_3536,N_2370,N_2374);
nor U3537 (N_3537,N_2223,N_796);
or U3538 (N_3538,N_2214,N_941);
or U3539 (N_3539,N_204,N_2004);
xor U3540 (N_3540,N_40,N_1435);
or U3541 (N_3541,N_194,N_1590);
xnor U3542 (N_3542,N_1682,N_2493);
xnor U3543 (N_3543,N_2158,N_2353);
or U3544 (N_3544,N_13,N_99);
xnor U3545 (N_3545,N_470,N_585);
xnor U3546 (N_3546,N_1974,N_168);
xnor U3547 (N_3547,N_1316,N_28);
nor U3548 (N_3548,N_2095,N_560);
nor U3549 (N_3549,N_1290,N_1853);
or U3550 (N_3550,N_1725,N_18);
and U3551 (N_3551,N_2195,N_777);
nand U3552 (N_3552,N_2317,N_2497);
xor U3553 (N_3553,N_1378,N_1177);
nor U3554 (N_3554,N_1862,N_1194);
or U3555 (N_3555,N_604,N_260);
xor U3556 (N_3556,N_797,N_654);
or U3557 (N_3557,N_359,N_1000);
and U3558 (N_3558,N_2184,N_150);
nand U3559 (N_3559,N_1893,N_2212);
and U3560 (N_3560,N_2378,N_744);
or U3561 (N_3561,N_452,N_1980);
nor U3562 (N_3562,N_1883,N_1674);
or U3563 (N_3563,N_2078,N_1291);
and U3564 (N_3564,N_905,N_93);
or U3565 (N_3565,N_2224,N_1287);
or U3566 (N_3566,N_1371,N_537);
nand U3567 (N_3567,N_468,N_788);
and U3568 (N_3568,N_2017,N_83);
nor U3569 (N_3569,N_2385,N_830);
nor U3570 (N_3570,N_1771,N_1903);
and U3571 (N_3571,N_856,N_129);
and U3572 (N_3572,N_1833,N_1224);
and U3573 (N_3573,N_2478,N_2077);
nor U3574 (N_3574,N_1042,N_2243);
and U3575 (N_3575,N_957,N_545);
nor U3576 (N_3576,N_900,N_852);
xor U3577 (N_3577,N_1706,N_1275);
or U3578 (N_3578,N_1584,N_107);
xnor U3579 (N_3579,N_872,N_1016);
and U3580 (N_3580,N_711,N_1927);
nand U3581 (N_3581,N_2164,N_276);
nand U3582 (N_3582,N_1923,N_1422);
xnor U3583 (N_3583,N_1458,N_2117);
or U3584 (N_3584,N_523,N_39);
xor U3585 (N_3585,N_285,N_536);
xor U3586 (N_3586,N_1983,N_1531);
or U3587 (N_3587,N_1353,N_1696);
xnor U3588 (N_3588,N_2422,N_196);
xnor U3589 (N_3589,N_551,N_1060);
nor U3590 (N_3590,N_355,N_1805);
nor U3591 (N_3591,N_952,N_1767);
nor U3592 (N_3592,N_2439,N_185);
nor U3593 (N_3593,N_2367,N_924);
nand U3594 (N_3594,N_127,N_1372);
and U3595 (N_3595,N_1802,N_2386);
xor U3596 (N_3596,N_1918,N_1587);
or U3597 (N_3597,N_2293,N_1021);
or U3598 (N_3598,N_417,N_145);
xnor U3599 (N_3599,N_692,N_1517);
nor U3600 (N_3600,N_977,N_1335);
and U3601 (N_3601,N_1300,N_811);
or U3602 (N_3602,N_1734,N_685);
xor U3603 (N_3603,N_2171,N_488);
or U3604 (N_3604,N_1418,N_379);
and U3605 (N_3605,N_2205,N_2325);
and U3606 (N_3606,N_691,N_1204);
nand U3607 (N_3607,N_652,N_2270);
nor U3608 (N_3608,N_1778,N_992);
nand U3609 (N_3609,N_139,N_2186);
nand U3610 (N_3610,N_1497,N_846);
and U3611 (N_3611,N_2274,N_66);
xor U3612 (N_3612,N_2402,N_2286);
nand U3613 (N_3613,N_2477,N_1878);
nand U3614 (N_3614,N_1888,N_2322);
and U3615 (N_3615,N_1541,N_257);
nand U3616 (N_3616,N_89,N_2103);
and U3617 (N_3617,N_1623,N_1774);
and U3618 (N_3618,N_1382,N_270);
nand U3619 (N_3619,N_819,N_1470);
and U3620 (N_3620,N_2350,N_450);
and U3621 (N_3621,N_2393,N_934);
nor U3622 (N_3622,N_1049,N_1479);
or U3623 (N_3623,N_656,N_17);
or U3624 (N_3624,N_369,N_803);
and U3625 (N_3625,N_723,N_2483);
nand U3626 (N_3626,N_1501,N_2245);
and U3627 (N_3627,N_1924,N_1301);
and U3628 (N_3628,N_1436,N_115);
xnor U3629 (N_3629,N_2211,N_1957);
nand U3630 (N_3630,N_843,N_1284);
and U3631 (N_3631,N_35,N_286);
and U3632 (N_3632,N_102,N_505);
nor U3633 (N_3633,N_2145,N_1288);
nand U3634 (N_3634,N_1005,N_1628);
xnor U3635 (N_3635,N_1669,N_1379);
nand U3636 (N_3636,N_1002,N_496);
nor U3637 (N_3637,N_1507,N_1821);
nor U3638 (N_3638,N_2420,N_382);
nand U3639 (N_3639,N_847,N_540);
xor U3640 (N_3640,N_698,N_1376);
nor U3641 (N_3641,N_776,N_1510);
nor U3642 (N_3642,N_1363,N_2490);
nor U3643 (N_3643,N_85,N_768);
nor U3644 (N_3644,N_1228,N_2430);
or U3645 (N_3645,N_2296,N_1314);
or U3646 (N_3646,N_1285,N_841);
nor U3647 (N_3647,N_1506,N_1009);
and U3648 (N_3648,N_2341,N_2476);
nor U3649 (N_3649,N_2234,N_1581);
and U3650 (N_3650,N_1812,N_546);
or U3651 (N_3651,N_1612,N_2281);
xor U3652 (N_3652,N_554,N_2174);
and U3653 (N_3653,N_19,N_1388);
and U3654 (N_3654,N_202,N_354);
and U3655 (N_3655,N_1747,N_2482);
nand U3656 (N_3656,N_805,N_1859);
nor U3657 (N_3657,N_1642,N_1480);
nor U3658 (N_3658,N_1901,N_1135);
nand U3659 (N_3659,N_1717,N_1059);
nand U3660 (N_3660,N_2054,N_2108);
xnor U3661 (N_3661,N_1952,N_2129);
and U3662 (N_3662,N_1894,N_833);
nor U3663 (N_3663,N_1277,N_222);
and U3664 (N_3664,N_1943,N_956);
and U3665 (N_3665,N_2401,N_2495);
xor U3666 (N_3666,N_364,N_1139);
nand U3667 (N_3667,N_1430,N_1475);
nor U3668 (N_3668,N_1516,N_228);
or U3669 (N_3669,N_2347,N_733);
or U3670 (N_3670,N_207,N_1247);
or U3671 (N_3671,N_620,N_1242);
xor U3672 (N_3672,N_212,N_2324);
or U3673 (N_3673,N_1072,N_985);
xor U3674 (N_3674,N_1665,N_729);
or U3675 (N_3675,N_1323,N_1910);
and U3676 (N_3676,N_110,N_1209);
xor U3677 (N_3677,N_75,N_909);
xor U3678 (N_3678,N_2396,N_592);
nand U3679 (N_3679,N_860,N_1513);
nor U3680 (N_3680,N_31,N_97);
xnor U3681 (N_3681,N_767,N_1712);
and U3682 (N_3682,N_43,N_2298);
or U3683 (N_3683,N_1077,N_1126);
xnor U3684 (N_3684,N_1474,N_553);
and U3685 (N_3685,N_201,N_1262);
or U3686 (N_3686,N_283,N_2473);
nand U3687 (N_3687,N_2240,N_2007);
nor U3688 (N_3688,N_2358,N_1472);
xnor U3689 (N_3689,N_1071,N_1134);
or U3690 (N_3690,N_702,N_1657);
or U3691 (N_3691,N_1790,N_1996);
and U3692 (N_3692,N_869,N_1057);
nand U3693 (N_3693,N_565,N_2257);
nand U3694 (N_3694,N_2244,N_2188);
or U3695 (N_3695,N_884,N_2474);
nor U3696 (N_3696,N_1999,N_1197);
and U3697 (N_3697,N_1604,N_1985);
or U3698 (N_3698,N_1630,N_135);
and U3699 (N_3699,N_389,N_914);
xnor U3700 (N_3700,N_1142,N_1634);
or U3701 (N_3701,N_108,N_945);
nor U3702 (N_3702,N_1711,N_176);
or U3703 (N_3703,N_1708,N_1227);
xor U3704 (N_3704,N_2360,N_1235);
or U3705 (N_3705,N_1737,N_2301);
xnor U3706 (N_3706,N_1701,N_775);
xnor U3707 (N_3707,N_1083,N_182);
nor U3708 (N_3708,N_1780,N_1417);
or U3709 (N_3709,N_2292,N_1700);
nand U3710 (N_3710,N_199,N_1255);
nor U3711 (N_3711,N_892,N_1672);
or U3712 (N_3712,N_273,N_1094);
or U3713 (N_3713,N_1954,N_365);
or U3714 (N_3714,N_1160,N_1874);
nand U3715 (N_3715,N_1222,N_1103);
xnor U3716 (N_3716,N_170,N_1477);
or U3717 (N_3717,N_1369,N_298);
xor U3718 (N_3718,N_1536,N_1831);
nor U3719 (N_3719,N_1293,N_522);
xor U3720 (N_3720,N_104,N_925);
nand U3721 (N_3721,N_969,N_527);
xnor U3722 (N_3722,N_2204,N_880);
and U3723 (N_3723,N_1982,N_773);
or U3724 (N_3724,N_1555,N_1887);
nor U3725 (N_3725,N_2379,N_544);
nor U3726 (N_3726,N_1014,N_183);
and U3727 (N_3727,N_2329,N_1120);
nor U3728 (N_3728,N_1012,N_879);
and U3729 (N_3729,N_111,N_1055);
xor U3730 (N_3730,N_984,N_1534);
and U3731 (N_3731,N_2437,N_927);
xnor U3732 (N_3732,N_789,N_1920);
xor U3733 (N_3733,N_1240,N_1520);
and U3734 (N_3734,N_2024,N_2213);
or U3735 (N_3735,N_1803,N_1560);
nand U3736 (N_3736,N_1212,N_1437);
xor U3737 (N_3737,N_1762,N_503);
or U3738 (N_3738,N_862,N_1882);
xnor U3739 (N_3739,N_1545,N_1415);
and U3740 (N_3740,N_2148,N_2051);
nand U3741 (N_3741,N_907,N_1129);
nand U3742 (N_3742,N_22,N_1946);
and U3743 (N_3743,N_1041,N_2068);
or U3744 (N_3744,N_1362,N_2143);
or U3745 (N_3745,N_2388,N_440);
and U3746 (N_3746,N_2182,N_898);
nand U3747 (N_3747,N_2452,N_827);
and U3748 (N_3748,N_77,N_926);
and U3749 (N_3749,N_1618,N_425);
and U3750 (N_3750,N_1302,N_67);
and U3751 (N_3751,N_17,N_776);
nor U3752 (N_3752,N_446,N_1972);
xor U3753 (N_3753,N_73,N_1923);
or U3754 (N_3754,N_1738,N_612);
nor U3755 (N_3755,N_1442,N_520);
or U3756 (N_3756,N_2387,N_1183);
xnor U3757 (N_3757,N_1809,N_658);
and U3758 (N_3758,N_1874,N_30);
and U3759 (N_3759,N_758,N_138);
and U3760 (N_3760,N_127,N_1991);
xnor U3761 (N_3761,N_318,N_968);
or U3762 (N_3762,N_448,N_2235);
or U3763 (N_3763,N_278,N_1130);
xor U3764 (N_3764,N_798,N_797);
nand U3765 (N_3765,N_1534,N_2066);
nand U3766 (N_3766,N_1929,N_1373);
nand U3767 (N_3767,N_2454,N_2087);
or U3768 (N_3768,N_587,N_1852);
and U3769 (N_3769,N_1489,N_885);
xnor U3770 (N_3770,N_585,N_185);
xnor U3771 (N_3771,N_2099,N_2453);
nand U3772 (N_3772,N_2457,N_455);
nand U3773 (N_3773,N_1086,N_936);
nor U3774 (N_3774,N_1040,N_1324);
nand U3775 (N_3775,N_2158,N_1202);
xor U3776 (N_3776,N_266,N_250);
or U3777 (N_3777,N_2444,N_45);
nor U3778 (N_3778,N_635,N_2045);
and U3779 (N_3779,N_396,N_58);
nand U3780 (N_3780,N_543,N_2147);
nor U3781 (N_3781,N_993,N_1182);
and U3782 (N_3782,N_2003,N_1634);
or U3783 (N_3783,N_1276,N_1536);
and U3784 (N_3784,N_1331,N_2179);
and U3785 (N_3785,N_239,N_2356);
nor U3786 (N_3786,N_2056,N_2489);
nor U3787 (N_3787,N_1492,N_1052);
xor U3788 (N_3788,N_822,N_111);
nand U3789 (N_3789,N_671,N_2443);
xor U3790 (N_3790,N_635,N_1808);
or U3791 (N_3791,N_564,N_410);
and U3792 (N_3792,N_417,N_1732);
and U3793 (N_3793,N_774,N_1263);
nand U3794 (N_3794,N_713,N_1676);
and U3795 (N_3795,N_715,N_1947);
nor U3796 (N_3796,N_1787,N_2100);
and U3797 (N_3797,N_2171,N_1997);
nand U3798 (N_3798,N_1094,N_2492);
nor U3799 (N_3799,N_2097,N_1269);
nand U3800 (N_3800,N_185,N_337);
and U3801 (N_3801,N_1695,N_1181);
or U3802 (N_3802,N_1266,N_1891);
or U3803 (N_3803,N_1067,N_1335);
nand U3804 (N_3804,N_1268,N_218);
or U3805 (N_3805,N_285,N_955);
nand U3806 (N_3806,N_1315,N_66);
nand U3807 (N_3807,N_419,N_363);
xnor U3808 (N_3808,N_513,N_1942);
nand U3809 (N_3809,N_1073,N_1667);
nor U3810 (N_3810,N_2150,N_319);
or U3811 (N_3811,N_502,N_942);
nand U3812 (N_3812,N_101,N_1048);
xor U3813 (N_3813,N_1915,N_941);
nand U3814 (N_3814,N_102,N_178);
nor U3815 (N_3815,N_827,N_724);
nand U3816 (N_3816,N_1571,N_1863);
nor U3817 (N_3817,N_348,N_881);
nand U3818 (N_3818,N_2265,N_1424);
and U3819 (N_3819,N_1983,N_22);
or U3820 (N_3820,N_2389,N_1518);
nand U3821 (N_3821,N_1123,N_1753);
xor U3822 (N_3822,N_327,N_1291);
nor U3823 (N_3823,N_937,N_431);
nand U3824 (N_3824,N_435,N_633);
xor U3825 (N_3825,N_1637,N_2042);
and U3826 (N_3826,N_1039,N_1783);
nor U3827 (N_3827,N_375,N_898);
xnor U3828 (N_3828,N_1280,N_1166);
or U3829 (N_3829,N_598,N_196);
xnor U3830 (N_3830,N_2205,N_354);
or U3831 (N_3831,N_2123,N_39);
xor U3832 (N_3832,N_1330,N_1032);
and U3833 (N_3833,N_1016,N_688);
or U3834 (N_3834,N_349,N_391);
nor U3835 (N_3835,N_2322,N_2180);
nor U3836 (N_3836,N_1418,N_729);
and U3837 (N_3837,N_781,N_2);
nand U3838 (N_3838,N_1475,N_221);
nor U3839 (N_3839,N_1992,N_1786);
or U3840 (N_3840,N_915,N_1895);
xnor U3841 (N_3841,N_309,N_1053);
nand U3842 (N_3842,N_378,N_1554);
and U3843 (N_3843,N_381,N_789);
and U3844 (N_3844,N_2378,N_125);
nor U3845 (N_3845,N_1081,N_1969);
nor U3846 (N_3846,N_1463,N_2084);
xnor U3847 (N_3847,N_641,N_351);
or U3848 (N_3848,N_1788,N_2283);
xnor U3849 (N_3849,N_931,N_724);
or U3850 (N_3850,N_1210,N_187);
and U3851 (N_3851,N_679,N_637);
nor U3852 (N_3852,N_1609,N_800);
nand U3853 (N_3853,N_1524,N_2292);
nor U3854 (N_3854,N_599,N_1922);
xor U3855 (N_3855,N_1989,N_1594);
and U3856 (N_3856,N_1872,N_1142);
and U3857 (N_3857,N_1955,N_200);
or U3858 (N_3858,N_92,N_1470);
nor U3859 (N_3859,N_2066,N_303);
and U3860 (N_3860,N_1372,N_1666);
nand U3861 (N_3861,N_1286,N_1688);
and U3862 (N_3862,N_1971,N_1035);
nor U3863 (N_3863,N_2089,N_300);
or U3864 (N_3864,N_916,N_2224);
or U3865 (N_3865,N_587,N_996);
nor U3866 (N_3866,N_86,N_1099);
and U3867 (N_3867,N_828,N_1911);
or U3868 (N_3868,N_557,N_29);
xnor U3869 (N_3869,N_1451,N_1974);
or U3870 (N_3870,N_2173,N_574);
or U3871 (N_3871,N_717,N_2106);
or U3872 (N_3872,N_2194,N_1009);
nand U3873 (N_3873,N_72,N_1168);
and U3874 (N_3874,N_1010,N_856);
or U3875 (N_3875,N_2367,N_2004);
xor U3876 (N_3876,N_1015,N_2051);
and U3877 (N_3877,N_532,N_2072);
xor U3878 (N_3878,N_1612,N_1062);
nor U3879 (N_3879,N_1486,N_1718);
nand U3880 (N_3880,N_525,N_632);
nand U3881 (N_3881,N_2272,N_561);
nor U3882 (N_3882,N_1941,N_1269);
and U3883 (N_3883,N_2490,N_165);
xnor U3884 (N_3884,N_618,N_327);
xnor U3885 (N_3885,N_2107,N_2255);
nand U3886 (N_3886,N_878,N_1814);
nand U3887 (N_3887,N_2142,N_192);
or U3888 (N_3888,N_505,N_499);
xor U3889 (N_3889,N_1593,N_576);
xnor U3890 (N_3890,N_1975,N_1021);
xnor U3891 (N_3891,N_1409,N_1084);
nand U3892 (N_3892,N_1848,N_1780);
nand U3893 (N_3893,N_1492,N_240);
or U3894 (N_3894,N_212,N_371);
nor U3895 (N_3895,N_927,N_1947);
and U3896 (N_3896,N_929,N_2194);
or U3897 (N_3897,N_462,N_2007);
xor U3898 (N_3898,N_2156,N_173);
nand U3899 (N_3899,N_1301,N_1393);
and U3900 (N_3900,N_114,N_1902);
nand U3901 (N_3901,N_1421,N_1892);
nand U3902 (N_3902,N_1325,N_1295);
nand U3903 (N_3903,N_1989,N_10);
or U3904 (N_3904,N_2226,N_384);
nor U3905 (N_3905,N_817,N_234);
or U3906 (N_3906,N_1192,N_1925);
xor U3907 (N_3907,N_903,N_1688);
and U3908 (N_3908,N_1417,N_2471);
nor U3909 (N_3909,N_147,N_1204);
nor U3910 (N_3910,N_801,N_2494);
xnor U3911 (N_3911,N_1667,N_39);
or U3912 (N_3912,N_2265,N_1597);
or U3913 (N_3913,N_2364,N_83);
or U3914 (N_3914,N_1747,N_328);
nor U3915 (N_3915,N_641,N_2417);
and U3916 (N_3916,N_186,N_2343);
and U3917 (N_3917,N_161,N_454);
and U3918 (N_3918,N_2210,N_717);
nand U3919 (N_3919,N_2474,N_945);
nand U3920 (N_3920,N_37,N_2244);
and U3921 (N_3921,N_1712,N_902);
nor U3922 (N_3922,N_1736,N_2334);
and U3923 (N_3923,N_2262,N_10);
nand U3924 (N_3924,N_53,N_1604);
and U3925 (N_3925,N_355,N_2366);
and U3926 (N_3926,N_1395,N_1418);
xnor U3927 (N_3927,N_2163,N_2193);
nor U3928 (N_3928,N_1619,N_836);
nand U3929 (N_3929,N_1486,N_1682);
or U3930 (N_3930,N_922,N_527);
nor U3931 (N_3931,N_1787,N_2025);
nand U3932 (N_3932,N_1144,N_1207);
and U3933 (N_3933,N_1898,N_855);
and U3934 (N_3934,N_1825,N_1646);
and U3935 (N_3935,N_2069,N_832);
nor U3936 (N_3936,N_1056,N_2385);
nor U3937 (N_3937,N_1541,N_1948);
nor U3938 (N_3938,N_150,N_789);
nand U3939 (N_3939,N_2414,N_975);
xnor U3940 (N_3940,N_2473,N_787);
nor U3941 (N_3941,N_63,N_1008);
xnor U3942 (N_3942,N_404,N_772);
or U3943 (N_3943,N_1199,N_1136);
nand U3944 (N_3944,N_1748,N_1965);
nand U3945 (N_3945,N_1943,N_367);
nand U3946 (N_3946,N_1016,N_1209);
xnor U3947 (N_3947,N_981,N_2299);
nor U3948 (N_3948,N_1044,N_1342);
xnor U3949 (N_3949,N_667,N_1745);
xor U3950 (N_3950,N_1120,N_1553);
nor U3951 (N_3951,N_292,N_586);
nor U3952 (N_3952,N_1615,N_1380);
and U3953 (N_3953,N_1757,N_1281);
xor U3954 (N_3954,N_2437,N_1369);
xor U3955 (N_3955,N_305,N_948);
nor U3956 (N_3956,N_2125,N_1960);
and U3957 (N_3957,N_1603,N_2207);
or U3958 (N_3958,N_2071,N_1471);
nor U3959 (N_3959,N_612,N_538);
nor U3960 (N_3960,N_1589,N_1833);
xnor U3961 (N_3961,N_771,N_1739);
xor U3962 (N_3962,N_433,N_1131);
or U3963 (N_3963,N_2347,N_167);
nor U3964 (N_3964,N_1384,N_2336);
nand U3965 (N_3965,N_1679,N_2064);
and U3966 (N_3966,N_2290,N_254);
nor U3967 (N_3967,N_418,N_1924);
xor U3968 (N_3968,N_1385,N_1604);
and U3969 (N_3969,N_949,N_1768);
nand U3970 (N_3970,N_1800,N_1593);
and U3971 (N_3971,N_302,N_2365);
nand U3972 (N_3972,N_933,N_1844);
nor U3973 (N_3973,N_1077,N_1976);
xor U3974 (N_3974,N_868,N_925);
nor U3975 (N_3975,N_377,N_205);
xor U3976 (N_3976,N_1106,N_1423);
nor U3977 (N_3977,N_2487,N_2111);
nand U3978 (N_3978,N_690,N_1327);
and U3979 (N_3979,N_916,N_539);
nor U3980 (N_3980,N_1012,N_2004);
and U3981 (N_3981,N_1288,N_975);
and U3982 (N_3982,N_277,N_1947);
nand U3983 (N_3983,N_403,N_275);
xor U3984 (N_3984,N_1365,N_2115);
or U3985 (N_3985,N_926,N_1955);
and U3986 (N_3986,N_1971,N_1473);
xnor U3987 (N_3987,N_1596,N_1801);
or U3988 (N_3988,N_914,N_58);
or U3989 (N_3989,N_2035,N_1418);
xor U3990 (N_3990,N_633,N_1581);
xnor U3991 (N_3991,N_2235,N_697);
xor U3992 (N_3992,N_1849,N_848);
or U3993 (N_3993,N_1741,N_1596);
and U3994 (N_3994,N_1013,N_734);
nand U3995 (N_3995,N_2185,N_2039);
nor U3996 (N_3996,N_1207,N_1281);
and U3997 (N_3997,N_1048,N_92);
and U3998 (N_3998,N_2037,N_2418);
or U3999 (N_3999,N_1654,N_2034);
and U4000 (N_4000,N_1924,N_1397);
and U4001 (N_4001,N_2075,N_2252);
xor U4002 (N_4002,N_1974,N_465);
nand U4003 (N_4003,N_1039,N_753);
and U4004 (N_4004,N_78,N_428);
and U4005 (N_4005,N_1706,N_651);
or U4006 (N_4006,N_52,N_1914);
nor U4007 (N_4007,N_708,N_1199);
or U4008 (N_4008,N_812,N_392);
or U4009 (N_4009,N_537,N_581);
nor U4010 (N_4010,N_1787,N_1349);
and U4011 (N_4011,N_2063,N_2106);
xor U4012 (N_4012,N_833,N_655);
xor U4013 (N_4013,N_435,N_1948);
nor U4014 (N_4014,N_921,N_1300);
and U4015 (N_4015,N_2066,N_241);
xor U4016 (N_4016,N_1295,N_1553);
nand U4017 (N_4017,N_2116,N_1542);
nor U4018 (N_4018,N_529,N_1106);
xor U4019 (N_4019,N_331,N_1350);
or U4020 (N_4020,N_1030,N_170);
and U4021 (N_4021,N_2282,N_1017);
or U4022 (N_4022,N_2474,N_237);
nand U4023 (N_4023,N_2389,N_1665);
xnor U4024 (N_4024,N_487,N_878);
nand U4025 (N_4025,N_1668,N_736);
and U4026 (N_4026,N_592,N_960);
xnor U4027 (N_4027,N_748,N_1680);
xor U4028 (N_4028,N_166,N_1661);
nand U4029 (N_4029,N_1533,N_255);
and U4030 (N_4030,N_1747,N_2252);
or U4031 (N_4031,N_1222,N_1145);
and U4032 (N_4032,N_337,N_730);
nor U4033 (N_4033,N_2055,N_526);
xor U4034 (N_4034,N_1586,N_562);
or U4035 (N_4035,N_1990,N_2043);
xnor U4036 (N_4036,N_1186,N_1517);
or U4037 (N_4037,N_2162,N_1457);
or U4038 (N_4038,N_1651,N_1558);
nor U4039 (N_4039,N_1653,N_1651);
and U4040 (N_4040,N_1044,N_257);
or U4041 (N_4041,N_2422,N_1888);
xor U4042 (N_4042,N_1056,N_311);
or U4043 (N_4043,N_1353,N_1652);
xor U4044 (N_4044,N_1765,N_927);
or U4045 (N_4045,N_343,N_1706);
nor U4046 (N_4046,N_1846,N_2218);
or U4047 (N_4047,N_1238,N_2283);
nor U4048 (N_4048,N_2343,N_2428);
nor U4049 (N_4049,N_2066,N_586);
nand U4050 (N_4050,N_143,N_183);
and U4051 (N_4051,N_765,N_1668);
or U4052 (N_4052,N_1283,N_1855);
nand U4053 (N_4053,N_1435,N_300);
xnor U4054 (N_4054,N_108,N_2368);
nor U4055 (N_4055,N_1584,N_1850);
nor U4056 (N_4056,N_812,N_781);
and U4057 (N_4057,N_283,N_1527);
xor U4058 (N_4058,N_1826,N_1496);
or U4059 (N_4059,N_410,N_879);
xor U4060 (N_4060,N_2146,N_2288);
or U4061 (N_4061,N_1850,N_1054);
nor U4062 (N_4062,N_2152,N_47);
or U4063 (N_4063,N_1042,N_2376);
xor U4064 (N_4064,N_2434,N_1508);
or U4065 (N_4065,N_1843,N_2171);
nor U4066 (N_4066,N_1839,N_2179);
nor U4067 (N_4067,N_2173,N_415);
nand U4068 (N_4068,N_1549,N_551);
nand U4069 (N_4069,N_311,N_1683);
nor U4070 (N_4070,N_1297,N_625);
and U4071 (N_4071,N_344,N_211);
or U4072 (N_4072,N_2099,N_1285);
nor U4073 (N_4073,N_1934,N_230);
or U4074 (N_4074,N_1083,N_2190);
nand U4075 (N_4075,N_791,N_1465);
nand U4076 (N_4076,N_1249,N_1818);
nor U4077 (N_4077,N_1079,N_2467);
xor U4078 (N_4078,N_127,N_1633);
and U4079 (N_4079,N_2350,N_814);
xnor U4080 (N_4080,N_1072,N_164);
xor U4081 (N_4081,N_664,N_2372);
xor U4082 (N_4082,N_2030,N_1206);
and U4083 (N_4083,N_2443,N_495);
nand U4084 (N_4084,N_1080,N_2307);
nor U4085 (N_4085,N_1574,N_2262);
and U4086 (N_4086,N_2250,N_1597);
nor U4087 (N_4087,N_1571,N_2277);
or U4088 (N_4088,N_1041,N_2491);
xnor U4089 (N_4089,N_386,N_907);
nor U4090 (N_4090,N_2254,N_1576);
xor U4091 (N_4091,N_2432,N_1418);
nand U4092 (N_4092,N_1341,N_1756);
nand U4093 (N_4093,N_2439,N_1516);
nand U4094 (N_4094,N_1869,N_259);
nand U4095 (N_4095,N_1444,N_2422);
xor U4096 (N_4096,N_124,N_516);
nand U4097 (N_4097,N_2428,N_1113);
xnor U4098 (N_4098,N_1649,N_660);
or U4099 (N_4099,N_1446,N_2327);
or U4100 (N_4100,N_2285,N_1318);
or U4101 (N_4101,N_1547,N_157);
nand U4102 (N_4102,N_2470,N_1334);
nor U4103 (N_4103,N_284,N_1665);
nand U4104 (N_4104,N_2089,N_33);
xor U4105 (N_4105,N_293,N_2432);
nand U4106 (N_4106,N_125,N_1377);
and U4107 (N_4107,N_989,N_1940);
nor U4108 (N_4108,N_320,N_708);
nand U4109 (N_4109,N_1280,N_150);
nand U4110 (N_4110,N_316,N_1292);
nand U4111 (N_4111,N_1528,N_1697);
xor U4112 (N_4112,N_2071,N_932);
nand U4113 (N_4113,N_734,N_2045);
nor U4114 (N_4114,N_1663,N_809);
or U4115 (N_4115,N_644,N_1029);
nand U4116 (N_4116,N_1079,N_265);
or U4117 (N_4117,N_1792,N_1075);
or U4118 (N_4118,N_895,N_1961);
nand U4119 (N_4119,N_1591,N_884);
xor U4120 (N_4120,N_1247,N_274);
nand U4121 (N_4121,N_1337,N_1685);
nand U4122 (N_4122,N_2204,N_1167);
xnor U4123 (N_4123,N_2412,N_1583);
nand U4124 (N_4124,N_167,N_203);
and U4125 (N_4125,N_2471,N_1919);
and U4126 (N_4126,N_563,N_2094);
nor U4127 (N_4127,N_457,N_364);
nor U4128 (N_4128,N_2191,N_467);
xnor U4129 (N_4129,N_555,N_2080);
nand U4130 (N_4130,N_246,N_1503);
nor U4131 (N_4131,N_878,N_1536);
and U4132 (N_4132,N_55,N_2166);
or U4133 (N_4133,N_86,N_558);
nand U4134 (N_4134,N_623,N_987);
xor U4135 (N_4135,N_138,N_153);
or U4136 (N_4136,N_1779,N_1249);
nand U4137 (N_4137,N_1586,N_1488);
or U4138 (N_4138,N_1692,N_1628);
xor U4139 (N_4139,N_2112,N_1166);
nand U4140 (N_4140,N_1436,N_2065);
or U4141 (N_4141,N_184,N_1170);
or U4142 (N_4142,N_2436,N_2378);
xnor U4143 (N_4143,N_1173,N_804);
and U4144 (N_4144,N_715,N_1986);
xnor U4145 (N_4145,N_200,N_1986);
nand U4146 (N_4146,N_1787,N_2213);
nor U4147 (N_4147,N_1429,N_1536);
nand U4148 (N_4148,N_1542,N_494);
and U4149 (N_4149,N_2462,N_1489);
and U4150 (N_4150,N_348,N_2392);
xor U4151 (N_4151,N_2289,N_2327);
or U4152 (N_4152,N_1338,N_2436);
nand U4153 (N_4153,N_808,N_64);
or U4154 (N_4154,N_2248,N_1732);
xor U4155 (N_4155,N_2033,N_2431);
nand U4156 (N_4156,N_1382,N_1506);
or U4157 (N_4157,N_554,N_1404);
nor U4158 (N_4158,N_1754,N_223);
nor U4159 (N_4159,N_1675,N_896);
or U4160 (N_4160,N_997,N_1868);
and U4161 (N_4161,N_893,N_1910);
xnor U4162 (N_4162,N_1574,N_147);
or U4163 (N_4163,N_2434,N_2103);
or U4164 (N_4164,N_960,N_2305);
or U4165 (N_4165,N_851,N_22);
or U4166 (N_4166,N_512,N_848);
nor U4167 (N_4167,N_519,N_1826);
nand U4168 (N_4168,N_1289,N_1373);
xnor U4169 (N_4169,N_1450,N_2094);
nor U4170 (N_4170,N_1412,N_2311);
and U4171 (N_4171,N_896,N_2199);
or U4172 (N_4172,N_389,N_1489);
nor U4173 (N_4173,N_1568,N_2269);
or U4174 (N_4174,N_1529,N_1695);
or U4175 (N_4175,N_507,N_2203);
nor U4176 (N_4176,N_443,N_1174);
nor U4177 (N_4177,N_951,N_1109);
xnor U4178 (N_4178,N_59,N_1944);
xnor U4179 (N_4179,N_444,N_20);
and U4180 (N_4180,N_2476,N_2321);
or U4181 (N_4181,N_2461,N_1569);
or U4182 (N_4182,N_1167,N_582);
nor U4183 (N_4183,N_938,N_896);
nor U4184 (N_4184,N_480,N_623);
nand U4185 (N_4185,N_1567,N_630);
nand U4186 (N_4186,N_1275,N_2272);
nor U4187 (N_4187,N_1359,N_1845);
nand U4188 (N_4188,N_2031,N_18);
or U4189 (N_4189,N_1261,N_2443);
xnor U4190 (N_4190,N_526,N_637);
nand U4191 (N_4191,N_1207,N_551);
and U4192 (N_4192,N_999,N_1015);
or U4193 (N_4193,N_434,N_739);
nor U4194 (N_4194,N_1395,N_1467);
nand U4195 (N_4195,N_2338,N_1563);
nand U4196 (N_4196,N_1228,N_1281);
and U4197 (N_4197,N_1584,N_2148);
and U4198 (N_4198,N_439,N_1532);
nand U4199 (N_4199,N_22,N_1116);
or U4200 (N_4200,N_902,N_2241);
or U4201 (N_4201,N_1220,N_2348);
nor U4202 (N_4202,N_1033,N_634);
nand U4203 (N_4203,N_946,N_879);
and U4204 (N_4204,N_78,N_2335);
nand U4205 (N_4205,N_2148,N_856);
and U4206 (N_4206,N_1920,N_150);
nand U4207 (N_4207,N_35,N_569);
xor U4208 (N_4208,N_1945,N_121);
nor U4209 (N_4209,N_2193,N_2196);
xor U4210 (N_4210,N_1587,N_956);
nor U4211 (N_4211,N_214,N_1676);
nand U4212 (N_4212,N_1856,N_1118);
nor U4213 (N_4213,N_2336,N_1859);
nand U4214 (N_4214,N_2326,N_1226);
nor U4215 (N_4215,N_2476,N_1480);
nand U4216 (N_4216,N_249,N_2336);
xor U4217 (N_4217,N_2287,N_10);
xor U4218 (N_4218,N_164,N_212);
and U4219 (N_4219,N_429,N_1708);
or U4220 (N_4220,N_2216,N_1768);
and U4221 (N_4221,N_2198,N_1891);
and U4222 (N_4222,N_2269,N_2211);
and U4223 (N_4223,N_790,N_489);
or U4224 (N_4224,N_1800,N_1672);
xor U4225 (N_4225,N_1069,N_1856);
and U4226 (N_4226,N_2051,N_18);
xor U4227 (N_4227,N_34,N_618);
xor U4228 (N_4228,N_548,N_1549);
and U4229 (N_4229,N_476,N_232);
xor U4230 (N_4230,N_1362,N_1864);
and U4231 (N_4231,N_1399,N_2084);
xor U4232 (N_4232,N_1515,N_1711);
and U4233 (N_4233,N_996,N_919);
or U4234 (N_4234,N_910,N_849);
and U4235 (N_4235,N_1471,N_406);
nand U4236 (N_4236,N_1420,N_898);
nand U4237 (N_4237,N_2298,N_2320);
nand U4238 (N_4238,N_998,N_364);
nand U4239 (N_4239,N_386,N_2104);
and U4240 (N_4240,N_1385,N_1611);
or U4241 (N_4241,N_1016,N_2178);
xor U4242 (N_4242,N_867,N_2397);
nor U4243 (N_4243,N_951,N_367);
nand U4244 (N_4244,N_465,N_842);
and U4245 (N_4245,N_117,N_2329);
or U4246 (N_4246,N_1820,N_2323);
or U4247 (N_4247,N_762,N_401);
or U4248 (N_4248,N_1085,N_1905);
nor U4249 (N_4249,N_996,N_1917);
xor U4250 (N_4250,N_1574,N_1953);
nand U4251 (N_4251,N_1458,N_1649);
and U4252 (N_4252,N_1610,N_619);
nand U4253 (N_4253,N_989,N_805);
or U4254 (N_4254,N_1174,N_2479);
nor U4255 (N_4255,N_34,N_1381);
nor U4256 (N_4256,N_389,N_2124);
nor U4257 (N_4257,N_982,N_1473);
or U4258 (N_4258,N_54,N_1038);
and U4259 (N_4259,N_822,N_1908);
and U4260 (N_4260,N_904,N_2150);
nand U4261 (N_4261,N_891,N_1906);
xnor U4262 (N_4262,N_1331,N_581);
nand U4263 (N_4263,N_233,N_1012);
and U4264 (N_4264,N_2390,N_1664);
nand U4265 (N_4265,N_2215,N_1575);
xnor U4266 (N_4266,N_2028,N_1817);
xnor U4267 (N_4267,N_229,N_313);
nand U4268 (N_4268,N_1450,N_1526);
nand U4269 (N_4269,N_1081,N_1024);
or U4270 (N_4270,N_676,N_1371);
and U4271 (N_4271,N_2161,N_34);
nor U4272 (N_4272,N_57,N_1127);
and U4273 (N_4273,N_1663,N_1058);
and U4274 (N_4274,N_2331,N_1514);
nor U4275 (N_4275,N_273,N_132);
and U4276 (N_4276,N_1500,N_938);
or U4277 (N_4277,N_352,N_476);
and U4278 (N_4278,N_852,N_1888);
and U4279 (N_4279,N_640,N_796);
xor U4280 (N_4280,N_256,N_170);
xnor U4281 (N_4281,N_2138,N_2479);
xnor U4282 (N_4282,N_1624,N_1929);
nor U4283 (N_4283,N_2139,N_1383);
nand U4284 (N_4284,N_329,N_1014);
nor U4285 (N_4285,N_971,N_1136);
or U4286 (N_4286,N_166,N_1533);
nor U4287 (N_4287,N_73,N_442);
or U4288 (N_4288,N_1808,N_836);
nand U4289 (N_4289,N_1813,N_423);
and U4290 (N_4290,N_597,N_2078);
xor U4291 (N_4291,N_2139,N_2339);
nand U4292 (N_4292,N_1359,N_253);
and U4293 (N_4293,N_334,N_789);
and U4294 (N_4294,N_2108,N_904);
nand U4295 (N_4295,N_1779,N_1063);
xnor U4296 (N_4296,N_529,N_1496);
or U4297 (N_4297,N_1790,N_1059);
xnor U4298 (N_4298,N_805,N_31);
or U4299 (N_4299,N_2153,N_1791);
xnor U4300 (N_4300,N_903,N_164);
and U4301 (N_4301,N_1102,N_2324);
nand U4302 (N_4302,N_55,N_338);
xnor U4303 (N_4303,N_1511,N_1482);
or U4304 (N_4304,N_306,N_2171);
or U4305 (N_4305,N_1581,N_1133);
xor U4306 (N_4306,N_1614,N_1202);
nor U4307 (N_4307,N_131,N_1258);
xnor U4308 (N_4308,N_2203,N_1163);
xor U4309 (N_4309,N_177,N_2352);
nor U4310 (N_4310,N_2147,N_1542);
nand U4311 (N_4311,N_1901,N_302);
and U4312 (N_4312,N_1470,N_1765);
or U4313 (N_4313,N_1481,N_1200);
nor U4314 (N_4314,N_2069,N_427);
xnor U4315 (N_4315,N_1493,N_848);
xor U4316 (N_4316,N_706,N_1755);
nand U4317 (N_4317,N_1680,N_1075);
nand U4318 (N_4318,N_1066,N_286);
nand U4319 (N_4319,N_7,N_2341);
and U4320 (N_4320,N_1768,N_1863);
and U4321 (N_4321,N_1476,N_735);
or U4322 (N_4322,N_1140,N_729);
nand U4323 (N_4323,N_435,N_1202);
or U4324 (N_4324,N_1819,N_2297);
xor U4325 (N_4325,N_2001,N_1956);
xor U4326 (N_4326,N_297,N_1267);
or U4327 (N_4327,N_1364,N_1975);
nand U4328 (N_4328,N_614,N_928);
nor U4329 (N_4329,N_1163,N_583);
or U4330 (N_4330,N_1610,N_272);
nand U4331 (N_4331,N_1471,N_1855);
or U4332 (N_4332,N_1043,N_866);
nand U4333 (N_4333,N_737,N_1759);
xor U4334 (N_4334,N_307,N_1710);
or U4335 (N_4335,N_2312,N_1802);
xor U4336 (N_4336,N_2496,N_1183);
or U4337 (N_4337,N_2330,N_1439);
and U4338 (N_4338,N_1960,N_731);
nor U4339 (N_4339,N_1744,N_248);
and U4340 (N_4340,N_685,N_1658);
nor U4341 (N_4341,N_1130,N_1398);
nand U4342 (N_4342,N_1257,N_2236);
nor U4343 (N_4343,N_1001,N_2324);
and U4344 (N_4344,N_1668,N_2490);
or U4345 (N_4345,N_812,N_620);
or U4346 (N_4346,N_2155,N_930);
nor U4347 (N_4347,N_2173,N_674);
nor U4348 (N_4348,N_1902,N_2146);
or U4349 (N_4349,N_1544,N_597);
xor U4350 (N_4350,N_528,N_401);
nand U4351 (N_4351,N_1254,N_905);
xor U4352 (N_4352,N_1660,N_580);
xor U4353 (N_4353,N_1979,N_127);
nand U4354 (N_4354,N_952,N_135);
nor U4355 (N_4355,N_2335,N_1619);
xnor U4356 (N_4356,N_547,N_1181);
nand U4357 (N_4357,N_258,N_1965);
nand U4358 (N_4358,N_1245,N_2040);
and U4359 (N_4359,N_1508,N_16);
or U4360 (N_4360,N_2339,N_854);
nor U4361 (N_4361,N_1017,N_2194);
and U4362 (N_4362,N_1556,N_378);
or U4363 (N_4363,N_417,N_1092);
and U4364 (N_4364,N_808,N_799);
or U4365 (N_4365,N_632,N_1337);
and U4366 (N_4366,N_1643,N_758);
xor U4367 (N_4367,N_22,N_1170);
or U4368 (N_4368,N_2095,N_1650);
nor U4369 (N_4369,N_2474,N_1279);
nand U4370 (N_4370,N_2491,N_117);
nor U4371 (N_4371,N_1156,N_1999);
or U4372 (N_4372,N_356,N_1877);
xor U4373 (N_4373,N_437,N_2482);
or U4374 (N_4374,N_66,N_42);
or U4375 (N_4375,N_934,N_2291);
xor U4376 (N_4376,N_196,N_1216);
or U4377 (N_4377,N_577,N_233);
nand U4378 (N_4378,N_1129,N_563);
or U4379 (N_4379,N_1825,N_1853);
and U4380 (N_4380,N_1560,N_2257);
nand U4381 (N_4381,N_1116,N_26);
nor U4382 (N_4382,N_348,N_152);
and U4383 (N_4383,N_2430,N_1982);
and U4384 (N_4384,N_889,N_984);
nand U4385 (N_4385,N_2179,N_2028);
xnor U4386 (N_4386,N_796,N_865);
nor U4387 (N_4387,N_856,N_273);
or U4388 (N_4388,N_1692,N_650);
nor U4389 (N_4389,N_827,N_1056);
nand U4390 (N_4390,N_845,N_1734);
nor U4391 (N_4391,N_1538,N_1167);
or U4392 (N_4392,N_948,N_105);
xor U4393 (N_4393,N_1449,N_2183);
nand U4394 (N_4394,N_1514,N_1895);
or U4395 (N_4395,N_1499,N_11);
nand U4396 (N_4396,N_917,N_1120);
and U4397 (N_4397,N_1270,N_291);
nor U4398 (N_4398,N_833,N_699);
nor U4399 (N_4399,N_1849,N_1040);
nor U4400 (N_4400,N_1064,N_1528);
or U4401 (N_4401,N_2466,N_1842);
and U4402 (N_4402,N_1394,N_1679);
or U4403 (N_4403,N_2417,N_879);
or U4404 (N_4404,N_1221,N_170);
or U4405 (N_4405,N_939,N_74);
nor U4406 (N_4406,N_234,N_1314);
or U4407 (N_4407,N_188,N_1982);
and U4408 (N_4408,N_1547,N_1249);
or U4409 (N_4409,N_441,N_1086);
nand U4410 (N_4410,N_365,N_186);
xor U4411 (N_4411,N_303,N_1772);
and U4412 (N_4412,N_743,N_1254);
nand U4413 (N_4413,N_1335,N_1297);
xor U4414 (N_4414,N_17,N_1867);
nand U4415 (N_4415,N_409,N_54);
and U4416 (N_4416,N_1017,N_1917);
nand U4417 (N_4417,N_2305,N_1024);
nand U4418 (N_4418,N_1177,N_2155);
and U4419 (N_4419,N_718,N_2176);
nor U4420 (N_4420,N_1599,N_1138);
or U4421 (N_4421,N_1290,N_234);
or U4422 (N_4422,N_1723,N_1823);
xnor U4423 (N_4423,N_1385,N_601);
or U4424 (N_4424,N_2378,N_1057);
and U4425 (N_4425,N_1486,N_1430);
and U4426 (N_4426,N_1894,N_1143);
nand U4427 (N_4427,N_634,N_1478);
and U4428 (N_4428,N_1078,N_2176);
or U4429 (N_4429,N_438,N_2145);
and U4430 (N_4430,N_1562,N_1583);
nor U4431 (N_4431,N_1116,N_2165);
xor U4432 (N_4432,N_1865,N_1171);
nor U4433 (N_4433,N_1271,N_466);
xor U4434 (N_4434,N_602,N_2365);
or U4435 (N_4435,N_692,N_854);
nand U4436 (N_4436,N_1812,N_2108);
nor U4437 (N_4437,N_1712,N_1907);
or U4438 (N_4438,N_843,N_435);
xnor U4439 (N_4439,N_1211,N_2248);
or U4440 (N_4440,N_962,N_1149);
xor U4441 (N_4441,N_132,N_1463);
nand U4442 (N_4442,N_866,N_404);
or U4443 (N_4443,N_2349,N_1684);
and U4444 (N_4444,N_456,N_814);
nor U4445 (N_4445,N_1796,N_821);
xnor U4446 (N_4446,N_1311,N_1546);
and U4447 (N_4447,N_284,N_2406);
nor U4448 (N_4448,N_1831,N_1102);
and U4449 (N_4449,N_2230,N_2492);
and U4450 (N_4450,N_721,N_2358);
xnor U4451 (N_4451,N_1466,N_2133);
nor U4452 (N_4452,N_1372,N_546);
nor U4453 (N_4453,N_2339,N_1425);
nand U4454 (N_4454,N_223,N_432);
or U4455 (N_4455,N_986,N_227);
or U4456 (N_4456,N_96,N_1168);
nand U4457 (N_4457,N_1352,N_119);
nor U4458 (N_4458,N_1132,N_665);
or U4459 (N_4459,N_1006,N_118);
or U4460 (N_4460,N_2436,N_1525);
xnor U4461 (N_4461,N_624,N_2491);
and U4462 (N_4462,N_2,N_1695);
nor U4463 (N_4463,N_525,N_972);
or U4464 (N_4464,N_2178,N_1935);
xor U4465 (N_4465,N_57,N_699);
nor U4466 (N_4466,N_1558,N_851);
nor U4467 (N_4467,N_1490,N_1711);
nand U4468 (N_4468,N_517,N_27);
nand U4469 (N_4469,N_16,N_746);
nand U4470 (N_4470,N_1359,N_1585);
nand U4471 (N_4471,N_1446,N_1357);
and U4472 (N_4472,N_497,N_2253);
xnor U4473 (N_4473,N_512,N_217);
or U4474 (N_4474,N_1593,N_600);
nor U4475 (N_4475,N_864,N_303);
nor U4476 (N_4476,N_1550,N_86);
nand U4477 (N_4477,N_674,N_1832);
or U4478 (N_4478,N_538,N_2487);
nand U4479 (N_4479,N_1266,N_525);
nor U4480 (N_4480,N_708,N_1129);
nor U4481 (N_4481,N_2065,N_2059);
or U4482 (N_4482,N_311,N_2381);
nand U4483 (N_4483,N_1485,N_672);
nand U4484 (N_4484,N_539,N_1748);
or U4485 (N_4485,N_1871,N_1396);
xnor U4486 (N_4486,N_2113,N_454);
nor U4487 (N_4487,N_874,N_195);
xnor U4488 (N_4488,N_2362,N_107);
xor U4489 (N_4489,N_439,N_1071);
or U4490 (N_4490,N_971,N_1893);
nor U4491 (N_4491,N_1670,N_1291);
or U4492 (N_4492,N_1693,N_1277);
nand U4493 (N_4493,N_601,N_1205);
nor U4494 (N_4494,N_1573,N_1992);
or U4495 (N_4495,N_1461,N_56);
nor U4496 (N_4496,N_1993,N_2369);
xnor U4497 (N_4497,N_1227,N_1448);
xnor U4498 (N_4498,N_1493,N_60);
nor U4499 (N_4499,N_2390,N_1910);
and U4500 (N_4500,N_68,N_959);
and U4501 (N_4501,N_1044,N_265);
or U4502 (N_4502,N_1176,N_675);
and U4503 (N_4503,N_559,N_1964);
xor U4504 (N_4504,N_81,N_330);
and U4505 (N_4505,N_2303,N_543);
and U4506 (N_4506,N_2189,N_125);
and U4507 (N_4507,N_1076,N_1033);
xnor U4508 (N_4508,N_1162,N_879);
nand U4509 (N_4509,N_2403,N_253);
and U4510 (N_4510,N_636,N_2325);
and U4511 (N_4511,N_1761,N_2137);
nand U4512 (N_4512,N_1524,N_1653);
xnor U4513 (N_4513,N_1840,N_1143);
nand U4514 (N_4514,N_1105,N_517);
xor U4515 (N_4515,N_2175,N_956);
xnor U4516 (N_4516,N_2023,N_1923);
or U4517 (N_4517,N_334,N_2131);
nor U4518 (N_4518,N_785,N_1773);
xor U4519 (N_4519,N_1017,N_1753);
nor U4520 (N_4520,N_657,N_1746);
or U4521 (N_4521,N_530,N_568);
nor U4522 (N_4522,N_2357,N_1779);
nor U4523 (N_4523,N_87,N_1626);
or U4524 (N_4524,N_2472,N_394);
or U4525 (N_4525,N_2071,N_1449);
nand U4526 (N_4526,N_100,N_2481);
or U4527 (N_4527,N_215,N_967);
nor U4528 (N_4528,N_2197,N_2460);
nand U4529 (N_4529,N_1770,N_504);
nor U4530 (N_4530,N_2382,N_1898);
and U4531 (N_4531,N_2005,N_56);
or U4532 (N_4532,N_1816,N_1439);
and U4533 (N_4533,N_1234,N_2087);
and U4534 (N_4534,N_305,N_762);
nand U4535 (N_4535,N_142,N_671);
or U4536 (N_4536,N_1682,N_17);
or U4537 (N_4537,N_1985,N_1248);
xnor U4538 (N_4538,N_1210,N_1061);
or U4539 (N_4539,N_1339,N_2380);
or U4540 (N_4540,N_247,N_719);
and U4541 (N_4541,N_860,N_536);
and U4542 (N_4542,N_642,N_1373);
nand U4543 (N_4543,N_1505,N_1500);
nand U4544 (N_4544,N_1627,N_1478);
nor U4545 (N_4545,N_12,N_1749);
xor U4546 (N_4546,N_1601,N_1454);
nor U4547 (N_4547,N_785,N_849);
xnor U4548 (N_4548,N_642,N_1134);
and U4549 (N_4549,N_41,N_1226);
xor U4550 (N_4550,N_1329,N_1550);
or U4551 (N_4551,N_1879,N_1601);
nor U4552 (N_4552,N_1424,N_28);
or U4553 (N_4553,N_890,N_797);
and U4554 (N_4554,N_2409,N_1009);
or U4555 (N_4555,N_575,N_273);
nor U4556 (N_4556,N_318,N_1150);
or U4557 (N_4557,N_1353,N_1812);
nor U4558 (N_4558,N_2309,N_1227);
or U4559 (N_4559,N_1543,N_782);
and U4560 (N_4560,N_2353,N_2418);
nand U4561 (N_4561,N_1584,N_2449);
nor U4562 (N_4562,N_406,N_1041);
xnor U4563 (N_4563,N_1742,N_1186);
or U4564 (N_4564,N_873,N_1545);
xor U4565 (N_4565,N_407,N_1141);
xor U4566 (N_4566,N_1057,N_2249);
xnor U4567 (N_4567,N_751,N_1310);
and U4568 (N_4568,N_2404,N_1762);
nor U4569 (N_4569,N_587,N_526);
nand U4570 (N_4570,N_542,N_523);
or U4571 (N_4571,N_1332,N_1881);
xor U4572 (N_4572,N_28,N_1375);
nand U4573 (N_4573,N_1715,N_1033);
or U4574 (N_4574,N_1725,N_1477);
nor U4575 (N_4575,N_1782,N_1019);
xor U4576 (N_4576,N_1711,N_290);
nand U4577 (N_4577,N_237,N_592);
nor U4578 (N_4578,N_2189,N_2358);
xnor U4579 (N_4579,N_1455,N_331);
or U4580 (N_4580,N_365,N_1933);
xor U4581 (N_4581,N_1764,N_2075);
and U4582 (N_4582,N_1062,N_570);
xor U4583 (N_4583,N_2474,N_325);
and U4584 (N_4584,N_1083,N_2446);
or U4585 (N_4585,N_643,N_2218);
or U4586 (N_4586,N_148,N_114);
nor U4587 (N_4587,N_1271,N_1274);
nand U4588 (N_4588,N_210,N_1633);
nor U4589 (N_4589,N_1614,N_429);
nor U4590 (N_4590,N_1911,N_1367);
and U4591 (N_4591,N_2283,N_662);
nor U4592 (N_4592,N_191,N_491);
xor U4593 (N_4593,N_2389,N_1946);
and U4594 (N_4594,N_312,N_489);
and U4595 (N_4595,N_1286,N_1574);
or U4596 (N_4596,N_1844,N_1015);
nand U4597 (N_4597,N_2051,N_843);
nand U4598 (N_4598,N_1186,N_1541);
xnor U4599 (N_4599,N_522,N_983);
xnor U4600 (N_4600,N_1810,N_261);
nand U4601 (N_4601,N_1239,N_1063);
nand U4602 (N_4602,N_2131,N_1877);
nand U4603 (N_4603,N_940,N_1568);
or U4604 (N_4604,N_427,N_1130);
xor U4605 (N_4605,N_154,N_1934);
nand U4606 (N_4606,N_2406,N_1119);
xor U4607 (N_4607,N_1078,N_1055);
and U4608 (N_4608,N_1262,N_598);
nand U4609 (N_4609,N_1586,N_1167);
nor U4610 (N_4610,N_398,N_379);
or U4611 (N_4611,N_1668,N_2096);
xor U4612 (N_4612,N_1426,N_1964);
nand U4613 (N_4613,N_1974,N_190);
or U4614 (N_4614,N_302,N_2071);
nor U4615 (N_4615,N_1387,N_1321);
or U4616 (N_4616,N_258,N_977);
nor U4617 (N_4617,N_1421,N_452);
nor U4618 (N_4618,N_1233,N_889);
nor U4619 (N_4619,N_1017,N_465);
xor U4620 (N_4620,N_772,N_1842);
nand U4621 (N_4621,N_1641,N_1527);
xor U4622 (N_4622,N_1327,N_532);
nand U4623 (N_4623,N_1414,N_1350);
or U4624 (N_4624,N_35,N_2314);
nand U4625 (N_4625,N_2235,N_1240);
and U4626 (N_4626,N_541,N_1804);
or U4627 (N_4627,N_855,N_1296);
nor U4628 (N_4628,N_1744,N_2179);
nand U4629 (N_4629,N_7,N_689);
xnor U4630 (N_4630,N_1395,N_1095);
or U4631 (N_4631,N_2161,N_525);
nand U4632 (N_4632,N_2461,N_553);
xnor U4633 (N_4633,N_1583,N_2022);
nand U4634 (N_4634,N_1286,N_1021);
nor U4635 (N_4635,N_472,N_2386);
or U4636 (N_4636,N_1299,N_200);
nand U4637 (N_4637,N_531,N_1334);
xnor U4638 (N_4638,N_667,N_1236);
or U4639 (N_4639,N_1668,N_1298);
or U4640 (N_4640,N_685,N_2002);
or U4641 (N_4641,N_2364,N_2463);
nor U4642 (N_4642,N_1079,N_1731);
and U4643 (N_4643,N_1581,N_1381);
xor U4644 (N_4644,N_1705,N_1293);
and U4645 (N_4645,N_1563,N_2485);
nand U4646 (N_4646,N_827,N_2371);
and U4647 (N_4647,N_2216,N_2393);
or U4648 (N_4648,N_1622,N_1973);
and U4649 (N_4649,N_1751,N_2345);
nand U4650 (N_4650,N_2149,N_2433);
xnor U4651 (N_4651,N_1673,N_20);
and U4652 (N_4652,N_461,N_2076);
nor U4653 (N_4653,N_250,N_1839);
and U4654 (N_4654,N_2093,N_1373);
nor U4655 (N_4655,N_2412,N_424);
or U4656 (N_4656,N_1902,N_1231);
and U4657 (N_4657,N_1828,N_182);
and U4658 (N_4658,N_1818,N_2019);
nand U4659 (N_4659,N_1481,N_1578);
and U4660 (N_4660,N_689,N_2262);
xnor U4661 (N_4661,N_1075,N_371);
xor U4662 (N_4662,N_38,N_1061);
nor U4663 (N_4663,N_312,N_546);
and U4664 (N_4664,N_1054,N_1624);
or U4665 (N_4665,N_2046,N_1819);
or U4666 (N_4666,N_906,N_1943);
or U4667 (N_4667,N_1960,N_458);
or U4668 (N_4668,N_1822,N_908);
and U4669 (N_4669,N_1623,N_1364);
nand U4670 (N_4670,N_55,N_139);
nand U4671 (N_4671,N_2112,N_896);
nand U4672 (N_4672,N_1417,N_2043);
or U4673 (N_4673,N_1661,N_1971);
nor U4674 (N_4674,N_1643,N_1783);
nand U4675 (N_4675,N_1032,N_2462);
nor U4676 (N_4676,N_1926,N_1408);
or U4677 (N_4677,N_2128,N_2299);
or U4678 (N_4678,N_748,N_2298);
or U4679 (N_4679,N_11,N_1926);
and U4680 (N_4680,N_2401,N_1252);
or U4681 (N_4681,N_2018,N_1641);
nand U4682 (N_4682,N_632,N_2038);
nand U4683 (N_4683,N_637,N_275);
or U4684 (N_4684,N_986,N_1971);
xor U4685 (N_4685,N_1278,N_922);
nor U4686 (N_4686,N_1860,N_980);
or U4687 (N_4687,N_376,N_692);
nand U4688 (N_4688,N_75,N_1196);
nand U4689 (N_4689,N_1258,N_1290);
xor U4690 (N_4690,N_936,N_774);
and U4691 (N_4691,N_30,N_767);
nor U4692 (N_4692,N_1572,N_2055);
and U4693 (N_4693,N_1894,N_2489);
nand U4694 (N_4694,N_81,N_1264);
nand U4695 (N_4695,N_1881,N_217);
nand U4696 (N_4696,N_222,N_551);
nand U4697 (N_4697,N_370,N_523);
nand U4698 (N_4698,N_1894,N_2347);
or U4699 (N_4699,N_763,N_993);
xor U4700 (N_4700,N_2213,N_1869);
and U4701 (N_4701,N_1864,N_57);
and U4702 (N_4702,N_682,N_2447);
and U4703 (N_4703,N_1317,N_2041);
or U4704 (N_4704,N_8,N_724);
nand U4705 (N_4705,N_1720,N_1566);
nor U4706 (N_4706,N_1176,N_370);
and U4707 (N_4707,N_2205,N_384);
nand U4708 (N_4708,N_1201,N_281);
and U4709 (N_4709,N_2095,N_1186);
and U4710 (N_4710,N_609,N_1552);
nor U4711 (N_4711,N_1559,N_1342);
and U4712 (N_4712,N_389,N_1418);
nor U4713 (N_4713,N_722,N_1993);
and U4714 (N_4714,N_500,N_429);
or U4715 (N_4715,N_1522,N_2081);
or U4716 (N_4716,N_1357,N_465);
nand U4717 (N_4717,N_774,N_1156);
nor U4718 (N_4718,N_1257,N_1115);
nand U4719 (N_4719,N_2197,N_227);
or U4720 (N_4720,N_827,N_1034);
or U4721 (N_4721,N_1158,N_2448);
and U4722 (N_4722,N_573,N_265);
or U4723 (N_4723,N_742,N_358);
and U4724 (N_4724,N_355,N_370);
or U4725 (N_4725,N_880,N_2188);
or U4726 (N_4726,N_677,N_1749);
or U4727 (N_4727,N_1755,N_961);
xnor U4728 (N_4728,N_1283,N_695);
xor U4729 (N_4729,N_1533,N_2226);
and U4730 (N_4730,N_1116,N_679);
and U4731 (N_4731,N_1107,N_1063);
or U4732 (N_4732,N_460,N_1868);
nand U4733 (N_4733,N_465,N_9);
or U4734 (N_4734,N_2015,N_1932);
or U4735 (N_4735,N_1120,N_2007);
or U4736 (N_4736,N_589,N_1383);
nand U4737 (N_4737,N_679,N_1968);
and U4738 (N_4738,N_1666,N_54);
xor U4739 (N_4739,N_912,N_1998);
xor U4740 (N_4740,N_1710,N_1588);
nand U4741 (N_4741,N_727,N_601);
nor U4742 (N_4742,N_1038,N_2268);
xnor U4743 (N_4743,N_287,N_390);
nor U4744 (N_4744,N_498,N_1356);
and U4745 (N_4745,N_2472,N_1733);
nand U4746 (N_4746,N_951,N_387);
and U4747 (N_4747,N_697,N_1931);
nor U4748 (N_4748,N_779,N_1085);
nand U4749 (N_4749,N_714,N_499);
and U4750 (N_4750,N_1142,N_2297);
nand U4751 (N_4751,N_1065,N_51);
and U4752 (N_4752,N_1488,N_781);
or U4753 (N_4753,N_1897,N_226);
and U4754 (N_4754,N_1469,N_1949);
nor U4755 (N_4755,N_620,N_1528);
and U4756 (N_4756,N_2128,N_2448);
xor U4757 (N_4757,N_810,N_98);
nand U4758 (N_4758,N_716,N_2138);
nand U4759 (N_4759,N_1468,N_1637);
xnor U4760 (N_4760,N_422,N_1664);
nand U4761 (N_4761,N_202,N_1671);
nand U4762 (N_4762,N_927,N_44);
or U4763 (N_4763,N_254,N_1676);
and U4764 (N_4764,N_1172,N_1403);
and U4765 (N_4765,N_2458,N_1689);
nor U4766 (N_4766,N_767,N_191);
nor U4767 (N_4767,N_465,N_2372);
or U4768 (N_4768,N_1053,N_2198);
nor U4769 (N_4769,N_965,N_1387);
and U4770 (N_4770,N_961,N_1641);
or U4771 (N_4771,N_2392,N_78);
nand U4772 (N_4772,N_417,N_861);
nand U4773 (N_4773,N_726,N_1165);
nand U4774 (N_4774,N_529,N_1231);
xor U4775 (N_4775,N_2341,N_1442);
xor U4776 (N_4776,N_2244,N_830);
nand U4777 (N_4777,N_2254,N_689);
or U4778 (N_4778,N_165,N_518);
nand U4779 (N_4779,N_910,N_351);
xnor U4780 (N_4780,N_2364,N_1967);
and U4781 (N_4781,N_542,N_639);
nand U4782 (N_4782,N_539,N_1135);
and U4783 (N_4783,N_1164,N_139);
nand U4784 (N_4784,N_877,N_1817);
and U4785 (N_4785,N_941,N_809);
and U4786 (N_4786,N_582,N_1936);
and U4787 (N_4787,N_2204,N_1614);
or U4788 (N_4788,N_2435,N_2081);
nor U4789 (N_4789,N_205,N_752);
and U4790 (N_4790,N_704,N_71);
or U4791 (N_4791,N_1007,N_694);
nand U4792 (N_4792,N_1660,N_212);
xnor U4793 (N_4793,N_792,N_40);
or U4794 (N_4794,N_1185,N_100);
nor U4795 (N_4795,N_1096,N_1353);
and U4796 (N_4796,N_692,N_528);
xor U4797 (N_4797,N_838,N_1422);
nand U4798 (N_4798,N_16,N_2432);
and U4799 (N_4799,N_686,N_750);
xor U4800 (N_4800,N_2454,N_1183);
and U4801 (N_4801,N_210,N_1493);
nand U4802 (N_4802,N_1851,N_2303);
or U4803 (N_4803,N_1671,N_1136);
nor U4804 (N_4804,N_1022,N_631);
or U4805 (N_4805,N_309,N_1670);
nand U4806 (N_4806,N_1512,N_767);
and U4807 (N_4807,N_1617,N_1608);
xnor U4808 (N_4808,N_551,N_2276);
and U4809 (N_4809,N_328,N_2173);
and U4810 (N_4810,N_785,N_1017);
and U4811 (N_4811,N_1274,N_825);
nor U4812 (N_4812,N_1031,N_467);
xnor U4813 (N_4813,N_1497,N_501);
nor U4814 (N_4814,N_1356,N_905);
or U4815 (N_4815,N_1341,N_1496);
nor U4816 (N_4816,N_493,N_1857);
xor U4817 (N_4817,N_258,N_17);
xor U4818 (N_4818,N_851,N_1990);
or U4819 (N_4819,N_1862,N_2442);
or U4820 (N_4820,N_2437,N_509);
nor U4821 (N_4821,N_1726,N_2363);
or U4822 (N_4822,N_1073,N_2453);
xnor U4823 (N_4823,N_44,N_305);
or U4824 (N_4824,N_157,N_1187);
nor U4825 (N_4825,N_703,N_1361);
nor U4826 (N_4826,N_2279,N_1615);
or U4827 (N_4827,N_1559,N_2438);
or U4828 (N_4828,N_1246,N_1027);
and U4829 (N_4829,N_1859,N_421);
and U4830 (N_4830,N_258,N_746);
nand U4831 (N_4831,N_1412,N_2269);
or U4832 (N_4832,N_1341,N_553);
and U4833 (N_4833,N_1730,N_1824);
nor U4834 (N_4834,N_1686,N_437);
xnor U4835 (N_4835,N_1042,N_362);
or U4836 (N_4836,N_1590,N_2331);
xor U4837 (N_4837,N_1964,N_77);
xor U4838 (N_4838,N_1292,N_1454);
xnor U4839 (N_4839,N_1546,N_957);
xnor U4840 (N_4840,N_1121,N_1704);
or U4841 (N_4841,N_964,N_1047);
nand U4842 (N_4842,N_910,N_2174);
or U4843 (N_4843,N_387,N_1092);
nor U4844 (N_4844,N_2394,N_1153);
and U4845 (N_4845,N_107,N_2307);
xor U4846 (N_4846,N_816,N_285);
and U4847 (N_4847,N_62,N_2041);
nand U4848 (N_4848,N_1508,N_201);
nor U4849 (N_4849,N_1311,N_400);
and U4850 (N_4850,N_778,N_1093);
nor U4851 (N_4851,N_2112,N_1028);
and U4852 (N_4852,N_1848,N_1502);
nor U4853 (N_4853,N_2453,N_2145);
or U4854 (N_4854,N_1194,N_598);
nor U4855 (N_4855,N_596,N_1679);
nand U4856 (N_4856,N_820,N_284);
or U4857 (N_4857,N_2374,N_1286);
xnor U4858 (N_4858,N_1620,N_510);
nand U4859 (N_4859,N_1449,N_825);
xnor U4860 (N_4860,N_1750,N_2271);
or U4861 (N_4861,N_2242,N_742);
nor U4862 (N_4862,N_1718,N_194);
nor U4863 (N_4863,N_1898,N_778);
nand U4864 (N_4864,N_741,N_2047);
nand U4865 (N_4865,N_1181,N_1100);
and U4866 (N_4866,N_1616,N_1910);
nand U4867 (N_4867,N_2156,N_798);
nand U4868 (N_4868,N_757,N_570);
nor U4869 (N_4869,N_157,N_316);
or U4870 (N_4870,N_1440,N_888);
nand U4871 (N_4871,N_1621,N_385);
and U4872 (N_4872,N_1802,N_723);
nand U4873 (N_4873,N_38,N_715);
and U4874 (N_4874,N_377,N_1096);
or U4875 (N_4875,N_251,N_883);
nor U4876 (N_4876,N_1396,N_728);
and U4877 (N_4877,N_492,N_1126);
or U4878 (N_4878,N_1125,N_2462);
and U4879 (N_4879,N_241,N_1784);
or U4880 (N_4880,N_350,N_256);
nand U4881 (N_4881,N_75,N_2193);
nor U4882 (N_4882,N_2322,N_308);
or U4883 (N_4883,N_1794,N_1493);
nor U4884 (N_4884,N_1605,N_2324);
xnor U4885 (N_4885,N_1602,N_1865);
xor U4886 (N_4886,N_2214,N_2026);
nand U4887 (N_4887,N_268,N_2276);
xor U4888 (N_4888,N_1833,N_2008);
xnor U4889 (N_4889,N_1973,N_1053);
nand U4890 (N_4890,N_1755,N_364);
nand U4891 (N_4891,N_2466,N_1625);
or U4892 (N_4892,N_1135,N_1574);
xor U4893 (N_4893,N_936,N_192);
nand U4894 (N_4894,N_233,N_2204);
nor U4895 (N_4895,N_874,N_450);
xor U4896 (N_4896,N_306,N_1188);
or U4897 (N_4897,N_55,N_2294);
nand U4898 (N_4898,N_1426,N_654);
nor U4899 (N_4899,N_1666,N_2097);
nand U4900 (N_4900,N_2413,N_495);
nand U4901 (N_4901,N_2370,N_1575);
or U4902 (N_4902,N_949,N_368);
or U4903 (N_4903,N_1494,N_611);
xnor U4904 (N_4904,N_1566,N_199);
or U4905 (N_4905,N_1229,N_1858);
or U4906 (N_4906,N_1088,N_2396);
or U4907 (N_4907,N_575,N_2181);
nand U4908 (N_4908,N_1936,N_1674);
xor U4909 (N_4909,N_1853,N_2058);
xor U4910 (N_4910,N_929,N_1234);
or U4911 (N_4911,N_1734,N_6);
nand U4912 (N_4912,N_2445,N_1233);
and U4913 (N_4913,N_1823,N_1301);
xor U4914 (N_4914,N_716,N_404);
and U4915 (N_4915,N_1333,N_1441);
xnor U4916 (N_4916,N_2288,N_1618);
nor U4917 (N_4917,N_2388,N_741);
and U4918 (N_4918,N_406,N_2263);
nor U4919 (N_4919,N_2116,N_2372);
nor U4920 (N_4920,N_359,N_2223);
and U4921 (N_4921,N_1785,N_1131);
and U4922 (N_4922,N_1239,N_2061);
xor U4923 (N_4923,N_647,N_2280);
nor U4924 (N_4924,N_1263,N_2482);
or U4925 (N_4925,N_961,N_1445);
nand U4926 (N_4926,N_947,N_2217);
and U4927 (N_4927,N_1546,N_224);
and U4928 (N_4928,N_2413,N_1893);
and U4929 (N_4929,N_39,N_883);
and U4930 (N_4930,N_1350,N_2443);
nand U4931 (N_4931,N_2384,N_1060);
nand U4932 (N_4932,N_414,N_714);
nand U4933 (N_4933,N_1223,N_125);
xnor U4934 (N_4934,N_441,N_1801);
and U4935 (N_4935,N_1926,N_965);
nand U4936 (N_4936,N_740,N_688);
xnor U4937 (N_4937,N_2020,N_1617);
nand U4938 (N_4938,N_2048,N_19);
nor U4939 (N_4939,N_1579,N_1290);
nand U4940 (N_4940,N_1367,N_626);
nor U4941 (N_4941,N_2173,N_716);
nor U4942 (N_4942,N_359,N_1161);
nor U4943 (N_4943,N_1533,N_1514);
nand U4944 (N_4944,N_2084,N_2364);
xor U4945 (N_4945,N_286,N_267);
nor U4946 (N_4946,N_2377,N_2415);
and U4947 (N_4947,N_2341,N_1970);
and U4948 (N_4948,N_637,N_1135);
and U4949 (N_4949,N_1134,N_1935);
nand U4950 (N_4950,N_2154,N_1214);
xnor U4951 (N_4951,N_29,N_1897);
and U4952 (N_4952,N_1268,N_768);
nor U4953 (N_4953,N_384,N_1063);
nor U4954 (N_4954,N_835,N_1841);
nand U4955 (N_4955,N_123,N_1768);
and U4956 (N_4956,N_967,N_1701);
nand U4957 (N_4957,N_508,N_361);
and U4958 (N_4958,N_2194,N_1013);
xor U4959 (N_4959,N_1998,N_732);
or U4960 (N_4960,N_590,N_694);
nor U4961 (N_4961,N_2351,N_111);
or U4962 (N_4962,N_1061,N_1757);
and U4963 (N_4963,N_1362,N_505);
xor U4964 (N_4964,N_803,N_237);
and U4965 (N_4965,N_1120,N_2456);
xnor U4966 (N_4966,N_1951,N_1979);
xnor U4967 (N_4967,N_378,N_2042);
xor U4968 (N_4968,N_1036,N_885);
xor U4969 (N_4969,N_445,N_1615);
and U4970 (N_4970,N_957,N_1291);
or U4971 (N_4971,N_389,N_618);
or U4972 (N_4972,N_541,N_571);
xnor U4973 (N_4973,N_1226,N_2089);
xor U4974 (N_4974,N_1597,N_928);
and U4975 (N_4975,N_1561,N_1603);
and U4976 (N_4976,N_633,N_300);
or U4977 (N_4977,N_2246,N_2111);
xnor U4978 (N_4978,N_582,N_714);
nor U4979 (N_4979,N_1622,N_1970);
nor U4980 (N_4980,N_431,N_2363);
nand U4981 (N_4981,N_8,N_2372);
nand U4982 (N_4982,N_602,N_1687);
nor U4983 (N_4983,N_1074,N_1330);
or U4984 (N_4984,N_1857,N_121);
nor U4985 (N_4985,N_347,N_2083);
xor U4986 (N_4986,N_1480,N_1212);
or U4987 (N_4987,N_1502,N_1556);
nor U4988 (N_4988,N_507,N_1734);
and U4989 (N_4989,N_30,N_1605);
or U4990 (N_4990,N_301,N_180);
and U4991 (N_4991,N_2129,N_470);
nor U4992 (N_4992,N_2304,N_909);
or U4993 (N_4993,N_2185,N_799);
nand U4994 (N_4994,N_791,N_1079);
and U4995 (N_4995,N_1851,N_1495);
and U4996 (N_4996,N_858,N_1651);
nand U4997 (N_4997,N_833,N_832);
or U4998 (N_4998,N_293,N_1824);
xnor U4999 (N_4999,N_565,N_341);
nand U5000 (N_5000,N_3840,N_2740);
and U5001 (N_5001,N_4799,N_3868);
nor U5002 (N_5002,N_2937,N_4712);
and U5003 (N_5003,N_4377,N_4468);
and U5004 (N_5004,N_4032,N_2862);
nor U5005 (N_5005,N_3589,N_4551);
nand U5006 (N_5006,N_4317,N_2883);
nor U5007 (N_5007,N_3978,N_4252);
nor U5008 (N_5008,N_2500,N_3258);
xnor U5009 (N_5009,N_3878,N_2729);
and U5010 (N_5010,N_4295,N_3770);
nor U5011 (N_5011,N_3246,N_3271);
nor U5012 (N_5012,N_4862,N_4091);
xnor U5013 (N_5013,N_2953,N_3910);
nand U5014 (N_5014,N_2938,N_4274);
nor U5015 (N_5015,N_3094,N_2537);
xor U5016 (N_5016,N_4577,N_3233);
or U5017 (N_5017,N_3270,N_4963);
nor U5018 (N_5018,N_4266,N_3937);
or U5019 (N_5019,N_3632,N_3342);
nand U5020 (N_5020,N_2545,N_4339);
xor U5021 (N_5021,N_4123,N_3154);
xnor U5022 (N_5022,N_3443,N_4459);
nor U5023 (N_5023,N_2534,N_3564);
nor U5024 (N_5024,N_4867,N_3595);
and U5025 (N_5025,N_3244,N_3002);
nor U5026 (N_5026,N_4897,N_2579);
or U5027 (N_5027,N_4375,N_3252);
and U5028 (N_5028,N_4848,N_2673);
and U5029 (N_5029,N_3839,N_3427);
nor U5030 (N_5030,N_3179,N_4492);
or U5031 (N_5031,N_3268,N_2564);
nor U5032 (N_5032,N_3349,N_2886);
nor U5033 (N_5033,N_4303,N_4803);
xor U5034 (N_5034,N_3764,N_3054);
and U5035 (N_5035,N_3475,N_3621);
and U5036 (N_5036,N_2657,N_3191);
xor U5037 (N_5037,N_3896,N_3486);
and U5038 (N_5038,N_3834,N_2565);
nor U5039 (N_5039,N_3719,N_2758);
and U5040 (N_5040,N_4210,N_4697);
and U5041 (N_5041,N_2645,N_2833);
or U5042 (N_5042,N_3231,N_4659);
nor U5043 (N_5043,N_3590,N_4720);
xnor U5044 (N_5044,N_4034,N_3630);
nand U5045 (N_5045,N_2697,N_4398);
nand U5046 (N_5046,N_3056,N_4545);
or U5047 (N_5047,N_4967,N_2675);
or U5048 (N_5048,N_4631,N_3112);
or U5049 (N_5049,N_3106,N_2686);
nor U5050 (N_5050,N_2829,N_4902);
or U5051 (N_5051,N_2837,N_2629);
nor U5052 (N_5052,N_4953,N_3298);
nand U5053 (N_5053,N_2956,N_4774);
or U5054 (N_5054,N_3105,N_4448);
or U5055 (N_5055,N_2583,N_4784);
xnor U5056 (N_5056,N_3129,N_3286);
and U5057 (N_5057,N_3123,N_2572);
xor U5058 (N_5058,N_4479,N_2547);
nand U5059 (N_5059,N_2672,N_2617);
nor U5060 (N_5060,N_3795,N_4980);
nor U5061 (N_5061,N_4601,N_3777);
or U5062 (N_5062,N_3666,N_3961);
xnor U5063 (N_5063,N_4998,N_3249);
nand U5064 (N_5064,N_4877,N_4363);
nand U5065 (N_5065,N_3197,N_4357);
or U5066 (N_5066,N_4160,N_3012);
nand U5067 (N_5067,N_4191,N_3288);
and U5068 (N_5068,N_3053,N_4837);
nor U5069 (N_5069,N_3874,N_4595);
or U5070 (N_5070,N_2989,N_3391);
xor U5071 (N_5071,N_2985,N_3411);
and U5072 (N_5072,N_3732,N_4331);
and U5073 (N_5073,N_3453,N_3651);
or U5074 (N_5074,N_3459,N_4383);
or U5075 (N_5075,N_3623,N_4237);
nand U5076 (N_5076,N_3706,N_2850);
nor U5077 (N_5077,N_4189,N_3846);
and U5078 (N_5078,N_2561,N_2846);
or U5079 (N_5079,N_3726,N_2549);
xor U5080 (N_5080,N_3801,N_2794);
nand U5081 (N_5081,N_4567,N_4236);
nor U5082 (N_5082,N_4334,N_2524);
and U5083 (N_5083,N_4040,N_3034);
xor U5084 (N_5084,N_3552,N_4914);
nand U5085 (N_5085,N_4858,N_3346);
nor U5086 (N_5086,N_4006,N_2805);
and U5087 (N_5087,N_3194,N_4855);
nor U5088 (N_5088,N_4834,N_4322);
nand U5089 (N_5089,N_4192,N_4195);
or U5090 (N_5090,N_4606,N_4395);
and U5091 (N_5091,N_2822,N_3320);
xor U5092 (N_5092,N_4095,N_4482);
xnor U5093 (N_5093,N_3082,N_4800);
and U5094 (N_5094,N_4526,N_3926);
xnor U5095 (N_5095,N_4932,N_4602);
and U5096 (N_5096,N_2655,N_3300);
nor U5097 (N_5097,N_4872,N_3296);
and U5098 (N_5098,N_2900,N_3240);
nor U5099 (N_5099,N_4136,N_4106);
xnor U5100 (N_5100,N_2571,N_4318);
and U5101 (N_5101,N_4950,N_3955);
or U5102 (N_5102,N_4374,N_3963);
nor U5103 (N_5103,N_3287,N_2706);
nand U5104 (N_5104,N_4805,N_3501);
nor U5105 (N_5105,N_2825,N_2540);
nand U5106 (N_5106,N_3267,N_3304);
nand U5107 (N_5107,N_3783,N_4974);
and U5108 (N_5108,N_3709,N_2926);
and U5109 (N_5109,N_4386,N_4080);
or U5110 (N_5110,N_4639,N_4047);
and U5111 (N_5111,N_3638,N_4497);
nand U5112 (N_5112,N_4504,N_4137);
xnor U5113 (N_5113,N_3462,N_2548);
nand U5114 (N_5114,N_3370,N_2855);
and U5115 (N_5115,N_2993,N_4089);
nand U5116 (N_5116,N_3163,N_2935);
or U5117 (N_5117,N_3114,N_2509);
or U5118 (N_5118,N_4409,N_4821);
and U5119 (N_5119,N_2960,N_4391);
nand U5120 (N_5120,N_3156,N_3852);
xor U5121 (N_5121,N_3535,N_3489);
nor U5122 (N_5122,N_4970,N_4445);
and U5123 (N_5123,N_3352,N_3151);
and U5124 (N_5124,N_3561,N_4696);
or U5125 (N_5125,N_4128,N_3090);
or U5126 (N_5126,N_3161,N_3598);
or U5127 (N_5127,N_2711,N_2893);
and U5128 (N_5128,N_3769,N_3134);
or U5129 (N_5129,N_4640,N_4478);
nand U5130 (N_5130,N_4686,N_3518);
nor U5131 (N_5131,N_4926,N_3182);
nand U5132 (N_5132,N_3964,N_3160);
nand U5133 (N_5133,N_3418,N_3136);
or U5134 (N_5134,N_3866,N_4271);
nor U5135 (N_5135,N_2601,N_3409);
xnor U5136 (N_5136,N_2618,N_4532);
xnor U5137 (N_5137,N_4026,N_4023);
or U5138 (N_5138,N_4874,N_4093);
xnor U5139 (N_5139,N_4178,N_4001);
nor U5140 (N_5140,N_2745,N_3139);
xnor U5141 (N_5141,N_3897,N_4279);
nand U5142 (N_5142,N_4224,N_2649);
or U5143 (N_5143,N_3525,N_4273);
or U5144 (N_5144,N_3325,N_4947);
or U5145 (N_5145,N_3004,N_4965);
or U5146 (N_5146,N_3399,N_3347);
xor U5147 (N_5147,N_4972,N_3005);
xnor U5148 (N_5148,N_2585,N_2691);
and U5149 (N_5149,N_4798,N_4120);
or U5150 (N_5150,N_3626,N_3850);
and U5151 (N_5151,N_4773,N_2936);
nor U5152 (N_5152,N_4957,N_4441);
nand U5153 (N_5153,N_3966,N_3417);
or U5154 (N_5154,N_4043,N_4718);
and U5155 (N_5155,N_4153,N_4045);
or U5156 (N_5156,N_2785,N_4215);
xnor U5157 (N_5157,N_3178,N_4309);
or U5158 (N_5158,N_3150,N_2523);
nor U5159 (N_5159,N_3691,N_3784);
nand U5160 (N_5160,N_3655,N_4263);
nand U5161 (N_5161,N_3956,N_4999);
xnor U5162 (N_5162,N_2831,N_3541);
xor U5163 (N_5163,N_3951,N_2780);
xnor U5164 (N_5164,N_3071,N_2727);
and U5165 (N_5165,N_3928,N_4529);
xnor U5166 (N_5166,N_4098,N_3921);
nand U5167 (N_5167,N_2597,N_4115);
and U5168 (N_5168,N_4973,N_4846);
nand U5169 (N_5169,N_4025,N_4766);
and U5170 (N_5170,N_3624,N_4525);
xnor U5171 (N_5171,N_2662,N_4477);
or U5172 (N_5172,N_2841,N_3587);
xnor U5173 (N_5173,N_4246,N_3339);
nor U5174 (N_5174,N_4096,N_3898);
nand U5175 (N_5175,N_4355,N_4683);
nand U5176 (N_5176,N_3037,N_4891);
nor U5177 (N_5177,N_2994,N_2615);
xor U5178 (N_5178,N_3100,N_2820);
nand U5179 (N_5179,N_2586,N_2828);
xnor U5180 (N_5180,N_4907,N_3254);
or U5181 (N_5181,N_2668,N_4730);
xor U5182 (N_5182,N_3842,N_2764);
and U5183 (N_5183,N_4767,N_3140);
xnor U5184 (N_5184,N_4397,N_2622);
and U5185 (N_5185,N_3656,N_3488);
or U5186 (N_5186,N_3751,N_3575);
and U5187 (N_5187,N_4996,N_3000);
xnor U5188 (N_5188,N_4533,N_3173);
xnor U5189 (N_5189,N_3434,N_4049);
or U5190 (N_5190,N_4473,N_3207);
nor U5191 (N_5191,N_2684,N_4134);
xnor U5192 (N_5192,N_3241,N_4489);
and U5193 (N_5193,N_4241,N_3953);
nor U5194 (N_5194,N_3622,N_2603);
xor U5195 (N_5195,N_4732,N_4495);
or U5196 (N_5196,N_4248,N_3545);
nand U5197 (N_5197,N_4351,N_3516);
or U5198 (N_5198,N_3102,N_4251);
nand U5199 (N_5199,N_3028,N_3245);
nand U5200 (N_5200,N_4937,N_2760);
nand U5201 (N_5201,N_3804,N_3600);
xnor U5202 (N_5202,N_3819,N_2942);
and U5203 (N_5203,N_3925,N_3932);
nand U5204 (N_5204,N_3558,N_4180);
xor U5205 (N_5205,N_3393,N_3234);
or U5206 (N_5206,N_3455,N_2701);
and U5207 (N_5207,N_3208,N_2640);
and U5208 (N_5208,N_4312,N_2527);
and U5209 (N_5209,N_4324,N_4822);
nand U5210 (N_5210,N_3413,N_2536);
nand U5211 (N_5211,N_3894,N_2884);
or U5212 (N_5212,N_4721,N_4889);
nand U5213 (N_5213,N_4503,N_4335);
xor U5214 (N_5214,N_3774,N_4181);
or U5215 (N_5215,N_4536,N_4223);
or U5216 (N_5216,N_4483,N_4208);
nand U5217 (N_5217,N_3506,N_3566);
xnor U5218 (N_5218,N_4265,N_3731);
nand U5219 (N_5219,N_2719,N_3767);
nand U5220 (N_5220,N_3923,N_3532);
xnor U5221 (N_5221,N_4596,N_4158);
nor U5222 (N_5222,N_3204,N_4658);
nor U5223 (N_5223,N_3505,N_3067);
or U5224 (N_5224,N_2860,N_4861);
nand U5225 (N_5225,N_4761,N_3788);
xnor U5226 (N_5226,N_2856,N_3072);
nand U5227 (N_5227,N_2660,N_3350);
or U5228 (N_5228,N_3849,N_4460);
and U5229 (N_5229,N_2703,N_4133);
nand U5230 (N_5230,N_3911,N_3493);
nand U5231 (N_5231,N_2984,N_4842);
nand U5232 (N_5232,N_2971,N_3760);
nor U5233 (N_5233,N_3196,N_2735);
xor U5234 (N_5234,N_4665,N_4036);
and U5235 (N_5235,N_4358,N_4175);
or U5236 (N_5236,N_2864,N_2897);
nor U5237 (N_5237,N_4188,N_3318);
xnor U5238 (N_5238,N_4446,N_4264);
or U5239 (N_5239,N_3713,N_3971);
xor U5240 (N_5240,N_4387,N_3825);
and U5241 (N_5241,N_2791,N_4003);
and U5242 (N_5242,N_3216,N_2742);
nor U5243 (N_5243,N_4808,N_3909);
nand U5244 (N_5244,N_3467,N_3107);
or U5245 (N_5245,N_3721,N_3968);
nor U5246 (N_5246,N_4756,N_3975);
nand U5247 (N_5247,N_2923,N_3480);
and U5248 (N_5248,N_2774,N_3883);
nor U5249 (N_5249,N_4486,N_2683);
xor U5250 (N_5250,N_4332,N_4813);
nand U5251 (N_5251,N_2685,N_2606);
xor U5252 (N_5252,N_4276,N_3021);
nor U5253 (N_5253,N_4587,N_4002);
or U5254 (N_5254,N_4961,N_4894);
or U5255 (N_5255,N_3727,N_4809);
and U5256 (N_5256,N_3328,N_3214);
xor U5257 (N_5257,N_4754,N_3935);
nor U5258 (N_5258,N_4305,N_2747);
xor U5259 (N_5259,N_3914,N_4788);
and U5260 (N_5260,N_2577,N_4917);
xnor U5261 (N_5261,N_3073,N_4421);
and U5262 (N_5262,N_2582,N_4228);
or U5263 (N_5263,N_3401,N_4909);
xnor U5264 (N_5264,N_2990,N_4690);
and U5265 (N_5265,N_4660,N_4102);
and U5266 (N_5266,N_3563,N_3510);
and U5267 (N_5267,N_3403,N_3987);
or U5268 (N_5268,N_4161,N_3994);
and U5269 (N_5269,N_4050,N_3415);
and U5270 (N_5270,N_3591,N_3712);
and U5271 (N_5271,N_3336,N_4267);
nor U5272 (N_5272,N_3165,N_3331);
nor U5273 (N_5273,N_2642,N_3038);
or U5274 (N_5274,N_4099,N_4182);
or U5275 (N_5275,N_2503,N_4183);
xor U5276 (N_5276,N_3250,N_4203);
and U5277 (N_5277,N_4428,N_2988);
xnor U5278 (N_5278,N_4240,N_2978);
xor U5279 (N_5279,N_4173,N_4513);
nor U5280 (N_5280,N_2717,N_4635);
nand U5281 (N_5281,N_3891,N_4649);
nand U5282 (N_5282,N_2551,N_3939);
xnor U5283 (N_5283,N_4143,N_4519);
xor U5284 (N_5284,N_3931,N_3431);
and U5285 (N_5285,N_4673,N_2975);
nand U5286 (N_5286,N_3618,N_4593);
and U5287 (N_5287,N_3084,N_2946);
nor U5288 (N_5288,N_3841,N_4878);
or U5289 (N_5289,N_2783,N_3612);
nor U5290 (N_5290,N_3686,N_3737);
or U5291 (N_5291,N_4594,N_3681);
nor U5292 (N_5292,N_3607,N_2819);
and U5293 (N_5293,N_2873,N_3663);
xnor U5294 (N_5294,N_2839,N_2612);
and U5295 (N_5295,N_4611,N_3035);
or U5296 (N_5296,N_3310,N_3020);
and U5297 (N_5297,N_2932,N_3863);
xnor U5298 (N_5298,N_2734,N_3809);
xor U5299 (N_5299,N_3211,N_4619);
xnor U5300 (N_5300,N_4242,N_4681);
or U5301 (N_5301,N_4575,N_4354);
and U5302 (N_5302,N_4652,N_4313);
nor U5303 (N_5303,N_4555,N_3006);
xor U5304 (N_5304,N_2705,N_4770);
nor U5305 (N_5305,N_4650,N_3451);
nor U5306 (N_5306,N_2714,N_4940);
and U5307 (N_5307,N_2656,N_4147);
and U5308 (N_5308,N_3908,N_2562);
nand U5309 (N_5309,N_4869,N_4527);
nand U5310 (N_5310,N_2777,N_2931);
nor U5311 (N_5311,N_4782,N_3083);
and U5312 (N_5312,N_3746,N_4287);
and U5313 (N_5313,N_3554,N_3902);
nor U5314 (N_5314,N_3135,N_4130);
xor U5315 (N_5315,N_4458,N_3147);
xnor U5316 (N_5316,N_4376,N_3168);
or U5317 (N_5317,N_4249,N_3571);
xnor U5318 (N_5318,N_2972,N_4943);
nor U5319 (N_5319,N_2575,N_4112);
nor U5320 (N_5320,N_4648,N_3755);
nand U5321 (N_5321,N_3494,N_2816);
nor U5322 (N_5322,N_3553,N_4368);
nor U5323 (N_5323,N_4843,N_3466);
nor U5324 (N_5324,N_2826,N_3423);
or U5325 (N_5325,N_2674,N_2599);
xor U5326 (N_5326,N_3110,N_3750);
nand U5327 (N_5327,N_3174,N_3456);
nor U5328 (N_5328,N_3177,N_4170);
nand U5329 (N_5329,N_4461,N_4912);
and U5330 (N_5330,N_3164,N_3301);
nor U5331 (N_5331,N_3040,N_4270);
xor U5332 (N_5332,N_4330,N_3967);
and U5333 (N_5333,N_3611,N_2743);
and U5334 (N_5334,N_3029,N_3924);
nor U5335 (N_5335,N_3594,N_4920);
or U5336 (N_5336,N_3522,N_4316);
nor U5337 (N_5337,N_3089,N_4085);
nand U5338 (N_5338,N_3620,N_3232);
and U5339 (N_5339,N_4742,N_4284);
or U5340 (N_5340,N_3887,N_3285);
and U5341 (N_5341,N_2632,N_3324);
nor U5342 (N_5342,N_4674,N_2687);
xnor U5343 (N_5343,N_2621,N_4992);
nor U5344 (N_5344,N_3458,N_3337);
and U5345 (N_5345,N_3775,N_3047);
or U5346 (N_5346,N_3912,N_2913);
nor U5347 (N_5347,N_3625,N_3273);
nor U5348 (N_5348,N_2614,N_2600);
or U5349 (N_5349,N_4360,N_3855);
or U5350 (N_5350,N_4925,N_2941);
nand U5351 (N_5351,N_4653,N_3817);
xnor U5352 (N_5352,N_3375,N_3380);
nand U5353 (N_5353,N_3400,N_3646);
or U5354 (N_5354,N_4282,N_3224);
nand U5355 (N_5355,N_4515,N_2689);
and U5356 (N_5356,N_3113,N_3429);
nor U5357 (N_5357,N_3687,N_4928);
xnor U5358 (N_5358,N_3441,N_4308);
nor U5359 (N_5359,N_3942,N_4453);
and U5360 (N_5360,N_2602,N_2918);
nand U5361 (N_5361,N_2584,N_3131);
or U5362 (N_5362,N_2637,N_3711);
or U5363 (N_5363,N_4576,N_2814);
and U5364 (N_5364,N_4201,N_2811);
nand U5365 (N_5365,N_4984,N_3816);
or U5366 (N_5366,N_3859,N_2793);
and U5367 (N_5367,N_4571,N_4977);
nand U5368 (N_5368,N_3395,N_3381);
xnor U5369 (N_5369,N_3017,N_3198);
xnor U5370 (N_5370,N_4910,N_3596);
and U5371 (N_5371,N_3291,N_2952);
and U5372 (N_5372,N_4481,N_4281);
xnor U5373 (N_5373,N_3997,N_4278);
nand U5374 (N_5374,N_2647,N_3226);
xor U5375 (N_5375,N_2535,N_3302);
nor U5376 (N_5376,N_3885,N_4845);
nand U5377 (N_5377,N_3972,N_3416);
nand U5378 (N_5378,N_3661,N_3531);
or U5379 (N_5379,N_2863,N_4678);
nand U5380 (N_5380,N_4618,N_4230);
nor U5381 (N_5381,N_3504,N_4654);
nor U5382 (N_5382,N_2636,N_3345);
xnor U5383 (N_5383,N_3761,N_4793);
and U5384 (N_5384,N_3837,N_4951);
nand U5385 (N_5385,N_4559,N_3445);
xnor U5386 (N_5386,N_2964,N_3469);
xor U5387 (N_5387,N_2766,N_4514);
and U5388 (N_5388,N_4218,N_4854);
or U5389 (N_5389,N_4087,N_4413);
and U5390 (N_5390,N_3754,N_3631);
nand U5391 (N_5391,N_2849,N_4423);
and U5392 (N_5392,N_3830,N_2519);
nor U5393 (N_5393,N_4027,N_3412);
xnor U5394 (N_5394,N_3452,N_4626);
nor U5395 (N_5395,N_3311,N_2707);
or U5396 (N_5396,N_2810,N_3474);
nand U5397 (N_5397,N_4008,N_4918);
or U5398 (N_5398,N_3022,N_3348);
nor U5399 (N_5399,N_4152,N_4488);
nand U5400 (N_5400,N_2933,N_3141);
and U5401 (N_5401,N_3387,N_3333);
nor U5402 (N_5402,N_4463,N_4820);
and U5403 (N_5403,N_3982,N_2501);
nand U5404 (N_5404,N_4150,N_3703);
nand U5405 (N_5405,N_2772,N_4729);
nor U5406 (N_5406,N_2916,N_3664);
xor U5407 (N_5407,N_4709,N_3463);
nand U5408 (N_5408,N_3604,N_4901);
and U5409 (N_5409,N_4662,N_2998);
and U5410 (N_5410,N_3890,N_3668);
and U5411 (N_5411,N_3540,N_3111);
nor U5412 (N_5412,N_2950,N_4562);
xnor U5413 (N_5413,N_2610,N_4728);
and U5414 (N_5414,N_3881,N_3895);
nand U5415 (N_5415,N_3952,N_3785);
and U5416 (N_5416,N_3776,N_4352);
or U5417 (N_5417,N_3326,N_3351);
xor U5418 (N_5418,N_4954,N_4088);
nand U5419 (N_5419,N_3503,N_3335);
nor U5420 (N_5420,N_4680,N_4939);
nand U5421 (N_5421,N_3122,N_4627);
or U5422 (N_5422,N_3359,N_4356);
nand U5423 (N_5423,N_3799,N_4944);
and U5424 (N_5424,N_2776,N_4927);
or U5425 (N_5425,N_3606,N_4864);
nor U5426 (N_5426,N_3689,N_4895);
and U5427 (N_5427,N_4046,N_3460);
and U5428 (N_5428,N_4824,N_3229);
and U5429 (N_5429,N_3752,N_4487);
nand U5430 (N_5430,N_2526,N_4698);
xnor U5431 (N_5431,N_2715,N_3421);
nor U5432 (N_5432,N_4149,N_4898);
or U5433 (N_5433,N_3379,N_3962);
or U5434 (N_5434,N_3950,N_3645);
or U5435 (N_5435,N_4879,N_2903);
and U5436 (N_5436,N_3907,N_3747);
xnor U5437 (N_5437,N_3448,N_3694);
nand U5438 (N_5438,N_4830,N_2695);
nand U5439 (N_5439,N_4056,N_4746);
or U5440 (N_5440,N_3547,N_3438);
or U5441 (N_5441,N_2559,N_3309);
or U5442 (N_5442,N_4253,N_4233);
nand U5443 (N_5443,N_4836,N_4625);
nand U5444 (N_5444,N_3414,N_2723);
and U5445 (N_5445,N_4315,N_3449);
or U5446 (N_5446,N_3092,N_3702);
xor U5447 (N_5447,N_4962,N_2521);
nor U5448 (N_5448,N_2895,N_3722);
xor U5449 (N_5449,N_4159,N_2716);
and U5450 (N_5450,N_3180,N_4005);
or U5451 (N_5451,N_2999,N_3739);
nor U5452 (N_5452,N_4296,N_3495);
nor U5453 (N_5453,N_3422,N_4131);
and U5454 (N_5454,N_3628,N_4531);
and U5455 (N_5455,N_3610,N_4748);
nor U5456 (N_5456,N_4780,N_4876);
nand U5457 (N_5457,N_4071,N_4058);
or U5458 (N_5458,N_4107,N_4818);
xnor U5459 (N_5459,N_2852,N_4232);
nor U5460 (N_5460,N_2563,N_4817);
or U5461 (N_5461,N_4676,N_4327);
nand U5462 (N_5462,N_2771,N_2851);
xnor U5463 (N_5463,N_4403,N_4715);
and U5464 (N_5464,N_3430,N_3853);
or U5465 (N_5465,N_4066,N_3748);
xor U5466 (N_5466,N_4077,N_2940);
xor U5467 (N_5467,N_3544,N_4190);
and U5468 (N_5468,N_4311,N_4638);
nand U5469 (N_5469,N_4537,N_4372);
nor U5470 (N_5470,N_3261,N_4866);
nand U5471 (N_5471,N_3292,N_4092);
or U5472 (N_5472,N_4044,N_3015);
nor U5473 (N_5473,N_3844,N_2506);
xnor U5474 (N_5474,N_4582,N_3314);
xor U5475 (N_5475,N_3189,N_4364);
and U5476 (N_5476,N_4506,N_3639);
and U5477 (N_5477,N_4140,N_3813);
xor U5478 (N_5478,N_3263,N_3779);
or U5479 (N_5479,N_4760,N_4166);
nor U5480 (N_5480,N_3201,N_4651);
or U5481 (N_5481,N_3382,N_2915);
and U5482 (N_5482,N_4451,N_2576);
xnor U5483 (N_5483,N_2678,N_3649);
nand U5484 (N_5484,N_3979,N_3652);
and U5485 (N_5485,N_4167,N_4052);
xnor U5486 (N_5486,N_3526,N_2808);
nand U5487 (N_5487,N_3410,N_4553);
nor U5488 (N_5488,N_3091,N_3678);
and U5489 (N_5489,N_4695,N_2904);
and U5490 (N_5490,N_3353,N_2867);
and U5491 (N_5491,N_3500,N_4404);
and U5492 (N_5492,N_4713,N_4717);
xnor U5493 (N_5493,N_3185,N_3036);
xnor U5494 (N_5494,N_4081,N_3172);
xor U5495 (N_5495,N_4369,N_4361);
or U5496 (N_5496,N_4226,N_4620);
nand U5497 (N_5497,N_3619,N_2955);
xnor U5498 (N_5498,N_4379,N_3127);
xor U5499 (N_5499,N_4393,N_4707);
nand U5500 (N_5500,N_2779,N_4510);
nand U5501 (N_5501,N_4930,N_3272);
nor U5502 (N_5502,N_3829,N_3426);
xor U5503 (N_5503,N_3152,N_2987);
nor U5504 (N_5504,N_4156,N_4518);
and U5505 (N_5505,N_3812,N_2670);
nand U5506 (N_5506,N_3823,N_3742);
and U5507 (N_5507,N_3990,N_4769);
xor U5508 (N_5508,N_4806,N_4524);
or U5509 (N_5509,N_2830,N_3059);
and U5510 (N_5510,N_2504,N_2677);
nor U5511 (N_5511,N_3960,N_3509);
and U5512 (N_5512,N_4275,N_4238);
nor U5513 (N_5513,N_3117,N_3052);
or U5514 (N_5514,N_4541,N_3593);
and U5515 (N_5515,N_3293,N_2898);
nand U5516 (N_5516,N_2721,N_3851);
nand U5517 (N_5517,N_2997,N_3366);
xnor U5518 (N_5518,N_2638,N_4857);
nor U5519 (N_5519,N_2694,N_3190);
nand U5520 (N_5520,N_3097,N_4629);
xor U5521 (N_5521,N_4015,N_3904);
nand U5522 (N_5522,N_2966,N_3384);
nand U5523 (N_5523,N_3585,N_3104);
xnor U5524 (N_5524,N_3132,N_4849);
nor U5525 (N_5525,N_3069,N_3943);
xnor U5526 (N_5526,N_2553,N_2891);
or U5527 (N_5527,N_2976,N_4304);
and U5528 (N_5528,N_3791,N_3714);
xor U5529 (N_5529,N_4724,N_4454);
nand U5530 (N_5530,N_4462,N_3376);
and U5531 (N_5531,N_3468,N_3903);
xnor U5532 (N_5532,N_3256,N_3394);
nand U5533 (N_5533,N_3317,N_3202);
and U5534 (N_5534,N_2626,N_3969);
or U5535 (N_5535,N_3843,N_2573);
nand U5536 (N_5536,N_3369,N_4222);
xor U5537 (N_5537,N_4781,N_3454);
and U5538 (N_5538,N_3723,N_3579);
and U5539 (N_5539,N_4657,N_2920);
xor U5540 (N_5540,N_4710,N_3371);
xor U5541 (N_5541,N_4388,N_2896);
nand U5542 (N_5542,N_2595,N_4646);
and U5543 (N_5543,N_3014,N_4528);
nor U5544 (N_5544,N_3698,N_4913);
nor U5545 (N_5545,N_4444,N_4757);
or U5546 (N_5546,N_3701,N_3444);
xor U5547 (N_5547,N_3856,N_4777);
and U5548 (N_5548,N_4125,N_3313);
nand U5549 (N_5549,N_2882,N_3944);
and U5550 (N_5550,N_2765,N_3567);
or U5551 (N_5551,N_3329,N_4342);
and U5552 (N_5552,N_4682,N_4135);
xor U5553 (N_5553,N_4018,N_4500);
xor U5554 (N_5554,N_3778,N_3278);
nor U5555 (N_5555,N_4438,N_2528);
and U5556 (N_5556,N_4948,N_4811);
nor U5557 (N_5557,N_3683,N_4888);
and U5558 (N_5558,N_2789,N_3936);
nand U5559 (N_5559,N_2639,N_3433);
or U5560 (N_5560,N_3039,N_3917);
nand U5561 (N_5561,N_3282,N_3995);
nand U5562 (N_5562,N_2731,N_2644);
or U5563 (N_5563,N_4637,N_4966);
or U5564 (N_5564,N_2604,N_4563);
and U5565 (N_5565,N_3133,N_4790);
xnor U5566 (N_5566,N_3577,N_2786);
and U5567 (N_5567,N_3338,N_4733);
or U5568 (N_5568,N_4412,N_4968);
nand U5569 (N_5569,N_3357,N_4073);
nor U5570 (N_5570,N_4250,N_4775);
and U5571 (N_5571,N_4589,N_4569);
xor U5572 (N_5572,N_3916,N_2741);
or U5573 (N_5573,N_2818,N_3109);
and U5574 (N_5574,N_4029,N_2651);
xnor U5575 (N_5575,N_4675,N_4430);
and U5576 (N_5576,N_4865,N_4185);
or U5577 (N_5577,N_3481,N_3186);
xnor U5578 (N_5578,N_4139,N_3633);
and U5579 (N_5579,N_4084,N_3636);
nor U5580 (N_5580,N_3574,N_3847);
nor U5581 (N_5581,N_4471,N_2804);
or U5582 (N_5582,N_4955,N_3170);
and U5583 (N_5583,N_4826,N_4320);
or U5584 (N_5584,N_4568,N_2821);
nor U5585 (N_5585,N_4416,N_4326);
nand U5586 (N_5586,N_3397,N_2557);
xnor U5587 (N_5587,N_4076,N_4988);
and U5588 (N_5588,N_4871,N_4007);
nor U5589 (N_5589,N_3334,N_2962);
or U5590 (N_5590,N_3279,N_3524);
nor U5591 (N_5591,N_3697,N_4346);
xor U5592 (N_5592,N_3062,N_2959);
or U5593 (N_5593,N_3557,N_3148);
nor U5594 (N_5594,N_3815,N_2505);
nand U5595 (N_5595,N_3848,N_3061);
nand U5596 (N_5596,N_3074,N_2661);
and U5597 (N_5597,N_2756,N_3992);
nor U5598 (N_5598,N_3762,N_4743);
nor U5599 (N_5599,N_2877,N_2623);
and U5600 (N_5600,N_3125,N_3653);
or U5601 (N_5601,N_3247,N_2543);
nand U5602 (N_5602,N_4692,N_4155);
or U5603 (N_5603,N_4039,N_4205);
or U5604 (N_5604,N_3832,N_3674);
nor U5605 (N_5605,N_2755,N_4814);
and U5606 (N_5606,N_4981,N_4011);
nand U5607 (N_5607,N_4225,N_2712);
nor U5608 (N_5608,N_3404,N_4905);
or U5609 (N_5609,N_3756,N_3704);
nand U5610 (N_5610,N_2538,N_2643);
xnor U5611 (N_5611,N_4070,N_3941);
or U5612 (N_5612,N_4666,N_3044);
nor U5613 (N_5613,N_4062,N_2592);
xor U5614 (N_5614,N_4366,N_4101);
nor U5615 (N_5615,N_2866,N_4938);
or U5616 (N_5616,N_4547,N_3613);
nand U5617 (N_5617,N_4856,N_2681);
or U5618 (N_5618,N_3305,N_2948);
xor U5619 (N_5619,N_4716,N_4405);
xor U5620 (N_5620,N_4197,N_3601);
nor U5621 (N_5621,N_3257,N_4259);
or U5622 (N_5622,N_3362,N_2663);
and U5623 (N_5623,N_3096,N_4186);
nand U5624 (N_5624,N_4432,N_2722);
nand U5625 (N_5625,N_3055,N_4329);
or U5626 (N_5626,N_3502,N_4176);
nand U5627 (N_5627,N_2633,N_3396);
and U5628 (N_5628,N_3991,N_2580);
or U5629 (N_5629,N_3306,N_4588);
or U5630 (N_5630,N_4945,N_2847);
or U5631 (N_5631,N_4127,N_3724);
xor U5632 (N_5632,N_4941,N_2951);
xor U5633 (N_5633,N_3368,N_3892);
nand U5634 (N_5634,N_3389,N_4427);
nand U5635 (N_5635,N_2525,N_3192);
nand U5636 (N_5636,N_4319,N_2546);
nor U5637 (N_5637,N_2919,N_3205);
nor U5638 (N_5638,N_4933,N_3818);
or U5639 (N_5639,N_4199,N_2620);
nand U5640 (N_5640,N_3507,N_3957);
and U5641 (N_5641,N_3277,N_3882);
nor U5642 (N_5642,N_2625,N_2510);
or U5643 (N_5643,N_4490,N_3116);
nor U5644 (N_5644,N_3641,N_4505);
nand U5645 (N_5645,N_4344,N_3374);
or U5646 (N_5646,N_4051,N_3070);
xnor U5647 (N_5647,N_4108,N_4020);
and U5648 (N_5648,N_4810,N_4893);
or U5649 (N_5649,N_3280,N_4566);
nor U5650 (N_5650,N_3559,N_4254);
or U5651 (N_5651,N_2619,N_4990);
nand U5652 (N_5652,N_3080,N_3341);
nor U5653 (N_5653,N_2871,N_4985);
and U5654 (N_5654,N_3741,N_3753);
or U5655 (N_5655,N_3568,N_4745);
or U5656 (N_5656,N_4494,N_4394);
or U5657 (N_5657,N_3523,N_4838);
nand U5658 (N_5658,N_4522,N_2667);
nor U5659 (N_5659,N_3659,N_4323);
xor U5660 (N_5660,N_4063,N_4801);
nand U5661 (N_5661,N_4169,N_3810);
xor U5662 (N_5662,N_3940,N_2749);
or U5663 (N_5663,N_3087,N_2763);
and U5664 (N_5664,N_2539,N_2874);
and U5665 (N_5665,N_3970,N_4994);
or U5666 (N_5666,N_3768,N_4310);
nand U5667 (N_5667,N_2533,N_4739);
nand U5668 (N_5668,N_3835,N_2634);
or U5669 (N_5669,N_4065,N_4472);
and U5670 (N_5670,N_3484,N_3520);
xnor U5671 (N_5671,N_3046,N_3048);
or U5672 (N_5672,N_3473,N_3243);
and U5673 (N_5673,N_4353,N_4455);
xnor U5674 (N_5674,N_3735,N_4916);
and U5675 (N_5675,N_4221,N_3521);
or U5676 (N_5676,N_4142,N_2507);
xnor U5677 (N_5677,N_4258,N_4164);
nand U5678 (N_5678,N_3435,N_4642);
xor U5679 (N_5679,N_4019,N_4535);
xor U5680 (N_5680,N_4960,N_2590);
nor U5681 (N_5681,N_2574,N_4105);
xnor U5682 (N_5682,N_4174,N_3730);
or U5683 (N_5683,N_4373,N_3432);
and U5684 (N_5684,N_3424,N_2781);
xor U5685 (N_5685,N_3215,N_4517);
nor U5686 (N_5686,N_4072,N_3548);
nand U5687 (N_5687,N_2885,N_4641);
nand U5688 (N_5688,N_3169,N_3041);
nand U5689 (N_5689,N_3260,N_2567);
xnor U5690 (N_5690,N_3699,N_3665);
or U5691 (N_5691,N_2554,N_3977);
nand U5692 (N_5692,N_3974,N_3390);
and U5693 (N_5693,N_4771,N_4672);
nor U5694 (N_5694,N_4367,N_3312);
or U5695 (N_5695,N_2890,N_3582);
nand U5696 (N_5696,N_2878,N_3385);
or U5697 (N_5697,N_3586,N_3378);
nand U5698 (N_5698,N_4550,N_3749);
and U5699 (N_5699,N_3230,N_2792);
nor U5700 (N_5700,N_2664,N_2550);
xnor U5701 (N_5701,N_4860,N_3705);
and U5702 (N_5702,N_3828,N_2702);
nor U5703 (N_5703,N_3508,N_4288);
and U5704 (N_5704,N_4949,N_3077);
nand U5705 (N_5705,N_4979,N_4964);
nor U5706 (N_5706,N_4887,N_3680);
and U5707 (N_5707,N_3529,N_4184);
or U5708 (N_5708,N_3343,N_4772);
xor U5709 (N_5709,N_4827,N_3537);
nand U5710 (N_5710,N_4982,N_4829);
nand U5711 (N_5711,N_3407,N_4663);
or U5712 (N_5712,N_3862,N_4217);
nor U5713 (N_5713,N_2875,N_4883);
xnor U5714 (N_5714,N_3796,N_2531);
and U5715 (N_5715,N_3218,N_4787);
xnor U5716 (N_5716,N_3806,N_4890);
and U5717 (N_5717,N_2911,N_4442);
nand U5718 (N_5718,N_3986,N_4163);
or U5719 (N_5719,N_3715,N_4750);
xnor U5720 (N_5720,N_3988,N_3672);
or U5721 (N_5721,N_2762,N_4591);
nand U5722 (N_5722,N_3228,N_4297);
or U5723 (N_5723,N_3906,N_3248);
and U5724 (N_5724,N_2778,N_3938);
or U5725 (N_5725,N_2532,N_3803);
and U5726 (N_5726,N_3845,N_2917);
xnor U5727 (N_5727,N_2888,N_3781);
nor U5728 (N_5728,N_3330,N_4452);
nor U5729 (N_5729,N_4198,N_4103);
and U5730 (N_5730,N_2815,N_4382);
nor U5731 (N_5731,N_3927,N_3128);
nor U5732 (N_5732,N_3888,N_3146);
and U5733 (N_5733,N_2568,N_2944);
nor U5734 (N_5734,N_2861,N_3792);
or U5735 (N_5735,N_2844,N_3085);
and U5736 (N_5736,N_2607,N_2653);
xnor U5737 (N_5737,N_3490,N_2799);
nor U5738 (N_5738,N_4614,N_4384);
or U5739 (N_5739,N_4693,N_3720);
and U5740 (N_5740,N_2876,N_3831);
or U5741 (N_5741,N_3143,N_4469);
or U5742 (N_5742,N_4751,N_3738);
or U5743 (N_5743,N_4090,N_3099);
xnor U5744 (N_5744,N_3790,N_4211);
and U5745 (N_5745,N_3303,N_3327);
nor U5746 (N_5746,N_4350,N_3536);
or U5747 (N_5747,N_4796,N_4704);
xnor U5748 (N_5748,N_3556,N_3063);
nand U5749 (N_5749,N_2704,N_2854);
xnor U5750 (N_5750,N_2710,N_3437);
nor U5751 (N_5751,N_3513,N_4923);
or U5752 (N_5752,N_4607,N_4285);
nand U5753 (N_5753,N_3981,N_3733);
xnor U5754 (N_5754,N_4307,N_4425);
or U5755 (N_5755,N_4196,N_4549);
or U5756 (N_5756,N_4752,N_3299);
and U5757 (N_5757,N_3918,N_4711);
or U5758 (N_5758,N_3934,N_2635);
or U5759 (N_5759,N_4243,N_3095);
and U5760 (N_5760,N_2542,N_4509);
xnor U5761 (N_5761,N_3833,N_3003);
xor U5762 (N_5762,N_3187,N_3615);
nor U5763 (N_5763,N_2843,N_2801);
or U5764 (N_5764,N_4321,N_4723);
xor U5765 (N_5765,N_4936,N_3743);
nor U5766 (N_5766,N_3031,N_3498);
nand U5767 (N_5767,N_2986,N_3479);
or U5768 (N_5768,N_4502,N_4162);
nor U5769 (N_5769,N_2517,N_3491);
and U5770 (N_5770,N_4338,N_2970);
xnor U5771 (N_5771,N_3142,N_4496);
and U5772 (N_5772,N_3654,N_2508);
nand U5773 (N_5773,N_3946,N_2693);
and U5774 (N_5774,N_2824,N_4560);
nand U5775 (N_5775,N_4035,N_3959);
or U5776 (N_5776,N_2654,N_2591);
nor U5777 (N_5777,N_4699,N_2530);
nor U5778 (N_5778,N_4257,N_2922);
nor U5779 (N_5779,N_2631,N_2757);
xnor U5780 (N_5780,N_3773,N_2737);
nor U5781 (N_5781,N_3865,N_3115);
nand U5782 (N_5782,N_3209,N_3482);
and U5783 (N_5783,N_4440,N_4655);
nor U5784 (N_5784,N_2902,N_4586);
nand U5785 (N_5785,N_2973,N_3629);
nor U5786 (N_5786,N_3569,N_3771);
and U5787 (N_5787,N_4079,N_3081);
or U5788 (N_5788,N_4260,N_3644);
xnor U5789 (N_5789,N_2823,N_2669);
xor U5790 (N_5790,N_2812,N_4903);
and U5791 (N_5791,N_3045,N_2608);
nor U5792 (N_5792,N_3637,N_3871);
nor U5793 (N_5793,N_4298,N_2981);
nand U5794 (N_5794,N_2840,N_3647);
nor U5795 (N_5795,N_3578,N_3176);
or U5796 (N_5796,N_3033,N_3728);
nand U5797 (N_5797,N_3064,N_4038);
and U5798 (N_5798,N_4705,N_2544);
or U5799 (N_5799,N_2813,N_3614);
xnor U5800 (N_5800,N_4873,N_3024);
nand U5801 (N_5801,N_3838,N_4293);
nor U5802 (N_5802,N_4419,N_3101);
nor U5803 (N_5803,N_3057,N_4832);
or U5804 (N_5804,N_4859,N_3984);
xnor U5805 (N_5805,N_3450,N_2899);
nor U5806 (N_5806,N_3093,N_4516);
nor U5807 (N_5807,N_4578,N_3565);
and U5808 (N_5808,N_4000,N_4573);
nor U5809 (N_5809,N_3693,N_4815);
nand U5810 (N_5810,N_3236,N_2982);
and U5811 (N_5811,N_2680,N_4231);
and U5812 (N_5812,N_3671,N_2859);
xnor U5813 (N_5813,N_4986,N_4082);
or U5814 (N_5814,N_2630,N_3667);
or U5815 (N_5815,N_2515,N_4969);
nor U5816 (N_5816,N_3253,N_2648);
nor U5817 (N_5817,N_3442,N_4068);
nand U5818 (N_5818,N_4359,N_4564);
nand U5819 (N_5819,N_4370,N_4117);
and U5820 (N_5820,N_3477,N_2797);
and U5821 (N_5821,N_4899,N_3319);
nand U5822 (N_5822,N_4255,N_2796);
xor U5823 (N_5823,N_3643,N_3220);
or U5824 (N_5824,N_3576,N_4691);
xnor U5825 (N_5825,N_2516,N_4802);
and U5826 (N_5826,N_3573,N_2939);
nand U5827 (N_5827,N_4734,N_2736);
and U5828 (N_5828,N_4570,N_4484);
xnor U5829 (N_5829,N_3259,N_4235);
nor U5830 (N_5830,N_4389,N_4280);
or U5831 (N_5831,N_2949,N_3239);
nor U5832 (N_5832,N_3602,N_4269);
nand U5833 (N_5833,N_4054,N_4449);
nand U5834 (N_5834,N_4671,N_2502);
xnor U5835 (N_5835,N_4789,N_3708);
nand U5836 (N_5836,N_4385,N_4501);
or U5837 (N_5837,N_3948,N_4314);
xnor U5838 (N_5838,N_3001,N_4292);
nand U5839 (N_5839,N_3905,N_4609);
nand U5840 (N_5840,N_3876,N_4753);
xnor U5841 (N_5841,N_4165,N_4580);
and U5842 (N_5842,N_3076,N_4679);
xnor U5843 (N_5843,N_3088,N_3406);
and U5844 (N_5844,N_4435,N_3470);
or U5845 (N_5845,N_4436,N_4333);
nand U5846 (N_5846,N_4929,N_4983);
or U5847 (N_5847,N_4261,N_4171);
nor U5848 (N_5848,N_3235,N_2541);
xnor U5849 (N_5849,N_4443,N_3275);
and U5850 (N_5850,N_4819,N_3605);
nor U5851 (N_5851,N_4840,N_4216);
or U5852 (N_5852,N_4083,N_4993);
and U5853 (N_5853,N_4031,N_3608);
or U5854 (N_5854,N_2782,N_3673);
or U5855 (N_5855,N_3213,N_2696);
or U5856 (N_5856,N_3583,N_4470);
nand U5857 (N_5857,N_2848,N_3157);
or U5858 (N_5858,N_4644,N_4557);
and U5859 (N_5859,N_2968,N_2969);
nor U5860 (N_5860,N_4126,N_2806);
nand U5861 (N_5861,N_3740,N_2767);
and U5862 (N_5862,N_3242,N_4778);
nand U5863 (N_5863,N_3289,N_4604);
or U5864 (N_5864,N_4465,N_4086);
and U5865 (N_5865,N_3922,N_2761);
nand U5866 (N_5866,N_4114,N_4202);
xor U5867 (N_5867,N_4612,N_4735);
or U5868 (N_5868,N_2943,N_4886);
or U5869 (N_5869,N_4615,N_4055);
nor U5870 (N_5870,N_2713,N_3332);
nand U5871 (N_5871,N_4302,N_3402);
nand U5872 (N_5872,N_4779,N_2754);
nor U5873 (N_5873,N_4213,N_4572);
nor U5874 (N_5874,N_2724,N_4493);
xor U5875 (N_5875,N_2725,N_4247);
or U5876 (N_5876,N_3323,N_4229);
nand U5877 (N_5877,N_4600,N_4429);
and U5878 (N_5878,N_2817,N_3255);
nor U5879 (N_5879,N_3913,N_3827);
or U5880 (N_5880,N_4349,N_3786);
xnor U5881 (N_5881,N_4530,N_4121);
xor U5882 (N_5882,N_3405,N_4100);
nor U5883 (N_5883,N_2977,N_4786);
xnor U5884 (N_5884,N_4783,N_4908);
nand U5885 (N_5885,N_4558,N_3546);
nand U5886 (N_5886,N_3820,N_4220);
xnor U5887 (N_5887,N_3124,N_4997);
and U5888 (N_5888,N_4340,N_2511);
and U5889 (N_5889,N_2892,N_2753);
xnor U5890 (N_5890,N_3870,N_4538);
xor U5891 (N_5891,N_2905,N_3016);
xor U5892 (N_5892,N_3465,N_3677);
xor U5893 (N_5893,N_3153,N_4727);
nand U5894 (N_5894,N_3126,N_3408);
and U5895 (N_5895,N_2961,N_4511);
and U5896 (N_5896,N_3707,N_3949);
nand U5897 (N_5897,N_3763,N_3050);
and U5898 (N_5898,N_3766,N_2730);
or U5899 (N_5899,N_3985,N_4244);
nand U5900 (N_5900,N_3222,N_3447);
xor U5901 (N_5901,N_3042,N_3199);
nand U5902 (N_5902,N_4823,N_4017);
or U5903 (N_5903,N_3262,N_4380);
nor U5904 (N_5904,N_3420,N_3428);
nor U5905 (N_5905,N_4119,N_3517);
xor U5906 (N_5906,N_2907,N_4885);
or U5907 (N_5907,N_4870,N_4059);
nand U5908 (N_5908,N_2512,N_3307);
nor U5909 (N_5909,N_3066,N_3032);
nand U5910 (N_5910,N_4978,N_3527);
nand U5911 (N_5911,N_3026,N_4294);
xor U5912 (N_5912,N_2679,N_3836);
and U5913 (N_5913,N_3499,N_4643);
nand U5914 (N_5914,N_3562,N_2858);
nor U5915 (N_5915,N_2593,N_4392);
nor U5916 (N_5916,N_4109,N_2739);
and U5917 (N_5917,N_3007,N_2522);
nand U5918 (N_5918,N_3717,N_4911);
nand U5919 (N_5919,N_3184,N_4022);
nand U5920 (N_5920,N_3363,N_4736);
nand U5921 (N_5921,N_4491,N_3805);
nand U5922 (N_5922,N_4546,N_4956);
xor U5923 (N_5923,N_4057,N_2979);
xor U5924 (N_5924,N_3120,N_4154);
nand U5925 (N_5925,N_3993,N_4623);
nand U5926 (N_5926,N_3162,N_4747);
or U5927 (N_5927,N_3539,N_4138);
nand U5928 (N_5928,N_2889,N_3538);
xor U5929 (N_5929,N_3800,N_4212);
or U5930 (N_5930,N_2750,N_4924);
nor U5931 (N_5931,N_4371,N_4552);
or U5932 (N_5932,N_4401,N_4976);
xor U5933 (N_5933,N_4033,N_3609);
nor U5934 (N_5934,N_4396,N_3485);
xnor U5935 (N_5935,N_2827,N_3534);
and U5936 (N_5936,N_3634,N_3492);
nand U5937 (N_5937,N_4958,N_3893);
and U5938 (N_5938,N_3210,N_4132);
nor U5939 (N_5939,N_4415,N_3919);
nand U5940 (N_5940,N_2556,N_4337);
and U5941 (N_5941,N_4656,N_2992);
or U5942 (N_5942,N_4113,N_4433);
and U5943 (N_5943,N_3149,N_3983);
nor U5944 (N_5944,N_2751,N_4485);
nor U5945 (N_5945,N_3237,N_4534);
nor U5946 (N_5946,N_3058,N_4613);
nor U5947 (N_5947,N_2513,N_2802);
nand U5948 (N_5948,N_4882,N_2784);
or U5949 (N_5949,N_3757,N_3284);
and U5950 (N_5950,N_4590,N_2666);
nand U5951 (N_5951,N_3873,N_3884);
and U5952 (N_5952,N_4622,N_4378);
xor U5953 (N_5953,N_4677,N_4239);
nand U5954 (N_5954,N_3372,N_2945);
or U5955 (N_5955,N_4991,N_4474);
and U5956 (N_5956,N_4014,N_3716);
and U5957 (N_5957,N_4475,N_2594);
nor U5958 (N_5958,N_2790,N_3798);
and U5959 (N_5959,N_4804,N_3684);
and U5960 (N_5960,N_4122,N_4447);
and U5961 (N_5961,N_3294,N_4701);
nor U5962 (N_5962,N_4365,N_2652);
or U5963 (N_5963,N_3879,N_3745);
nand U5964 (N_5964,N_4410,N_4042);
xnor U5965 (N_5965,N_4794,N_4041);
and U5966 (N_5966,N_4407,N_4706);
or U5967 (N_5967,N_4521,N_4325);
xor U5968 (N_5968,N_4256,N_3660);
nor U5969 (N_5969,N_3688,N_4540);
xnor U5970 (N_5970,N_4341,N_3340);
or U5971 (N_5971,N_3297,N_3976);
nand U5972 (N_5972,N_2838,N_4758);
or U5973 (N_5973,N_4884,N_4875);
and U5974 (N_5974,N_4016,N_3808);
xnor U5975 (N_5975,N_4048,N_2869);
and U5976 (N_5976,N_4931,N_4880);
nand U5977 (N_5977,N_3542,N_4585);
and U5978 (N_5978,N_2611,N_3386);
and U5979 (N_5979,N_3782,N_4118);
and U5980 (N_5980,N_4097,N_2752);
xnor U5981 (N_5981,N_3603,N_4381);
and U5982 (N_5982,N_3025,N_4290);
or U5983 (N_5983,N_4896,N_3360);
xnor U5984 (N_5984,N_2928,N_4694);
nor U5985 (N_5985,N_4703,N_3560);
and U5986 (N_5986,N_4919,N_4124);
and U5987 (N_5987,N_3079,N_3794);
nor U5988 (N_5988,N_3274,N_3290);
or U5989 (N_5989,N_2894,N_2881);
and U5990 (N_5990,N_3592,N_2947);
or U5991 (N_5991,N_4012,N_3367);
and U5992 (N_5992,N_3018,N_4610);
and U5993 (N_5993,N_4069,N_3789);
or U5994 (N_5994,N_4645,N_4157);
and U5995 (N_5995,N_4512,N_3251);
nand U5996 (N_5996,N_4708,N_4194);
or U5997 (N_5997,N_4850,N_4306);
and U5998 (N_5998,N_4630,N_4647);
nor U5999 (N_5999,N_2718,N_2906);
nor U6000 (N_6000,N_3354,N_3497);
nor U6001 (N_6001,N_2974,N_2676);
xnor U6002 (N_6002,N_2514,N_4457);
and U6003 (N_6003,N_2598,N_4868);
xnor U6004 (N_6004,N_2996,N_4347);
and U6005 (N_6005,N_3171,N_4300);
or U6006 (N_6006,N_4111,N_4688);
or U6007 (N_6007,N_3206,N_3635);
and U6008 (N_6008,N_3780,N_4476);
and U6009 (N_6009,N_3869,N_3315);
and U6010 (N_6010,N_4853,N_4634);
nand U6011 (N_6011,N_2868,N_4765);
nor U6012 (N_6012,N_4971,N_2518);
nand U6013 (N_6013,N_4299,N_2795);
nand U6014 (N_6014,N_3580,N_3690);
nand U6015 (N_6015,N_4599,N_4464);
and U6016 (N_6016,N_3188,N_2800);
nand U6017 (N_6017,N_4565,N_3864);
or U6018 (N_6018,N_3858,N_3512);
or U6019 (N_6019,N_2700,N_3200);
nand U6020 (N_6020,N_3483,N_2759);
nand U6021 (N_6021,N_3640,N_4336);
or U6022 (N_6022,N_3227,N_4234);
nand U6023 (N_6023,N_4934,N_2787);
xor U6024 (N_6024,N_4328,N_4851);
nor U6025 (N_6025,N_3597,N_3759);
nand U6026 (N_6026,N_2587,N_4807);
nor U6027 (N_6027,N_4825,N_3533);
nor U6028 (N_6028,N_2788,N_2914);
nor U6029 (N_6029,N_3158,N_4738);
nand U6030 (N_6030,N_4785,N_4915);
xor U6031 (N_6031,N_3514,N_4207);
nand U6032 (N_6032,N_4791,N_4277);
nor U6033 (N_6033,N_4797,N_4343);
xor U6034 (N_6034,N_4922,N_4831);
nand U6035 (N_6035,N_3419,N_4146);
nor U6036 (N_6036,N_4064,N_3383);
or U6037 (N_6037,N_3772,N_2720);
or U6038 (N_6038,N_3648,N_3103);
or U6039 (N_6039,N_3945,N_2887);
or U6040 (N_6040,N_4200,N_4574);
nor U6041 (N_6041,N_4556,N_4592);
xnor U6042 (N_6042,N_3725,N_2613);
nor U6043 (N_6043,N_4544,N_4792);
nand U6044 (N_6044,N_4104,N_4844);
nor U6045 (N_6045,N_4621,N_3221);
and U6046 (N_6046,N_4624,N_3344);
xor U6047 (N_6047,N_4740,N_4881);
or U6048 (N_6048,N_3439,N_2967);
and U6049 (N_6049,N_2520,N_4776);
nor U6050 (N_6050,N_3049,N_3822);
or U6051 (N_6051,N_4959,N_3364);
nand U6052 (N_6052,N_4543,N_4508);
nor U6053 (N_6053,N_4434,N_4204);
and U6054 (N_6054,N_4816,N_4668);
nor U6055 (N_6055,N_4633,N_3999);
nor U6056 (N_6056,N_4579,N_4636);
nor U6057 (N_6057,N_4053,N_2909);
nand U6058 (N_6058,N_2798,N_4145);
nand U6059 (N_6059,N_2835,N_4289);
or U6060 (N_6060,N_3078,N_4116);
and U6061 (N_6061,N_3388,N_3857);
xnor U6062 (N_6062,N_3930,N_4193);
and U6063 (N_6063,N_4689,N_3138);
and U6064 (N_6064,N_4841,N_2628);
nor U6065 (N_6065,N_4847,N_4702);
nand U6066 (N_6066,N_2853,N_4010);
nand U6067 (N_6067,N_3797,N_2641);
nor U6068 (N_6068,N_3662,N_3996);
nand U6069 (N_6069,N_3860,N_4021);
and U6070 (N_6070,N_2529,N_4437);
nand U6071 (N_6071,N_3175,N_3098);
nor U6072 (N_6072,N_2560,N_2930);
nor U6073 (N_6073,N_2732,N_3900);
nor U6074 (N_6074,N_3679,N_4078);
or U6075 (N_6075,N_4605,N_3676);
or U6076 (N_6076,N_4722,N_4661);
xnor U6077 (N_6077,N_3958,N_4616);
and U6078 (N_6078,N_4060,N_2566);
and U6079 (N_6079,N_2958,N_4542);
xnor U6080 (N_6080,N_4177,N_2596);
and U6081 (N_6081,N_4399,N_3617);
nor U6082 (N_6082,N_3358,N_3710);
xor U6083 (N_6083,N_3166,N_4168);
nand U6084 (N_6084,N_2746,N_4466);
nor U6085 (N_6085,N_4406,N_3487);
xor U6086 (N_6086,N_3308,N_4737);
nor U6087 (N_6087,N_4684,N_4719);
xor U6088 (N_6088,N_3219,N_2658);
nor U6089 (N_6089,N_4554,N_2699);
and U6090 (N_6090,N_3446,N_2698);
and U6091 (N_6091,N_4144,N_3392);
or U6092 (N_6092,N_3519,N_3658);
nand U6093 (N_6093,N_4523,N_3886);
nand U6094 (N_6094,N_3824,N_2934);
and U6095 (N_6095,N_4268,N_3130);
and U6096 (N_6096,N_3181,N_3599);
nand U6097 (N_6097,N_4061,N_4214);
nand U6098 (N_6098,N_3060,N_2872);
xor U6099 (N_6099,N_3889,N_4987);
or U6100 (N_6100,N_4759,N_2908);
xnor U6101 (N_6101,N_2690,N_4584);
xor U6102 (N_6102,N_3899,N_3321);
nand U6103 (N_6103,N_4744,N_4839);
or U6104 (N_6104,N_2671,N_4219);
nor U6105 (N_6105,N_3193,N_4725);
nand U6106 (N_6106,N_3043,N_2991);
xor U6107 (N_6107,N_3973,N_3023);
nor U6108 (N_6108,N_4670,N_4024);
nand U6109 (N_6109,N_3030,N_4067);
and U6110 (N_6110,N_2857,N_3814);
xnor U6111 (N_6111,N_3065,N_2809);
nand U6112 (N_6112,N_4141,N_3195);
and U6113 (N_6113,N_4632,N_4262);
nand U6114 (N_6114,N_4548,N_4700);
and U6115 (N_6115,N_4037,N_4714);
nand U6116 (N_6116,N_4764,N_3657);
xnor U6117 (N_6117,N_3642,N_3811);
nor U6118 (N_6118,N_3266,N_3121);
nand U6119 (N_6119,N_4414,N_3075);
nand U6120 (N_6120,N_3119,N_2589);
and U6121 (N_6121,N_4424,N_3802);
and U6122 (N_6122,N_4598,N_4074);
xnor U6123 (N_6123,N_2609,N_4148);
nor U6124 (N_6124,N_3316,N_2769);
xnor U6125 (N_6125,N_2659,N_3398);
nor U6126 (N_6126,N_4935,N_4946);
nor U6127 (N_6127,N_2624,N_4094);
xor U6128 (N_6128,N_3915,N_4499);
nand U6129 (N_6129,N_2901,N_3807);
nor U6130 (N_6130,N_4151,N_2957);
nand U6131 (N_6131,N_4975,N_4301);
xor U6132 (N_6132,N_4009,N_2682);
and U6133 (N_6133,N_3471,N_4608);
xor U6134 (N_6134,N_3373,N_3027);
xor U6135 (N_6135,N_4408,N_3880);
xor U6136 (N_6136,N_3322,N_4348);
or U6137 (N_6137,N_4617,N_4755);
or U6138 (N_6138,N_2726,N_4411);
nand U6139 (N_6139,N_4402,N_3223);
nor U6140 (N_6140,N_2834,N_3212);
or U6141 (N_6141,N_3478,N_3068);
or U6142 (N_6142,N_3765,N_4906);
and U6143 (N_6143,N_3675,N_3555);
and U6144 (N_6144,N_3682,N_3826);
and U6145 (N_6145,N_3627,N_2927);
xnor U6146 (N_6146,N_3550,N_4507);
xnor U6147 (N_6147,N_4989,N_3265);
and U6148 (N_6148,N_2842,N_3572);
nor U6149 (N_6149,N_4995,N_4687);
nand U6150 (N_6150,N_3549,N_4450);
nand U6151 (N_6151,N_3821,N_4628);
nor U6152 (N_6152,N_2570,N_4520);
nand U6153 (N_6153,N_3019,N_3225);
xor U6154 (N_6154,N_3496,N_3269);
and U6155 (N_6155,N_2688,N_3877);
or U6156 (N_6156,N_4749,N_4952);
xor U6157 (N_6157,N_4835,N_4852);
or U6158 (N_6158,N_3947,N_3581);
or U6159 (N_6159,N_4828,N_3744);
and U6160 (N_6160,N_2646,N_3588);
nor U6161 (N_6161,N_3528,N_3159);
and U6162 (N_6162,N_4480,N_3145);
or U6163 (N_6163,N_3009,N_3203);
and U6164 (N_6164,N_2692,N_3118);
or U6165 (N_6165,N_4272,N_4345);
or U6166 (N_6166,N_3616,N_3051);
nor U6167 (N_6167,N_3472,N_2588);
nand U6168 (N_6168,N_2709,N_3734);
nand U6169 (N_6169,N_2845,N_3108);
nor U6170 (N_6170,N_2803,N_4731);
xor U6171 (N_6171,N_2738,N_4795);
nand U6172 (N_6172,N_4597,N_4900);
nor U6173 (N_6173,N_4004,N_4439);
and U6174 (N_6174,N_4286,N_3695);
xor U6175 (N_6175,N_3276,N_3530);
nand U6176 (N_6176,N_4030,N_2770);
and U6177 (N_6177,N_4431,N_3283);
xor U6178 (N_6178,N_3718,N_4921);
and U6179 (N_6179,N_3361,N_2728);
xor U6180 (N_6180,N_4075,N_2708);
nor U6181 (N_6181,N_3692,N_3144);
nand U6182 (N_6182,N_2925,N_3086);
nor U6183 (N_6183,N_3670,N_2748);
and U6184 (N_6184,N_2616,N_3793);
nor U6185 (N_6185,N_3700,N_4904);
xor U6186 (N_6186,N_2965,N_3365);
nand U6187 (N_6187,N_3013,N_2744);
and U6188 (N_6188,N_3137,N_2921);
or U6189 (N_6189,N_4110,N_4417);
and U6190 (N_6190,N_3551,N_3901);
nor U6191 (N_6191,N_3440,N_2912);
or U6192 (N_6192,N_3954,N_2555);
xor U6193 (N_6193,N_3264,N_4741);
xor U6194 (N_6194,N_4028,N_4426);
xor U6195 (N_6195,N_4669,N_3736);
or U6196 (N_6196,N_3281,N_3476);
nand U6197 (N_6197,N_4942,N_2879);
or U6198 (N_6198,N_4420,N_2552);
xor U6199 (N_6199,N_2807,N_2963);
xnor U6200 (N_6200,N_4726,N_4129);
nor U6201 (N_6201,N_2650,N_4561);
nand U6202 (N_6202,N_4206,N_3685);
nand U6203 (N_6203,N_4763,N_2627);
or U6204 (N_6204,N_2910,N_3217);
xnor U6205 (N_6205,N_3669,N_4603);
nand U6206 (N_6206,N_3238,N_4833);
nor U6207 (N_6207,N_3425,N_4209);
xor U6208 (N_6208,N_2775,N_3758);
or U6209 (N_6209,N_4498,N_3011);
xnor U6210 (N_6210,N_3515,N_4685);
or U6211 (N_6211,N_2832,N_4418);
nand U6212 (N_6212,N_3008,N_3010);
xor U6213 (N_6213,N_3875,N_4172);
nor U6214 (N_6214,N_3989,N_3998);
or U6215 (N_6215,N_2870,N_4422);
or U6216 (N_6216,N_3167,N_3729);
or U6217 (N_6217,N_3854,N_3867);
nor U6218 (N_6218,N_3543,N_2954);
nand U6219 (N_6219,N_2605,N_2558);
or U6220 (N_6220,N_3861,N_3155);
nor U6221 (N_6221,N_4291,N_4581);
and U6222 (N_6222,N_2995,N_4467);
nor U6223 (N_6223,N_4892,N_3872);
xnor U6224 (N_6224,N_3570,N_4539);
nand U6225 (N_6225,N_2733,N_4227);
and U6226 (N_6226,N_2569,N_2768);
nor U6227 (N_6227,N_3511,N_4283);
and U6228 (N_6228,N_2865,N_3355);
or U6229 (N_6229,N_2836,N_4362);
and U6230 (N_6230,N_3183,N_2578);
or U6231 (N_6231,N_2929,N_3436);
or U6232 (N_6232,N_4667,N_3377);
and U6233 (N_6233,N_2924,N_4400);
and U6234 (N_6234,N_3933,N_4762);
and U6235 (N_6235,N_4456,N_4390);
or U6236 (N_6236,N_3650,N_2581);
xnor U6237 (N_6237,N_4179,N_3457);
xnor U6238 (N_6238,N_4583,N_4013);
xnor U6239 (N_6239,N_4812,N_3787);
and U6240 (N_6240,N_3965,N_4768);
xor U6241 (N_6241,N_2880,N_3696);
and U6242 (N_6242,N_2665,N_4245);
nor U6243 (N_6243,N_3929,N_3464);
xnor U6244 (N_6244,N_4664,N_3920);
and U6245 (N_6245,N_4187,N_3980);
nor U6246 (N_6246,N_3461,N_3584);
xor U6247 (N_6247,N_4863,N_3295);
nand U6248 (N_6248,N_2773,N_2983);
nor U6249 (N_6249,N_2980,N_3356);
xor U6250 (N_6250,N_3884,N_3231);
xor U6251 (N_6251,N_4803,N_3504);
and U6252 (N_6252,N_3874,N_3983);
nand U6253 (N_6253,N_2948,N_4429);
xnor U6254 (N_6254,N_2719,N_2944);
and U6255 (N_6255,N_3859,N_4548);
or U6256 (N_6256,N_3513,N_3279);
nor U6257 (N_6257,N_4886,N_2505);
and U6258 (N_6258,N_2670,N_3539);
and U6259 (N_6259,N_2634,N_3753);
nor U6260 (N_6260,N_4115,N_3226);
and U6261 (N_6261,N_4188,N_2848);
or U6262 (N_6262,N_3635,N_3289);
and U6263 (N_6263,N_4177,N_3663);
or U6264 (N_6264,N_4581,N_2648);
or U6265 (N_6265,N_4520,N_3357);
nand U6266 (N_6266,N_4774,N_4596);
nor U6267 (N_6267,N_3938,N_3754);
nand U6268 (N_6268,N_3501,N_4370);
or U6269 (N_6269,N_3519,N_3360);
xnor U6270 (N_6270,N_4519,N_4814);
or U6271 (N_6271,N_3917,N_3209);
and U6272 (N_6272,N_3001,N_3033);
xor U6273 (N_6273,N_2725,N_4365);
and U6274 (N_6274,N_2833,N_3006);
or U6275 (N_6275,N_3968,N_2598);
xor U6276 (N_6276,N_4173,N_4835);
or U6277 (N_6277,N_3799,N_3139);
nor U6278 (N_6278,N_3773,N_4347);
nand U6279 (N_6279,N_2783,N_3519);
or U6280 (N_6280,N_4022,N_2764);
or U6281 (N_6281,N_2758,N_4836);
and U6282 (N_6282,N_3910,N_4833);
xnor U6283 (N_6283,N_4677,N_4178);
and U6284 (N_6284,N_4419,N_2542);
or U6285 (N_6285,N_3632,N_2956);
xor U6286 (N_6286,N_4324,N_4526);
nor U6287 (N_6287,N_2641,N_3011);
xnor U6288 (N_6288,N_3221,N_3265);
or U6289 (N_6289,N_4674,N_4534);
nand U6290 (N_6290,N_3553,N_3614);
nand U6291 (N_6291,N_3710,N_3315);
nor U6292 (N_6292,N_3322,N_2711);
nand U6293 (N_6293,N_4588,N_4980);
or U6294 (N_6294,N_4880,N_3953);
nand U6295 (N_6295,N_3658,N_4188);
xor U6296 (N_6296,N_3156,N_3666);
xnor U6297 (N_6297,N_4892,N_3891);
and U6298 (N_6298,N_3248,N_4047);
nor U6299 (N_6299,N_4844,N_2946);
and U6300 (N_6300,N_3147,N_3027);
or U6301 (N_6301,N_4884,N_3098);
xnor U6302 (N_6302,N_4458,N_4335);
and U6303 (N_6303,N_4000,N_2932);
xnor U6304 (N_6304,N_4224,N_4877);
and U6305 (N_6305,N_4287,N_3386);
and U6306 (N_6306,N_3247,N_2689);
nand U6307 (N_6307,N_4141,N_3081);
nor U6308 (N_6308,N_2919,N_3262);
xnor U6309 (N_6309,N_4419,N_3737);
nor U6310 (N_6310,N_3550,N_4392);
and U6311 (N_6311,N_4739,N_4566);
nand U6312 (N_6312,N_4643,N_3155);
or U6313 (N_6313,N_4948,N_2856);
xnor U6314 (N_6314,N_3988,N_4785);
and U6315 (N_6315,N_4577,N_3892);
or U6316 (N_6316,N_3755,N_3488);
or U6317 (N_6317,N_3928,N_3961);
and U6318 (N_6318,N_3538,N_4353);
nand U6319 (N_6319,N_4310,N_3229);
or U6320 (N_6320,N_4490,N_4515);
and U6321 (N_6321,N_2501,N_2666);
and U6322 (N_6322,N_3095,N_3988);
nand U6323 (N_6323,N_3419,N_3130);
xnor U6324 (N_6324,N_3521,N_4351);
and U6325 (N_6325,N_4859,N_4429);
and U6326 (N_6326,N_4400,N_4240);
nor U6327 (N_6327,N_4648,N_4534);
or U6328 (N_6328,N_4628,N_4550);
xor U6329 (N_6329,N_4982,N_3340);
or U6330 (N_6330,N_2578,N_2918);
xnor U6331 (N_6331,N_3171,N_4634);
or U6332 (N_6332,N_4004,N_2691);
and U6333 (N_6333,N_4960,N_3282);
nand U6334 (N_6334,N_4755,N_3904);
xor U6335 (N_6335,N_2667,N_2878);
or U6336 (N_6336,N_4788,N_2792);
nand U6337 (N_6337,N_2853,N_4847);
and U6338 (N_6338,N_4020,N_4568);
xor U6339 (N_6339,N_4842,N_2525);
xor U6340 (N_6340,N_4747,N_3613);
xnor U6341 (N_6341,N_2787,N_3470);
or U6342 (N_6342,N_3591,N_3927);
or U6343 (N_6343,N_4099,N_3197);
and U6344 (N_6344,N_3643,N_3031);
or U6345 (N_6345,N_2875,N_4974);
nor U6346 (N_6346,N_2798,N_4765);
and U6347 (N_6347,N_3941,N_3427);
or U6348 (N_6348,N_3552,N_2864);
xor U6349 (N_6349,N_2993,N_3877);
nand U6350 (N_6350,N_3912,N_2505);
or U6351 (N_6351,N_3515,N_2554);
nor U6352 (N_6352,N_4262,N_3803);
nand U6353 (N_6353,N_4092,N_4208);
nand U6354 (N_6354,N_2516,N_3657);
xor U6355 (N_6355,N_3389,N_4724);
and U6356 (N_6356,N_2817,N_3890);
xor U6357 (N_6357,N_4969,N_2759);
or U6358 (N_6358,N_4102,N_4375);
or U6359 (N_6359,N_4054,N_2953);
xnor U6360 (N_6360,N_4377,N_2530);
nand U6361 (N_6361,N_3301,N_4471);
or U6362 (N_6362,N_3220,N_3813);
nand U6363 (N_6363,N_4062,N_3915);
and U6364 (N_6364,N_4860,N_3377);
nor U6365 (N_6365,N_3656,N_4788);
nand U6366 (N_6366,N_4166,N_4298);
and U6367 (N_6367,N_3229,N_3047);
or U6368 (N_6368,N_4866,N_4799);
xnor U6369 (N_6369,N_4566,N_3237);
xor U6370 (N_6370,N_3129,N_2612);
xor U6371 (N_6371,N_3014,N_4080);
nor U6372 (N_6372,N_3215,N_4444);
nand U6373 (N_6373,N_4426,N_4092);
or U6374 (N_6374,N_3279,N_3347);
or U6375 (N_6375,N_3889,N_4290);
xor U6376 (N_6376,N_4071,N_4097);
or U6377 (N_6377,N_3416,N_2558);
or U6378 (N_6378,N_3610,N_4419);
or U6379 (N_6379,N_4619,N_2733);
nand U6380 (N_6380,N_3160,N_3921);
nor U6381 (N_6381,N_2977,N_4606);
xnor U6382 (N_6382,N_4258,N_3055);
or U6383 (N_6383,N_3029,N_2532);
nor U6384 (N_6384,N_3185,N_4474);
or U6385 (N_6385,N_4971,N_3511);
or U6386 (N_6386,N_4748,N_3084);
xor U6387 (N_6387,N_3251,N_4610);
and U6388 (N_6388,N_4953,N_4924);
nand U6389 (N_6389,N_3360,N_4558);
nand U6390 (N_6390,N_4617,N_4781);
xnor U6391 (N_6391,N_4128,N_4842);
xnor U6392 (N_6392,N_3361,N_3649);
nor U6393 (N_6393,N_4095,N_2709);
nand U6394 (N_6394,N_2979,N_4609);
nor U6395 (N_6395,N_3829,N_4586);
or U6396 (N_6396,N_4765,N_4124);
nand U6397 (N_6397,N_2759,N_3481);
or U6398 (N_6398,N_3022,N_4245);
nor U6399 (N_6399,N_2696,N_4800);
nor U6400 (N_6400,N_4725,N_4654);
and U6401 (N_6401,N_4119,N_3548);
nor U6402 (N_6402,N_4512,N_3092);
nand U6403 (N_6403,N_3593,N_3667);
or U6404 (N_6404,N_3986,N_4243);
nand U6405 (N_6405,N_2817,N_4827);
xnor U6406 (N_6406,N_2889,N_4724);
xnor U6407 (N_6407,N_3438,N_3312);
nand U6408 (N_6408,N_3013,N_4776);
xnor U6409 (N_6409,N_4150,N_3794);
or U6410 (N_6410,N_2806,N_4853);
and U6411 (N_6411,N_4160,N_4384);
nand U6412 (N_6412,N_3191,N_2538);
xnor U6413 (N_6413,N_4667,N_3961);
nand U6414 (N_6414,N_4734,N_4749);
nand U6415 (N_6415,N_4491,N_3457);
nor U6416 (N_6416,N_4824,N_3197);
nand U6417 (N_6417,N_3555,N_2589);
nor U6418 (N_6418,N_4658,N_2818);
and U6419 (N_6419,N_2790,N_3968);
nor U6420 (N_6420,N_3873,N_4654);
xor U6421 (N_6421,N_2702,N_4784);
nor U6422 (N_6422,N_3404,N_4880);
xnor U6423 (N_6423,N_4113,N_3157);
nand U6424 (N_6424,N_3345,N_4726);
nor U6425 (N_6425,N_2773,N_4205);
xor U6426 (N_6426,N_2550,N_4248);
xor U6427 (N_6427,N_4122,N_4634);
nor U6428 (N_6428,N_3845,N_4301);
nor U6429 (N_6429,N_4808,N_4576);
or U6430 (N_6430,N_4144,N_2858);
or U6431 (N_6431,N_3942,N_3634);
xnor U6432 (N_6432,N_3075,N_4472);
nor U6433 (N_6433,N_4814,N_4340);
nor U6434 (N_6434,N_2727,N_3345);
or U6435 (N_6435,N_2791,N_4092);
nand U6436 (N_6436,N_2827,N_3642);
xor U6437 (N_6437,N_3279,N_3491);
or U6438 (N_6438,N_3527,N_4705);
nand U6439 (N_6439,N_4738,N_2910);
nor U6440 (N_6440,N_2954,N_3914);
and U6441 (N_6441,N_2607,N_3448);
nand U6442 (N_6442,N_2562,N_4605);
and U6443 (N_6443,N_2598,N_4757);
nand U6444 (N_6444,N_4102,N_2933);
or U6445 (N_6445,N_4354,N_4737);
nand U6446 (N_6446,N_3800,N_3290);
or U6447 (N_6447,N_2620,N_4634);
and U6448 (N_6448,N_4257,N_3044);
or U6449 (N_6449,N_2923,N_4048);
nor U6450 (N_6450,N_4979,N_4469);
and U6451 (N_6451,N_4464,N_3309);
xor U6452 (N_6452,N_3632,N_4855);
and U6453 (N_6453,N_3009,N_4143);
and U6454 (N_6454,N_4549,N_3383);
nand U6455 (N_6455,N_4752,N_3825);
xnor U6456 (N_6456,N_4595,N_4153);
or U6457 (N_6457,N_3313,N_4591);
nand U6458 (N_6458,N_2589,N_4792);
or U6459 (N_6459,N_4782,N_3807);
xor U6460 (N_6460,N_4074,N_2794);
xnor U6461 (N_6461,N_4582,N_3260);
or U6462 (N_6462,N_3250,N_3949);
or U6463 (N_6463,N_2931,N_3312);
xnor U6464 (N_6464,N_4718,N_3561);
and U6465 (N_6465,N_4593,N_4442);
xnor U6466 (N_6466,N_4481,N_3679);
nand U6467 (N_6467,N_4944,N_3150);
nand U6468 (N_6468,N_3835,N_2664);
or U6469 (N_6469,N_3871,N_2595);
nand U6470 (N_6470,N_2963,N_4917);
nor U6471 (N_6471,N_4877,N_4957);
nor U6472 (N_6472,N_4313,N_3984);
xor U6473 (N_6473,N_3998,N_4561);
or U6474 (N_6474,N_3256,N_3349);
and U6475 (N_6475,N_3741,N_3516);
and U6476 (N_6476,N_4768,N_4618);
or U6477 (N_6477,N_4721,N_3817);
nand U6478 (N_6478,N_3851,N_2884);
xor U6479 (N_6479,N_3933,N_2591);
nor U6480 (N_6480,N_4725,N_4598);
and U6481 (N_6481,N_4721,N_3087);
xnor U6482 (N_6482,N_4759,N_3922);
xor U6483 (N_6483,N_4229,N_3150);
xor U6484 (N_6484,N_3998,N_4806);
or U6485 (N_6485,N_2963,N_3026);
nor U6486 (N_6486,N_4992,N_4427);
xnor U6487 (N_6487,N_2875,N_2981);
nand U6488 (N_6488,N_2968,N_4119);
and U6489 (N_6489,N_2648,N_4378);
xnor U6490 (N_6490,N_4694,N_4804);
nand U6491 (N_6491,N_2741,N_3191);
or U6492 (N_6492,N_3556,N_2829);
xor U6493 (N_6493,N_3153,N_4218);
nor U6494 (N_6494,N_3397,N_3128);
nor U6495 (N_6495,N_3722,N_2968);
nand U6496 (N_6496,N_2923,N_3645);
nor U6497 (N_6497,N_3984,N_4229);
and U6498 (N_6498,N_3046,N_3389);
nand U6499 (N_6499,N_4149,N_4135);
nor U6500 (N_6500,N_2710,N_3594);
and U6501 (N_6501,N_4550,N_3665);
nand U6502 (N_6502,N_3635,N_4708);
or U6503 (N_6503,N_3874,N_4322);
and U6504 (N_6504,N_4440,N_4580);
nand U6505 (N_6505,N_4546,N_4173);
nand U6506 (N_6506,N_4727,N_4068);
nand U6507 (N_6507,N_4232,N_3582);
or U6508 (N_6508,N_4494,N_2589);
and U6509 (N_6509,N_4423,N_2748);
or U6510 (N_6510,N_3337,N_2641);
and U6511 (N_6511,N_4262,N_3045);
or U6512 (N_6512,N_2875,N_4277);
xnor U6513 (N_6513,N_4473,N_4623);
xor U6514 (N_6514,N_2829,N_3171);
nand U6515 (N_6515,N_4854,N_4948);
nor U6516 (N_6516,N_3904,N_3099);
or U6517 (N_6517,N_4866,N_2639);
nand U6518 (N_6518,N_4138,N_4093);
and U6519 (N_6519,N_4446,N_4088);
or U6520 (N_6520,N_2617,N_3039);
nand U6521 (N_6521,N_4247,N_4364);
nand U6522 (N_6522,N_4368,N_2810);
nor U6523 (N_6523,N_3686,N_3085);
and U6524 (N_6524,N_4693,N_3152);
and U6525 (N_6525,N_3968,N_4078);
nand U6526 (N_6526,N_2886,N_3045);
xnor U6527 (N_6527,N_4778,N_2975);
nor U6528 (N_6528,N_3111,N_3074);
nor U6529 (N_6529,N_4158,N_4887);
xor U6530 (N_6530,N_4596,N_4530);
xor U6531 (N_6531,N_4455,N_4974);
xnor U6532 (N_6532,N_4397,N_3523);
nand U6533 (N_6533,N_3101,N_3708);
nor U6534 (N_6534,N_2735,N_2977);
or U6535 (N_6535,N_4346,N_3578);
nand U6536 (N_6536,N_3000,N_2652);
or U6537 (N_6537,N_3623,N_4579);
xnor U6538 (N_6538,N_2567,N_4129);
and U6539 (N_6539,N_4733,N_3981);
and U6540 (N_6540,N_3406,N_4912);
nand U6541 (N_6541,N_4823,N_2926);
or U6542 (N_6542,N_3649,N_4570);
nand U6543 (N_6543,N_4470,N_3325);
and U6544 (N_6544,N_4995,N_3910);
xnor U6545 (N_6545,N_2975,N_2951);
nor U6546 (N_6546,N_3797,N_4014);
and U6547 (N_6547,N_4271,N_4470);
and U6548 (N_6548,N_2641,N_4570);
xor U6549 (N_6549,N_4723,N_3790);
or U6550 (N_6550,N_4760,N_2715);
xnor U6551 (N_6551,N_4252,N_4213);
nor U6552 (N_6552,N_2682,N_3432);
nand U6553 (N_6553,N_4378,N_2960);
nor U6554 (N_6554,N_3564,N_4575);
nand U6555 (N_6555,N_4145,N_3261);
nand U6556 (N_6556,N_4020,N_4569);
xor U6557 (N_6557,N_4838,N_4489);
xor U6558 (N_6558,N_3178,N_4818);
or U6559 (N_6559,N_4405,N_3896);
xor U6560 (N_6560,N_4638,N_2745);
nand U6561 (N_6561,N_3608,N_2928);
xor U6562 (N_6562,N_3637,N_4633);
nor U6563 (N_6563,N_4017,N_3921);
xnor U6564 (N_6564,N_2652,N_3945);
nand U6565 (N_6565,N_4194,N_4297);
and U6566 (N_6566,N_3281,N_4630);
nor U6567 (N_6567,N_3388,N_2680);
nor U6568 (N_6568,N_3407,N_4648);
or U6569 (N_6569,N_3889,N_2699);
nor U6570 (N_6570,N_2866,N_2575);
nand U6571 (N_6571,N_3558,N_4114);
xnor U6572 (N_6572,N_4666,N_2810);
or U6573 (N_6573,N_2744,N_3183);
or U6574 (N_6574,N_4558,N_2648);
xnor U6575 (N_6575,N_3966,N_4297);
nor U6576 (N_6576,N_4552,N_4768);
nand U6577 (N_6577,N_2770,N_3013);
xnor U6578 (N_6578,N_3603,N_4718);
or U6579 (N_6579,N_3947,N_4171);
or U6580 (N_6580,N_3418,N_3395);
nor U6581 (N_6581,N_3303,N_2816);
xnor U6582 (N_6582,N_4069,N_3097);
nand U6583 (N_6583,N_3312,N_3192);
and U6584 (N_6584,N_3932,N_3953);
xnor U6585 (N_6585,N_4106,N_4795);
or U6586 (N_6586,N_3302,N_3576);
xor U6587 (N_6587,N_4652,N_4163);
and U6588 (N_6588,N_3392,N_3554);
xnor U6589 (N_6589,N_4960,N_4283);
or U6590 (N_6590,N_3702,N_3249);
and U6591 (N_6591,N_4235,N_2985);
nand U6592 (N_6592,N_2529,N_2771);
nand U6593 (N_6593,N_4888,N_4867);
xnor U6594 (N_6594,N_4356,N_3226);
nor U6595 (N_6595,N_4969,N_3352);
nand U6596 (N_6596,N_3279,N_2720);
and U6597 (N_6597,N_4321,N_4682);
nor U6598 (N_6598,N_3809,N_2564);
nor U6599 (N_6599,N_3298,N_4077);
xnor U6600 (N_6600,N_2874,N_2519);
nor U6601 (N_6601,N_3380,N_4157);
nand U6602 (N_6602,N_2697,N_2792);
nand U6603 (N_6603,N_2628,N_2587);
xor U6604 (N_6604,N_4784,N_2670);
nand U6605 (N_6605,N_3189,N_4296);
nand U6606 (N_6606,N_2579,N_4183);
nor U6607 (N_6607,N_2936,N_4388);
and U6608 (N_6608,N_4867,N_4157);
and U6609 (N_6609,N_2839,N_4751);
or U6610 (N_6610,N_4162,N_3181);
nand U6611 (N_6611,N_2615,N_4693);
and U6612 (N_6612,N_4232,N_4530);
or U6613 (N_6613,N_4834,N_2512);
or U6614 (N_6614,N_4712,N_2954);
or U6615 (N_6615,N_3115,N_2618);
and U6616 (N_6616,N_3643,N_4387);
nand U6617 (N_6617,N_4737,N_4771);
nand U6618 (N_6618,N_4722,N_4109);
xor U6619 (N_6619,N_4309,N_2988);
nor U6620 (N_6620,N_2931,N_2730);
nand U6621 (N_6621,N_4647,N_3393);
xnor U6622 (N_6622,N_4204,N_4620);
or U6623 (N_6623,N_3438,N_3590);
and U6624 (N_6624,N_4205,N_3106);
nand U6625 (N_6625,N_4063,N_2668);
nor U6626 (N_6626,N_2587,N_3785);
and U6627 (N_6627,N_2828,N_4074);
or U6628 (N_6628,N_4264,N_3432);
xor U6629 (N_6629,N_4733,N_3698);
nor U6630 (N_6630,N_3408,N_4648);
and U6631 (N_6631,N_2782,N_4426);
nand U6632 (N_6632,N_4092,N_4704);
or U6633 (N_6633,N_3547,N_2586);
or U6634 (N_6634,N_3088,N_4421);
nand U6635 (N_6635,N_4780,N_4178);
nor U6636 (N_6636,N_3376,N_4149);
and U6637 (N_6637,N_4015,N_3057);
xnor U6638 (N_6638,N_2727,N_4681);
nor U6639 (N_6639,N_3087,N_3853);
nand U6640 (N_6640,N_4937,N_4268);
nand U6641 (N_6641,N_3876,N_2512);
nand U6642 (N_6642,N_3620,N_2999);
nor U6643 (N_6643,N_3527,N_4750);
or U6644 (N_6644,N_2658,N_4712);
nand U6645 (N_6645,N_4613,N_3924);
and U6646 (N_6646,N_3627,N_2728);
or U6647 (N_6647,N_2707,N_4416);
and U6648 (N_6648,N_2935,N_4515);
nand U6649 (N_6649,N_4820,N_2714);
or U6650 (N_6650,N_3372,N_3258);
nor U6651 (N_6651,N_4957,N_4624);
or U6652 (N_6652,N_3562,N_4209);
nor U6653 (N_6653,N_4733,N_2832);
and U6654 (N_6654,N_2520,N_3791);
or U6655 (N_6655,N_2626,N_2818);
nand U6656 (N_6656,N_2754,N_2644);
and U6657 (N_6657,N_3800,N_2703);
and U6658 (N_6658,N_3511,N_4968);
or U6659 (N_6659,N_4471,N_4130);
nor U6660 (N_6660,N_4025,N_3556);
or U6661 (N_6661,N_3556,N_3266);
and U6662 (N_6662,N_3434,N_3241);
nand U6663 (N_6663,N_4271,N_3605);
xnor U6664 (N_6664,N_2906,N_4102);
nand U6665 (N_6665,N_3026,N_2520);
xnor U6666 (N_6666,N_3863,N_3438);
and U6667 (N_6667,N_3600,N_4127);
and U6668 (N_6668,N_3757,N_4630);
or U6669 (N_6669,N_2533,N_4709);
nand U6670 (N_6670,N_4579,N_3009);
and U6671 (N_6671,N_2900,N_4368);
nand U6672 (N_6672,N_4703,N_4399);
nor U6673 (N_6673,N_2700,N_2569);
nor U6674 (N_6674,N_3092,N_2964);
xor U6675 (N_6675,N_4486,N_3392);
nand U6676 (N_6676,N_4670,N_3803);
xnor U6677 (N_6677,N_4111,N_4093);
and U6678 (N_6678,N_3406,N_4085);
or U6679 (N_6679,N_4765,N_3043);
or U6680 (N_6680,N_3818,N_3091);
nand U6681 (N_6681,N_3628,N_3586);
and U6682 (N_6682,N_2865,N_2534);
and U6683 (N_6683,N_3468,N_4394);
and U6684 (N_6684,N_4130,N_4038);
nor U6685 (N_6685,N_2935,N_3048);
xor U6686 (N_6686,N_3773,N_3091);
nand U6687 (N_6687,N_3711,N_3562);
nor U6688 (N_6688,N_3264,N_4175);
nand U6689 (N_6689,N_3832,N_2937);
nand U6690 (N_6690,N_3543,N_3233);
nand U6691 (N_6691,N_2936,N_4501);
nor U6692 (N_6692,N_3497,N_3057);
and U6693 (N_6693,N_4468,N_4397);
and U6694 (N_6694,N_3435,N_3587);
and U6695 (N_6695,N_4866,N_3980);
nand U6696 (N_6696,N_2698,N_3492);
and U6697 (N_6697,N_4647,N_3670);
nor U6698 (N_6698,N_3519,N_3514);
and U6699 (N_6699,N_3277,N_3045);
nand U6700 (N_6700,N_4369,N_4521);
or U6701 (N_6701,N_4498,N_2936);
or U6702 (N_6702,N_3601,N_2549);
xor U6703 (N_6703,N_4500,N_4104);
xnor U6704 (N_6704,N_2995,N_2553);
xnor U6705 (N_6705,N_4035,N_2705);
nor U6706 (N_6706,N_3227,N_2601);
nand U6707 (N_6707,N_4804,N_3489);
or U6708 (N_6708,N_4098,N_3966);
xnor U6709 (N_6709,N_3912,N_3113);
xnor U6710 (N_6710,N_4879,N_2875);
or U6711 (N_6711,N_4396,N_2709);
nor U6712 (N_6712,N_4480,N_4157);
nand U6713 (N_6713,N_4149,N_3467);
or U6714 (N_6714,N_4529,N_3353);
nand U6715 (N_6715,N_3961,N_4499);
xor U6716 (N_6716,N_4374,N_2523);
nor U6717 (N_6717,N_4471,N_2985);
nor U6718 (N_6718,N_4390,N_3870);
nand U6719 (N_6719,N_4144,N_4267);
nand U6720 (N_6720,N_2600,N_2772);
nor U6721 (N_6721,N_3141,N_4579);
nand U6722 (N_6722,N_2735,N_4882);
or U6723 (N_6723,N_2525,N_3791);
and U6724 (N_6724,N_4791,N_3324);
nand U6725 (N_6725,N_2834,N_2912);
xor U6726 (N_6726,N_3148,N_4573);
xnor U6727 (N_6727,N_3804,N_4236);
nor U6728 (N_6728,N_2685,N_2578);
or U6729 (N_6729,N_4183,N_2702);
xnor U6730 (N_6730,N_3984,N_2723);
and U6731 (N_6731,N_2558,N_4473);
and U6732 (N_6732,N_4822,N_4761);
xor U6733 (N_6733,N_4056,N_2695);
or U6734 (N_6734,N_3911,N_2609);
xnor U6735 (N_6735,N_2610,N_4743);
and U6736 (N_6736,N_2655,N_2951);
xnor U6737 (N_6737,N_3084,N_3332);
nand U6738 (N_6738,N_3514,N_2967);
and U6739 (N_6739,N_3411,N_4898);
or U6740 (N_6740,N_3884,N_3692);
or U6741 (N_6741,N_2676,N_3678);
xnor U6742 (N_6742,N_4754,N_4788);
nand U6743 (N_6743,N_3892,N_2500);
nor U6744 (N_6744,N_3189,N_3179);
and U6745 (N_6745,N_4324,N_3648);
nor U6746 (N_6746,N_4440,N_3446);
or U6747 (N_6747,N_3465,N_4404);
and U6748 (N_6748,N_4132,N_2987);
xor U6749 (N_6749,N_4246,N_4016);
xnor U6750 (N_6750,N_4085,N_4551);
nor U6751 (N_6751,N_4483,N_3456);
nand U6752 (N_6752,N_2629,N_4270);
or U6753 (N_6753,N_4531,N_4945);
xor U6754 (N_6754,N_3983,N_3118);
nand U6755 (N_6755,N_4900,N_2642);
nor U6756 (N_6756,N_3703,N_2888);
nand U6757 (N_6757,N_3846,N_2663);
or U6758 (N_6758,N_3484,N_4845);
and U6759 (N_6759,N_3212,N_4832);
nor U6760 (N_6760,N_4687,N_3969);
xnor U6761 (N_6761,N_3018,N_2608);
xnor U6762 (N_6762,N_3673,N_2691);
nand U6763 (N_6763,N_3762,N_4327);
or U6764 (N_6764,N_2557,N_3167);
nor U6765 (N_6765,N_4059,N_3168);
nor U6766 (N_6766,N_2791,N_2822);
or U6767 (N_6767,N_4140,N_4011);
nor U6768 (N_6768,N_4983,N_3565);
xnor U6769 (N_6769,N_4933,N_4227);
nand U6770 (N_6770,N_2541,N_2910);
or U6771 (N_6771,N_3804,N_2832);
and U6772 (N_6772,N_3173,N_3354);
or U6773 (N_6773,N_3424,N_3188);
nor U6774 (N_6774,N_4305,N_3278);
or U6775 (N_6775,N_2858,N_3646);
or U6776 (N_6776,N_3396,N_3457);
or U6777 (N_6777,N_4260,N_3243);
nand U6778 (N_6778,N_3741,N_4591);
nor U6779 (N_6779,N_3574,N_3300);
xor U6780 (N_6780,N_4059,N_2580);
and U6781 (N_6781,N_3539,N_3165);
or U6782 (N_6782,N_4697,N_3097);
xor U6783 (N_6783,N_4761,N_3190);
xor U6784 (N_6784,N_3395,N_3639);
and U6785 (N_6785,N_2785,N_3239);
nand U6786 (N_6786,N_2849,N_4325);
and U6787 (N_6787,N_3709,N_3058);
and U6788 (N_6788,N_2519,N_3038);
or U6789 (N_6789,N_3551,N_4045);
nor U6790 (N_6790,N_3653,N_3219);
or U6791 (N_6791,N_4060,N_3705);
nand U6792 (N_6792,N_3183,N_3275);
xor U6793 (N_6793,N_4884,N_4352);
and U6794 (N_6794,N_3461,N_2869);
nor U6795 (N_6795,N_2599,N_4286);
or U6796 (N_6796,N_4334,N_2683);
nor U6797 (N_6797,N_2895,N_3906);
or U6798 (N_6798,N_4613,N_4369);
or U6799 (N_6799,N_3111,N_2723);
xor U6800 (N_6800,N_4351,N_3462);
or U6801 (N_6801,N_2904,N_3901);
nor U6802 (N_6802,N_3460,N_3148);
xnor U6803 (N_6803,N_4685,N_4186);
xnor U6804 (N_6804,N_4382,N_2701);
or U6805 (N_6805,N_3108,N_3051);
nor U6806 (N_6806,N_3109,N_4743);
nand U6807 (N_6807,N_3758,N_4751);
and U6808 (N_6808,N_4678,N_3561);
xor U6809 (N_6809,N_3592,N_4268);
and U6810 (N_6810,N_4474,N_4367);
or U6811 (N_6811,N_3256,N_4130);
xnor U6812 (N_6812,N_2546,N_3599);
xor U6813 (N_6813,N_3094,N_3689);
nand U6814 (N_6814,N_2628,N_3327);
and U6815 (N_6815,N_4250,N_3949);
or U6816 (N_6816,N_4942,N_3507);
nor U6817 (N_6817,N_4035,N_4881);
nand U6818 (N_6818,N_2807,N_2646);
or U6819 (N_6819,N_4330,N_4510);
and U6820 (N_6820,N_2946,N_3106);
or U6821 (N_6821,N_2809,N_4575);
xor U6822 (N_6822,N_4715,N_4104);
nor U6823 (N_6823,N_3671,N_2979);
nand U6824 (N_6824,N_4887,N_4807);
or U6825 (N_6825,N_4348,N_3129);
xnor U6826 (N_6826,N_4476,N_3212);
xor U6827 (N_6827,N_3567,N_4963);
xnor U6828 (N_6828,N_3343,N_2706);
and U6829 (N_6829,N_3505,N_2532);
or U6830 (N_6830,N_2978,N_4316);
nand U6831 (N_6831,N_3706,N_3021);
nand U6832 (N_6832,N_2659,N_4373);
or U6833 (N_6833,N_3266,N_3936);
nor U6834 (N_6834,N_4995,N_4640);
nand U6835 (N_6835,N_3766,N_2748);
nand U6836 (N_6836,N_4395,N_3718);
nand U6837 (N_6837,N_3367,N_2644);
or U6838 (N_6838,N_4890,N_3641);
nand U6839 (N_6839,N_4366,N_3595);
nor U6840 (N_6840,N_4567,N_3872);
nand U6841 (N_6841,N_3329,N_2539);
nand U6842 (N_6842,N_3223,N_4125);
and U6843 (N_6843,N_4051,N_4103);
xnor U6844 (N_6844,N_3470,N_3545);
nand U6845 (N_6845,N_3843,N_3753);
nor U6846 (N_6846,N_4255,N_2535);
xor U6847 (N_6847,N_2817,N_2732);
nand U6848 (N_6848,N_2731,N_4791);
nor U6849 (N_6849,N_3517,N_2989);
and U6850 (N_6850,N_2733,N_3112);
or U6851 (N_6851,N_4016,N_4153);
nand U6852 (N_6852,N_2996,N_4975);
nand U6853 (N_6853,N_3018,N_2917);
or U6854 (N_6854,N_3747,N_2929);
or U6855 (N_6855,N_2905,N_2566);
nor U6856 (N_6856,N_4147,N_4912);
or U6857 (N_6857,N_4659,N_4580);
nand U6858 (N_6858,N_4517,N_2623);
nand U6859 (N_6859,N_4728,N_2619);
or U6860 (N_6860,N_2976,N_3571);
and U6861 (N_6861,N_3888,N_4976);
nand U6862 (N_6862,N_3732,N_4024);
nor U6863 (N_6863,N_4042,N_3962);
xnor U6864 (N_6864,N_3987,N_4350);
nor U6865 (N_6865,N_2704,N_4045);
or U6866 (N_6866,N_3673,N_3314);
nor U6867 (N_6867,N_2946,N_3484);
xnor U6868 (N_6868,N_3123,N_2761);
and U6869 (N_6869,N_4195,N_2559);
nand U6870 (N_6870,N_3775,N_2942);
nor U6871 (N_6871,N_4293,N_2948);
nand U6872 (N_6872,N_3478,N_2932);
and U6873 (N_6873,N_2840,N_4033);
nand U6874 (N_6874,N_4341,N_2626);
or U6875 (N_6875,N_4410,N_4223);
and U6876 (N_6876,N_3988,N_3324);
nand U6877 (N_6877,N_3099,N_3511);
nor U6878 (N_6878,N_3985,N_2976);
xor U6879 (N_6879,N_2633,N_4070);
xor U6880 (N_6880,N_3007,N_3866);
nor U6881 (N_6881,N_4136,N_4993);
xor U6882 (N_6882,N_3786,N_3986);
nand U6883 (N_6883,N_2757,N_3878);
nand U6884 (N_6884,N_3106,N_3673);
and U6885 (N_6885,N_3695,N_3970);
xnor U6886 (N_6886,N_2803,N_4138);
xor U6887 (N_6887,N_3526,N_3711);
and U6888 (N_6888,N_4090,N_4256);
nor U6889 (N_6889,N_4461,N_3913);
xor U6890 (N_6890,N_3770,N_2953);
or U6891 (N_6891,N_3760,N_2554);
or U6892 (N_6892,N_2953,N_3569);
xnor U6893 (N_6893,N_3376,N_4814);
and U6894 (N_6894,N_3817,N_3856);
xor U6895 (N_6895,N_4989,N_3211);
or U6896 (N_6896,N_2990,N_3243);
and U6897 (N_6897,N_4531,N_3090);
nor U6898 (N_6898,N_3644,N_4886);
xnor U6899 (N_6899,N_2889,N_2902);
nor U6900 (N_6900,N_2866,N_3438);
nand U6901 (N_6901,N_2900,N_4173);
nand U6902 (N_6902,N_3387,N_4044);
xor U6903 (N_6903,N_4160,N_3004);
or U6904 (N_6904,N_3201,N_4037);
or U6905 (N_6905,N_2812,N_4354);
or U6906 (N_6906,N_4075,N_3238);
or U6907 (N_6907,N_4874,N_4906);
or U6908 (N_6908,N_4790,N_3402);
nor U6909 (N_6909,N_2914,N_4233);
nor U6910 (N_6910,N_3970,N_4834);
nor U6911 (N_6911,N_4310,N_3024);
nor U6912 (N_6912,N_4790,N_3520);
or U6913 (N_6913,N_4399,N_4535);
nand U6914 (N_6914,N_4508,N_4372);
xnor U6915 (N_6915,N_4697,N_4195);
nand U6916 (N_6916,N_4320,N_4323);
nand U6917 (N_6917,N_3076,N_2718);
nand U6918 (N_6918,N_4844,N_4166);
or U6919 (N_6919,N_3515,N_3788);
or U6920 (N_6920,N_2702,N_3843);
xor U6921 (N_6921,N_3766,N_3460);
nand U6922 (N_6922,N_3084,N_3499);
nor U6923 (N_6923,N_4978,N_3800);
xnor U6924 (N_6924,N_4452,N_4928);
nor U6925 (N_6925,N_3210,N_4578);
xnor U6926 (N_6926,N_3218,N_3986);
or U6927 (N_6927,N_4829,N_2888);
and U6928 (N_6928,N_4625,N_2855);
xor U6929 (N_6929,N_3462,N_3600);
nand U6930 (N_6930,N_4222,N_3368);
nand U6931 (N_6931,N_3696,N_2860);
nor U6932 (N_6932,N_3384,N_4197);
nor U6933 (N_6933,N_3507,N_3164);
and U6934 (N_6934,N_3620,N_4097);
and U6935 (N_6935,N_2718,N_3336);
and U6936 (N_6936,N_4926,N_4111);
nor U6937 (N_6937,N_2572,N_3248);
xor U6938 (N_6938,N_4687,N_4534);
or U6939 (N_6939,N_2529,N_3407);
xnor U6940 (N_6940,N_3733,N_4319);
or U6941 (N_6941,N_4006,N_3396);
nor U6942 (N_6942,N_3702,N_2531);
nor U6943 (N_6943,N_4577,N_3092);
or U6944 (N_6944,N_3258,N_2652);
nand U6945 (N_6945,N_4133,N_4511);
and U6946 (N_6946,N_3752,N_3130);
nor U6947 (N_6947,N_4325,N_4310);
and U6948 (N_6948,N_2745,N_4092);
or U6949 (N_6949,N_4377,N_3182);
or U6950 (N_6950,N_2643,N_2838);
nor U6951 (N_6951,N_3529,N_4929);
nand U6952 (N_6952,N_3824,N_3977);
xor U6953 (N_6953,N_3698,N_3560);
and U6954 (N_6954,N_4842,N_3671);
nand U6955 (N_6955,N_4450,N_3544);
xnor U6956 (N_6956,N_3910,N_3599);
nor U6957 (N_6957,N_3191,N_4721);
nand U6958 (N_6958,N_2827,N_4951);
nor U6959 (N_6959,N_4178,N_3867);
nor U6960 (N_6960,N_3661,N_4180);
nand U6961 (N_6961,N_2948,N_2755);
or U6962 (N_6962,N_3851,N_4876);
nand U6963 (N_6963,N_4511,N_2521);
nor U6964 (N_6964,N_2571,N_2985);
and U6965 (N_6965,N_4547,N_3089);
or U6966 (N_6966,N_3234,N_3423);
nor U6967 (N_6967,N_2981,N_3140);
or U6968 (N_6968,N_3803,N_4460);
or U6969 (N_6969,N_4709,N_2642);
xnor U6970 (N_6970,N_3416,N_4681);
or U6971 (N_6971,N_4582,N_4471);
nand U6972 (N_6972,N_4531,N_4330);
nand U6973 (N_6973,N_3503,N_2609);
xor U6974 (N_6974,N_4607,N_4442);
nor U6975 (N_6975,N_3540,N_3857);
or U6976 (N_6976,N_4417,N_4006);
or U6977 (N_6977,N_2727,N_3748);
or U6978 (N_6978,N_3684,N_4724);
nand U6979 (N_6979,N_4277,N_4969);
xor U6980 (N_6980,N_4373,N_3069);
xor U6981 (N_6981,N_3387,N_3544);
xor U6982 (N_6982,N_3213,N_4412);
nor U6983 (N_6983,N_4293,N_4484);
or U6984 (N_6984,N_3384,N_2577);
and U6985 (N_6985,N_2748,N_4546);
or U6986 (N_6986,N_4412,N_4857);
nor U6987 (N_6987,N_3383,N_3013);
xor U6988 (N_6988,N_4077,N_4164);
nor U6989 (N_6989,N_4543,N_3887);
and U6990 (N_6990,N_3878,N_2739);
or U6991 (N_6991,N_3215,N_3727);
or U6992 (N_6992,N_4158,N_3117);
xnor U6993 (N_6993,N_4367,N_3295);
and U6994 (N_6994,N_3634,N_2611);
xor U6995 (N_6995,N_3508,N_2725);
nor U6996 (N_6996,N_4735,N_4361);
xor U6997 (N_6997,N_4839,N_3341);
or U6998 (N_6998,N_3670,N_2666);
xnor U6999 (N_6999,N_4012,N_4682);
and U7000 (N_7000,N_3258,N_3621);
and U7001 (N_7001,N_3775,N_4848);
nand U7002 (N_7002,N_3206,N_3074);
and U7003 (N_7003,N_2703,N_4671);
nor U7004 (N_7004,N_2664,N_3277);
and U7005 (N_7005,N_4838,N_4165);
or U7006 (N_7006,N_4503,N_4447);
or U7007 (N_7007,N_2960,N_3389);
or U7008 (N_7008,N_3810,N_3934);
and U7009 (N_7009,N_4162,N_4786);
nor U7010 (N_7010,N_2729,N_3080);
or U7011 (N_7011,N_4203,N_3548);
or U7012 (N_7012,N_4041,N_3099);
nand U7013 (N_7013,N_4112,N_4453);
or U7014 (N_7014,N_2828,N_2574);
and U7015 (N_7015,N_3748,N_2654);
and U7016 (N_7016,N_4282,N_4319);
or U7017 (N_7017,N_4064,N_4683);
or U7018 (N_7018,N_2857,N_3243);
nor U7019 (N_7019,N_2784,N_4313);
nand U7020 (N_7020,N_4473,N_4021);
or U7021 (N_7021,N_2665,N_4028);
nor U7022 (N_7022,N_4844,N_4201);
and U7023 (N_7023,N_2935,N_2517);
nor U7024 (N_7024,N_3135,N_4592);
and U7025 (N_7025,N_2672,N_3219);
xor U7026 (N_7026,N_4392,N_3758);
xor U7027 (N_7027,N_4353,N_4790);
and U7028 (N_7028,N_4193,N_3569);
or U7029 (N_7029,N_3935,N_3190);
nand U7030 (N_7030,N_3841,N_2984);
xor U7031 (N_7031,N_4389,N_3917);
or U7032 (N_7032,N_4898,N_4817);
and U7033 (N_7033,N_4247,N_4892);
nand U7034 (N_7034,N_3720,N_4925);
nand U7035 (N_7035,N_3913,N_4185);
or U7036 (N_7036,N_2945,N_4025);
or U7037 (N_7037,N_4372,N_4515);
or U7038 (N_7038,N_3313,N_4956);
nand U7039 (N_7039,N_4624,N_3837);
nand U7040 (N_7040,N_4649,N_3466);
xnor U7041 (N_7041,N_4996,N_4891);
or U7042 (N_7042,N_2717,N_4258);
nor U7043 (N_7043,N_3308,N_3968);
nand U7044 (N_7044,N_4771,N_4024);
nand U7045 (N_7045,N_2553,N_4483);
xnor U7046 (N_7046,N_3305,N_4594);
nor U7047 (N_7047,N_3245,N_2798);
nand U7048 (N_7048,N_3598,N_4426);
nand U7049 (N_7049,N_4414,N_4593);
xnor U7050 (N_7050,N_3758,N_2990);
or U7051 (N_7051,N_2828,N_2723);
nor U7052 (N_7052,N_2629,N_4203);
xor U7053 (N_7053,N_2804,N_3930);
nor U7054 (N_7054,N_3952,N_4834);
or U7055 (N_7055,N_4268,N_2623);
nand U7056 (N_7056,N_2507,N_3662);
nand U7057 (N_7057,N_4085,N_2792);
and U7058 (N_7058,N_3762,N_4613);
or U7059 (N_7059,N_4481,N_3462);
and U7060 (N_7060,N_2693,N_4677);
nor U7061 (N_7061,N_4321,N_2739);
nand U7062 (N_7062,N_4776,N_3602);
nand U7063 (N_7063,N_2928,N_3053);
nor U7064 (N_7064,N_3162,N_3201);
and U7065 (N_7065,N_4397,N_2909);
or U7066 (N_7066,N_2551,N_3437);
nand U7067 (N_7067,N_2580,N_3880);
nand U7068 (N_7068,N_3325,N_4506);
nor U7069 (N_7069,N_2755,N_4224);
and U7070 (N_7070,N_3289,N_2926);
xnor U7071 (N_7071,N_3787,N_3885);
and U7072 (N_7072,N_4793,N_4295);
nand U7073 (N_7073,N_2975,N_4217);
nand U7074 (N_7074,N_3336,N_4352);
nand U7075 (N_7075,N_3995,N_2642);
or U7076 (N_7076,N_3071,N_3922);
nor U7077 (N_7077,N_2796,N_3726);
nand U7078 (N_7078,N_3131,N_3245);
xor U7079 (N_7079,N_4751,N_3096);
xor U7080 (N_7080,N_3368,N_4883);
and U7081 (N_7081,N_2610,N_4265);
nand U7082 (N_7082,N_4460,N_3067);
nand U7083 (N_7083,N_3196,N_3019);
and U7084 (N_7084,N_4897,N_3919);
and U7085 (N_7085,N_3329,N_4557);
or U7086 (N_7086,N_4092,N_4231);
nand U7087 (N_7087,N_3643,N_4570);
or U7088 (N_7088,N_2559,N_3200);
or U7089 (N_7089,N_2997,N_3030);
nor U7090 (N_7090,N_4113,N_4675);
and U7091 (N_7091,N_2511,N_4929);
or U7092 (N_7092,N_3173,N_3943);
xor U7093 (N_7093,N_4423,N_2943);
nand U7094 (N_7094,N_2868,N_3053);
nand U7095 (N_7095,N_4622,N_4823);
xnor U7096 (N_7096,N_2926,N_4209);
xor U7097 (N_7097,N_2502,N_3637);
and U7098 (N_7098,N_4265,N_4960);
nor U7099 (N_7099,N_3258,N_3800);
and U7100 (N_7100,N_4572,N_2568);
and U7101 (N_7101,N_4282,N_2943);
and U7102 (N_7102,N_4299,N_3200);
and U7103 (N_7103,N_2527,N_4374);
nand U7104 (N_7104,N_4593,N_3476);
nand U7105 (N_7105,N_3223,N_3709);
nor U7106 (N_7106,N_3741,N_3961);
or U7107 (N_7107,N_3317,N_3275);
or U7108 (N_7108,N_4246,N_3896);
or U7109 (N_7109,N_3425,N_4145);
xnor U7110 (N_7110,N_3556,N_4235);
and U7111 (N_7111,N_4554,N_4460);
nor U7112 (N_7112,N_3550,N_4990);
xor U7113 (N_7113,N_4960,N_4143);
nand U7114 (N_7114,N_4873,N_4498);
xnor U7115 (N_7115,N_2565,N_2518);
xor U7116 (N_7116,N_3649,N_2758);
nor U7117 (N_7117,N_3889,N_4183);
and U7118 (N_7118,N_4523,N_3275);
and U7119 (N_7119,N_4799,N_3948);
nand U7120 (N_7120,N_4320,N_4613);
nand U7121 (N_7121,N_4716,N_4133);
nand U7122 (N_7122,N_3335,N_2612);
or U7123 (N_7123,N_3011,N_4764);
nor U7124 (N_7124,N_2922,N_2967);
or U7125 (N_7125,N_2979,N_3809);
nor U7126 (N_7126,N_2660,N_3929);
nor U7127 (N_7127,N_2915,N_3514);
xnor U7128 (N_7128,N_2774,N_4649);
or U7129 (N_7129,N_3605,N_3188);
nand U7130 (N_7130,N_3026,N_3037);
nand U7131 (N_7131,N_4638,N_3872);
xnor U7132 (N_7132,N_3754,N_2720);
nand U7133 (N_7133,N_4637,N_4103);
nor U7134 (N_7134,N_4078,N_2815);
xor U7135 (N_7135,N_4374,N_4513);
nor U7136 (N_7136,N_2558,N_3110);
and U7137 (N_7137,N_2567,N_4093);
nor U7138 (N_7138,N_4156,N_3392);
nor U7139 (N_7139,N_4931,N_3110);
and U7140 (N_7140,N_4098,N_4603);
and U7141 (N_7141,N_3390,N_3590);
xnor U7142 (N_7142,N_3204,N_3437);
or U7143 (N_7143,N_4555,N_4223);
xor U7144 (N_7144,N_3703,N_3589);
nand U7145 (N_7145,N_3490,N_2560);
and U7146 (N_7146,N_4576,N_4912);
or U7147 (N_7147,N_2524,N_4523);
and U7148 (N_7148,N_4093,N_3184);
nor U7149 (N_7149,N_4740,N_4893);
or U7150 (N_7150,N_3079,N_4779);
nor U7151 (N_7151,N_4272,N_4861);
and U7152 (N_7152,N_3505,N_4880);
or U7153 (N_7153,N_2953,N_3659);
nor U7154 (N_7154,N_3556,N_3530);
or U7155 (N_7155,N_4655,N_3071);
nor U7156 (N_7156,N_4759,N_2640);
or U7157 (N_7157,N_4461,N_4597);
nand U7158 (N_7158,N_4675,N_4728);
xnor U7159 (N_7159,N_4232,N_2889);
nor U7160 (N_7160,N_4816,N_3538);
or U7161 (N_7161,N_2542,N_4485);
nand U7162 (N_7162,N_4990,N_3968);
nand U7163 (N_7163,N_4731,N_3823);
and U7164 (N_7164,N_3723,N_4557);
xnor U7165 (N_7165,N_2787,N_3543);
nor U7166 (N_7166,N_3426,N_3359);
nand U7167 (N_7167,N_3956,N_3048);
and U7168 (N_7168,N_4322,N_2571);
xnor U7169 (N_7169,N_3387,N_3701);
nor U7170 (N_7170,N_4745,N_4333);
xor U7171 (N_7171,N_4877,N_4369);
nor U7172 (N_7172,N_3362,N_3444);
xnor U7173 (N_7173,N_4445,N_4262);
nor U7174 (N_7174,N_4925,N_3461);
and U7175 (N_7175,N_3690,N_3284);
and U7176 (N_7176,N_3538,N_4898);
nor U7177 (N_7177,N_4802,N_2995);
nor U7178 (N_7178,N_3921,N_2577);
and U7179 (N_7179,N_3490,N_2699);
or U7180 (N_7180,N_4010,N_3107);
xnor U7181 (N_7181,N_3631,N_4816);
and U7182 (N_7182,N_4476,N_2993);
or U7183 (N_7183,N_2837,N_3043);
nand U7184 (N_7184,N_4889,N_4677);
nand U7185 (N_7185,N_3902,N_3839);
and U7186 (N_7186,N_2573,N_4094);
or U7187 (N_7187,N_4643,N_3565);
or U7188 (N_7188,N_3213,N_2705);
or U7189 (N_7189,N_3794,N_2763);
or U7190 (N_7190,N_4611,N_4168);
and U7191 (N_7191,N_2606,N_3160);
or U7192 (N_7192,N_4145,N_4008);
nand U7193 (N_7193,N_2857,N_4783);
nor U7194 (N_7194,N_3754,N_4897);
and U7195 (N_7195,N_4927,N_4463);
or U7196 (N_7196,N_4583,N_3172);
and U7197 (N_7197,N_3569,N_2745);
or U7198 (N_7198,N_4091,N_3372);
or U7199 (N_7199,N_3211,N_4149);
or U7200 (N_7200,N_4390,N_4175);
nand U7201 (N_7201,N_4471,N_4954);
or U7202 (N_7202,N_3441,N_4854);
and U7203 (N_7203,N_4066,N_4084);
nand U7204 (N_7204,N_4699,N_2554);
and U7205 (N_7205,N_3974,N_3040);
xnor U7206 (N_7206,N_3314,N_3596);
xor U7207 (N_7207,N_2657,N_3805);
xor U7208 (N_7208,N_3506,N_2570);
or U7209 (N_7209,N_4225,N_4054);
nor U7210 (N_7210,N_4696,N_2745);
nand U7211 (N_7211,N_3029,N_3690);
nor U7212 (N_7212,N_3162,N_4130);
and U7213 (N_7213,N_3978,N_3653);
or U7214 (N_7214,N_3653,N_2668);
xnor U7215 (N_7215,N_3432,N_2985);
nand U7216 (N_7216,N_4126,N_4591);
nand U7217 (N_7217,N_4347,N_4304);
nand U7218 (N_7218,N_2836,N_4109);
nand U7219 (N_7219,N_3719,N_4275);
or U7220 (N_7220,N_4717,N_4757);
nor U7221 (N_7221,N_4808,N_2844);
nand U7222 (N_7222,N_4493,N_2625);
xnor U7223 (N_7223,N_2533,N_3258);
xnor U7224 (N_7224,N_4622,N_3532);
and U7225 (N_7225,N_4737,N_3616);
nor U7226 (N_7226,N_2611,N_3694);
nor U7227 (N_7227,N_4379,N_3479);
xnor U7228 (N_7228,N_2947,N_3110);
xnor U7229 (N_7229,N_4015,N_4601);
nor U7230 (N_7230,N_2709,N_4695);
and U7231 (N_7231,N_4000,N_4533);
or U7232 (N_7232,N_4823,N_4741);
nor U7233 (N_7233,N_3098,N_2706);
or U7234 (N_7234,N_4463,N_2610);
or U7235 (N_7235,N_2958,N_4338);
or U7236 (N_7236,N_4851,N_2651);
xor U7237 (N_7237,N_3606,N_3689);
nand U7238 (N_7238,N_4946,N_3506);
and U7239 (N_7239,N_2870,N_3638);
and U7240 (N_7240,N_3752,N_3558);
xor U7241 (N_7241,N_3256,N_4328);
nor U7242 (N_7242,N_3531,N_2613);
and U7243 (N_7243,N_3965,N_3108);
nor U7244 (N_7244,N_4102,N_2707);
and U7245 (N_7245,N_3562,N_4206);
xor U7246 (N_7246,N_4721,N_4748);
xor U7247 (N_7247,N_3800,N_3445);
nand U7248 (N_7248,N_3269,N_4250);
xnor U7249 (N_7249,N_4348,N_2773);
xor U7250 (N_7250,N_4798,N_2582);
or U7251 (N_7251,N_4811,N_3333);
nand U7252 (N_7252,N_2569,N_2672);
and U7253 (N_7253,N_3764,N_4056);
xnor U7254 (N_7254,N_3460,N_3042);
or U7255 (N_7255,N_3636,N_3971);
and U7256 (N_7256,N_2760,N_4793);
nor U7257 (N_7257,N_4410,N_4763);
and U7258 (N_7258,N_2913,N_3984);
nor U7259 (N_7259,N_3360,N_3016);
or U7260 (N_7260,N_4438,N_3373);
or U7261 (N_7261,N_3861,N_3276);
or U7262 (N_7262,N_2886,N_3309);
nor U7263 (N_7263,N_3697,N_4717);
nor U7264 (N_7264,N_4384,N_3337);
or U7265 (N_7265,N_3232,N_3703);
and U7266 (N_7266,N_3015,N_4742);
nor U7267 (N_7267,N_3492,N_4702);
nand U7268 (N_7268,N_4373,N_3598);
nor U7269 (N_7269,N_3741,N_4005);
nand U7270 (N_7270,N_4086,N_2928);
nand U7271 (N_7271,N_4338,N_4675);
nand U7272 (N_7272,N_4888,N_4353);
xor U7273 (N_7273,N_3350,N_4946);
nand U7274 (N_7274,N_4605,N_3350);
nor U7275 (N_7275,N_4609,N_2649);
and U7276 (N_7276,N_2768,N_2666);
nor U7277 (N_7277,N_3225,N_4734);
xnor U7278 (N_7278,N_3779,N_4563);
nand U7279 (N_7279,N_2795,N_4448);
nor U7280 (N_7280,N_4813,N_3641);
nand U7281 (N_7281,N_3741,N_4994);
nor U7282 (N_7282,N_3879,N_3329);
nand U7283 (N_7283,N_4532,N_2718);
and U7284 (N_7284,N_3071,N_4939);
or U7285 (N_7285,N_2804,N_3946);
nor U7286 (N_7286,N_3530,N_3475);
nor U7287 (N_7287,N_4146,N_3009);
nor U7288 (N_7288,N_4120,N_4514);
and U7289 (N_7289,N_4662,N_4845);
xor U7290 (N_7290,N_4275,N_2582);
xnor U7291 (N_7291,N_3724,N_4882);
and U7292 (N_7292,N_2540,N_3078);
and U7293 (N_7293,N_3614,N_2718);
nand U7294 (N_7294,N_3933,N_3979);
and U7295 (N_7295,N_4259,N_3151);
xnor U7296 (N_7296,N_3883,N_2982);
nand U7297 (N_7297,N_3568,N_4094);
nand U7298 (N_7298,N_3535,N_4601);
or U7299 (N_7299,N_3445,N_2625);
xor U7300 (N_7300,N_3886,N_4533);
and U7301 (N_7301,N_3306,N_4082);
xor U7302 (N_7302,N_3136,N_2958);
nand U7303 (N_7303,N_3497,N_3495);
xnor U7304 (N_7304,N_2579,N_3692);
or U7305 (N_7305,N_4672,N_2871);
nor U7306 (N_7306,N_3548,N_2738);
and U7307 (N_7307,N_4735,N_4995);
xnor U7308 (N_7308,N_4105,N_3190);
nand U7309 (N_7309,N_4075,N_4225);
or U7310 (N_7310,N_3888,N_4958);
or U7311 (N_7311,N_4134,N_2863);
nor U7312 (N_7312,N_2669,N_3744);
and U7313 (N_7313,N_2608,N_4634);
xnor U7314 (N_7314,N_4439,N_2800);
or U7315 (N_7315,N_4333,N_4503);
nand U7316 (N_7316,N_2801,N_4165);
and U7317 (N_7317,N_3083,N_3026);
nor U7318 (N_7318,N_4106,N_3290);
and U7319 (N_7319,N_2991,N_3905);
nand U7320 (N_7320,N_4382,N_2543);
nor U7321 (N_7321,N_4657,N_2630);
nand U7322 (N_7322,N_3915,N_3636);
nor U7323 (N_7323,N_2981,N_4416);
nand U7324 (N_7324,N_3006,N_3212);
and U7325 (N_7325,N_4801,N_3024);
nand U7326 (N_7326,N_3148,N_4542);
nor U7327 (N_7327,N_2707,N_4740);
or U7328 (N_7328,N_2936,N_4294);
or U7329 (N_7329,N_2706,N_2997);
or U7330 (N_7330,N_4436,N_2704);
xor U7331 (N_7331,N_4086,N_3439);
or U7332 (N_7332,N_4570,N_4022);
xnor U7333 (N_7333,N_3556,N_2558);
or U7334 (N_7334,N_4765,N_3806);
or U7335 (N_7335,N_2816,N_4839);
or U7336 (N_7336,N_4346,N_4137);
or U7337 (N_7337,N_4492,N_4655);
or U7338 (N_7338,N_3308,N_4788);
or U7339 (N_7339,N_4949,N_4006);
nor U7340 (N_7340,N_4032,N_3784);
nor U7341 (N_7341,N_2724,N_4311);
xnor U7342 (N_7342,N_3449,N_4906);
and U7343 (N_7343,N_4560,N_3577);
nor U7344 (N_7344,N_3514,N_3505);
or U7345 (N_7345,N_4245,N_4373);
xor U7346 (N_7346,N_4728,N_3559);
nor U7347 (N_7347,N_4750,N_3566);
xor U7348 (N_7348,N_2526,N_3200);
xnor U7349 (N_7349,N_4379,N_4656);
and U7350 (N_7350,N_4474,N_3739);
nor U7351 (N_7351,N_4406,N_3580);
and U7352 (N_7352,N_3096,N_3929);
xnor U7353 (N_7353,N_4288,N_4361);
nor U7354 (N_7354,N_3475,N_4826);
and U7355 (N_7355,N_4628,N_3951);
xor U7356 (N_7356,N_3572,N_4433);
xor U7357 (N_7357,N_4380,N_3536);
nor U7358 (N_7358,N_3809,N_2545);
nand U7359 (N_7359,N_4211,N_3481);
nand U7360 (N_7360,N_4562,N_2984);
and U7361 (N_7361,N_2576,N_4720);
nor U7362 (N_7362,N_2933,N_3216);
and U7363 (N_7363,N_3881,N_2832);
xor U7364 (N_7364,N_3962,N_3922);
and U7365 (N_7365,N_4921,N_3338);
and U7366 (N_7366,N_2609,N_4498);
and U7367 (N_7367,N_3039,N_3844);
or U7368 (N_7368,N_2961,N_2676);
nand U7369 (N_7369,N_3288,N_2586);
and U7370 (N_7370,N_4779,N_4942);
xnor U7371 (N_7371,N_3133,N_4319);
nor U7372 (N_7372,N_4479,N_2913);
and U7373 (N_7373,N_4157,N_3103);
xor U7374 (N_7374,N_3289,N_3576);
and U7375 (N_7375,N_3993,N_2982);
and U7376 (N_7376,N_3447,N_3205);
and U7377 (N_7377,N_4303,N_3947);
xnor U7378 (N_7378,N_3303,N_4531);
nor U7379 (N_7379,N_2817,N_4722);
nor U7380 (N_7380,N_3960,N_2549);
or U7381 (N_7381,N_4212,N_4943);
and U7382 (N_7382,N_3597,N_2718);
xor U7383 (N_7383,N_4179,N_2733);
or U7384 (N_7384,N_4211,N_4937);
nand U7385 (N_7385,N_2867,N_2671);
xnor U7386 (N_7386,N_4899,N_2961);
or U7387 (N_7387,N_2753,N_2620);
nor U7388 (N_7388,N_2872,N_2594);
or U7389 (N_7389,N_4401,N_4147);
nand U7390 (N_7390,N_3966,N_3404);
xor U7391 (N_7391,N_3363,N_3899);
and U7392 (N_7392,N_3791,N_3535);
xor U7393 (N_7393,N_4541,N_2734);
or U7394 (N_7394,N_2999,N_4956);
or U7395 (N_7395,N_2876,N_2868);
and U7396 (N_7396,N_4298,N_4174);
and U7397 (N_7397,N_4067,N_4983);
xor U7398 (N_7398,N_3972,N_2984);
and U7399 (N_7399,N_4902,N_3745);
nor U7400 (N_7400,N_3044,N_4195);
nor U7401 (N_7401,N_3471,N_3717);
nand U7402 (N_7402,N_4403,N_4806);
nand U7403 (N_7403,N_4326,N_4294);
xor U7404 (N_7404,N_4796,N_3347);
xnor U7405 (N_7405,N_2673,N_4015);
nand U7406 (N_7406,N_3916,N_4396);
nor U7407 (N_7407,N_3642,N_2733);
or U7408 (N_7408,N_3205,N_2767);
and U7409 (N_7409,N_4393,N_4143);
nor U7410 (N_7410,N_3938,N_3263);
or U7411 (N_7411,N_4709,N_2866);
and U7412 (N_7412,N_4264,N_4738);
nor U7413 (N_7413,N_4908,N_4960);
and U7414 (N_7414,N_4164,N_4509);
nor U7415 (N_7415,N_4912,N_4262);
and U7416 (N_7416,N_3294,N_2796);
xnor U7417 (N_7417,N_2689,N_4165);
or U7418 (N_7418,N_4088,N_4098);
xor U7419 (N_7419,N_2857,N_3450);
xor U7420 (N_7420,N_4812,N_4320);
and U7421 (N_7421,N_3773,N_2666);
xnor U7422 (N_7422,N_3492,N_4001);
nand U7423 (N_7423,N_3250,N_4823);
nor U7424 (N_7424,N_3098,N_3662);
or U7425 (N_7425,N_4220,N_4371);
nand U7426 (N_7426,N_3633,N_3621);
nor U7427 (N_7427,N_3441,N_3747);
xor U7428 (N_7428,N_4377,N_2710);
or U7429 (N_7429,N_4457,N_2907);
nand U7430 (N_7430,N_3103,N_4778);
nor U7431 (N_7431,N_4419,N_4333);
nand U7432 (N_7432,N_3826,N_3688);
or U7433 (N_7433,N_3045,N_2920);
nor U7434 (N_7434,N_3211,N_2934);
or U7435 (N_7435,N_3776,N_4689);
and U7436 (N_7436,N_4322,N_3108);
or U7437 (N_7437,N_3312,N_4270);
and U7438 (N_7438,N_4162,N_2687);
xnor U7439 (N_7439,N_3972,N_4537);
nor U7440 (N_7440,N_4796,N_3428);
nand U7441 (N_7441,N_4255,N_4960);
nand U7442 (N_7442,N_2937,N_2527);
and U7443 (N_7443,N_4115,N_3259);
and U7444 (N_7444,N_3525,N_4365);
nand U7445 (N_7445,N_4611,N_4420);
nand U7446 (N_7446,N_3509,N_3865);
xnor U7447 (N_7447,N_2854,N_3283);
nand U7448 (N_7448,N_3245,N_3414);
and U7449 (N_7449,N_3243,N_2789);
or U7450 (N_7450,N_2725,N_3724);
nor U7451 (N_7451,N_4217,N_4675);
or U7452 (N_7452,N_3601,N_4216);
xor U7453 (N_7453,N_3282,N_4457);
nor U7454 (N_7454,N_3231,N_4894);
or U7455 (N_7455,N_3607,N_4139);
nand U7456 (N_7456,N_4925,N_4197);
nor U7457 (N_7457,N_4486,N_3372);
or U7458 (N_7458,N_4031,N_3309);
nor U7459 (N_7459,N_4730,N_3748);
nor U7460 (N_7460,N_2987,N_2752);
or U7461 (N_7461,N_3970,N_4890);
and U7462 (N_7462,N_4156,N_4176);
and U7463 (N_7463,N_3259,N_4129);
xor U7464 (N_7464,N_4553,N_3576);
or U7465 (N_7465,N_4228,N_3807);
nand U7466 (N_7466,N_3950,N_4776);
xnor U7467 (N_7467,N_2714,N_3592);
nand U7468 (N_7468,N_2602,N_3063);
or U7469 (N_7469,N_3468,N_4117);
or U7470 (N_7470,N_3879,N_2797);
and U7471 (N_7471,N_4098,N_2952);
nand U7472 (N_7472,N_4443,N_2542);
nand U7473 (N_7473,N_3106,N_4820);
nor U7474 (N_7474,N_4823,N_2989);
nand U7475 (N_7475,N_4556,N_3374);
and U7476 (N_7476,N_3829,N_2970);
or U7477 (N_7477,N_3058,N_4577);
xor U7478 (N_7478,N_4309,N_2670);
nor U7479 (N_7479,N_3019,N_4362);
nor U7480 (N_7480,N_3438,N_2657);
and U7481 (N_7481,N_2670,N_3183);
nor U7482 (N_7482,N_4688,N_3465);
nor U7483 (N_7483,N_2610,N_4682);
nor U7484 (N_7484,N_2813,N_4186);
or U7485 (N_7485,N_4293,N_3521);
and U7486 (N_7486,N_3219,N_4374);
nor U7487 (N_7487,N_3742,N_3231);
or U7488 (N_7488,N_4275,N_3686);
nand U7489 (N_7489,N_4901,N_2501);
nand U7490 (N_7490,N_3891,N_3018);
nor U7491 (N_7491,N_3191,N_4399);
nor U7492 (N_7492,N_4707,N_3876);
or U7493 (N_7493,N_4868,N_3573);
nand U7494 (N_7494,N_3841,N_4620);
xor U7495 (N_7495,N_4683,N_3151);
or U7496 (N_7496,N_2771,N_4273);
or U7497 (N_7497,N_3444,N_2745);
and U7498 (N_7498,N_3273,N_4090);
nand U7499 (N_7499,N_4498,N_2587);
or U7500 (N_7500,N_7390,N_6349);
or U7501 (N_7501,N_5530,N_5772);
xnor U7502 (N_7502,N_6447,N_6511);
nand U7503 (N_7503,N_6508,N_7457);
xnor U7504 (N_7504,N_5705,N_5189);
nand U7505 (N_7505,N_5792,N_5216);
xor U7506 (N_7506,N_5934,N_6072);
and U7507 (N_7507,N_6970,N_5817);
nand U7508 (N_7508,N_6356,N_6293);
nand U7509 (N_7509,N_5857,N_6085);
and U7510 (N_7510,N_5135,N_5402);
nand U7511 (N_7511,N_5725,N_7415);
or U7512 (N_7512,N_5999,N_7095);
xnor U7513 (N_7513,N_6324,N_6055);
and U7514 (N_7514,N_5200,N_6022);
xnor U7515 (N_7515,N_6229,N_6272);
and U7516 (N_7516,N_6310,N_7492);
nand U7517 (N_7517,N_5115,N_5472);
nor U7518 (N_7518,N_6778,N_7302);
or U7519 (N_7519,N_7349,N_5665);
nor U7520 (N_7520,N_5034,N_7294);
nand U7521 (N_7521,N_5796,N_5214);
or U7522 (N_7522,N_7073,N_5460);
and U7523 (N_7523,N_6953,N_6692);
nor U7524 (N_7524,N_7091,N_6120);
xnor U7525 (N_7525,N_5848,N_5639);
nor U7526 (N_7526,N_5161,N_6737);
nand U7527 (N_7527,N_7358,N_6122);
xor U7528 (N_7528,N_7374,N_6113);
or U7529 (N_7529,N_6541,N_6433);
nor U7530 (N_7530,N_5106,N_7029);
and U7531 (N_7531,N_6018,N_6769);
or U7532 (N_7532,N_5950,N_5112);
nand U7533 (N_7533,N_5630,N_5248);
and U7534 (N_7534,N_5465,N_6593);
nor U7535 (N_7535,N_5127,N_5209);
and U7536 (N_7536,N_6030,N_7327);
or U7537 (N_7537,N_5096,N_6691);
xnor U7538 (N_7538,N_5610,N_6994);
nand U7539 (N_7539,N_5253,N_7317);
or U7540 (N_7540,N_7257,N_6276);
xnor U7541 (N_7541,N_6024,N_5450);
nor U7542 (N_7542,N_6532,N_6282);
xor U7543 (N_7543,N_7168,N_6884);
xnor U7544 (N_7544,N_6245,N_6173);
nand U7545 (N_7545,N_7410,N_5063);
or U7546 (N_7546,N_5957,N_6244);
or U7547 (N_7547,N_6971,N_7241);
nand U7548 (N_7548,N_6452,N_6852);
nand U7549 (N_7549,N_7036,N_7391);
nor U7550 (N_7550,N_6557,N_6649);
nor U7551 (N_7551,N_5653,N_6608);
nor U7552 (N_7552,N_5418,N_5692);
nand U7553 (N_7553,N_5607,N_5855);
xnor U7554 (N_7554,N_7218,N_5880);
and U7555 (N_7555,N_5844,N_6596);
and U7556 (N_7556,N_6257,N_7493);
xnor U7557 (N_7557,N_5237,N_6377);
and U7558 (N_7558,N_6958,N_5094);
xor U7559 (N_7559,N_6800,N_5730);
or U7560 (N_7560,N_5286,N_7201);
nor U7561 (N_7561,N_7476,N_7392);
and U7562 (N_7562,N_6683,N_7301);
xnor U7563 (N_7563,N_6715,N_5419);
and U7564 (N_7564,N_7446,N_5411);
xnor U7565 (N_7565,N_6560,N_7086);
or U7566 (N_7566,N_6001,N_6076);
nand U7567 (N_7567,N_6662,N_7396);
and U7568 (N_7568,N_6862,N_7094);
nand U7569 (N_7569,N_5138,N_5350);
or U7570 (N_7570,N_6496,N_7130);
xor U7571 (N_7571,N_6809,N_6960);
or U7572 (N_7572,N_6627,N_6540);
or U7573 (N_7573,N_6318,N_5806);
nand U7574 (N_7574,N_5697,N_7092);
nand U7575 (N_7575,N_5318,N_5433);
nor U7576 (N_7576,N_6652,N_5375);
xor U7577 (N_7577,N_5654,N_6527);
and U7578 (N_7578,N_6198,N_6071);
xor U7579 (N_7579,N_7107,N_5833);
nor U7580 (N_7580,N_6039,N_7019);
nand U7581 (N_7581,N_6822,N_6591);
or U7582 (N_7582,N_5882,N_7297);
xnor U7583 (N_7583,N_6690,N_5786);
or U7584 (N_7584,N_6562,N_5232);
and U7585 (N_7585,N_5013,N_5660);
and U7586 (N_7586,N_6297,N_6668);
xor U7587 (N_7587,N_5552,N_5159);
nor U7588 (N_7588,N_6184,N_5977);
nor U7589 (N_7589,N_5005,N_5525);
or U7590 (N_7590,N_6028,N_7269);
and U7591 (N_7591,N_6736,N_5073);
or U7592 (N_7592,N_6456,N_7346);
nand U7593 (N_7593,N_6416,N_6760);
nand U7594 (N_7594,N_5881,N_6016);
nand U7595 (N_7595,N_5603,N_7286);
or U7596 (N_7596,N_5533,N_7287);
xor U7597 (N_7597,N_6892,N_7261);
xnor U7598 (N_7598,N_5541,N_6674);
or U7599 (N_7599,N_5695,N_6186);
and U7600 (N_7600,N_5234,N_6873);
nand U7601 (N_7601,N_5694,N_5685);
and U7602 (N_7602,N_5536,N_5688);
xnor U7603 (N_7603,N_6929,N_6187);
and U7604 (N_7604,N_5324,N_5733);
nand U7605 (N_7605,N_6576,N_6483);
nor U7606 (N_7606,N_5279,N_5929);
nand U7607 (N_7607,N_6740,N_6226);
nand U7608 (N_7608,N_6175,N_6107);
or U7609 (N_7609,N_6845,N_5345);
xor U7610 (N_7610,N_7025,N_6921);
xnor U7611 (N_7611,N_7109,N_6969);
nor U7612 (N_7612,N_6987,N_5343);
nand U7613 (N_7613,N_5262,N_6831);
or U7614 (N_7614,N_6756,N_5722);
nand U7615 (N_7615,N_5176,N_6752);
nand U7616 (N_7616,N_5462,N_6328);
xnor U7617 (N_7617,N_5192,N_5739);
xor U7618 (N_7618,N_5782,N_5947);
or U7619 (N_7619,N_7401,N_7122);
nand U7620 (N_7620,N_7311,N_7322);
or U7621 (N_7621,N_5898,N_7223);
or U7622 (N_7622,N_5829,N_5937);
and U7623 (N_7623,N_7151,N_5001);
nand U7624 (N_7624,N_5217,N_5448);
or U7625 (N_7625,N_6636,N_7234);
and U7626 (N_7626,N_5308,N_6474);
nor U7627 (N_7627,N_5342,N_6991);
and U7628 (N_7628,N_5471,N_7451);
nor U7629 (N_7629,N_6457,N_6200);
nor U7630 (N_7630,N_6743,N_5015);
or U7631 (N_7631,N_7207,N_6855);
nand U7632 (N_7632,N_6367,N_5229);
nand U7633 (N_7633,N_7440,N_5596);
and U7634 (N_7634,N_5781,N_7146);
nor U7635 (N_7635,N_7143,N_6643);
and U7636 (N_7636,N_6926,N_6035);
xnor U7637 (N_7637,N_7368,N_6777);
nor U7638 (N_7638,N_5434,N_5316);
and U7639 (N_7639,N_7382,N_6336);
nor U7640 (N_7640,N_7189,N_7418);
and U7641 (N_7641,N_5297,N_6753);
or U7642 (N_7642,N_6426,N_6125);
xnor U7643 (N_7643,N_6917,N_5128);
nand U7644 (N_7644,N_5206,N_5687);
and U7645 (N_7645,N_7467,N_7357);
nand U7646 (N_7646,N_6091,N_5900);
nor U7647 (N_7647,N_7149,N_6597);
and U7648 (N_7648,N_5721,N_6667);
and U7649 (N_7649,N_5632,N_6555);
nor U7650 (N_7650,N_5803,N_5720);
nor U7651 (N_7651,N_6682,N_7360);
xnor U7652 (N_7652,N_6017,N_7370);
nand U7653 (N_7653,N_7147,N_7248);
nor U7654 (N_7654,N_6203,N_5018);
nor U7655 (N_7655,N_6007,N_6536);
xor U7656 (N_7656,N_6851,N_7246);
nor U7657 (N_7657,N_6195,N_5989);
or U7658 (N_7658,N_5769,N_5897);
nor U7659 (N_7659,N_6906,N_7075);
or U7660 (N_7660,N_6403,N_5995);
nand U7661 (N_7661,N_7059,N_6083);
and U7662 (N_7662,N_6946,N_7018);
or U7663 (N_7663,N_5489,N_5033);
xnor U7664 (N_7664,N_5809,N_5502);
nand U7665 (N_7665,N_5435,N_5506);
nor U7666 (N_7666,N_5913,N_5355);
or U7667 (N_7667,N_5773,N_7238);
nand U7668 (N_7668,N_6032,N_6810);
or U7669 (N_7669,N_6728,N_5028);
or U7670 (N_7670,N_6641,N_7138);
nand U7671 (N_7671,N_6115,N_6241);
xor U7672 (N_7672,N_7131,N_5668);
nor U7673 (N_7673,N_6653,N_6348);
xnor U7674 (N_7674,N_5710,N_6242);
nand U7675 (N_7675,N_7343,N_5540);
nor U7676 (N_7676,N_6407,N_6026);
or U7677 (N_7677,N_5867,N_7008);
nand U7678 (N_7678,N_5284,N_5495);
nor U7679 (N_7679,N_5949,N_7173);
nand U7680 (N_7680,N_5129,N_5246);
xnor U7681 (N_7681,N_5859,N_6044);
xor U7682 (N_7682,N_5119,N_7152);
xnor U7683 (N_7683,N_7288,N_5439);
nand U7684 (N_7684,N_6650,N_5706);
or U7685 (N_7685,N_5932,N_5547);
or U7686 (N_7686,N_5992,N_5481);
or U7687 (N_7687,N_6706,N_5320);
xnor U7688 (N_7688,N_5601,N_5340);
and U7689 (N_7689,N_7264,N_6751);
and U7690 (N_7690,N_6366,N_5312);
nand U7691 (N_7691,N_6931,N_5738);
nor U7692 (N_7692,N_6069,N_5838);
nand U7693 (N_7693,N_5363,N_5716);
xnor U7694 (N_7694,N_6219,N_6619);
nor U7695 (N_7695,N_5445,N_7193);
xnor U7696 (N_7696,N_6135,N_7011);
nand U7697 (N_7697,N_6982,N_6110);
and U7698 (N_7698,N_7273,N_5178);
nor U7699 (N_7699,N_6501,N_6616);
nor U7700 (N_7700,N_6043,N_5538);
xor U7701 (N_7701,N_5917,N_6793);
xor U7702 (N_7702,N_7045,N_5130);
and U7703 (N_7703,N_6867,N_6856);
xnor U7704 (N_7704,N_5628,N_5226);
and U7705 (N_7705,N_7290,N_6734);
nand U7706 (N_7706,N_6615,N_5595);
and U7707 (N_7707,N_7206,N_5605);
or U7708 (N_7708,N_6334,N_6630);
and U7709 (N_7709,N_5650,N_5008);
nand U7710 (N_7710,N_5975,N_5671);
nor U7711 (N_7711,N_5633,N_5746);
nor U7712 (N_7712,N_5409,N_5466);
or U7713 (N_7713,N_6454,N_6701);
nor U7714 (N_7714,N_5948,N_5441);
nor U7715 (N_7715,N_5927,N_6123);
and U7716 (N_7716,N_6546,N_5459);
nand U7717 (N_7717,N_7432,N_6677);
and U7718 (N_7718,N_6640,N_6181);
xor U7719 (N_7719,N_7425,N_6573);
nor U7720 (N_7720,N_6111,N_5485);
and U7721 (N_7721,N_6236,N_5800);
or U7722 (N_7722,N_6357,N_5813);
nor U7723 (N_7723,N_6484,N_7190);
xnor U7724 (N_7724,N_6844,N_5099);
nand U7725 (N_7725,N_7420,N_7466);
nand U7726 (N_7726,N_5449,N_5087);
nand U7727 (N_7727,N_5114,N_5606);
and U7728 (N_7728,N_6581,N_5236);
xnor U7729 (N_7729,N_6171,N_7030);
nand U7730 (N_7730,N_6725,N_7461);
nand U7731 (N_7731,N_6149,N_6933);
nand U7732 (N_7732,N_6054,N_7389);
xnor U7733 (N_7733,N_6232,N_6658);
nor U7734 (N_7734,N_7009,N_6977);
and U7735 (N_7735,N_6185,N_6827);
and U7736 (N_7736,N_6666,N_6141);
nand U7737 (N_7737,N_5560,N_6839);
xor U7738 (N_7738,N_5887,N_5821);
nand U7739 (N_7739,N_6162,N_6216);
or U7740 (N_7740,N_6944,N_6466);
nand U7741 (N_7741,N_6595,N_5615);
nand U7742 (N_7742,N_7385,N_6296);
nor U7743 (N_7743,N_5689,N_6673);
nor U7744 (N_7744,N_5251,N_7077);
nor U7745 (N_7745,N_5580,N_6579);
nor U7746 (N_7746,N_7039,N_5837);
nand U7747 (N_7747,N_7178,N_5670);
nor U7748 (N_7748,N_5858,N_5583);
or U7749 (N_7749,N_7135,N_7249);
or U7750 (N_7750,N_5933,N_5860);
and U7751 (N_7751,N_5699,N_6190);
and U7752 (N_7752,N_5609,N_6240);
nand U7753 (N_7753,N_6235,N_5469);
and U7754 (N_7754,N_6518,N_5923);
nand U7755 (N_7755,N_6699,N_5420);
or U7756 (N_7756,N_6303,N_5513);
nand U7757 (N_7757,N_6369,N_6380);
nand U7758 (N_7758,N_5959,N_5338);
nand U7759 (N_7759,N_5458,N_7049);
or U7760 (N_7760,N_5600,N_5511);
nor U7761 (N_7761,N_6470,N_6872);
xnor U7762 (N_7762,N_5684,N_5423);
xor U7763 (N_7763,N_5354,N_5719);
or U7764 (N_7764,N_5916,N_6217);
nand U7765 (N_7765,N_7215,N_6770);
nor U7766 (N_7766,N_6840,N_7139);
nor U7767 (N_7767,N_7335,N_7012);
nor U7768 (N_7768,N_5870,N_7277);
and U7769 (N_7769,N_5282,N_6811);
and U7770 (N_7770,N_5010,N_7427);
and U7771 (N_7771,N_5840,N_6212);
and U7772 (N_7772,N_7491,N_5543);
nand U7773 (N_7773,N_5035,N_7235);
and U7774 (N_7774,N_5404,N_7081);
and U7775 (N_7775,N_5007,N_7226);
nand U7776 (N_7776,N_5118,N_6823);
nand U7777 (N_7777,N_5962,N_6813);
and U7778 (N_7778,N_5056,N_5673);
or U7779 (N_7779,N_7419,N_7462);
or U7780 (N_7780,N_6904,N_7089);
xnor U7781 (N_7781,N_6014,N_6819);
nand U7782 (N_7782,N_5197,N_6561);
and U7783 (N_7783,N_6340,N_5331);
or U7784 (N_7784,N_5539,N_6847);
xnor U7785 (N_7785,N_5845,N_5339);
and U7786 (N_7786,N_5698,N_5535);
xor U7787 (N_7787,N_7098,N_6460);
nor U7788 (N_7788,N_6126,N_6264);
and U7789 (N_7789,N_6776,N_5184);
xor U7790 (N_7790,N_5271,N_5915);
or U7791 (N_7791,N_5059,N_5785);
and U7792 (N_7792,N_5604,N_5202);
nor U7793 (N_7793,N_7123,N_5139);
nand U7794 (N_7794,N_5240,N_6271);
nand U7795 (N_7795,N_7478,N_5017);
or U7796 (N_7796,N_6693,N_7097);
nor U7797 (N_7797,N_5274,N_6721);
xor U7798 (N_7798,N_6999,N_5378);
or U7799 (N_7799,N_5478,N_7268);
nand U7800 (N_7800,N_6464,N_6785);
nand U7801 (N_7801,N_6758,N_7198);
xor U7802 (N_7802,N_5242,N_6495);
nand U7803 (N_7803,N_7101,N_6140);
or U7804 (N_7804,N_6473,N_6559);
nor U7805 (N_7805,N_6385,N_5476);
and U7806 (N_7806,N_6624,N_7371);
xor U7807 (N_7807,N_5238,N_6422);
or U7808 (N_7808,N_5473,N_6459);
or U7809 (N_7809,N_5333,N_6611);
xnor U7810 (N_7810,N_6409,N_7027);
nor U7811 (N_7811,N_6489,N_5815);
xor U7812 (N_7812,N_6976,N_5198);
xnor U7813 (N_7813,N_5620,N_6723);
and U7814 (N_7814,N_5662,N_5255);
nand U7815 (N_7815,N_6830,N_6879);
and U7816 (N_7816,N_7166,N_5527);
and U7817 (N_7817,N_5199,N_6520);
nor U7818 (N_7818,N_5122,N_5045);
or U7819 (N_7819,N_5414,N_7158);
nor U7820 (N_7820,N_6764,N_5515);
nor U7821 (N_7821,N_5092,N_6121);
and U7822 (N_7822,N_6246,N_5145);
xnor U7823 (N_7823,N_5040,N_7085);
and U7824 (N_7824,N_5407,N_7087);
nand U7825 (N_7825,N_5613,N_5143);
and U7826 (N_7826,N_7284,N_7006);
or U7827 (N_7827,N_5847,N_6912);
and U7828 (N_7828,N_5336,N_6471);
nor U7829 (N_7829,N_5006,N_5967);
nor U7830 (N_7830,N_7378,N_5366);
or U7831 (N_7831,N_5589,N_5842);
and U7832 (N_7832,N_6942,N_6494);
xnor U7833 (N_7833,N_7079,N_7154);
or U7834 (N_7834,N_6535,N_7452);
and U7835 (N_7835,N_5546,N_6761);
or U7836 (N_7836,N_5287,N_6712);
xnor U7837 (N_7837,N_5759,N_6045);
nand U7838 (N_7838,N_5454,N_6599);
or U7839 (N_7839,N_5621,N_5909);
or U7840 (N_7840,N_5531,N_5283);
nand U7841 (N_7841,N_6739,N_5510);
xor U7842 (N_7842,N_5966,N_6945);
xnor U7843 (N_7843,N_7066,N_6100);
nand U7844 (N_7844,N_6503,N_6763);
nor U7845 (N_7845,N_6364,N_6963);
nor U7846 (N_7846,N_5497,N_7195);
or U7847 (N_7847,N_5368,N_7416);
or U7848 (N_7848,N_6803,N_7369);
and U7849 (N_7849,N_6021,N_7340);
and U7850 (N_7850,N_5003,N_5883);
nor U7851 (N_7851,N_6694,N_6404);
nand U7852 (N_7852,N_5463,N_5179);
nor U7853 (N_7853,N_7342,N_5252);
and U7854 (N_7854,N_6439,N_7103);
xnor U7855 (N_7855,N_5386,N_5791);
and U7856 (N_7856,N_5461,N_6675);
or U7857 (N_7857,N_6394,N_7188);
nand U7858 (N_7858,N_5727,N_5464);
xor U7859 (N_7859,N_6702,N_5911);
xor U7860 (N_7860,N_6345,N_5623);
or U7861 (N_7861,N_6808,N_7161);
or U7862 (N_7862,N_5765,N_5853);
xnor U7863 (N_7863,N_6986,N_6932);
or U7864 (N_7864,N_7219,N_5379);
or U7865 (N_7865,N_7316,N_5154);
and U7866 (N_7866,N_7240,N_6850);
xnor U7867 (N_7867,N_7080,N_5961);
nor U7868 (N_7868,N_5222,N_6934);
and U7869 (N_7869,N_6388,N_5270);
and U7870 (N_7870,N_6883,N_5009);
and U7871 (N_7871,N_6151,N_7351);
nand U7872 (N_7872,N_7397,N_5690);
or U7873 (N_7873,N_7383,N_6622);
and U7874 (N_7874,N_6773,N_5888);
nor U7875 (N_7875,N_7324,N_7328);
and U7876 (N_7876,N_5349,N_6664);
or U7877 (N_7877,N_5146,N_5227);
nand U7878 (N_7878,N_5292,N_7084);
xor U7879 (N_7879,N_6603,N_6697);
nand U7880 (N_7880,N_5072,N_5212);
nand U7881 (N_7881,N_6335,N_6886);
or U7882 (N_7882,N_7388,N_5125);
xor U7883 (N_7883,N_5616,N_5669);
nor U7884 (N_7884,N_5475,N_5327);
nor U7885 (N_7885,N_6825,N_6317);
and U7886 (N_7886,N_6256,N_7184);
xnor U7887 (N_7887,N_7165,N_5239);
nor U7888 (N_7888,N_5295,N_6263);
xor U7889 (N_7889,N_5259,N_5208);
xor U7890 (N_7890,N_5281,N_5373);
xor U7891 (N_7891,N_5391,N_7118);
nand U7892 (N_7892,N_5869,N_7162);
xnor U7893 (N_7893,N_6368,N_5732);
nand U7894 (N_7894,N_6829,N_7472);
and U7895 (N_7895,N_5424,N_6424);
or U7896 (N_7896,N_5528,N_6027);
nor U7897 (N_7897,N_6646,N_5401);
or U7898 (N_7898,N_6136,N_6020);
or U7899 (N_7899,N_5807,N_5862);
nor U7900 (N_7900,N_5814,N_5770);
xnor U7901 (N_7901,N_6314,N_7229);
nor U7902 (N_7902,N_6259,N_6635);
nand U7903 (N_7903,N_6634,N_5737);
nand U7904 (N_7904,N_7475,N_6922);
or U7905 (N_7905,N_7377,N_7498);
nand U7906 (N_7906,N_7295,N_7348);
or U7907 (N_7907,N_6613,N_5592);
and U7908 (N_7908,N_5885,N_5672);
nand U7909 (N_7909,N_7453,N_6997);
xor U7910 (N_7910,N_6057,N_6589);
or U7911 (N_7911,N_6300,N_5392);
nor U7912 (N_7912,N_6247,N_5181);
xnor U7913 (N_7913,N_6949,N_5574);
nand U7914 (N_7914,N_6871,N_5228);
and U7915 (N_7915,N_7037,N_5514);
xor U7916 (N_7916,N_6816,N_7034);
nor U7917 (N_7917,N_5451,N_5661);
nand U7918 (N_7918,N_6291,N_5643);
xor U7919 (N_7919,N_6907,N_5652);
or U7920 (N_7920,N_5123,N_6323);
or U7921 (N_7921,N_6313,N_6669);
xnor U7922 (N_7922,N_7259,N_6432);
and U7923 (N_7923,N_5500,N_6476);
xor U7924 (N_7924,N_5309,N_7291);
nor U7925 (N_7925,N_7445,N_5030);
or U7926 (N_7926,N_5986,N_5522);
or U7927 (N_7927,N_6552,N_6529);
and U7928 (N_7928,N_6610,N_6009);
nor U7929 (N_7929,N_7347,N_6801);
nand U7930 (N_7930,N_6465,N_6802);
or U7931 (N_7931,N_7014,N_5376);
nor U7932 (N_7932,N_6360,N_7244);
and U7933 (N_7933,N_7366,N_6787);
and U7934 (N_7934,N_5693,N_5337);
nor U7935 (N_7935,N_5841,N_7058);
nand U7936 (N_7936,N_6746,N_5098);
nor U7937 (N_7937,N_5958,N_6854);
nand U7938 (N_7938,N_6431,N_5456);
or U7939 (N_7939,N_7265,N_5077);
and U7940 (N_7940,N_5026,N_5306);
and U7941 (N_7941,N_6866,N_5415);
xor U7942 (N_7942,N_7127,N_5873);
nand U7943 (N_7943,N_6420,N_6563);
or U7944 (N_7944,N_7454,N_5205);
xnor U7945 (N_7945,N_7171,N_6642);
and U7946 (N_7946,N_7434,N_6250);
and U7947 (N_7947,N_5682,N_5677);
or U7948 (N_7948,N_6889,N_6860);
nor U7949 (N_7949,N_5120,N_5365);
xnor U7950 (N_7950,N_6428,N_5194);
nor U7951 (N_7951,N_7145,N_5074);
nand U7952 (N_7952,N_6004,N_5593);
or U7953 (N_7953,N_6477,N_5261);
or U7954 (N_7954,N_7481,N_5755);
nor U7955 (N_7955,N_7289,N_6909);
xnor U7956 (N_7956,N_5707,N_6099);
nor U7957 (N_7957,N_6713,N_6647);
and U7958 (N_7958,N_6755,N_6209);
or U7959 (N_7959,N_6170,N_7033);
nor U7960 (N_7960,N_5753,N_5488);
nand U7961 (N_7961,N_5884,N_7444);
and U7962 (N_7962,N_5784,N_7280);
nor U7963 (N_7963,N_5068,N_7004);
and U7964 (N_7964,N_6019,N_5575);
and U7965 (N_7965,N_7069,N_6047);
and U7966 (N_7966,N_6089,N_7140);
or U7967 (N_7967,N_5381,N_7242);
and U7968 (N_7968,N_6502,N_5047);
nand U7969 (N_7969,N_6178,N_6657);
nand U7970 (N_7970,N_5190,N_7499);
nand U7971 (N_7971,N_5905,N_5997);
nor U7972 (N_7972,N_7022,N_5468);
or U7973 (N_7973,N_5969,N_6578);
or U7974 (N_7974,N_6362,N_6878);
nor U7975 (N_7975,N_6485,N_6700);
or U7976 (N_7976,N_7251,N_6981);
or U7977 (N_7977,N_7353,N_5490);
nor U7978 (N_7978,N_5083,N_6530);
nor U7979 (N_7979,N_5132,N_5484);
nand U7980 (N_7980,N_7225,N_5301);
and U7981 (N_7981,N_6451,N_6900);
nand U7982 (N_7982,N_6343,N_5117);
or U7983 (N_7983,N_6423,N_7061);
and U7984 (N_7984,N_5608,N_6732);
xnor U7985 (N_7985,N_7001,N_5830);
or U7986 (N_7986,N_7394,N_7088);
or U7987 (N_7987,N_6567,N_5091);
or U7988 (N_7988,N_6183,N_6771);
nand U7989 (N_7989,N_6533,N_6584);
nand U7990 (N_7990,N_7344,N_5496);
xor U7991 (N_7991,N_7482,N_6188);
xnor U7992 (N_7992,N_6880,N_5012);
nand U7993 (N_7993,N_7200,N_7417);
nor U7994 (N_7994,N_5902,N_5076);
xor U7995 (N_7995,N_5836,N_6637);
nand U7996 (N_7996,N_6227,N_5799);
nor U7997 (N_7997,N_6143,N_7495);
xor U7998 (N_7998,N_6056,N_6097);
nand U7999 (N_7999,N_5517,N_5914);
and U8000 (N_8000,N_6923,N_6656);
and U8001 (N_8001,N_6168,N_7187);
and U8002 (N_8002,N_7469,N_5300);
nor U8003 (N_8003,N_5055,N_5988);
nand U8004 (N_8004,N_5219,N_7477);
nor U8005 (N_8005,N_5935,N_6620);
and U8006 (N_8006,N_7384,N_5417);
nand U8007 (N_8007,N_6260,N_7026);
and U8008 (N_8008,N_7448,N_6008);
or U8009 (N_8009,N_5371,N_5372);
nor U8010 (N_8010,N_6663,N_5569);
nor U8011 (N_8011,N_6425,N_6305);
nand U8012 (N_8012,N_5597,N_5649);
nand U8013 (N_8013,N_7456,N_6671);
nand U8014 (N_8014,N_6606,N_5747);
or U8015 (N_8015,N_7192,N_7422);
and U8016 (N_8016,N_6445,N_6835);
nor U8017 (N_8017,N_7015,N_5131);
nor U8018 (N_8018,N_6436,N_5731);
nand U8019 (N_8019,N_6547,N_7279);
nor U8020 (N_8020,N_7313,N_6458);
nor U8021 (N_8021,N_5060,N_7055);
nand U8022 (N_8022,N_5922,N_6449);
xor U8023 (N_8023,N_7338,N_7310);
and U8024 (N_8024,N_7038,N_5944);
or U8025 (N_8025,N_5571,N_5573);
or U8026 (N_8026,N_5851,N_6077);
or U8027 (N_8027,N_5408,N_6719);
or U8028 (N_8028,N_5344,N_7157);
nor U8029 (N_8029,N_5648,N_5195);
nor U8030 (N_8030,N_6644,N_5942);
nor U8031 (N_8031,N_5004,N_6538);
xor U8032 (N_8032,N_7175,N_7380);
nor U8033 (N_8033,N_7325,N_6196);
or U8034 (N_8034,N_7413,N_5256);
or U8035 (N_8035,N_6843,N_5728);
and U8036 (N_8036,N_6228,N_7044);
nor U8037 (N_8037,N_6583,N_7428);
and U8038 (N_8038,N_5903,N_5827);
and U8039 (N_8039,N_5069,N_6002);
xnor U8040 (N_8040,N_6182,N_5526);
or U8041 (N_8041,N_6029,N_7115);
and U8042 (N_8042,N_5912,N_6602);
or U8043 (N_8043,N_5360,N_6116);
or U8044 (N_8044,N_5824,N_7485);
xor U8045 (N_8045,N_5941,N_6522);
nand U8046 (N_8046,N_6096,N_6372);
xor U8047 (N_8047,N_7105,N_7308);
and U8048 (N_8048,N_7455,N_6497);
nor U8049 (N_8049,N_5521,N_6478);
or U8050 (N_8050,N_6322,N_5021);
nor U8051 (N_8051,N_7468,N_5704);
xor U8052 (N_8052,N_6223,N_5266);
and U8053 (N_8053,N_6079,N_6448);
or U8054 (N_8054,N_7064,N_6939);
nand U8055 (N_8055,N_6499,N_7116);
and U8056 (N_8056,N_6782,N_6796);
nor U8057 (N_8057,N_6230,N_6134);
nand U8058 (N_8058,N_7159,N_5825);
nand U8059 (N_8059,N_5764,N_7156);
xor U8060 (N_8060,N_5152,N_6972);
and U8061 (N_8061,N_6309,N_5024);
nand U8062 (N_8062,N_6011,N_7437);
and U8063 (N_8063,N_6440,N_7020);
xor U8064 (N_8064,N_6393,N_7365);
xor U8065 (N_8065,N_5160,N_5136);
xor U8066 (N_8066,N_5503,N_5751);
xnor U8067 (N_8067,N_6166,N_5249);
and U8068 (N_8068,N_6234,N_5879);
nand U8069 (N_8069,N_5230,N_6101);
and U8070 (N_8070,N_5524,N_6475);
and U8071 (N_8071,N_6070,N_5019);
nand U8072 (N_8072,N_6119,N_6543);
xor U8073 (N_8073,N_5137,N_6549);
or U8074 (N_8074,N_7023,N_5567);
nor U8075 (N_8075,N_6491,N_6869);
or U8076 (N_8076,N_5919,N_7275);
nand U8077 (N_8077,N_6676,N_6975);
nand U8078 (N_8078,N_7395,N_5637);
or U8079 (N_8079,N_6379,N_6859);
xnor U8080 (N_8080,N_5691,N_6531);
or U8081 (N_8081,N_7362,N_6651);
nand U8082 (N_8082,N_5663,N_6565);
nand U8083 (N_8083,N_6383,N_5241);
nand U8084 (N_8084,N_5029,N_6818);
nand U8085 (N_8085,N_5871,N_6537);
and U8086 (N_8086,N_5162,N_5054);
nor U8087 (N_8087,N_6148,N_6127);
nor U8088 (N_8088,N_5834,N_6320);
or U8089 (N_8089,N_6361,N_5895);
nand U8090 (N_8090,N_6853,N_5067);
and U8091 (N_8091,N_6709,N_6073);
nand U8092 (N_8092,N_5619,N_5482);
or U8093 (N_8093,N_6680,N_6574);
nand U8094 (N_8094,N_7212,N_6150);
xor U8095 (N_8095,N_5714,N_5713);
nor U8096 (N_8096,N_5452,N_6251);
nor U8097 (N_8097,N_7120,N_6005);
xor U8098 (N_8098,N_5956,N_5794);
and U8099 (N_8099,N_6015,N_5431);
nand U8100 (N_8100,N_5244,N_6744);
and U8101 (N_8101,N_6881,N_6792);
nor U8102 (N_8102,N_5037,N_7332);
nor U8103 (N_8103,N_7398,N_6211);
xor U8104 (N_8104,N_7307,N_6078);
nand U8105 (N_8105,N_7443,N_5544);
nand U8106 (N_8106,N_5474,N_7114);
nand U8107 (N_8107,N_5416,N_6930);
and U8108 (N_8108,N_5171,N_6888);
or U8109 (N_8109,N_5812,N_6075);
or U8110 (N_8110,N_5723,N_7488);
xor U8111 (N_8111,N_7104,N_6633);
nand U8112 (N_8112,N_5470,N_7035);
and U8113 (N_8113,N_7387,N_5101);
xor U8114 (N_8114,N_6902,N_6920);
and U8115 (N_8115,N_5598,N_7341);
or U8116 (N_8116,N_7426,N_6290);
and U8117 (N_8117,N_5886,N_5718);
nor U8118 (N_8118,N_5954,N_5974);
nor U8119 (N_8119,N_5981,N_5724);
or U8120 (N_8120,N_6176,N_6312);
or U8121 (N_8121,N_7272,N_6927);
nand U8122 (N_8122,N_5865,N_6566);
and U8123 (N_8123,N_7232,N_5290);
xor U8124 (N_8124,N_6998,N_5675);
xor U8125 (N_8125,N_6940,N_6731);
nor U8126 (N_8126,N_7208,N_7048);
nor U8127 (N_8127,N_5210,N_6842);
nor U8128 (N_8128,N_5715,N_6947);
nor U8129 (N_8129,N_5108,N_6411);
nor U8130 (N_8130,N_7227,N_5749);
xor U8131 (N_8131,N_6500,N_5636);
xnor U8132 (N_8132,N_5635,N_5810);
nand U8133 (N_8133,N_7202,N_7439);
nor U8134 (N_8134,N_7172,N_7017);
or U8135 (N_8135,N_7355,N_5711);
and U8136 (N_8136,N_6687,N_7211);
nor U8137 (N_8137,N_5061,N_7068);
xnor U8138 (N_8138,N_6806,N_6040);
nand U8139 (N_8139,N_6544,N_7442);
xor U8140 (N_8140,N_5382,N_7032);
xnor U8141 (N_8141,N_6479,N_6749);
and U8142 (N_8142,N_5166,N_6951);
or U8143 (N_8143,N_5776,N_6267);
and U8144 (N_8144,N_7361,N_5611);
nor U8145 (N_8145,N_5686,N_6220);
xnor U8146 (N_8146,N_5020,N_6539);
nand U8147 (N_8147,N_7250,N_6252);
xor U8148 (N_8148,N_7431,N_6086);
xor U8149 (N_8149,N_6556,N_5651);
or U8150 (N_8150,N_7209,N_6068);
nor U8151 (N_8151,N_5618,N_7067);
nor U8152 (N_8152,N_7155,N_7237);
nor U8153 (N_8153,N_5788,N_6003);
nor U8154 (N_8154,N_7356,N_5972);
nand U8155 (N_8155,N_7352,N_5549);
nand U8156 (N_8156,N_7222,N_6553);
or U8157 (N_8157,N_5756,N_7196);
nor U8158 (N_8158,N_5089,N_5388);
nor U8159 (N_8159,N_6598,N_5196);
and U8160 (N_8160,N_6206,N_5483);
nand U8161 (N_8161,N_6983,N_5736);
and U8162 (N_8162,N_5518,N_6254);
or U8163 (N_8163,N_7489,N_6468);
nor U8164 (N_8164,N_7065,N_5863);
nor U8165 (N_8165,N_7405,N_5752);
and U8166 (N_8166,N_5664,N_6164);
or U8167 (N_8167,N_5667,N_5116);
and U8168 (N_8168,N_5779,N_5385);
xor U8169 (N_8169,N_6661,N_5310);
nand U8170 (N_8170,N_5626,N_6600);
xor U8171 (N_8171,N_6799,N_5215);
nand U8172 (N_8172,N_5828,N_5529);
or U8173 (N_8173,N_6858,N_5348);
and U8174 (N_8174,N_6618,N_7194);
xnor U8175 (N_8175,N_5787,N_7412);
nor U8176 (N_8176,N_6194,N_5224);
and U8177 (N_8177,N_5141,N_5617);
nand U8178 (N_8178,N_5578,N_7197);
nor U8179 (N_8179,N_5278,N_7003);
nand U8180 (N_8180,N_6523,N_5398);
nor U8181 (N_8181,N_7247,N_6696);
or U8182 (N_8182,N_5313,N_5167);
xnor U8183 (N_8183,N_5432,N_5780);
nor U8184 (N_8184,N_6935,N_6490);
nor U8185 (N_8185,N_5314,N_5078);
xor U8186 (N_8186,N_7363,N_5394);
xor U8187 (N_8187,N_5920,N_6199);
nor U8188 (N_8188,N_6665,N_6304);
nand U8189 (N_8189,N_5823,N_6161);
nor U8190 (N_8190,N_5493,N_7174);
or U8191 (N_8191,N_6179,N_6132);
nand U8192 (N_8192,N_6978,N_5356);
and U8193 (N_8193,N_5326,N_7497);
nor U8194 (N_8194,N_5487,N_5629);
or U8195 (N_8195,N_6833,N_5579);
or U8196 (N_8196,N_5156,N_6506);
nand U8197 (N_8197,N_6570,N_6572);
or U8198 (N_8198,N_5861,N_6036);
nand U8199 (N_8199,N_5288,N_5086);
nor U8200 (N_8200,N_5247,N_6237);
or U8201 (N_8201,N_6326,N_6821);
or U8202 (N_8202,N_6472,N_5702);
xor U8203 (N_8203,N_5491,N_6836);
and U8204 (N_8204,N_5188,N_7047);
and U8205 (N_8205,N_6807,N_6046);
nand U8206 (N_8206,N_6392,N_5507);
nor U8207 (N_8207,N_6105,N_5039);
nand U8208 (N_8208,N_6759,N_5908);
nand U8209 (N_8209,N_6060,N_5332);
or U8210 (N_8210,N_6895,N_6401);
xor U8211 (N_8211,N_7013,N_5275);
nor U8212 (N_8212,N_5943,N_6726);
nand U8213 (N_8213,N_5646,N_6387);
and U8214 (N_8214,N_5890,N_5352);
and U8215 (N_8215,N_5254,N_5296);
nand U8216 (N_8216,N_6748,N_6093);
nor U8217 (N_8217,N_5025,N_5878);
nor U8218 (N_8218,N_7078,N_7271);
or U8219 (N_8219,N_7424,N_7256);
xor U8220 (N_8220,N_5852,N_5798);
nand U8221 (N_8221,N_6358,N_6757);
nor U8222 (N_8222,N_5708,N_6061);
xor U8223 (N_8223,N_5822,N_6885);
nand U8224 (N_8224,N_6985,N_7136);
nand U8225 (N_8225,N_6180,N_5811);
xnor U8226 (N_8226,N_6365,N_5323);
xnor U8227 (N_8227,N_6528,N_6331);
and U8228 (N_8228,N_6504,N_5447);
nand U8229 (N_8229,N_5058,N_7441);
and U8230 (N_8230,N_6418,N_5298);
or U8231 (N_8231,N_6767,N_6213);
or U8232 (N_8232,N_6315,N_5777);
xor U8233 (N_8233,N_6542,N_5548);
and U8234 (N_8234,N_6695,N_6189);
or U8235 (N_8235,N_5631,N_6204);
and U8236 (N_8236,N_7239,N_7057);
and U8237 (N_8237,N_5322,N_6412);
or U8238 (N_8238,N_6507,N_5429);
nor U8239 (N_8239,N_6289,N_6033);
and U8240 (N_8240,N_5519,N_5877);
nand U8241 (N_8241,N_5168,N_6386);
and U8242 (N_8242,N_5926,N_5557);
or U8243 (N_8243,N_6876,N_6302);
or U8244 (N_8244,N_7319,N_6167);
nand U8245 (N_8245,N_6727,N_5520);
nand U8246 (N_8246,N_5364,N_5624);
xor U8247 (N_8247,N_6221,N_5644);
or U8248 (N_8248,N_6812,N_6545);
nand U8249 (N_8249,N_6038,N_7262);
and U8250 (N_8250,N_6000,N_6612);
nand U8251 (N_8251,N_6258,N_6399);
xor U8252 (N_8252,N_7354,N_6679);
nand U8253 (N_8253,N_5124,N_6238);
xor U8254 (N_8254,N_5676,N_5816);
and U8255 (N_8255,N_5970,N_5896);
nor U8256 (N_8256,N_7305,N_7217);
and U8257 (N_8257,N_5022,N_5412);
nor U8258 (N_8258,N_7263,N_6266);
nor U8259 (N_8259,N_6861,N_5095);
or U8260 (N_8260,N_5370,N_7110);
xnor U8261 (N_8261,N_6395,N_5103);
nand U8262 (N_8262,N_5501,N_5551);
nand U8263 (N_8263,N_7278,N_7460);
and U8264 (N_8264,N_5889,N_6828);
xnor U8265 (N_8265,N_5754,N_5965);
and U8266 (N_8266,N_6655,N_5534);
nor U8267 (N_8267,N_5436,N_6405);
nor U8268 (N_8268,N_6996,N_5396);
nand U8269 (N_8269,N_5170,N_6384);
and U8270 (N_8270,N_6215,N_6925);
and U8271 (N_8271,N_5042,N_5940);
nand U8272 (N_8272,N_6789,N_5289);
xnor U8273 (N_8273,N_7333,N_7108);
nand U8274 (N_8274,N_6210,N_5032);
nand U8275 (N_8275,N_6512,N_6910);
xnor U8276 (N_8276,N_6762,N_5492);
xor U8277 (N_8277,N_5361,N_6074);
and U8278 (N_8278,N_6708,N_5735);
or U8279 (N_8279,N_5745,N_6898);
nor U8280 (N_8280,N_5771,N_5740);
and U8281 (N_8281,N_6049,N_6338);
or U8282 (N_8282,N_7314,N_5696);
nor U8283 (N_8283,N_6041,N_6438);
nor U8284 (N_8284,N_5438,N_6430);
nor U8285 (N_8285,N_6006,N_7167);
or U8286 (N_8286,N_7230,N_5325);
or U8287 (N_8287,N_7129,N_6887);
or U8288 (N_8288,N_6280,N_5050);
xor U8289 (N_8289,N_6577,N_6990);
nand U8290 (N_8290,N_5218,N_5031);
or U8291 (N_8291,N_6239,N_5572);
or U8292 (N_8292,N_6908,N_6730);
nor U8293 (N_8293,N_7414,N_5276);
and U8294 (N_8294,N_7490,N_5043);
and U8295 (N_8295,N_6592,N_7228);
nor U8296 (N_8296,N_5273,N_7076);
xor U8297 (N_8297,N_5084,N_7163);
xor U8298 (N_8298,N_7063,N_6979);
xor U8299 (N_8299,N_5987,N_6467);
nand U8300 (N_8300,N_6899,N_5577);
nand U8301 (N_8301,N_6558,N_5100);
xnor U8302 (N_8302,N_7283,N_7486);
nand U8303 (N_8303,N_7373,N_5051);
or U8304 (N_8304,N_6103,N_5964);
xor U8305 (N_8305,N_6112,N_7408);
nor U8306 (N_8306,N_5951,N_6059);
and U8307 (N_8307,N_5868,N_7320);
or U8308 (N_8308,N_5584,N_6421);
nand U8309 (N_8309,N_6865,N_5742);
nor U8310 (N_8310,N_6397,N_5918);
nand U8311 (N_8311,N_6901,N_5757);
nor U8312 (N_8312,N_7473,N_6916);
xnor U8313 (N_8313,N_6623,N_7180);
and U8314 (N_8314,N_7304,N_5155);
and U8315 (N_8315,N_5894,N_6964);
and U8316 (N_8316,N_7056,N_5268);
and U8317 (N_8317,N_5299,N_7203);
or U8318 (N_8318,N_6857,N_5679);
and U8319 (N_8319,N_5599,N_7031);
nand U8320 (N_8320,N_6875,N_5064);
nor U8321 (N_8321,N_6794,N_5768);
nor U8322 (N_8322,N_5395,N_6742);
xnor U8323 (N_8323,N_6724,N_5169);
nor U8324 (N_8324,N_6864,N_5400);
and U8325 (N_8325,N_5369,N_7224);
or U8326 (N_8326,N_7170,N_5991);
and U8327 (N_8327,N_5978,N_6109);
and U8328 (N_8328,N_5133,N_5142);
nand U8329 (N_8329,N_6950,N_6295);
or U8330 (N_8330,N_7306,N_5430);
and U8331 (N_8331,N_6973,N_6780);
nor U8332 (N_8332,N_6688,N_6129);
nor U8333 (N_8333,N_6158,N_5512);
and U8334 (N_8334,N_6745,N_6534);
nor U8335 (N_8335,N_5163,N_7128);
xor U8336 (N_8336,N_6952,N_6034);
nor U8337 (N_8337,N_5203,N_6571);
nand U8338 (N_8338,N_5389,N_5832);
nand U8339 (N_8339,N_6341,N_6434);
and U8340 (N_8340,N_7021,N_7150);
nor U8341 (N_8341,N_6098,N_6350);
nor U8342 (N_8342,N_6515,N_7375);
xnor U8343 (N_8343,N_6928,N_7113);
xor U8344 (N_8344,N_6482,N_7364);
or U8345 (N_8345,N_5187,N_6231);
and U8346 (N_8346,N_5647,N_6639);
nand U8347 (N_8347,N_6037,N_6294);
or U8348 (N_8348,N_6717,N_5048);
or U8349 (N_8349,N_7474,N_6890);
or U8350 (N_8350,N_6722,N_5437);
xor U8351 (N_8351,N_6897,N_7179);
nor U8352 (N_8352,N_5081,N_7465);
xor U8353 (N_8353,N_5453,N_5328);
and U8354 (N_8354,N_5778,N_6948);
and U8355 (N_8355,N_6645,N_5955);
nor U8356 (N_8356,N_6087,N_5330);
or U8357 (N_8357,N_7496,N_5570);
nor U8358 (N_8358,N_6124,N_5263);
nand U8359 (N_8359,N_5849,N_5107);
or U8360 (N_8360,N_6487,N_5892);
nor U8361 (N_8361,N_7204,N_6628);
nand U8362 (N_8362,N_6159,N_5204);
and U8363 (N_8363,N_6156,N_6957);
or U8364 (N_8364,N_5023,N_5269);
xnor U8365 (N_8365,N_5655,N_5563);
nor U8366 (N_8366,N_5839,N_5979);
or U8367 (N_8367,N_5576,N_6133);
and U8368 (N_8368,N_5582,N_7134);
nor U8369 (N_8369,N_6965,N_5831);
or U8370 (N_8370,N_5564,N_6720);
and U8371 (N_8371,N_5147,N_6492);
or U8372 (N_8372,N_6344,N_5658);
nor U8373 (N_8373,N_5614,N_6685);
and U8374 (N_8374,N_5993,N_6278);
xnor U8375 (N_8375,N_5426,N_5111);
nor U8376 (N_8376,N_5904,N_7483);
nand U8377 (N_8377,N_7402,N_7480);
or U8378 (N_8378,N_6268,N_5347);
xnor U8379 (N_8379,N_7329,N_6954);
or U8380 (N_8380,N_5113,N_5041);
and U8381 (N_8381,N_7210,N_6805);
and U8382 (N_8382,N_5568,N_7285);
nand U8383 (N_8383,N_7125,N_6672);
nand U8384 (N_8384,N_6153,N_6903);
nand U8385 (N_8385,N_6192,N_6131);
nor U8386 (N_8386,N_7334,N_5952);
nor U8387 (N_8387,N_6814,N_5835);
nor U8388 (N_8388,N_5052,N_6262);
xor U8389 (N_8389,N_6346,N_5383);
and U8390 (N_8390,N_7407,N_6373);
xor U8391 (N_8391,N_6788,N_5102);
and U8392 (N_8392,N_6408,N_5444);
nor U8393 (N_8393,N_6741,N_5591);
or U8394 (N_8394,N_5329,N_6498);
nor U8395 (N_8395,N_7433,N_7133);
xor U8396 (N_8396,N_5893,N_5446);
nand U8397 (N_8397,N_5294,N_5678);
and U8398 (N_8398,N_7216,N_6735);
nor U8399 (N_8399,N_7372,N_7220);
and U8400 (N_8400,N_6139,N_7185);
nand U8401 (N_8401,N_5413,N_7484);
and U8402 (N_8402,N_6172,N_6114);
nand U8403 (N_8403,N_6795,N_6363);
nand U8404 (N_8404,N_5265,N_5406);
xnor U8405 (N_8405,N_5760,N_6775);
nand U8406 (N_8406,N_6588,N_5443);
nand U8407 (N_8407,N_5627,N_7438);
xnor U8408 (N_8408,N_5766,N_6205);
nor U8409 (N_8409,N_6117,N_7336);
and U8410 (N_8410,N_5175,N_5057);
nand U8411 (N_8411,N_6147,N_5674);
xnor U8412 (N_8412,N_6410,N_5642);
nor U8413 (N_8413,N_6733,N_6450);
nand U8414 (N_8414,N_7323,N_6919);
and U8415 (N_8415,N_5442,N_6868);
nand U8416 (N_8416,N_6351,N_5223);
or U8417 (N_8417,N_6359,N_5494);
or U8418 (N_8418,N_6980,N_5357);
nand U8419 (N_8419,N_6768,N_5744);
or U8420 (N_8420,N_5808,N_6327);
xor U8421 (N_8421,N_7236,N_6582);
or U8422 (N_8422,N_6347,N_5985);
or U8423 (N_8423,N_6165,N_5856);
xnor U8424 (N_8424,N_7148,N_5554);
nand U8425 (N_8425,N_7050,N_5984);
nor U8426 (N_8426,N_7303,N_5201);
or U8427 (N_8427,N_6607,N_6993);
nor U8428 (N_8428,N_6992,N_5477);
or U8429 (N_8429,N_6265,N_6191);
xor U8430 (N_8430,N_6157,N_5182);
nor U8431 (N_8431,N_5153,N_6718);
nand U8432 (N_8432,N_6201,N_6747);
nor U8433 (N_8433,N_6396,N_7260);
and U8434 (N_8434,N_5990,N_6480);
nand U8435 (N_8435,N_5250,N_7339);
xnor U8436 (N_8436,N_7321,N_6137);
and U8437 (N_8437,N_5945,N_6288);
or U8438 (N_8438,N_5681,N_6065);
xnor U8439 (N_8439,N_7429,N_6617);
xnor U8440 (N_8440,N_6058,N_7010);
and U8441 (N_8441,N_5767,N_5174);
nor U8442 (N_8442,N_6848,N_6779);
nand U8443 (N_8443,N_7053,N_6064);
nor U8444 (N_8444,N_5960,N_7191);
nor U8445 (N_8445,N_7186,N_6193);
xor U8446 (N_8446,N_5109,N_6834);
nor U8447 (N_8447,N_5924,N_6568);
and U8448 (N_8448,N_5144,N_6585);
or U8449 (N_8449,N_7117,N_5207);
nor U8450 (N_8450,N_5532,N_6286);
and U8451 (N_8451,N_6067,N_6790);
nand U8452 (N_8452,N_6417,N_5264);
and U8453 (N_8453,N_7000,N_6678);
nor U8454 (N_8454,N_6052,N_5587);
or U8455 (N_8455,N_5774,N_6435);
nand U8456 (N_8456,N_5457,N_7090);
and U8457 (N_8457,N_5225,N_5038);
or U8458 (N_8458,N_5319,N_6774);
xor U8459 (N_8459,N_5387,N_6437);
xor U8460 (N_8460,N_5854,N_5105);
and U8461 (N_8461,N_5709,N_5090);
xnor U8462 (N_8462,N_6704,N_6516);
or U8463 (N_8463,N_6152,N_6031);
nor U8464 (N_8464,N_5080,N_7132);
nand U8465 (N_8465,N_5906,N_7096);
nor U8466 (N_8466,N_7376,N_5002);
or U8467 (N_8467,N_5211,N_6284);
or U8468 (N_8468,N_5891,N_5508);
nor U8469 (N_8469,N_6648,N_6815);
or U8470 (N_8470,N_7106,N_5701);
nor U8471 (N_8471,N_5523,N_5422);
xnor U8472 (N_8472,N_7142,N_6798);
nand U8473 (N_8473,N_6249,N_7470);
xnor U8474 (N_8474,N_5285,N_5983);
xnor U8475 (N_8475,N_6882,N_5380);
xor U8476 (N_8476,N_6292,N_7024);
nor U8477 (N_8477,N_6959,N_5036);
and U8478 (N_8478,N_5165,N_6924);
xor U8479 (N_8479,N_5561,N_6281);
and U8480 (N_8480,N_5930,N_5805);
nor U8481 (N_8481,N_6654,N_7312);
and U8482 (N_8482,N_5558,N_5410);
and U8483 (N_8483,N_6846,N_5645);
nor U8484 (N_8484,N_6750,N_7074);
and U8485 (N_8485,N_5151,N_6248);
xor U8486 (N_8486,N_6670,N_5866);
and U8487 (N_8487,N_7182,N_5998);
nor U8488 (N_8488,N_5763,N_7449);
xor U8489 (N_8489,N_6586,N_6804);
or U8490 (N_8490,N_5931,N_6943);
xnor U8491 (N_8491,N_5843,N_5351);
nand U8492 (N_8492,N_5044,N_6961);
and U8493 (N_8493,N_6453,N_7471);
nand U8494 (N_8494,N_5928,N_5625);
and U8495 (N_8495,N_6053,N_6488);
and U8496 (N_8496,N_6705,N_6080);
nand U8497 (N_8497,N_6956,N_6094);
and U8498 (N_8498,N_5467,N_5790);
or U8499 (N_8499,N_7326,N_7062);
nand U8500 (N_8500,N_5243,N_5793);
nor U8501 (N_8501,N_6301,N_6375);
nand U8502 (N_8502,N_7060,N_5820);
xor U8503 (N_8503,N_6224,N_7266);
nand U8504 (N_8504,N_5221,N_6781);
xnor U8505 (N_8505,N_5397,N_7112);
xor U8506 (N_8506,N_6051,N_6285);
nor U8507 (N_8507,N_5311,N_6629);
xnor U8508 (N_8508,N_6837,N_6108);
or U8509 (N_8509,N_5075,N_6510);
nand U8510 (N_8510,N_5304,N_5399);
nor U8511 (N_8511,N_7337,N_5353);
nand U8512 (N_8512,N_6023,N_7099);
and U8513 (N_8513,N_6374,N_6299);
xnor U8514 (N_8514,N_5700,N_6413);
nor U8515 (N_8515,N_5973,N_5053);
xor U8516 (N_8516,N_6505,N_5555);
xnor U8517 (N_8517,N_7400,N_5499);
nor U8518 (N_8518,N_6824,N_5065);
xor U8519 (N_8519,N_5826,N_6308);
and U8520 (N_8520,N_5110,N_5703);
and U8521 (N_8521,N_6548,N_6838);
nand U8522 (N_8522,N_7041,N_7040);
xor U8523 (N_8523,N_6088,N_6817);
nor U8524 (N_8524,N_5257,N_5157);
or U8525 (N_8525,N_6689,N_7421);
and U8526 (N_8526,N_6863,N_5939);
xor U8527 (N_8527,N_6968,N_5334);
or U8528 (N_8528,N_7435,N_6605);
nor U8529 (N_8529,N_6287,N_5659);
xor U8530 (N_8530,N_7052,N_6632);
xnor U8531 (N_8531,N_6826,N_7258);
xor U8532 (N_8532,N_5996,N_5748);
nor U8533 (N_8533,N_7233,N_6169);
and U8534 (N_8534,N_5641,N_6604);
or U8535 (N_8535,N_5946,N_6911);
or U8536 (N_8536,N_7007,N_6329);
and U8537 (N_8537,N_7464,N_6066);
nand U8538 (N_8538,N_6138,N_6390);
or U8539 (N_8539,N_6354,N_5818);
and U8540 (N_8540,N_6261,N_5302);
nor U8541 (N_8541,N_6106,N_5963);
nand U8542 (N_8542,N_5134,N_5797);
and U8543 (N_8543,N_6154,N_5071);
nor U8544 (N_8544,N_6988,N_5657);
xor U8545 (N_8545,N_6660,N_6524);
nor U8546 (N_8546,N_6275,N_5802);
or U8547 (N_8547,N_6325,N_6090);
nor U8548 (N_8548,N_5968,N_5588);
or U8549 (N_8549,N_6048,N_7051);
and U8550 (N_8550,N_5516,N_7160);
and U8551 (N_8551,N_6050,N_7459);
nand U8552 (N_8552,N_6594,N_6493);
and U8553 (N_8553,N_6062,N_5185);
xnor U8554 (N_8554,N_7411,N_5585);
nor U8555 (N_8555,N_5341,N_6376);
or U8556 (N_8556,N_6092,N_6877);
nand U8557 (N_8557,N_5245,N_6130);
or U8558 (N_8558,N_6277,N_7253);
xnor U8559 (N_8559,N_6918,N_6316);
nand U8560 (N_8560,N_5537,N_5088);
and U8561 (N_8561,N_5565,N_7144);
and U8562 (N_8562,N_6208,N_7213);
nand U8563 (N_8563,N_5743,N_5480);
xnor U8564 (N_8564,N_6514,N_6163);
nand U8565 (N_8565,N_5070,N_5213);
xor U8566 (N_8566,N_5594,N_6160);
and U8567 (N_8567,N_6698,N_6915);
xnor U8568 (N_8568,N_6214,N_6554);
xnor U8569 (N_8569,N_6707,N_7423);
or U8570 (N_8570,N_7345,N_6155);
or U8571 (N_8571,N_5427,N_7276);
and U8572 (N_8572,N_5804,N_6614);
and U8573 (N_8573,N_5622,N_6332);
nand U8574 (N_8574,N_6874,N_7296);
xor U8575 (N_8575,N_5027,N_5186);
and U8576 (N_8576,N_5590,N_7404);
or U8577 (N_8577,N_5267,N_5403);
nand U8578 (N_8578,N_7281,N_6681);
xor U8579 (N_8579,N_6711,N_5910);
and U8580 (N_8580,N_6896,N_6415);
nor U8581 (N_8581,N_5121,N_6174);
nor U8582 (N_8582,N_6870,N_6765);
and U8583 (N_8583,N_6995,N_5509);
or U8584 (N_8584,N_5062,N_6521);
nor U8585 (N_8585,N_6306,N_5158);
nand U8586 (N_8586,N_7330,N_6609);
xor U8587 (N_8587,N_6517,N_5321);
nand U8588 (N_8588,N_7100,N_6893);
and U8589 (N_8589,N_6269,N_6102);
nand U8590 (N_8590,N_6984,N_7393);
or U8591 (N_8591,N_6526,N_5864);
or U8592 (N_8592,N_5729,N_5761);
nand U8593 (N_8593,N_5783,N_7177);
or U8594 (N_8594,N_5634,N_5293);
xor U8595 (N_8595,N_5173,N_5359);
and U8596 (N_8596,N_5581,N_6402);
nand U8597 (N_8597,N_6279,N_5172);
nor U8598 (N_8598,N_5762,N_5260);
nand U8599 (N_8599,N_5358,N_6462);
nor U8600 (N_8600,N_6625,N_5220);
and U8601 (N_8601,N_5734,N_5272);
nor U8602 (N_8602,N_6936,N_6378);
nor U8603 (N_8603,N_5346,N_6626);
or U8604 (N_8604,N_6729,N_6307);
or U8605 (N_8605,N_6966,N_6081);
xnor U8606 (N_8606,N_5016,N_6754);
xor U8607 (N_8607,N_5612,N_5789);
and U8608 (N_8608,N_6955,N_7403);
nand U8609 (N_8609,N_5504,N_7231);
nand U8610 (N_8610,N_6519,N_6569);
nor U8611 (N_8611,N_5307,N_6382);
and U8612 (N_8612,N_7409,N_6025);
nand U8613 (N_8613,N_7331,N_6414);
and U8614 (N_8614,N_5980,N_6371);
and U8615 (N_8615,N_7274,N_6427);
and U8616 (N_8616,N_6461,N_6270);
or U8617 (N_8617,N_6177,N_5421);
nor U8618 (N_8618,N_6575,N_6914);
and U8619 (N_8619,N_5874,N_5149);
nor U8620 (N_8620,N_6444,N_7169);
nor U8621 (N_8621,N_7046,N_6342);
nor U8622 (N_8622,N_5280,N_5717);
nand U8623 (N_8623,N_6330,N_6938);
nand U8624 (N_8624,N_6391,N_5545);
and U8625 (N_8625,N_7267,N_5556);
xnor U8626 (N_8626,N_5562,N_7043);
nand U8627 (N_8627,N_5428,N_6042);
and U8628 (N_8628,N_5666,N_6659);
nor U8629 (N_8629,N_5148,N_7016);
nor U8630 (N_8630,N_6255,N_7137);
nor U8631 (N_8631,N_5850,N_5082);
or U8632 (N_8632,N_6989,N_6082);
xor U8633 (N_8633,N_7199,N_6621);
and U8634 (N_8634,N_6772,N_7350);
and U8635 (N_8635,N_6580,N_7111);
and U8636 (N_8636,N_5846,N_6370);
and U8637 (N_8637,N_5390,N_5683);
xnor U8638 (N_8638,N_6894,N_6710);
or U8639 (N_8639,N_5315,N_5335);
or U8640 (N_8640,N_6832,N_7252);
nor U8641 (N_8641,N_7436,N_6012);
or U8642 (N_8642,N_6233,N_6311);
nor U8643 (N_8643,N_6784,N_5656);
and U8644 (N_8644,N_7299,N_7359);
and U8645 (N_8645,N_5303,N_7487);
nor U8646 (N_8646,N_7183,N_5553);
nor U8647 (N_8647,N_7126,N_7164);
nand U8648 (N_8648,N_5953,N_7300);
or U8649 (N_8649,N_6222,N_6590);
and U8650 (N_8650,N_7315,N_5150);
nand U8651 (N_8651,N_5566,N_6419);
nor U8652 (N_8652,N_7406,N_6321);
xor U8653 (N_8653,N_7002,N_6243);
and U8654 (N_8654,N_6225,N_7292);
and U8655 (N_8655,N_7176,N_6974);
xnor U8656 (N_8656,N_5367,N_6797);
xnor U8657 (N_8657,N_6463,N_7386);
and U8658 (N_8658,N_5097,N_6443);
xor U8659 (N_8659,N_7054,N_5819);
and U8660 (N_8660,N_7072,N_5085);
nor U8661 (N_8661,N_6381,N_6891);
nand U8662 (N_8662,N_5638,N_7450);
and U8663 (N_8663,N_5505,N_6013);
xor U8664 (N_8664,N_6142,N_6941);
and U8665 (N_8665,N_6400,N_5140);
nand U8666 (N_8666,N_5049,N_5104);
nand U8667 (N_8667,N_5191,N_5542);
xor U8668 (N_8668,N_7463,N_5901);
nor U8669 (N_8669,N_7254,N_6339);
nor U8670 (N_8670,N_7270,N_5440);
nand U8671 (N_8671,N_5362,N_6095);
or U8672 (N_8672,N_7399,N_6509);
nor U8673 (N_8673,N_5602,N_7494);
nand U8674 (N_8674,N_7381,N_7102);
and U8675 (N_8675,N_5455,N_5907);
xor U8676 (N_8676,N_5640,N_6145);
or U8677 (N_8677,N_6849,N_5795);
xnor U8678 (N_8678,N_6937,N_6218);
nand U8679 (N_8679,N_7083,N_6686);
nand U8680 (N_8680,N_7028,N_6738);
nor U8681 (N_8681,N_6967,N_6551);
nor U8682 (N_8682,N_6791,N_6298);
or U8683 (N_8683,N_5277,N_6486);
xor U8684 (N_8684,N_6913,N_6104);
and U8685 (N_8685,N_5164,N_5726);
nand U8686 (N_8686,N_5374,N_6513);
nor U8687 (N_8687,N_5801,N_7181);
or U8688 (N_8688,N_6398,N_5014);
xor U8689 (N_8689,N_7141,N_7153);
xnor U8690 (N_8690,N_5011,N_5233);
and U8691 (N_8691,N_5393,N_7214);
nand U8692 (N_8692,N_5384,N_6638);
or U8693 (N_8693,N_7447,N_5193);
nand U8694 (N_8694,N_5872,N_7119);
and U8695 (N_8695,N_5559,N_5741);
xnor U8696 (N_8696,N_6283,N_6010);
or U8697 (N_8697,N_5486,N_7042);
nand U8698 (N_8698,N_5921,N_6962);
xor U8699 (N_8699,N_5291,N_6253);
xnor U8700 (N_8700,N_6352,N_7255);
nor U8701 (N_8701,N_6550,N_5876);
or U8702 (N_8702,N_7318,N_5750);
nor U8703 (N_8703,N_6406,N_5925);
or U8704 (N_8704,N_6197,N_5177);
nor U8705 (N_8705,N_6273,N_7221);
and U8706 (N_8706,N_6353,N_5258);
xor U8707 (N_8707,N_5994,N_6469);
or U8708 (N_8708,N_6455,N_7005);
and U8709 (N_8709,N_5079,N_5183);
nand U8710 (N_8710,N_5550,N_5976);
or U8711 (N_8711,N_5982,N_5758);
or U8712 (N_8712,N_5317,N_5875);
nor U8713 (N_8713,N_6841,N_7298);
xnor U8714 (N_8714,N_6319,N_6084);
nand U8715 (N_8715,N_5066,N_5046);
or U8716 (N_8716,N_6446,N_5938);
and U8717 (N_8717,N_7093,N_6564);
nand U8718 (N_8718,N_5093,N_7293);
nor U8719 (N_8719,N_5775,N_5180);
nor U8720 (N_8720,N_5425,N_6525);
and U8721 (N_8721,N_6128,N_5231);
xnor U8722 (N_8722,N_5899,N_7458);
nand U8723 (N_8723,N_7282,N_5586);
nor U8724 (N_8724,N_6601,N_7367);
nand U8725 (N_8725,N_7479,N_6389);
or U8726 (N_8726,N_7243,N_6207);
or U8727 (N_8727,N_6355,N_5126);
nor U8728 (N_8728,N_6202,N_5936);
xnor U8729 (N_8729,N_6703,N_6820);
or U8730 (N_8730,N_6442,N_7245);
nor U8731 (N_8731,N_6063,N_7205);
nand U8732 (N_8732,N_6783,N_6684);
and U8733 (N_8733,N_5712,N_5498);
nand U8734 (N_8734,N_5971,N_7082);
xor U8735 (N_8735,N_7121,N_6905);
xnor U8736 (N_8736,N_6274,N_6144);
nor U8737 (N_8737,N_7379,N_7430);
xor U8738 (N_8738,N_5377,N_5235);
nor U8739 (N_8739,N_7070,N_6337);
xnor U8740 (N_8740,N_6716,N_7071);
and U8741 (N_8741,N_6441,N_5000);
nand U8742 (N_8742,N_6766,N_6333);
nand U8743 (N_8743,N_5680,N_6481);
nor U8744 (N_8744,N_7124,N_6587);
and U8745 (N_8745,N_5405,N_5305);
nand U8746 (N_8746,N_6631,N_6786);
or U8747 (N_8747,N_6118,N_6429);
and U8748 (N_8748,N_6146,N_7309);
nand U8749 (N_8749,N_5479,N_6714);
and U8750 (N_8750,N_5092,N_7188);
nor U8751 (N_8751,N_5117,N_6958);
and U8752 (N_8752,N_6949,N_5567);
nand U8753 (N_8753,N_5372,N_5778);
nand U8754 (N_8754,N_5965,N_5098);
nor U8755 (N_8755,N_6079,N_5436);
and U8756 (N_8756,N_6366,N_6761);
or U8757 (N_8757,N_7177,N_5670);
xor U8758 (N_8758,N_7176,N_5351);
and U8759 (N_8759,N_6686,N_5745);
and U8760 (N_8760,N_5713,N_7027);
xor U8761 (N_8761,N_7361,N_6281);
or U8762 (N_8762,N_5522,N_5794);
nor U8763 (N_8763,N_6834,N_6720);
nor U8764 (N_8764,N_6552,N_5401);
and U8765 (N_8765,N_7386,N_6342);
nor U8766 (N_8766,N_6752,N_7419);
nand U8767 (N_8767,N_6342,N_6627);
and U8768 (N_8768,N_6965,N_5048);
nor U8769 (N_8769,N_5809,N_6897);
nand U8770 (N_8770,N_6413,N_6285);
nand U8771 (N_8771,N_6176,N_6819);
nand U8772 (N_8772,N_6148,N_5510);
or U8773 (N_8773,N_6342,N_6753);
or U8774 (N_8774,N_6859,N_6671);
xor U8775 (N_8775,N_6649,N_7316);
and U8776 (N_8776,N_5702,N_6758);
nand U8777 (N_8777,N_6268,N_7074);
xor U8778 (N_8778,N_5718,N_5166);
xor U8779 (N_8779,N_5484,N_5009);
nor U8780 (N_8780,N_7265,N_6318);
and U8781 (N_8781,N_6577,N_5634);
or U8782 (N_8782,N_5098,N_6016);
and U8783 (N_8783,N_7220,N_6981);
nor U8784 (N_8784,N_5806,N_7202);
or U8785 (N_8785,N_5404,N_5438);
nand U8786 (N_8786,N_5885,N_6661);
or U8787 (N_8787,N_7359,N_6412);
xnor U8788 (N_8788,N_5692,N_6233);
nor U8789 (N_8789,N_5713,N_5667);
nor U8790 (N_8790,N_5809,N_5777);
nand U8791 (N_8791,N_6389,N_5515);
nor U8792 (N_8792,N_5900,N_6412);
and U8793 (N_8793,N_7333,N_6602);
or U8794 (N_8794,N_7034,N_6113);
xor U8795 (N_8795,N_5232,N_6110);
nand U8796 (N_8796,N_5191,N_6568);
nor U8797 (N_8797,N_6613,N_6746);
and U8798 (N_8798,N_7354,N_6967);
or U8799 (N_8799,N_5490,N_6399);
xnor U8800 (N_8800,N_6435,N_5309);
and U8801 (N_8801,N_6478,N_5092);
and U8802 (N_8802,N_6269,N_6394);
xnor U8803 (N_8803,N_5345,N_6095);
nand U8804 (N_8804,N_5755,N_5237);
nor U8805 (N_8805,N_6499,N_6023);
and U8806 (N_8806,N_6852,N_7106);
or U8807 (N_8807,N_5988,N_7172);
and U8808 (N_8808,N_5185,N_6587);
or U8809 (N_8809,N_7091,N_5658);
and U8810 (N_8810,N_6639,N_5401);
nor U8811 (N_8811,N_6443,N_5244);
or U8812 (N_8812,N_5590,N_5430);
or U8813 (N_8813,N_6046,N_5207);
and U8814 (N_8814,N_5891,N_5170);
xor U8815 (N_8815,N_6458,N_5221);
nand U8816 (N_8816,N_5595,N_6386);
or U8817 (N_8817,N_5032,N_7436);
and U8818 (N_8818,N_5033,N_5361);
or U8819 (N_8819,N_7241,N_6957);
or U8820 (N_8820,N_6117,N_5076);
or U8821 (N_8821,N_6719,N_5638);
xnor U8822 (N_8822,N_7227,N_5653);
nand U8823 (N_8823,N_5911,N_6801);
nand U8824 (N_8824,N_5892,N_7052);
nand U8825 (N_8825,N_7394,N_7457);
and U8826 (N_8826,N_5533,N_6326);
nand U8827 (N_8827,N_7083,N_5577);
nor U8828 (N_8828,N_7272,N_6231);
nor U8829 (N_8829,N_6018,N_6288);
or U8830 (N_8830,N_5668,N_5713);
xnor U8831 (N_8831,N_6432,N_5117);
or U8832 (N_8832,N_6036,N_6606);
and U8833 (N_8833,N_5646,N_6312);
and U8834 (N_8834,N_6984,N_5652);
or U8835 (N_8835,N_5736,N_5371);
and U8836 (N_8836,N_5337,N_5161);
nor U8837 (N_8837,N_5565,N_5773);
nor U8838 (N_8838,N_6553,N_5574);
and U8839 (N_8839,N_5798,N_6811);
and U8840 (N_8840,N_6143,N_5857);
nor U8841 (N_8841,N_5583,N_5832);
and U8842 (N_8842,N_7406,N_6171);
or U8843 (N_8843,N_6782,N_5013);
nor U8844 (N_8844,N_6172,N_6909);
and U8845 (N_8845,N_7154,N_5708);
or U8846 (N_8846,N_7004,N_5044);
and U8847 (N_8847,N_6679,N_7249);
xor U8848 (N_8848,N_6601,N_6409);
xnor U8849 (N_8849,N_6810,N_5322);
or U8850 (N_8850,N_6289,N_5605);
or U8851 (N_8851,N_5504,N_5790);
nor U8852 (N_8852,N_5680,N_7204);
and U8853 (N_8853,N_5871,N_5212);
and U8854 (N_8854,N_5776,N_5862);
or U8855 (N_8855,N_5199,N_7181);
nand U8856 (N_8856,N_6991,N_5686);
or U8857 (N_8857,N_7497,N_6464);
nor U8858 (N_8858,N_7085,N_5260);
and U8859 (N_8859,N_6558,N_6670);
or U8860 (N_8860,N_6940,N_5315);
nand U8861 (N_8861,N_5159,N_5740);
nand U8862 (N_8862,N_6687,N_5148);
xnor U8863 (N_8863,N_7117,N_5549);
nor U8864 (N_8864,N_5646,N_5813);
nand U8865 (N_8865,N_5231,N_6708);
and U8866 (N_8866,N_7273,N_5515);
nand U8867 (N_8867,N_6896,N_6568);
and U8868 (N_8868,N_6322,N_7034);
nor U8869 (N_8869,N_6868,N_6203);
or U8870 (N_8870,N_5353,N_5263);
and U8871 (N_8871,N_5727,N_7039);
nand U8872 (N_8872,N_5544,N_5423);
nor U8873 (N_8873,N_6333,N_5570);
or U8874 (N_8874,N_7464,N_6944);
or U8875 (N_8875,N_6163,N_7377);
nand U8876 (N_8876,N_5817,N_6790);
nor U8877 (N_8877,N_7090,N_5529);
and U8878 (N_8878,N_5082,N_5319);
nor U8879 (N_8879,N_7204,N_6723);
or U8880 (N_8880,N_5314,N_6724);
nor U8881 (N_8881,N_5017,N_5274);
nand U8882 (N_8882,N_7318,N_7453);
nand U8883 (N_8883,N_5645,N_5347);
xor U8884 (N_8884,N_5144,N_7011);
or U8885 (N_8885,N_6479,N_6118);
nor U8886 (N_8886,N_6735,N_5270);
nand U8887 (N_8887,N_7029,N_7169);
or U8888 (N_8888,N_5352,N_5471);
nor U8889 (N_8889,N_6566,N_5447);
or U8890 (N_8890,N_5351,N_5102);
and U8891 (N_8891,N_6711,N_7387);
and U8892 (N_8892,N_5970,N_5034);
and U8893 (N_8893,N_5874,N_7174);
or U8894 (N_8894,N_5800,N_7173);
nand U8895 (N_8895,N_7343,N_6230);
nand U8896 (N_8896,N_5861,N_5624);
nor U8897 (N_8897,N_7260,N_7255);
nand U8898 (N_8898,N_6154,N_5051);
nand U8899 (N_8899,N_7324,N_7179);
nor U8900 (N_8900,N_5609,N_6111);
nand U8901 (N_8901,N_5556,N_7439);
nor U8902 (N_8902,N_6535,N_7138);
and U8903 (N_8903,N_6880,N_7002);
xnor U8904 (N_8904,N_6192,N_6148);
nand U8905 (N_8905,N_6411,N_6508);
or U8906 (N_8906,N_7434,N_5148);
or U8907 (N_8907,N_6631,N_6648);
or U8908 (N_8908,N_6878,N_6177);
xnor U8909 (N_8909,N_7464,N_5355);
or U8910 (N_8910,N_5837,N_5261);
xnor U8911 (N_8911,N_5196,N_5174);
nand U8912 (N_8912,N_5741,N_6759);
xnor U8913 (N_8913,N_7414,N_7119);
nor U8914 (N_8914,N_6938,N_6987);
nor U8915 (N_8915,N_7299,N_7018);
nor U8916 (N_8916,N_6332,N_6538);
nand U8917 (N_8917,N_6805,N_6197);
and U8918 (N_8918,N_6625,N_5530);
nor U8919 (N_8919,N_6033,N_7144);
xnor U8920 (N_8920,N_5579,N_6397);
or U8921 (N_8921,N_7211,N_5236);
xnor U8922 (N_8922,N_7240,N_5000);
or U8923 (N_8923,N_5929,N_6188);
nor U8924 (N_8924,N_5522,N_7044);
and U8925 (N_8925,N_7188,N_6782);
nand U8926 (N_8926,N_5715,N_6501);
and U8927 (N_8927,N_5512,N_7086);
nor U8928 (N_8928,N_6246,N_6124);
xnor U8929 (N_8929,N_6671,N_5257);
or U8930 (N_8930,N_5651,N_7050);
or U8931 (N_8931,N_6792,N_7039);
nand U8932 (N_8932,N_6273,N_7138);
or U8933 (N_8933,N_6247,N_6638);
and U8934 (N_8934,N_5286,N_5859);
and U8935 (N_8935,N_6555,N_5658);
or U8936 (N_8936,N_6910,N_5826);
nor U8937 (N_8937,N_6113,N_6410);
or U8938 (N_8938,N_6311,N_5295);
and U8939 (N_8939,N_6146,N_5245);
nand U8940 (N_8940,N_6359,N_5193);
nand U8941 (N_8941,N_6225,N_7326);
or U8942 (N_8942,N_6987,N_7149);
nand U8943 (N_8943,N_5240,N_6856);
and U8944 (N_8944,N_6677,N_7145);
or U8945 (N_8945,N_6461,N_5829);
nor U8946 (N_8946,N_5900,N_7385);
or U8947 (N_8947,N_7362,N_5267);
and U8948 (N_8948,N_6631,N_5991);
or U8949 (N_8949,N_6953,N_6134);
nand U8950 (N_8950,N_5781,N_5616);
nand U8951 (N_8951,N_6091,N_7175);
nand U8952 (N_8952,N_5243,N_6061);
xor U8953 (N_8953,N_5438,N_7236);
or U8954 (N_8954,N_6565,N_7064);
nor U8955 (N_8955,N_5656,N_6762);
and U8956 (N_8956,N_6817,N_5553);
nand U8957 (N_8957,N_5217,N_7290);
or U8958 (N_8958,N_7397,N_6168);
or U8959 (N_8959,N_6034,N_6202);
nand U8960 (N_8960,N_5427,N_6847);
and U8961 (N_8961,N_5400,N_7261);
nor U8962 (N_8962,N_7204,N_7114);
and U8963 (N_8963,N_5540,N_6675);
or U8964 (N_8964,N_5457,N_5977);
xnor U8965 (N_8965,N_6202,N_7408);
nand U8966 (N_8966,N_6075,N_6701);
nand U8967 (N_8967,N_6062,N_6801);
and U8968 (N_8968,N_5846,N_6028);
or U8969 (N_8969,N_6424,N_5401);
or U8970 (N_8970,N_6480,N_6043);
or U8971 (N_8971,N_7369,N_6115);
xor U8972 (N_8972,N_6231,N_7028);
or U8973 (N_8973,N_7174,N_5668);
and U8974 (N_8974,N_6288,N_7061);
and U8975 (N_8975,N_6325,N_6024);
xor U8976 (N_8976,N_5234,N_6009);
nand U8977 (N_8977,N_6739,N_6699);
nand U8978 (N_8978,N_7042,N_5751);
or U8979 (N_8979,N_6951,N_5844);
nand U8980 (N_8980,N_5589,N_5537);
nor U8981 (N_8981,N_5089,N_6783);
or U8982 (N_8982,N_5351,N_6079);
xor U8983 (N_8983,N_7261,N_5933);
and U8984 (N_8984,N_7344,N_5276);
or U8985 (N_8985,N_5329,N_6559);
nor U8986 (N_8986,N_6022,N_5143);
nor U8987 (N_8987,N_6534,N_6476);
xnor U8988 (N_8988,N_5112,N_5467);
nand U8989 (N_8989,N_6663,N_6462);
nor U8990 (N_8990,N_6560,N_5325);
nor U8991 (N_8991,N_6951,N_6744);
nand U8992 (N_8992,N_6680,N_6185);
xnor U8993 (N_8993,N_5244,N_6278);
xnor U8994 (N_8994,N_6008,N_5964);
or U8995 (N_8995,N_5965,N_6407);
nor U8996 (N_8996,N_5257,N_7365);
and U8997 (N_8997,N_5141,N_5830);
xor U8998 (N_8998,N_6624,N_5637);
nand U8999 (N_8999,N_6031,N_5542);
nor U9000 (N_9000,N_6720,N_6263);
nand U9001 (N_9001,N_5322,N_6720);
nand U9002 (N_9002,N_5349,N_5170);
nand U9003 (N_9003,N_6865,N_5402);
nand U9004 (N_9004,N_6806,N_5429);
or U9005 (N_9005,N_7318,N_6390);
xor U9006 (N_9006,N_6929,N_5313);
nand U9007 (N_9007,N_6379,N_5157);
nand U9008 (N_9008,N_6991,N_5223);
or U9009 (N_9009,N_6630,N_5598);
nor U9010 (N_9010,N_6526,N_5883);
or U9011 (N_9011,N_6544,N_6240);
and U9012 (N_9012,N_5833,N_6445);
or U9013 (N_9013,N_5316,N_5936);
or U9014 (N_9014,N_6518,N_7383);
nor U9015 (N_9015,N_5582,N_6697);
nor U9016 (N_9016,N_5559,N_5854);
nand U9017 (N_9017,N_5115,N_6686);
or U9018 (N_9018,N_6653,N_5762);
xor U9019 (N_9019,N_6345,N_5013);
xor U9020 (N_9020,N_5395,N_5761);
and U9021 (N_9021,N_5715,N_6981);
or U9022 (N_9022,N_5155,N_5756);
or U9023 (N_9023,N_7368,N_7222);
or U9024 (N_9024,N_7275,N_5979);
or U9025 (N_9025,N_6549,N_5333);
nor U9026 (N_9026,N_5844,N_7034);
xor U9027 (N_9027,N_6308,N_5604);
nor U9028 (N_9028,N_6650,N_5966);
nor U9029 (N_9029,N_5446,N_7010);
and U9030 (N_9030,N_6764,N_7498);
xor U9031 (N_9031,N_6185,N_5515);
xnor U9032 (N_9032,N_5667,N_5320);
nor U9033 (N_9033,N_6164,N_6900);
nand U9034 (N_9034,N_6637,N_6655);
xnor U9035 (N_9035,N_5755,N_7245);
and U9036 (N_9036,N_7420,N_6751);
or U9037 (N_9037,N_7270,N_5626);
xnor U9038 (N_9038,N_6990,N_5047);
nand U9039 (N_9039,N_6672,N_5086);
nor U9040 (N_9040,N_7281,N_6678);
nand U9041 (N_9041,N_5220,N_6588);
nand U9042 (N_9042,N_6198,N_6965);
nand U9043 (N_9043,N_5129,N_5836);
nand U9044 (N_9044,N_6487,N_5978);
and U9045 (N_9045,N_6555,N_6608);
nand U9046 (N_9046,N_5903,N_5739);
nand U9047 (N_9047,N_7312,N_5789);
and U9048 (N_9048,N_5298,N_5418);
nor U9049 (N_9049,N_6785,N_5999);
xnor U9050 (N_9050,N_7242,N_6297);
nand U9051 (N_9051,N_5929,N_7136);
xor U9052 (N_9052,N_6774,N_6826);
and U9053 (N_9053,N_6745,N_5323);
and U9054 (N_9054,N_5728,N_7433);
or U9055 (N_9055,N_6066,N_7062);
and U9056 (N_9056,N_5091,N_6202);
and U9057 (N_9057,N_6905,N_6649);
or U9058 (N_9058,N_5739,N_6318);
or U9059 (N_9059,N_5312,N_7377);
or U9060 (N_9060,N_7025,N_5979);
nor U9061 (N_9061,N_7159,N_7298);
xor U9062 (N_9062,N_5070,N_5943);
xnor U9063 (N_9063,N_6301,N_5329);
and U9064 (N_9064,N_5737,N_6505);
and U9065 (N_9065,N_6475,N_5418);
xor U9066 (N_9066,N_6740,N_6327);
nor U9067 (N_9067,N_7390,N_6602);
nor U9068 (N_9068,N_6372,N_5353);
or U9069 (N_9069,N_6442,N_6474);
or U9070 (N_9070,N_6519,N_6525);
xor U9071 (N_9071,N_5691,N_5750);
nand U9072 (N_9072,N_7126,N_6041);
or U9073 (N_9073,N_6423,N_6583);
nor U9074 (N_9074,N_6822,N_6968);
and U9075 (N_9075,N_7232,N_5876);
nand U9076 (N_9076,N_5994,N_6760);
and U9077 (N_9077,N_5024,N_5702);
nor U9078 (N_9078,N_7423,N_5145);
or U9079 (N_9079,N_7308,N_5015);
xor U9080 (N_9080,N_5516,N_5244);
xor U9081 (N_9081,N_7406,N_6187);
xor U9082 (N_9082,N_6294,N_6972);
and U9083 (N_9083,N_5812,N_6337);
nor U9084 (N_9084,N_6309,N_6018);
or U9085 (N_9085,N_5986,N_5151);
or U9086 (N_9086,N_5253,N_7484);
nand U9087 (N_9087,N_5407,N_5695);
xnor U9088 (N_9088,N_6850,N_5243);
or U9089 (N_9089,N_6063,N_6751);
and U9090 (N_9090,N_7058,N_6095);
xnor U9091 (N_9091,N_6773,N_7266);
and U9092 (N_9092,N_6551,N_7200);
nand U9093 (N_9093,N_7240,N_5156);
and U9094 (N_9094,N_5162,N_7275);
xnor U9095 (N_9095,N_5404,N_5265);
xnor U9096 (N_9096,N_5143,N_6455);
and U9097 (N_9097,N_6017,N_6382);
and U9098 (N_9098,N_7342,N_6333);
nand U9099 (N_9099,N_6716,N_6005);
nor U9100 (N_9100,N_5670,N_6821);
or U9101 (N_9101,N_5852,N_5573);
nor U9102 (N_9102,N_7204,N_6428);
xnor U9103 (N_9103,N_6751,N_5237);
and U9104 (N_9104,N_6558,N_7316);
nand U9105 (N_9105,N_5488,N_7124);
and U9106 (N_9106,N_6352,N_5469);
nor U9107 (N_9107,N_6169,N_6636);
xnor U9108 (N_9108,N_6489,N_6983);
and U9109 (N_9109,N_5695,N_6491);
nor U9110 (N_9110,N_6292,N_7331);
nand U9111 (N_9111,N_6650,N_6945);
nand U9112 (N_9112,N_6611,N_5867);
nand U9113 (N_9113,N_6741,N_5473);
xor U9114 (N_9114,N_5832,N_5064);
xor U9115 (N_9115,N_6856,N_6699);
nor U9116 (N_9116,N_7432,N_5276);
and U9117 (N_9117,N_7107,N_6780);
nand U9118 (N_9118,N_5119,N_7489);
nand U9119 (N_9119,N_7099,N_5049);
or U9120 (N_9120,N_6928,N_5208);
xor U9121 (N_9121,N_7419,N_6097);
or U9122 (N_9122,N_7035,N_5283);
or U9123 (N_9123,N_5120,N_5956);
nor U9124 (N_9124,N_5939,N_6898);
nand U9125 (N_9125,N_6487,N_6357);
nand U9126 (N_9126,N_6686,N_6261);
nor U9127 (N_9127,N_5827,N_6422);
or U9128 (N_9128,N_7233,N_6172);
xnor U9129 (N_9129,N_6585,N_6989);
or U9130 (N_9130,N_6261,N_7103);
xnor U9131 (N_9131,N_6110,N_5940);
or U9132 (N_9132,N_6788,N_6786);
nand U9133 (N_9133,N_6901,N_7391);
or U9134 (N_9134,N_7441,N_6131);
xor U9135 (N_9135,N_7238,N_5277);
xor U9136 (N_9136,N_6044,N_5571);
or U9137 (N_9137,N_5193,N_5984);
nor U9138 (N_9138,N_5227,N_5104);
nor U9139 (N_9139,N_5130,N_6004);
xor U9140 (N_9140,N_5426,N_5171);
and U9141 (N_9141,N_5771,N_7032);
nand U9142 (N_9142,N_6442,N_5887);
xor U9143 (N_9143,N_6313,N_5033);
and U9144 (N_9144,N_6895,N_5116);
nor U9145 (N_9145,N_6876,N_6409);
or U9146 (N_9146,N_5347,N_5193);
xnor U9147 (N_9147,N_5102,N_5243);
or U9148 (N_9148,N_6900,N_6982);
nand U9149 (N_9149,N_7042,N_6084);
or U9150 (N_9150,N_6890,N_5875);
nand U9151 (N_9151,N_7179,N_7268);
or U9152 (N_9152,N_6391,N_6919);
nor U9153 (N_9153,N_7045,N_6040);
or U9154 (N_9154,N_6095,N_5288);
and U9155 (N_9155,N_5974,N_5461);
nor U9156 (N_9156,N_5392,N_6255);
nand U9157 (N_9157,N_5886,N_6550);
nor U9158 (N_9158,N_5248,N_5801);
or U9159 (N_9159,N_5239,N_5057);
nand U9160 (N_9160,N_7411,N_5225);
nand U9161 (N_9161,N_6026,N_6053);
nand U9162 (N_9162,N_6636,N_5706);
and U9163 (N_9163,N_6341,N_7158);
nand U9164 (N_9164,N_6696,N_6551);
nor U9165 (N_9165,N_5658,N_6164);
xnor U9166 (N_9166,N_5245,N_6122);
or U9167 (N_9167,N_5484,N_6977);
or U9168 (N_9168,N_6308,N_6117);
or U9169 (N_9169,N_5455,N_6718);
xnor U9170 (N_9170,N_6480,N_6688);
nor U9171 (N_9171,N_6982,N_6446);
or U9172 (N_9172,N_6027,N_7238);
and U9173 (N_9173,N_5361,N_5836);
nor U9174 (N_9174,N_7369,N_6704);
nand U9175 (N_9175,N_5636,N_6711);
nor U9176 (N_9176,N_6082,N_6916);
nor U9177 (N_9177,N_5041,N_7213);
xor U9178 (N_9178,N_6855,N_5437);
nand U9179 (N_9179,N_5856,N_5582);
nand U9180 (N_9180,N_6227,N_6735);
nand U9181 (N_9181,N_6374,N_7125);
nor U9182 (N_9182,N_5585,N_5954);
xor U9183 (N_9183,N_7245,N_6970);
nand U9184 (N_9184,N_5470,N_6454);
nand U9185 (N_9185,N_7221,N_5497);
or U9186 (N_9186,N_7219,N_7206);
xor U9187 (N_9187,N_5039,N_5433);
or U9188 (N_9188,N_5527,N_5070);
or U9189 (N_9189,N_6851,N_6219);
nor U9190 (N_9190,N_5394,N_7301);
nor U9191 (N_9191,N_5085,N_6837);
xor U9192 (N_9192,N_6182,N_5845);
nor U9193 (N_9193,N_5081,N_5496);
and U9194 (N_9194,N_5366,N_6122);
and U9195 (N_9195,N_6353,N_6318);
xnor U9196 (N_9196,N_6668,N_5234);
nor U9197 (N_9197,N_6743,N_6578);
and U9198 (N_9198,N_6702,N_6562);
and U9199 (N_9199,N_5299,N_5956);
nand U9200 (N_9200,N_7075,N_5441);
or U9201 (N_9201,N_5929,N_7040);
xor U9202 (N_9202,N_5647,N_6815);
and U9203 (N_9203,N_6066,N_7048);
and U9204 (N_9204,N_6417,N_6859);
and U9205 (N_9205,N_5886,N_6252);
and U9206 (N_9206,N_5452,N_5678);
nor U9207 (N_9207,N_7031,N_5141);
nand U9208 (N_9208,N_5672,N_6818);
and U9209 (N_9209,N_6869,N_6794);
nor U9210 (N_9210,N_5912,N_6792);
and U9211 (N_9211,N_5357,N_6692);
nand U9212 (N_9212,N_7345,N_7442);
xnor U9213 (N_9213,N_6805,N_6160);
or U9214 (N_9214,N_5090,N_5365);
and U9215 (N_9215,N_6241,N_6610);
nand U9216 (N_9216,N_7112,N_6930);
nand U9217 (N_9217,N_6985,N_6132);
and U9218 (N_9218,N_6611,N_6574);
or U9219 (N_9219,N_6049,N_5171);
xor U9220 (N_9220,N_5568,N_6953);
nor U9221 (N_9221,N_6721,N_5903);
or U9222 (N_9222,N_5504,N_5179);
and U9223 (N_9223,N_7158,N_5313);
nor U9224 (N_9224,N_5973,N_5577);
nor U9225 (N_9225,N_5219,N_6332);
nor U9226 (N_9226,N_6450,N_6318);
nor U9227 (N_9227,N_5492,N_5881);
or U9228 (N_9228,N_5377,N_7094);
nand U9229 (N_9229,N_7259,N_5462);
and U9230 (N_9230,N_6669,N_7285);
nand U9231 (N_9231,N_5529,N_6254);
and U9232 (N_9232,N_5545,N_5684);
nand U9233 (N_9233,N_6623,N_7402);
or U9234 (N_9234,N_6486,N_6473);
nand U9235 (N_9235,N_5734,N_6612);
nor U9236 (N_9236,N_6015,N_5457);
nand U9237 (N_9237,N_6876,N_6022);
nand U9238 (N_9238,N_6331,N_5837);
xnor U9239 (N_9239,N_6888,N_5810);
and U9240 (N_9240,N_7470,N_6906);
or U9241 (N_9241,N_5068,N_5212);
or U9242 (N_9242,N_6451,N_6985);
and U9243 (N_9243,N_5639,N_5018);
nand U9244 (N_9244,N_5367,N_6272);
or U9245 (N_9245,N_5751,N_5907);
nand U9246 (N_9246,N_7194,N_5224);
and U9247 (N_9247,N_6159,N_5721);
nand U9248 (N_9248,N_7170,N_5603);
nand U9249 (N_9249,N_5929,N_5347);
or U9250 (N_9250,N_5477,N_5604);
and U9251 (N_9251,N_5257,N_6846);
or U9252 (N_9252,N_6894,N_7182);
nor U9253 (N_9253,N_5076,N_6872);
or U9254 (N_9254,N_7251,N_6064);
nor U9255 (N_9255,N_5921,N_6444);
nor U9256 (N_9256,N_6325,N_6172);
xor U9257 (N_9257,N_6594,N_6958);
nor U9258 (N_9258,N_6366,N_5406);
or U9259 (N_9259,N_6366,N_5241);
nand U9260 (N_9260,N_7072,N_6664);
and U9261 (N_9261,N_5352,N_7197);
nor U9262 (N_9262,N_5723,N_6005);
and U9263 (N_9263,N_6185,N_5047);
and U9264 (N_9264,N_7063,N_6330);
nand U9265 (N_9265,N_5782,N_6174);
nor U9266 (N_9266,N_7068,N_5165);
nand U9267 (N_9267,N_5683,N_6583);
and U9268 (N_9268,N_7102,N_6618);
and U9269 (N_9269,N_6607,N_7214);
and U9270 (N_9270,N_7254,N_7490);
nand U9271 (N_9271,N_5822,N_5717);
nand U9272 (N_9272,N_5456,N_7484);
and U9273 (N_9273,N_5970,N_6895);
nand U9274 (N_9274,N_6231,N_7494);
nor U9275 (N_9275,N_5732,N_7101);
or U9276 (N_9276,N_7007,N_5625);
xor U9277 (N_9277,N_6000,N_7323);
nand U9278 (N_9278,N_6096,N_5942);
nand U9279 (N_9279,N_6308,N_5077);
xnor U9280 (N_9280,N_6183,N_7083);
or U9281 (N_9281,N_6211,N_6962);
or U9282 (N_9282,N_6169,N_6173);
nand U9283 (N_9283,N_7134,N_6193);
nand U9284 (N_9284,N_5154,N_5590);
nor U9285 (N_9285,N_6645,N_5011);
xnor U9286 (N_9286,N_6523,N_7139);
xnor U9287 (N_9287,N_6149,N_6031);
nand U9288 (N_9288,N_5793,N_6827);
and U9289 (N_9289,N_5293,N_7261);
nand U9290 (N_9290,N_5836,N_5118);
nand U9291 (N_9291,N_6125,N_6069);
or U9292 (N_9292,N_7123,N_6506);
nor U9293 (N_9293,N_6917,N_5323);
nand U9294 (N_9294,N_5591,N_5674);
nand U9295 (N_9295,N_7198,N_6421);
or U9296 (N_9296,N_6174,N_6587);
nand U9297 (N_9297,N_7431,N_5647);
nor U9298 (N_9298,N_5898,N_7398);
nor U9299 (N_9299,N_5842,N_7110);
nor U9300 (N_9300,N_6381,N_7425);
xnor U9301 (N_9301,N_7490,N_7170);
and U9302 (N_9302,N_7297,N_5410);
or U9303 (N_9303,N_6100,N_7487);
or U9304 (N_9304,N_6448,N_6951);
nand U9305 (N_9305,N_6320,N_6220);
and U9306 (N_9306,N_5245,N_5184);
xor U9307 (N_9307,N_5418,N_5856);
and U9308 (N_9308,N_5609,N_6449);
or U9309 (N_9309,N_5310,N_5920);
nor U9310 (N_9310,N_5163,N_5857);
or U9311 (N_9311,N_5017,N_5478);
and U9312 (N_9312,N_6743,N_6018);
and U9313 (N_9313,N_6199,N_6124);
nand U9314 (N_9314,N_5047,N_6174);
or U9315 (N_9315,N_7126,N_5616);
and U9316 (N_9316,N_6403,N_7398);
nand U9317 (N_9317,N_7091,N_6307);
nand U9318 (N_9318,N_5122,N_6441);
or U9319 (N_9319,N_6734,N_6969);
or U9320 (N_9320,N_5903,N_7321);
nand U9321 (N_9321,N_6926,N_5485);
and U9322 (N_9322,N_5910,N_7397);
xnor U9323 (N_9323,N_7427,N_5364);
and U9324 (N_9324,N_5459,N_7359);
or U9325 (N_9325,N_7211,N_6156);
and U9326 (N_9326,N_7477,N_7276);
or U9327 (N_9327,N_7153,N_5370);
nor U9328 (N_9328,N_5925,N_5544);
or U9329 (N_9329,N_6077,N_5583);
nor U9330 (N_9330,N_6503,N_6990);
and U9331 (N_9331,N_5368,N_5804);
and U9332 (N_9332,N_5389,N_6960);
nand U9333 (N_9333,N_5400,N_5795);
and U9334 (N_9334,N_7319,N_5605);
or U9335 (N_9335,N_6504,N_5317);
nor U9336 (N_9336,N_7261,N_5708);
or U9337 (N_9337,N_6178,N_6527);
xnor U9338 (N_9338,N_6481,N_5453);
or U9339 (N_9339,N_7266,N_5485);
nor U9340 (N_9340,N_6721,N_7357);
or U9341 (N_9341,N_6971,N_7007);
nor U9342 (N_9342,N_7364,N_7031);
nor U9343 (N_9343,N_5385,N_6306);
nor U9344 (N_9344,N_6926,N_5827);
or U9345 (N_9345,N_5106,N_5414);
xor U9346 (N_9346,N_5903,N_6223);
or U9347 (N_9347,N_6767,N_5935);
or U9348 (N_9348,N_5888,N_5953);
or U9349 (N_9349,N_6344,N_6651);
nor U9350 (N_9350,N_6300,N_5070);
or U9351 (N_9351,N_7101,N_6814);
xnor U9352 (N_9352,N_5966,N_7195);
xnor U9353 (N_9353,N_7000,N_5657);
xor U9354 (N_9354,N_5571,N_5166);
and U9355 (N_9355,N_5309,N_6018);
xnor U9356 (N_9356,N_5524,N_5681);
nor U9357 (N_9357,N_6188,N_5864);
nand U9358 (N_9358,N_5050,N_6550);
nand U9359 (N_9359,N_7234,N_6948);
nor U9360 (N_9360,N_6305,N_5691);
or U9361 (N_9361,N_6745,N_6842);
and U9362 (N_9362,N_5435,N_6834);
and U9363 (N_9363,N_5177,N_7420);
nor U9364 (N_9364,N_7181,N_7013);
nor U9365 (N_9365,N_6967,N_6668);
and U9366 (N_9366,N_7426,N_6706);
and U9367 (N_9367,N_6494,N_5350);
nand U9368 (N_9368,N_5490,N_5997);
nand U9369 (N_9369,N_5046,N_7266);
nand U9370 (N_9370,N_5483,N_6786);
and U9371 (N_9371,N_6753,N_6241);
and U9372 (N_9372,N_6587,N_6542);
nand U9373 (N_9373,N_5368,N_5412);
nand U9374 (N_9374,N_6523,N_5367);
and U9375 (N_9375,N_6933,N_5446);
nand U9376 (N_9376,N_6880,N_5782);
nor U9377 (N_9377,N_6554,N_7272);
nor U9378 (N_9378,N_5419,N_5475);
nand U9379 (N_9379,N_6523,N_7424);
nand U9380 (N_9380,N_6420,N_6685);
or U9381 (N_9381,N_7257,N_7285);
or U9382 (N_9382,N_6496,N_6346);
and U9383 (N_9383,N_6041,N_5777);
xnor U9384 (N_9384,N_5446,N_7079);
nor U9385 (N_9385,N_6783,N_5354);
or U9386 (N_9386,N_5406,N_6490);
and U9387 (N_9387,N_6926,N_6718);
and U9388 (N_9388,N_5952,N_5078);
and U9389 (N_9389,N_7469,N_6464);
nor U9390 (N_9390,N_5364,N_6407);
nand U9391 (N_9391,N_5823,N_6611);
nor U9392 (N_9392,N_6624,N_7308);
and U9393 (N_9393,N_5823,N_6976);
xor U9394 (N_9394,N_7078,N_5018);
nor U9395 (N_9395,N_6130,N_7187);
nand U9396 (N_9396,N_6685,N_7463);
nor U9397 (N_9397,N_7105,N_6456);
xnor U9398 (N_9398,N_5091,N_6499);
nor U9399 (N_9399,N_5486,N_6106);
or U9400 (N_9400,N_5602,N_5992);
nor U9401 (N_9401,N_5050,N_6562);
nor U9402 (N_9402,N_5823,N_7071);
nor U9403 (N_9403,N_6050,N_7017);
nor U9404 (N_9404,N_6395,N_5076);
and U9405 (N_9405,N_5392,N_6945);
nand U9406 (N_9406,N_7364,N_5357);
xnor U9407 (N_9407,N_6456,N_6153);
nor U9408 (N_9408,N_6908,N_5525);
and U9409 (N_9409,N_6028,N_5147);
nor U9410 (N_9410,N_5067,N_6016);
and U9411 (N_9411,N_6085,N_5649);
xnor U9412 (N_9412,N_5709,N_5052);
xor U9413 (N_9413,N_5163,N_6109);
or U9414 (N_9414,N_6605,N_6322);
and U9415 (N_9415,N_5126,N_5184);
xnor U9416 (N_9416,N_5270,N_7298);
xor U9417 (N_9417,N_7345,N_5752);
or U9418 (N_9418,N_5196,N_5537);
nor U9419 (N_9419,N_5654,N_5027);
nor U9420 (N_9420,N_5962,N_5351);
nand U9421 (N_9421,N_6734,N_7025);
nand U9422 (N_9422,N_6720,N_5327);
xnor U9423 (N_9423,N_7115,N_5194);
nor U9424 (N_9424,N_5782,N_5466);
xor U9425 (N_9425,N_6566,N_5565);
or U9426 (N_9426,N_6487,N_5764);
and U9427 (N_9427,N_7136,N_5047);
nor U9428 (N_9428,N_7489,N_5889);
or U9429 (N_9429,N_5751,N_6672);
and U9430 (N_9430,N_5513,N_7265);
or U9431 (N_9431,N_6967,N_5019);
nand U9432 (N_9432,N_5712,N_6640);
xor U9433 (N_9433,N_6189,N_6768);
and U9434 (N_9434,N_5026,N_5932);
or U9435 (N_9435,N_6811,N_7420);
or U9436 (N_9436,N_5939,N_7254);
and U9437 (N_9437,N_5423,N_6104);
nand U9438 (N_9438,N_6178,N_5516);
nor U9439 (N_9439,N_7409,N_7469);
xor U9440 (N_9440,N_7120,N_5447);
nand U9441 (N_9441,N_7242,N_5583);
nand U9442 (N_9442,N_6379,N_5164);
or U9443 (N_9443,N_5219,N_6360);
nand U9444 (N_9444,N_5897,N_5002);
or U9445 (N_9445,N_5033,N_7489);
and U9446 (N_9446,N_6805,N_5150);
nor U9447 (N_9447,N_6878,N_6443);
nand U9448 (N_9448,N_7154,N_5428);
xor U9449 (N_9449,N_6508,N_5504);
and U9450 (N_9450,N_6378,N_7331);
nand U9451 (N_9451,N_7440,N_6801);
xnor U9452 (N_9452,N_6838,N_5756);
xnor U9453 (N_9453,N_5463,N_7059);
nand U9454 (N_9454,N_7158,N_7371);
and U9455 (N_9455,N_7076,N_6098);
or U9456 (N_9456,N_6350,N_7009);
nand U9457 (N_9457,N_5020,N_6777);
nor U9458 (N_9458,N_6068,N_6873);
xor U9459 (N_9459,N_6121,N_5461);
or U9460 (N_9460,N_7221,N_5684);
nor U9461 (N_9461,N_6111,N_5781);
or U9462 (N_9462,N_6338,N_7060);
xor U9463 (N_9463,N_6395,N_5890);
xnor U9464 (N_9464,N_6644,N_6926);
nor U9465 (N_9465,N_5096,N_5134);
nand U9466 (N_9466,N_6393,N_6523);
nor U9467 (N_9467,N_5778,N_5353);
xnor U9468 (N_9468,N_7134,N_5950);
xor U9469 (N_9469,N_5898,N_6169);
and U9470 (N_9470,N_6592,N_6006);
and U9471 (N_9471,N_7223,N_6258);
or U9472 (N_9472,N_6320,N_6922);
nor U9473 (N_9473,N_7359,N_5685);
and U9474 (N_9474,N_7022,N_6564);
xnor U9475 (N_9475,N_5264,N_5423);
and U9476 (N_9476,N_5418,N_6884);
nand U9477 (N_9477,N_5282,N_5522);
or U9478 (N_9478,N_6244,N_5113);
nor U9479 (N_9479,N_5257,N_5577);
xor U9480 (N_9480,N_6473,N_5294);
and U9481 (N_9481,N_6856,N_6420);
xor U9482 (N_9482,N_5647,N_7230);
nand U9483 (N_9483,N_5967,N_7314);
xnor U9484 (N_9484,N_5312,N_5264);
and U9485 (N_9485,N_5451,N_5593);
nand U9486 (N_9486,N_7338,N_5694);
nor U9487 (N_9487,N_5150,N_5250);
or U9488 (N_9488,N_5756,N_7414);
xnor U9489 (N_9489,N_6811,N_6675);
or U9490 (N_9490,N_7137,N_7166);
xor U9491 (N_9491,N_7106,N_7084);
xor U9492 (N_9492,N_7343,N_6394);
nor U9493 (N_9493,N_6579,N_6188);
xor U9494 (N_9494,N_5435,N_5298);
and U9495 (N_9495,N_5302,N_6390);
or U9496 (N_9496,N_5335,N_6991);
nand U9497 (N_9497,N_5168,N_6237);
nor U9498 (N_9498,N_7043,N_5672);
and U9499 (N_9499,N_7185,N_5472);
or U9500 (N_9500,N_5785,N_7388);
nor U9501 (N_9501,N_5551,N_6967);
nor U9502 (N_9502,N_5764,N_7166);
xnor U9503 (N_9503,N_6645,N_5511);
nor U9504 (N_9504,N_6258,N_7090);
and U9505 (N_9505,N_6830,N_7170);
nand U9506 (N_9506,N_5919,N_6829);
and U9507 (N_9507,N_5830,N_5486);
or U9508 (N_9508,N_6432,N_6473);
nand U9509 (N_9509,N_7131,N_6606);
or U9510 (N_9510,N_6266,N_5097);
nand U9511 (N_9511,N_5372,N_6588);
nor U9512 (N_9512,N_7064,N_7267);
nor U9513 (N_9513,N_7486,N_7074);
xnor U9514 (N_9514,N_5116,N_5118);
nor U9515 (N_9515,N_6384,N_7357);
and U9516 (N_9516,N_7125,N_5652);
xor U9517 (N_9517,N_7006,N_7213);
xor U9518 (N_9518,N_6411,N_5841);
xor U9519 (N_9519,N_7064,N_6984);
nand U9520 (N_9520,N_6907,N_6310);
and U9521 (N_9521,N_7202,N_6681);
or U9522 (N_9522,N_5656,N_6544);
or U9523 (N_9523,N_5743,N_6615);
xor U9524 (N_9524,N_7144,N_5161);
nand U9525 (N_9525,N_5741,N_6174);
nor U9526 (N_9526,N_6898,N_7211);
nor U9527 (N_9527,N_6552,N_6814);
or U9528 (N_9528,N_5471,N_6063);
or U9529 (N_9529,N_5476,N_5134);
or U9530 (N_9530,N_5743,N_6852);
nor U9531 (N_9531,N_6817,N_5848);
or U9532 (N_9532,N_7188,N_5812);
nand U9533 (N_9533,N_6194,N_5365);
and U9534 (N_9534,N_6224,N_6030);
nand U9535 (N_9535,N_5257,N_5759);
nor U9536 (N_9536,N_5000,N_5425);
nor U9537 (N_9537,N_5433,N_7487);
or U9538 (N_9538,N_5546,N_6331);
xnor U9539 (N_9539,N_5701,N_7229);
xnor U9540 (N_9540,N_5655,N_5262);
nand U9541 (N_9541,N_5005,N_5391);
nor U9542 (N_9542,N_5044,N_6393);
xor U9543 (N_9543,N_5599,N_5863);
or U9544 (N_9544,N_5205,N_7383);
or U9545 (N_9545,N_7197,N_7019);
nor U9546 (N_9546,N_6334,N_5112);
xor U9547 (N_9547,N_5766,N_7012);
and U9548 (N_9548,N_6200,N_6407);
or U9549 (N_9549,N_6624,N_5880);
and U9550 (N_9550,N_6028,N_5904);
or U9551 (N_9551,N_6175,N_5607);
or U9552 (N_9552,N_5992,N_5797);
nand U9553 (N_9553,N_5163,N_5823);
nand U9554 (N_9554,N_6022,N_5380);
nor U9555 (N_9555,N_5982,N_5898);
nor U9556 (N_9556,N_5744,N_7418);
xor U9557 (N_9557,N_5692,N_6200);
nand U9558 (N_9558,N_6418,N_7460);
xnor U9559 (N_9559,N_5722,N_5763);
nand U9560 (N_9560,N_7480,N_5073);
and U9561 (N_9561,N_7228,N_7171);
nand U9562 (N_9562,N_5464,N_6504);
xor U9563 (N_9563,N_7379,N_5945);
and U9564 (N_9564,N_6060,N_6922);
nand U9565 (N_9565,N_5322,N_5339);
and U9566 (N_9566,N_7013,N_6582);
nand U9567 (N_9567,N_5150,N_5623);
nand U9568 (N_9568,N_6979,N_5548);
nand U9569 (N_9569,N_5392,N_6622);
or U9570 (N_9570,N_5895,N_5085);
or U9571 (N_9571,N_5637,N_5271);
nand U9572 (N_9572,N_6075,N_6244);
or U9573 (N_9573,N_6919,N_5445);
or U9574 (N_9574,N_5206,N_7109);
nor U9575 (N_9575,N_6738,N_6827);
xor U9576 (N_9576,N_6975,N_5887);
nand U9577 (N_9577,N_7022,N_6098);
nor U9578 (N_9578,N_5073,N_5035);
and U9579 (N_9579,N_7050,N_7138);
and U9580 (N_9580,N_6587,N_6897);
nand U9581 (N_9581,N_6599,N_6074);
xnor U9582 (N_9582,N_5075,N_6697);
or U9583 (N_9583,N_5520,N_5538);
nor U9584 (N_9584,N_7339,N_6891);
xnor U9585 (N_9585,N_7271,N_5566);
and U9586 (N_9586,N_6052,N_5245);
nand U9587 (N_9587,N_7450,N_5226);
and U9588 (N_9588,N_6977,N_5439);
or U9589 (N_9589,N_6241,N_6545);
nor U9590 (N_9590,N_6564,N_7392);
and U9591 (N_9591,N_5360,N_6084);
nor U9592 (N_9592,N_5077,N_6973);
nand U9593 (N_9593,N_6775,N_7462);
xnor U9594 (N_9594,N_7475,N_7077);
nand U9595 (N_9595,N_6398,N_6022);
or U9596 (N_9596,N_5562,N_6109);
nand U9597 (N_9597,N_6828,N_7066);
or U9598 (N_9598,N_7000,N_7324);
xnor U9599 (N_9599,N_5062,N_5378);
and U9600 (N_9600,N_6132,N_6738);
xnor U9601 (N_9601,N_7192,N_5851);
or U9602 (N_9602,N_6065,N_6082);
and U9603 (N_9603,N_6975,N_7067);
nand U9604 (N_9604,N_5399,N_6525);
nand U9605 (N_9605,N_6159,N_6823);
nor U9606 (N_9606,N_5904,N_6353);
or U9607 (N_9607,N_6932,N_6686);
or U9608 (N_9608,N_6565,N_5303);
or U9609 (N_9609,N_5696,N_6127);
and U9610 (N_9610,N_5840,N_6498);
or U9611 (N_9611,N_6187,N_6934);
nor U9612 (N_9612,N_7283,N_7488);
nor U9613 (N_9613,N_5321,N_5539);
nor U9614 (N_9614,N_5514,N_5343);
and U9615 (N_9615,N_6275,N_5545);
nand U9616 (N_9616,N_7083,N_6922);
nand U9617 (N_9617,N_5044,N_5283);
and U9618 (N_9618,N_6131,N_5272);
nor U9619 (N_9619,N_6262,N_6519);
and U9620 (N_9620,N_6595,N_5392);
xnor U9621 (N_9621,N_7118,N_6936);
and U9622 (N_9622,N_6569,N_6773);
and U9623 (N_9623,N_6128,N_7146);
xor U9624 (N_9624,N_5622,N_6704);
and U9625 (N_9625,N_5547,N_7089);
xnor U9626 (N_9626,N_5122,N_7109);
and U9627 (N_9627,N_5537,N_6977);
or U9628 (N_9628,N_6269,N_6826);
or U9629 (N_9629,N_5497,N_6644);
and U9630 (N_9630,N_5564,N_6693);
and U9631 (N_9631,N_6967,N_7171);
or U9632 (N_9632,N_5327,N_6457);
or U9633 (N_9633,N_6667,N_7398);
nand U9634 (N_9634,N_7388,N_6245);
and U9635 (N_9635,N_6031,N_5300);
xor U9636 (N_9636,N_6958,N_6742);
nand U9637 (N_9637,N_6336,N_7394);
nor U9638 (N_9638,N_6771,N_6803);
and U9639 (N_9639,N_6313,N_5016);
xor U9640 (N_9640,N_6893,N_5462);
nand U9641 (N_9641,N_6225,N_6833);
and U9642 (N_9642,N_7185,N_5126);
nand U9643 (N_9643,N_5735,N_6735);
and U9644 (N_9644,N_6494,N_6342);
xor U9645 (N_9645,N_6574,N_6855);
or U9646 (N_9646,N_5320,N_6709);
or U9647 (N_9647,N_6814,N_6782);
or U9648 (N_9648,N_6330,N_6579);
nor U9649 (N_9649,N_5972,N_5577);
or U9650 (N_9650,N_6357,N_6935);
or U9651 (N_9651,N_7405,N_6159);
or U9652 (N_9652,N_5718,N_5013);
or U9653 (N_9653,N_6692,N_7291);
nor U9654 (N_9654,N_7219,N_5807);
and U9655 (N_9655,N_6183,N_6454);
nand U9656 (N_9656,N_5466,N_5379);
nand U9657 (N_9657,N_5172,N_5140);
and U9658 (N_9658,N_6169,N_5496);
and U9659 (N_9659,N_6733,N_5030);
nor U9660 (N_9660,N_7433,N_6439);
or U9661 (N_9661,N_7469,N_6801);
and U9662 (N_9662,N_5182,N_6100);
nor U9663 (N_9663,N_6453,N_5019);
and U9664 (N_9664,N_7081,N_5656);
and U9665 (N_9665,N_6487,N_7268);
xor U9666 (N_9666,N_7476,N_6335);
xnor U9667 (N_9667,N_5578,N_6843);
nand U9668 (N_9668,N_5485,N_6826);
nand U9669 (N_9669,N_7042,N_6071);
or U9670 (N_9670,N_6993,N_6716);
or U9671 (N_9671,N_7030,N_5868);
xnor U9672 (N_9672,N_6253,N_6519);
and U9673 (N_9673,N_6194,N_6234);
nand U9674 (N_9674,N_5370,N_7327);
nand U9675 (N_9675,N_5011,N_7202);
nand U9676 (N_9676,N_5376,N_7334);
nand U9677 (N_9677,N_7126,N_5950);
nand U9678 (N_9678,N_5227,N_5806);
or U9679 (N_9679,N_5530,N_5344);
nand U9680 (N_9680,N_7132,N_5190);
or U9681 (N_9681,N_6750,N_6725);
and U9682 (N_9682,N_7092,N_6165);
or U9683 (N_9683,N_5529,N_6206);
and U9684 (N_9684,N_6794,N_6687);
xor U9685 (N_9685,N_7197,N_5861);
xor U9686 (N_9686,N_6800,N_7213);
or U9687 (N_9687,N_7310,N_6658);
or U9688 (N_9688,N_7003,N_5423);
or U9689 (N_9689,N_5772,N_7449);
and U9690 (N_9690,N_7142,N_5128);
or U9691 (N_9691,N_6547,N_7485);
or U9692 (N_9692,N_6265,N_5078);
and U9693 (N_9693,N_7464,N_6232);
nand U9694 (N_9694,N_6199,N_6019);
xor U9695 (N_9695,N_6337,N_5578);
and U9696 (N_9696,N_6595,N_6908);
nand U9697 (N_9697,N_5518,N_5278);
nand U9698 (N_9698,N_5365,N_6064);
or U9699 (N_9699,N_5107,N_6889);
xor U9700 (N_9700,N_5127,N_6986);
xor U9701 (N_9701,N_7242,N_5514);
and U9702 (N_9702,N_6296,N_5053);
xor U9703 (N_9703,N_7368,N_6737);
nand U9704 (N_9704,N_6982,N_5329);
nor U9705 (N_9705,N_6233,N_6064);
xor U9706 (N_9706,N_6591,N_5477);
and U9707 (N_9707,N_7036,N_6868);
and U9708 (N_9708,N_6199,N_7270);
or U9709 (N_9709,N_5076,N_6864);
nand U9710 (N_9710,N_5793,N_6173);
nand U9711 (N_9711,N_5806,N_7014);
xnor U9712 (N_9712,N_7177,N_5837);
or U9713 (N_9713,N_5977,N_5058);
and U9714 (N_9714,N_5612,N_6251);
nor U9715 (N_9715,N_7072,N_5707);
xnor U9716 (N_9716,N_5654,N_5296);
or U9717 (N_9717,N_5119,N_6870);
nor U9718 (N_9718,N_5753,N_5151);
nand U9719 (N_9719,N_5072,N_5360);
nor U9720 (N_9720,N_5810,N_6437);
nor U9721 (N_9721,N_6103,N_6504);
and U9722 (N_9722,N_6464,N_6692);
nand U9723 (N_9723,N_6999,N_6680);
and U9724 (N_9724,N_7452,N_5692);
and U9725 (N_9725,N_6238,N_7090);
nor U9726 (N_9726,N_5237,N_6029);
nand U9727 (N_9727,N_6142,N_7459);
or U9728 (N_9728,N_6206,N_6656);
nor U9729 (N_9729,N_7330,N_5713);
nand U9730 (N_9730,N_6198,N_6914);
and U9731 (N_9731,N_5878,N_7165);
nor U9732 (N_9732,N_5643,N_5371);
xnor U9733 (N_9733,N_6171,N_5748);
nand U9734 (N_9734,N_6070,N_5456);
xor U9735 (N_9735,N_5902,N_6227);
nor U9736 (N_9736,N_6444,N_6715);
and U9737 (N_9737,N_7090,N_6535);
or U9738 (N_9738,N_5907,N_5943);
nand U9739 (N_9739,N_6077,N_6377);
nor U9740 (N_9740,N_7214,N_6025);
or U9741 (N_9741,N_6592,N_7270);
nand U9742 (N_9742,N_5383,N_7174);
nor U9743 (N_9743,N_6495,N_6108);
nor U9744 (N_9744,N_5968,N_6273);
xnor U9745 (N_9745,N_6397,N_6311);
nor U9746 (N_9746,N_5728,N_7123);
and U9747 (N_9747,N_7389,N_6365);
or U9748 (N_9748,N_5644,N_7102);
or U9749 (N_9749,N_5544,N_7468);
nor U9750 (N_9750,N_6709,N_6827);
and U9751 (N_9751,N_5392,N_5149);
nand U9752 (N_9752,N_6364,N_6717);
and U9753 (N_9753,N_5078,N_6138);
xnor U9754 (N_9754,N_6214,N_6676);
or U9755 (N_9755,N_6981,N_6592);
or U9756 (N_9756,N_6134,N_7211);
or U9757 (N_9757,N_7069,N_5455);
or U9758 (N_9758,N_5458,N_7165);
or U9759 (N_9759,N_6410,N_6162);
xor U9760 (N_9760,N_6282,N_7343);
nor U9761 (N_9761,N_5093,N_7141);
and U9762 (N_9762,N_6606,N_7371);
or U9763 (N_9763,N_7112,N_5636);
or U9764 (N_9764,N_6873,N_6381);
nor U9765 (N_9765,N_6045,N_6984);
nor U9766 (N_9766,N_7185,N_5526);
nand U9767 (N_9767,N_7380,N_6282);
xnor U9768 (N_9768,N_5083,N_6354);
or U9769 (N_9769,N_5155,N_7444);
nand U9770 (N_9770,N_7131,N_5721);
nand U9771 (N_9771,N_6997,N_7104);
nor U9772 (N_9772,N_5537,N_5766);
or U9773 (N_9773,N_7275,N_5825);
or U9774 (N_9774,N_6989,N_5967);
and U9775 (N_9775,N_7311,N_6845);
nand U9776 (N_9776,N_5785,N_7112);
and U9777 (N_9777,N_7086,N_5523);
and U9778 (N_9778,N_5589,N_5484);
and U9779 (N_9779,N_5171,N_5725);
nand U9780 (N_9780,N_7058,N_5988);
xnor U9781 (N_9781,N_7039,N_6629);
and U9782 (N_9782,N_7073,N_5171);
or U9783 (N_9783,N_6501,N_6273);
xor U9784 (N_9784,N_5289,N_5821);
or U9785 (N_9785,N_5964,N_5659);
nor U9786 (N_9786,N_5179,N_5360);
or U9787 (N_9787,N_5895,N_6312);
and U9788 (N_9788,N_7121,N_6384);
nor U9789 (N_9789,N_5952,N_5106);
nor U9790 (N_9790,N_6435,N_5290);
nor U9791 (N_9791,N_6152,N_5542);
nand U9792 (N_9792,N_5038,N_6711);
and U9793 (N_9793,N_5562,N_6875);
or U9794 (N_9794,N_6375,N_6953);
or U9795 (N_9795,N_6085,N_5732);
nand U9796 (N_9796,N_7154,N_6029);
or U9797 (N_9797,N_5749,N_7408);
nor U9798 (N_9798,N_6853,N_6625);
nor U9799 (N_9799,N_6959,N_6476);
xnor U9800 (N_9800,N_7426,N_6043);
or U9801 (N_9801,N_6667,N_5631);
and U9802 (N_9802,N_5782,N_5492);
xor U9803 (N_9803,N_5613,N_7492);
nor U9804 (N_9804,N_5024,N_5786);
nor U9805 (N_9805,N_6531,N_5351);
xnor U9806 (N_9806,N_7403,N_5113);
and U9807 (N_9807,N_5269,N_7261);
and U9808 (N_9808,N_5410,N_6498);
nand U9809 (N_9809,N_7306,N_6282);
nor U9810 (N_9810,N_5166,N_6458);
nand U9811 (N_9811,N_6542,N_6926);
xnor U9812 (N_9812,N_5594,N_7364);
nor U9813 (N_9813,N_6485,N_6195);
or U9814 (N_9814,N_6609,N_5023);
nand U9815 (N_9815,N_7238,N_6634);
xnor U9816 (N_9816,N_5697,N_7279);
nand U9817 (N_9817,N_6195,N_6475);
or U9818 (N_9818,N_5450,N_6045);
nand U9819 (N_9819,N_5657,N_6168);
xor U9820 (N_9820,N_5732,N_6471);
xor U9821 (N_9821,N_5280,N_7009);
nor U9822 (N_9822,N_5489,N_6652);
nor U9823 (N_9823,N_5789,N_7125);
or U9824 (N_9824,N_6266,N_6272);
xor U9825 (N_9825,N_5467,N_7164);
and U9826 (N_9826,N_5199,N_5919);
nand U9827 (N_9827,N_7244,N_5822);
and U9828 (N_9828,N_7112,N_5095);
or U9829 (N_9829,N_6672,N_6512);
and U9830 (N_9830,N_5745,N_5031);
nand U9831 (N_9831,N_6168,N_6186);
nand U9832 (N_9832,N_5949,N_5809);
nor U9833 (N_9833,N_5770,N_5797);
or U9834 (N_9834,N_6880,N_5061);
nand U9835 (N_9835,N_6600,N_5793);
nor U9836 (N_9836,N_5783,N_6963);
nor U9837 (N_9837,N_5885,N_6587);
nor U9838 (N_9838,N_5033,N_5915);
and U9839 (N_9839,N_5434,N_6503);
nor U9840 (N_9840,N_7468,N_6872);
nor U9841 (N_9841,N_5247,N_7337);
nor U9842 (N_9842,N_5556,N_6872);
nor U9843 (N_9843,N_7350,N_6941);
nor U9844 (N_9844,N_6447,N_6504);
or U9845 (N_9845,N_7139,N_5062);
or U9846 (N_9846,N_7164,N_5535);
nor U9847 (N_9847,N_6593,N_6961);
xnor U9848 (N_9848,N_6557,N_7019);
nand U9849 (N_9849,N_6406,N_5881);
and U9850 (N_9850,N_6582,N_5316);
nand U9851 (N_9851,N_5395,N_5298);
or U9852 (N_9852,N_5043,N_7145);
xor U9853 (N_9853,N_6400,N_7166);
or U9854 (N_9854,N_5000,N_7090);
nor U9855 (N_9855,N_7314,N_5298);
or U9856 (N_9856,N_5369,N_6983);
nor U9857 (N_9857,N_5810,N_6621);
nor U9858 (N_9858,N_5387,N_5110);
xnor U9859 (N_9859,N_5549,N_6887);
nand U9860 (N_9860,N_5132,N_6143);
or U9861 (N_9861,N_5840,N_7072);
nand U9862 (N_9862,N_6153,N_6213);
xnor U9863 (N_9863,N_6575,N_5785);
nand U9864 (N_9864,N_6690,N_5987);
nand U9865 (N_9865,N_6749,N_7020);
or U9866 (N_9866,N_5073,N_6130);
xnor U9867 (N_9867,N_5046,N_6112);
and U9868 (N_9868,N_5970,N_6276);
nand U9869 (N_9869,N_5118,N_7373);
nand U9870 (N_9870,N_6678,N_5738);
nand U9871 (N_9871,N_6282,N_6971);
xnor U9872 (N_9872,N_5714,N_6593);
or U9873 (N_9873,N_6186,N_5394);
or U9874 (N_9874,N_6326,N_6668);
or U9875 (N_9875,N_5729,N_6077);
nor U9876 (N_9876,N_5002,N_5379);
or U9877 (N_9877,N_6742,N_6911);
nor U9878 (N_9878,N_6566,N_5318);
nand U9879 (N_9879,N_6907,N_5346);
nor U9880 (N_9880,N_6501,N_6166);
xnor U9881 (N_9881,N_7275,N_6855);
nor U9882 (N_9882,N_5377,N_7343);
nor U9883 (N_9883,N_7153,N_5271);
nor U9884 (N_9884,N_7451,N_7345);
or U9885 (N_9885,N_7219,N_6426);
and U9886 (N_9886,N_7242,N_6319);
or U9887 (N_9887,N_5318,N_7282);
nand U9888 (N_9888,N_5250,N_5756);
or U9889 (N_9889,N_5928,N_7383);
and U9890 (N_9890,N_6574,N_7036);
or U9891 (N_9891,N_5604,N_5907);
nand U9892 (N_9892,N_7440,N_6698);
xor U9893 (N_9893,N_7167,N_5773);
nor U9894 (N_9894,N_5956,N_5389);
nor U9895 (N_9895,N_6231,N_6707);
nand U9896 (N_9896,N_5441,N_5942);
xnor U9897 (N_9897,N_5546,N_6322);
and U9898 (N_9898,N_5107,N_5410);
or U9899 (N_9899,N_6156,N_7277);
nand U9900 (N_9900,N_5183,N_6238);
nor U9901 (N_9901,N_6671,N_6568);
nor U9902 (N_9902,N_5865,N_5509);
nand U9903 (N_9903,N_5382,N_7130);
nor U9904 (N_9904,N_6067,N_7057);
or U9905 (N_9905,N_5659,N_5881);
and U9906 (N_9906,N_5154,N_5039);
xor U9907 (N_9907,N_5998,N_7490);
nor U9908 (N_9908,N_5510,N_5592);
and U9909 (N_9909,N_7425,N_6004);
xnor U9910 (N_9910,N_5262,N_6651);
and U9911 (N_9911,N_7111,N_5958);
nand U9912 (N_9912,N_7395,N_5019);
or U9913 (N_9913,N_7309,N_6859);
nor U9914 (N_9914,N_6751,N_6426);
or U9915 (N_9915,N_7484,N_5084);
or U9916 (N_9916,N_5311,N_7489);
xnor U9917 (N_9917,N_5816,N_5779);
and U9918 (N_9918,N_6442,N_5616);
or U9919 (N_9919,N_6485,N_5253);
and U9920 (N_9920,N_5092,N_5440);
nor U9921 (N_9921,N_5771,N_6608);
and U9922 (N_9922,N_6208,N_5975);
and U9923 (N_9923,N_6326,N_5449);
nor U9924 (N_9924,N_6587,N_5949);
xor U9925 (N_9925,N_5125,N_5777);
nand U9926 (N_9926,N_5168,N_7011);
or U9927 (N_9927,N_7192,N_6518);
nand U9928 (N_9928,N_6470,N_7340);
nand U9929 (N_9929,N_6825,N_6423);
nor U9930 (N_9930,N_7045,N_6501);
nor U9931 (N_9931,N_5708,N_6730);
and U9932 (N_9932,N_6777,N_7433);
nor U9933 (N_9933,N_5338,N_5348);
nand U9934 (N_9934,N_6714,N_5414);
nor U9935 (N_9935,N_5567,N_7464);
and U9936 (N_9936,N_6885,N_5877);
xnor U9937 (N_9937,N_6618,N_7272);
nor U9938 (N_9938,N_6237,N_7136);
or U9939 (N_9939,N_5716,N_5538);
or U9940 (N_9940,N_6678,N_6172);
and U9941 (N_9941,N_5803,N_6310);
xnor U9942 (N_9942,N_5489,N_5853);
and U9943 (N_9943,N_5917,N_5347);
and U9944 (N_9944,N_6024,N_5978);
nand U9945 (N_9945,N_5733,N_7011);
nor U9946 (N_9946,N_6149,N_6367);
nor U9947 (N_9947,N_5092,N_6652);
nand U9948 (N_9948,N_6327,N_6774);
or U9949 (N_9949,N_6059,N_5836);
nor U9950 (N_9950,N_5314,N_7113);
nand U9951 (N_9951,N_5003,N_5155);
and U9952 (N_9952,N_5148,N_7212);
nor U9953 (N_9953,N_6695,N_6696);
nor U9954 (N_9954,N_5180,N_5217);
nand U9955 (N_9955,N_6297,N_5793);
or U9956 (N_9956,N_5706,N_6790);
nand U9957 (N_9957,N_6838,N_6928);
xnor U9958 (N_9958,N_6386,N_6065);
xnor U9959 (N_9959,N_5279,N_7349);
and U9960 (N_9960,N_5947,N_5709);
xor U9961 (N_9961,N_7373,N_5176);
nand U9962 (N_9962,N_6881,N_5652);
nor U9963 (N_9963,N_6853,N_7426);
or U9964 (N_9964,N_7098,N_6629);
nand U9965 (N_9965,N_6447,N_6188);
nor U9966 (N_9966,N_7106,N_6337);
nor U9967 (N_9967,N_6222,N_7346);
nand U9968 (N_9968,N_5882,N_6673);
nor U9969 (N_9969,N_6650,N_6557);
xor U9970 (N_9970,N_5166,N_7120);
nand U9971 (N_9971,N_6018,N_5285);
nor U9972 (N_9972,N_7261,N_6411);
or U9973 (N_9973,N_6605,N_5624);
or U9974 (N_9974,N_6718,N_7351);
or U9975 (N_9975,N_6805,N_5067);
nor U9976 (N_9976,N_5545,N_5827);
nand U9977 (N_9977,N_5105,N_6024);
nand U9978 (N_9978,N_7071,N_5564);
or U9979 (N_9979,N_5813,N_6805);
xnor U9980 (N_9980,N_5938,N_6917);
or U9981 (N_9981,N_5571,N_5024);
xnor U9982 (N_9982,N_5262,N_6169);
nor U9983 (N_9983,N_5365,N_5872);
nand U9984 (N_9984,N_6709,N_7147);
xor U9985 (N_9985,N_6545,N_6317);
and U9986 (N_9986,N_6120,N_6070);
and U9987 (N_9987,N_5354,N_5787);
nor U9988 (N_9988,N_6167,N_6046);
nand U9989 (N_9989,N_7346,N_6426);
nor U9990 (N_9990,N_6719,N_5540);
nor U9991 (N_9991,N_6520,N_6505);
nand U9992 (N_9992,N_6846,N_5414);
nor U9993 (N_9993,N_6413,N_7155);
nand U9994 (N_9994,N_7245,N_6604);
nand U9995 (N_9995,N_7384,N_7240);
or U9996 (N_9996,N_7331,N_5687);
or U9997 (N_9997,N_5885,N_6688);
nand U9998 (N_9998,N_5785,N_5348);
xor U9999 (N_9999,N_5636,N_5015);
nand UO_0 (O_0,N_9744,N_9628);
nor UO_1 (O_1,N_7612,N_9674);
nor UO_2 (O_2,N_9240,N_9389);
xor UO_3 (O_3,N_9293,N_9680);
and UO_4 (O_4,N_9685,N_7508);
nor UO_5 (O_5,N_7956,N_9368);
nand UO_6 (O_6,N_9622,N_9113);
xor UO_7 (O_7,N_8719,N_8779);
nand UO_8 (O_8,N_9634,N_9983);
or UO_9 (O_9,N_9927,N_8252);
and UO_10 (O_10,N_8987,N_8793);
xnor UO_11 (O_11,N_7877,N_7908);
nand UO_12 (O_12,N_9866,N_9617);
nand UO_13 (O_13,N_7797,N_8760);
xor UO_14 (O_14,N_8137,N_9521);
and UO_15 (O_15,N_8458,N_7762);
or UO_16 (O_16,N_9449,N_8929);
xnor UO_17 (O_17,N_8228,N_9852);
and UO_18 (O_18,N_8715,N_9311);
nand UO_19 (O_19,N_9724,N_9097);
nand UO_20 (O_20,N_7750,N_9797);
xnor UO_21 (O_21,N_9402,N_9718);
or UO_22 (O_22,N_8275,N_7851);
nor UO_23 (O_23,N_9187,N_9826);
or UO_24 (O_24,N_9963,N_9078);
xnor UO_25 (O_25,N_8886,N_7689);
or UO_26 (O_26,N_7624,N_8396);
nand UO_27 (O_27,N_7619,N_8803);
and UO_28 (O_28,N_9992,N_8170);
nand UO_29 (O_29,N_7921,N_8849);
nand UO_30 (O_30,N_7969,N_7790);
nor UO_31 (O_31,N_8147,N_9639);
or UO_32 (O_32,N_8654,N_9986);
or UO_33 (O_33,N_8100,N_8066);
and UO_34 (O_34,N_8238,N_9928);
and UO_35 (O_35,N_9651,N_8500);
and UO_36 (O_36,N_8941,N_7606);
or UO_37 (O_37,N_9995,N_8885);
nor UO_38 (O_38,N_9609,N_8254);
and UO_39 (O_39,N_8272,N_9231);
nand UO_40 (O_40,N_7636,N_8414);
or UO_41 (O_41,N_9557,N_9728);
nor UO_42 (O_42,N_7869,N_9751);
or UO_43 (O_43,N_8707,N_9641);
and UO_44 (O_44,N_9978,N_8448);
and UO_45 (O_45,N_9530,N_8295);
and UO_46 (O_46,N_7661,N_9794);
or UO_47 (O_47,N_7557,N_7771);
nand UO_48 (O_48,N_9915,N_8980);
nor UO_49 (O_49,N_8278,N_7766);
nand UO_50 (O_50,N_8496,N_9920);
and UO_51 (O_51,N_9009,N_9971);
xnor UO_52 (O_52,N_8853,N_9583);
nand UO_53 (O_53,N_8319,N_8955);
nor UO_54 (O_54,N_8599,N_9525);
nor UO_55 (O_55,N_9711,N_8482);
nand UO_56 (O_56,N_8587,N_8423);
and UO_57 (O_57,N_8261,N_8576);
nor UO_58 (O_58,N_7964,N_9167);
xor UO_59 (O_59,N_9709,N_9734);
nand UO_60 (O_60,N_9904,N_9791);
nand UO_61 (O_61,N_9395,N_8361);
xnor UO_62 (O_62,N_7996,N_9966);
xor UO_63 (O_63,N_8995,N_8483);
or UO_64 (O_64,N_9569,N_9339);
or UO_65 (O_65,N_8026,N_9315);
xnor UO_66 (O_66,N_8809,N_9682);
nor UO_67 (O_67,N_8753,N_9754);
and UO_68 (O_68,N_7602,N_9343);
nand UO_69 (O_69,N_7706,N_9401);
xnor UO_70 (O_70,N_8472,N_8209);
nor UO_71 (O_71,N_8083,N_8766);
and UO_72 (O_72,N_9428,N_7922);
and UO_73 (O_73,N_7947,N_9917);
xnor UO_74 (O_74,N_8136,N_8233);
xor UO_75 (O_75,N_9790,N_9138);
and UO_76 (O_76,N_8893,N_7838);
xor UO_77 (O_77,N_9446,N_9829);
xnor UO_78 (O_78,N_8774,N_8836);
and UO_79 (O_79,N_7933,N_9417);
or UO_80 (O_80,N_9710,N_9391);
nor UO_81 (O_81,N_9721,N_9518);
xor UO_82 (O_82,N_7630,N_7920);
nand UO_83 (O_83,N_7957,N_9498);
or UO_84 (O_84,N_7569,N_7768);
xnor UO_85 (O_85,N_7783,N_9129);
nand UO_86 (O_86,N_8574,N_8968);
or UO_87 (O_87,N_7695,N_7543);
or UO_88 (O_88,N_9823,N_8276);
xnor UO_89 (O_89,N_7615,N_9548);
nand UO_90 (O_90,N_9454,N_9946);
nor UO_91 (O_91,N_7801,N_9363);
xnor UO_92 (O_92,N_9938,N_9541);
nand UO_93 (O_93,N_9566,N_9091);
xnor UO_94 (O_94,N_7726,N_9325);
nor UO_95 (O_95,N_8926,N_7659);
nand UO_96 (O_96,N_7798,N_8614);
nor UO_97 (O_97,N_8003,N_8530);
and UO_98 (O_98,N_9887,N_9032);
and UO_99 (O_99,N_8429,N_7611);
and UO_100 (O_100,N_8972,N_9044);
nor UO_101 (O_101,N_9783,N_9037);
nand UO_102 (O_102,N_8292,N_7911);
and UO_103 (O_103,N_9073,N_8901);
nor UO_104 (O_104,N_7539,N_7603);
nor UO_105 (O_105,N_9468,N_9051);
xnor UO_106 (O_106,N_9761,N_8314);
or UO_107 (O_107,N_8401,N_7931);
and UO_108 (O_108,N_8315,N_8438);
and UO_109 (O_109,N_7940,N_7562);
xor UO_110 (O_110,N_9623,N_7868);
nor UO_111 (O_111,N_9195,N_7573);
and UO_112 (O_112,N_9850,N_7503);
nand UO_113 (O_113,N_7909,N_8508);
and UO_114 (O_114,N_8864,N_9427);
or UO_115 (O_115,N_7679,N_7918);
nor UO_116 (O_116,N_9964,N_7667);
and UO_117 (O_117,N_7577,N_9178);
nor UO_118 (O_118,N_8203,N_9650);
nand UO_119 (O_119,N_7622,N_8873);
xor UO_120 (O_120,N_9683,N_8855);
nand UO_121 (O_121,N_8813,N_7678);
nor UO_122 (O_122,N_9506,N_7916);
nand UO_123 (O_123,N_7582,N_8287);
nor UO_124 (O_124,N_9227,N_9547);
or UO_125 (O_125,N_9045,N_8206);
or UO_126 (O_126,N_9221,N_9279);
nor UO_127 (O_127,N_7968,N_9869);
and UO_128 (O_128,N_7914,N_9840);
xnor UO_129 (O_129,N_9644,N_8101);
nor UO_130 (O_130,N_7684,N_9316);
xor UO_131 (O_131,N_9069,N_9372);
or UO_132 (O_132,N_9635,N_7997);
nor UO_133 (O_133,N_8207,N_7891);
or UO_134 (O_134,N_9041,N_9740);
nand UO_135 (O_135,N_9160,N_7613);
and UO_136 (O_136,N_8461,N_9262);
nand UO_137 (O_137,N_9871,N_8814);
xnor UO_138 (O_138,N_8397,N_9356);
and UO_139 (O_139,N_9726,N_9435);
or UO_140 (O_140,N_9245,N_9458);
or UO_141 (O_141,N_9592,N_8785);
nand UO_142 (O_142,N_7532,N_9234);
and UO_143 (O_143,N_9555,N_8568);
nand UO_144 (O_144,N_9573,N_8830);
nand UO_145 (O_145,N_9008,N_8918);
or UO_146 (O_146,N_8798,N_8143);
xnor UO_147 (O_147,N_9038,N_8718);
xnor UO_148 (O_148,N_7810,N_8708);
xor UO_149 (O_149,N_8964,N_9969);
nand UO_150 (O_150,N_8515,N_8600);
nor UO_151 (O_151,N_7520,N_9994);
or UO_152 (O_152,N_9911,N_7552);
and UO_153 (O_153,N_8132,N_8916);
nor UO_154 (O_154,N_9077,N_8581);
nand UO_155 (O_155,N_7887,N_7523);
nand UO_156 (O_156,N_9578,N_8925);
nor UO_157 (O_157,N_9590,N_9305);
nand UO_158 (O_158,N_7896,N_8265);
nor UO_159 (O_159,N_9903,N_9531);
and UO_160 (O_160,N_9588,N_9845);
or UO_161 (O_161,N_8250,N_8459);
and UO_162 (O_162,N_8106,N_8450);
nor UO_163 (O_163,N_7501,N_8210);
and UO_164 (O_164,N_8620,N_9342);
xnor UO_165 (O_165,N_9184,N_8741);
and UO_166 (O_166,N_7561,N_9649);
or UO_167 (O_167,N_9747,N_8200);
and UO_168 (O_168,N_7795,N_7820);
nand UO_169 (O_169,N_9941,N_8984);
or UO_170 (O_170,N_8366,N_9265);
xor UO_171 (O_171,N_8205,N_8591);
nand UO_172 (O_172,N_9460,N_9816);
nand UO_173 (O_173,N_8532,N_7811);
xor UO_174 (O_174,N_9593,N_8122);
nor UO_175 (O_175,N_9317,N_8175);
and UO_176 (O_176,N_9602,N_9165);
and UO_177 (O_177,N_9672,N_8764);
xor UO_178 (O_178,N_8196,N_9171);
and UO_179 (O_179,N_7741,N_8380);
and UO_180 (O_180,N_8037,N_8476);
xor UO_181 (O_181,N_9445,N_7510);
or UO_182 (O_182,N_8381,N_9143);
nand UO_183 (O_183,N_7821,N_9340);
or UO_184 (O_184,N_9450,N_9040);
nor UO_185 (O_185,N_8235,N_8298);
nand UO_186 (O_186,N_7785,N_9205);
nor UO_187 (O_187,N_8131,N_7961);
nor UO_188 (O_188,N_8327,N_9695);
xor UO_189 (O_189,N_8640,N_7595);
or UO_190 (O_190,N_9284,N_8477);
nand UO_191 (O_191,N_8602,N_9604);
or UO_192 (O_192,N_9615,N_9482);
or UO_193 (O_193,N_9601,N_9440);
xor UO_194 (O_194,N_9631,N_9083);
xor UO_195 (O_195,N_9459,N_9054);
xor UO_196 (O_196,N_7852,N_9875);
or UO_197 (O_197,N_8229,N_8068);
xnor UO_198 (O_198,N_8994,N_9485);
and UO_199 (O_199,N_8804,N_8788);
or UO_200 (O_200,N_8728,N_8892);
nor UO_201 (O_201,N_7675,N_9101);
xor UO_202 (O_202,N_8240,N_9970);
nand UO_203 (O_203,N_8952,N_9847);
and UO_204 (O_204,N_8484,N_7842);
nor UO_205 (O_205,N_8927,N_9164);
xor UO_206 (O_206,N_8535,N_9088);
nor UO_207 (O_207,N_9373,N_9627);
xnor UO_208 (O_208,N_9872,N_9412);
nand UO_209 (O_209,N_8466,N_8251);
or UO_210 (O_210,N_9965,N_8526);
nor UO_211 (O_211,N_8112,N_9287);
or UO_212 (O_212,N_8998,N_9330);
nor UO_213 (O_213,N_8110,N_8672);
or UO_214 (O_214,N_8040,N_8236);
and UO_215 (O_215,N_9586,N_7743);
nor UO_216 (O_216,N_9140,N_8491);
nand UO_217 (O_217,N_9860,N_7815);
nand UO_218 (O_218,N_9523,N_9224);
or UO_219 (O_219,N_8231,N_8969);
and UO_220 (O_220,N_7549,N_7625);
nand UO_221 (O_221,N_7696,N_9378);
nor UO_222 (O_222,N_8079,N_8870);
nand UO_223 (O_223,N_8379,N_8427);
and UO_224 (O_224,N_8595,N_9808);
xnor UO_225 (O_225,N_8214,N_7999);
nor UO_226 (O_226,N_9309,N_9406);
or UO_227 (O_227,N_7698,N_7749);
and UO_228 (O_228,N_7834,N_8027);
or UO_229 (O_229,N_9748,N_8481);
nand UO_230 (O_230,N_9087,N_7976);
nand UO_231 (O_231,N_8360,N_8345);
nor UO_232 (O_232,N_8019,N_7609);
and UO_233 (O_233,N_9658,N_9407);
nand UO_234 (O_234,N_9802,N_9849);
and UO_235 (O_235,N_7645,N_8406);
or UO_236 (O_236,N_8632,N_8844);
nand UO_237 (O_237,N_9151,N_9731);
nand UO_238 (O_238,N_9912,N_8978);
xnor UO_239 (O_239,N_8783,N_9777);
xor UO_240 (O_240,N_7502,N_9225);
and UO_241 (O_241,N_8597,N_7776);
or UO_242 (O_242,N_9246,N_9220);
or UO_243 (O_243,N_7949,N_9319);
nor UO_244 (O_244,N_9494,N_8557);
nand UO_245 (O_245,N_9800,N_9846);
xnor UO_246 (O_246,N_8316,N_9772);
xnor UO_247 (O_247,N_9824,N_9384);
and UO_248 (O_248,N_8422,N_8693);
or UO_249 (O_249,N_9335,N_9512);
xnor UO_250 (O_250,N_9688,N_8045);
nor UO_251 (O_251,N_8913,N_9139);
xnor UO_252 (O_252,N_8882,N_8069);
nor UO_253 (O_253,N_9410,N_7534);
nor UO_254 (O_254,N_7863,N_8243);
nor UO_255 (O_255,N_7690,N_8695);
and UO_256 (O_256,N_9441,N_8943);
nor UO_257 (O_257,N_9766,N_9544);
nand UO_258 (O_258,N_7945,N_8453);
xnor UO_259 (O_259,N_8359,N_8135);
nand UO_260 (O_260,N_9413,N_9629);
xor UO_261 (O_261,N_8042,N_7687);
nor UO_262 (O_262,N_8081,N_8290);
xor UO_263 (O_263,N_9306,N_9526);
or UO_264 (O_264,N_7703,N_8811);
and UO_265 (O_265,N_8773,N_8956);
nor UO_266 (O_266,N_9470,N_8879);
and UO_267 (O_267,N_9930,N_9393);
xor UO_268 (O_268,N_9414,N_8454);
or UO_269 (O_269,N_8226,N_8612);
nor UO_270 (O_270,N_7917,N_8981);
and UO_271 (O_271,N_7500,N_9795);
and UO_272 (O_272,N_8056,N_8058);
nor UO_273 (O_273,N_9758,N_8904);
and UO_274 (O_274,N_7751,N_9489);
xnor UO_275 (O_275,N_9807,N_8639);
and UO_276 (O_276,N_9700,N_7676);
and UO_277 (O_277,N_8220,N_9906);
nor UO_278 (O_278,N_9621,N_9955);
nand UO_279 (O_279,N_8108,N_7840);
nand UO_280 (O_280,N_9462,N_9580);
xnor UO_281 (O_281,N_8837,N_8677);
and UO_282 (O_282,N_8506,N_8687);
and UO_283 (O_283,N_7734,N_9565);
or UO_284 (O_284,N_9042,N_9606);
and UO_285 (O_285,N_9484,N_9191);
xnor UO_286 (O_286,N_9982,N_9355);
and UO_287 (O_287,N_8649,N_9023);
nand UO_288 (O_288,N_9898,N_8294);
and UO_289 (O_289,N_9273,N_9333);
nor UO_290 (O_290,N_9248,N_8513);
xnor UO_291 (O_291,N_9997,N_7725);
nor UO_292 (O_292,N_8141,N_7610);
and UO_293 (O_293,N_8098,N_9211);
or UO_294 (O_294,N_7867,N_9620);
and UO_295 (O_295,N_9331,N_7827);
xor UO_296 (O_296,N_9676,N_9338);
nor UO_297 (O_297,N_9519,N_8628);
xnor UO_298 (O_298,N_8709,N_7664);
and UO_299 (O_299,N_8221,N_7632);
and UO_300 (O_300,N_8159,N_8242);
or UO_301 (O_301,N_8311,N_9940);
xnor UO_302 (O_302,N_8195,N_8739);
nand UO_303 (O_303,N_8171,N_9960);
or UO_304 (O_304,N_7756,N_7585);
xor UO_305 (O_305,N_7589,N_8877);
and UO_306 (O_306,N_8665,N_9770);
or UO_307 (O_307,N_7928,N_8494);
xor UO_308 (O_308,N_7903,N_8761);
nand UO_309 (O_309,N_8103,N_9432);
or UO_310 (O_310,N_9361,N_8362);
xnor UO_311 (O_311,N_9998,N_9839);
or UO_312 (O_312,N_8645,N_8580);
or UO_313 (O_313,N_8704,N_8909);
or UO_314 (O_314,N_8288,N_9614);
nand UO_315 (O_315,N_9673,N_9568);
nor UO_316 (O_316,N_9229,N_8102);
nand UO_317 (O_317,N_8398,N_9297);
or UO_318 (O_318,N_8520,N_9351);
nand UO_319 (O_319,N_8551,N_8385);
xnor UO_320 (O_320,N_8237,N_8149);
and UO_321 (O_321,N_9300,N_9242);
and UO_322 (O_322,N_8938,N_8765);
and UO_323 (O_323,N_7980,N_7804);
nor UO_324 (O_324,N_7631,N_8902);
nor UO_325 (O_325,N_9065,N_8652);
and UO_326 (O_326,N_9295,N_8517);
xnor UO_327 (O_327,N_9831,N_8331);
nor UO_328 (O_328,N_8451,N_9874);
nor UO_329 (O_329,N_8178,N_8322);
and UO_330 (O_330,N_8321,N_9640);
nor UO_331 (O_331,N_9324,N_8138);
and UO_332 (O_332,N_9142,N_9163);
or UO_333 (O_333,N_8168,N_9691);
and UO_334 (O_334,N_8723,N_7818);
xnor UO_335 (O_335,N_8967,N_9301);
and UO_336 (O_336,N_9254,N_8320);
xnor UO_337 (O_337,N_7954,N_7878);
or UO_338 (O_338,N_8651,N_9843);
xnor UO_339 (O_339,N_8395,N_8184);
or UO_340 (O_340,N_8383,N_9514);
xnor UO_341 (O_341,N_7910,N_9561);
nor UO_342 (O_342,N_8786,N_9341);
or UO_343 (O_343,N_8562,N_9861);
xor UO_344 (O_344,N_8501,N_9382);
xor UO_345 (O_345,N_9947,N_8791);
nand UO_346 (O_346,N_9597,N_9553);
xnor UO_347 (O_347,N_8659,N_8795);
nand UO_348 (O_348,N_9499,N_8324);
nand UO_349 (O_349,N_8375,N_8618);
or UO_350 (O_350,N_8908,N_8441);
and UO_351 (O_351,N_8073,N_9024);
nor UO_352 (O_352,N_9334,N_8922);
or UO_353 (O_353,N_9067,N_7727);
and UO_354 (O_354,N_9697,N_9817);
or UO_355 (O_355,N_7707,N_8227);
or UO_356 (O_356,N_9785,N_8550);
nor UO_357 (O_357,N_8782,N_9642);
nand UO_358 (O_358,N_9689,N_8428);
and UO_359 (O_359,N_9477,N_8619);
and UO_360 (O_360,N_9675,N_8239);
nand UO_361 (O_361,N_8151,N_9663);
nand UO_362 (O_362,N_9177,N_8077);
and UO_363 (O_363,N_7959,N_9457);
and UO_364 (O_364,N_7568,N_8588);
nand UO_365 (O_365,N_8903,N_7651);
nor UO_366 (O_366,N_7871,N_8474);
or UO_367 (O_367,N_8216,N_8827);
nor UO_368 (O_368,N_8493,N_9660);
nor UO_369 (O_369,N_8875,N_8305);
xnor UO_370 (O_370,N_9172,N_8424);
or UO_371 (O_371,N_9764,N_9968);
nand UO_372 (O_372,N_8514,N_9865);
nand UO_373 (O_373,N_7740,N_8548);
or UO_374 (O_374,N_8394,N_9094);
and UO_375 (O_375,N_9421,N_7836);
and UO_376 (O_376,N_8626,N_8790);
and UO_377 (O_377,N_7854,N_8638);
nand UO_378 (O_378,N_8358,N_9611);
nor UO_379 (O_379,N_8062,N_8961);
and UO_380 (O_380,N_8558,N_9692);
or UO_381 (O_381,N_9259,N_8865);
and UO_382 (O_382,N_9288,N_9476);
or UO_383 (O_383,N_8607,N_8642);
nor UO_384 (O_384,N_8129,N_7662);
xor UO_385 (O_385,N_8009,N_7984);
nor UO_386 (O_386,N_7946,N_7833);
or UO_387 (O_387,N_7879,N_7773);
nand UO_388 (O_388,N_8650,N_7641);
xor UO_389 (O_389,N_7814,N_9626);
xor UO_390 (O_390,N_9844,N_7958);
and UO_391 (O_391,N_8720,N_8347);
nor UO_392 (O_392,N_9522,N_9769);
xnor UO_393 (O_393,N_7786,N_8933);
or UO_394 (O_394,N_9504,N_8144);
nand UO_395 (O_395,N_9099,N_8817);
nor UO_396 (O_396,N_8117,N_9922);
xnor UO_397 (O_397,N_7967,N_8312);
nor UO_398 (O_398,N_8637,N_9954);
xor UO_399 (O_399,N_7658,N_9895);
nand UO_400 (O_400,N_9020,N_9638);
and UO_401 (O_401,N_8653,N_9868);
or UO_402 (O_402,N_7809,N_7578);
and UO_403 (O_403,N_9048,N_9552);
nor UO_404 (O_404,N_9481,N_7711);
xor UO_405 (O_405,N_9505,N_7979);
nand UO_406 (O_406,N_9228,N_9618);
nand UO_407 (O_407,N_7799,N_7919);
and UO_408 (O_408,N_9612,N_9010);
nor UO_409 (O_409,N_9788,N_9186);
nor UO_410 (O_410,N_9174,N_8738);
xor UO_411 (O_411,N_9517,N_8094);
or UO_412 (O_412,N_9422,N_8076);
and UO_413 (O_413,N_8356,N_9249);
nor UO_414 (O_414,N_8133,N_7587);
and UO_415 (O_415,N_9116,N_9900);
or UO_416 (O_416,N_9131,N_8368);
nor UO_417 (O_417,N_8856,N_8928);
xor UO_418 (O_418,N_7699,N_9752);
nor UO_419 (O_419,N_9332,N_9092);
nor UO_420 (O_420,N_8286,N_9702);
or UO_421 (O_421,N_9365,N_9084);
or UO_422 (O_422,N_8165,N_8389);
nand UO_423 (O_423,N_9987,N_9803);
or UO_424 (O_424,N_9133,N_8572);
nand UO_425 (O_425,N_9155,N_7982);
and UO_426 (O_426,N_8057,N_9493);
and UO_427 (O_427,N_9813,N_9135);
and UO_428 (O_428,N_8338,N_8656);
nor UO_429 (O_429,N_8912,N_8946);
xor UO_430 (O_430,N_7538,N_8890);
xnor UO_431 (O_431,N_9774,N_8516);
and UO_432 (O_432,N_8683,N_7524);
or UO_433 (O_433,N_9239,N_9303);
xnor UO_434 (O_434,N_7880,N_8993);
and UO_435 (O_435,N_8148,N_9690);
or UO_436 (O_436,N_9028,N_7832);
or UO_437 (O_437,N_8266,N_9058);
and UO_438 (O_438,N_9878,N_7816);
xnor UO_439 (O_439,N_9423,N_9196);
nand UO_440 (O_440,N_8182,N_8512);
and UO_441 (O_441,N_8778,N_8940);
nand UO_442 (O_442,N_9532,N_8979);
nor UO_443 (O_443,N_9717,N_8378);
xnor UO_444 (O_444,N_8215,N_7823);
nand UO_445 (O_445,N_9773,N_8053);
and UO_446 (O_446,N_8464,N_7873);
nand UO_447 (O_447,N_8546,N_7835);
and UO_448 (O_448,N_8097,N_9496);
and UO_449 (O_449,N_8124,N_9511);
nor UO_450 (O_450,N_8431,N_9809);
nor UO_451 (O_451,N_8889,N_7974);
xnor UO_452 (O_452,N_8293,N_9775);
nor UO_453 (O_453,N_9200,N_8334);
xnor UO_454 (O_454,N_9294,N_9006);
and UO_455 (O_455,N_9562,N_8958);
or UO_456 (O_456,N_9409,N_9720);
or UO_457 (O_457,N_9107,N_7870);
xnor UO_458 (O_458,N_9359,N_7764);
and UO_459 (O_459,N_9148,N_7507);
and UO_460 (O_460,N_8012,N_8585);
or UO_461 (O_461,N_9607,N_9778);
nand UO_462 (O_462,N_9537,N_9579);
nand UO_463 (O_463,N_9576,N_7812);
nand UO_464 (O_464,N_9090,N_8049);
xor UO_465 (O_465,N_8852,N_8923);
and UO_466 (O_466,N_9812,N_9792);
xnor UO_467 (O_467,N_8644,N_9226);
or UO_468 (O_468,N_9197,N_8211);
xnor UO_469 (O_469,N_9833,N_9290);
and UO_470 (O_470,N_8816,N_8328);
xnor UO_471 (O_471,N_9034,N_7626);
or UO_472 (O_472,N_8470,N_8084);
and UO_473 (O_473,N_8539,N_7597);
nor UO_474 (O_474,N_8430,N_7864);
xnor UO_475 (O_475,N_8734,N_7738);
xnor UO_476 (O_476,N_7605,N_8996);
and UO_477 (O_477,N_9267,N_9924);
or UO_478 (O_478,N_8598,N_8480);
or UO_479 (O_479,N_9286,N_7729);
xnor UO_480 (O_480,N_9436,N_8681);
nor UO_481 (O_481,N_7767,N_8488);
nand UO_482 (O_482,N_7596,N_9320);
nand UO_483 (O_483,N_8408,N_8154);
nor UO_484 (O_484,N_8419,N_9012);
xor UO_485 (O_485,N_8035,N_8682);
nand UO_486 (O_486,N_9266,N_8744);
or UO_487 (O_487,N_7763,N_9513);
nand UO_488 (O_488,N_9729,N_8435);
and UO_489 (O_489,N_9071,N_8538);
and UO_490 (O_490,N_7781,N_8806);
or UO_491 (O_491,N_8655,N_8016);
nand UO_492 (O_492,N_9507,N_8861);
and UO_493 (O_493,N_8308,N_8573);
nor UO_494 (O_494,N_9275,N_8740);
nand UO_495 (O_495,N_8669,N_8365);
xor UO_496 (O_496,N_9182,N_7950);
or UO_497 (O_497,N_8868,N_9283);
nand UO_498 (O_498,N_8177,N_9694);
nand UO_499 (O_499,N_9349,N_8306);
or UO_500 (O_500,N_9781,N_8411);
nor UO_501 (O_501,N_9318,N_8421);
or UO_502 (O_502,N_9759,N_9201);
nand UO_503 (O_503,N_9358,N_9798);
nand UO_504 (O_504,N_7583,N_7653);
or UO_505 (O_505,N_7712,N_8567);
xnor UO_506 (O_506,N_8537,N_9789);
nor UO_507 (O_507,N_7761,N_8080);
nand UO_508 (O_508,N_9188,N_9973);
xnor UO_509 (O_509,N_9921,N_8088);
nor UO_510 (O_510,N_9072,N_7563);
nor UO_511 (O_511,N_7941,N_9509);
xnor UO_512 (O_512,N_9656,N_8030);
or UO_513 (O_513,N_7504,N_8763);
nand UO_514 (O_514,N_8099,N_9503);
nand UO_515 (O_515,N_8721,N_7813);
or UO_516 (O_516,N_8399,N_9857);
xor UO_517 (O_517,N_7888,N_9080);
nand UO_518 (O_518,N_8064,N_8982);
xor UO_519 (O_519,N_8452,N_9890);
xor UO_520 (O_520,N_8187,N_7544);
and UO_521 (O_521,N_9208,N_8256);
and UO_522 (O_522,N_8859,N_9003);
nor UO_523 (O_523,N_9913,N_7780);
nor UO_524 (O_524,N_9841,N_8444);
xnor UO_525 (O_525,N_9686,N_9419);
nor UO_526 (O_526,N_9433,N_8162);
or UO_527 (O_527,N_9806,N_7590);
or UO_528 (O_528,N_8199,N_9510);
nand UO_529 (O_529,N_9112,N_7521);
and UO_530 (O_530,N_8490,N_8770);
and UO_531 (O_531,N_8780,N_9238);
xnor UO_532 (O_532,N_9959,N_7607);
and UO_533 (O_533,N_8247,N_7844);
nor UO_534 (O_534,N_9264,N_8096);
or UO_535 (O_535,N_9661,N_8291);
nor UO_536 (O_536,N_9370,N_9705);
and UO_537 (O_537,N_9529,N_7998);
and UO_538 (O_538,N_8282,N_9070);
and UO_539 (O_539,N_8742,N_9957);
or UO_540 (O_540,N_8089,N_9241);
nand UO_541 (O_541,N_8161,N_8633);
xor UO_542 (O_542,N_9362,N_8412);
and UO_543 (O_543,N_7591,N_8953);
xor UO_544 (O_544,N_8285,N_8111);
nor UO_545 (O_545,N_7992,N_8437);
nor UO_546 (O_546,N_8751,N_9130);
nand UO_547 (O_547,N_8085,N_9154);
or UO_548 (O_548,N_8478,N_9589);
xnor UO_549 (O_549,N_7926,N_9452);
xor UO_550 (O_550,N_9085,N_8255);
xnor UO_551 (O_551,N_8340,N_8087);
xnor UO_552 (O_552,N_8336,N_8575);
xor UO_553 (O_553,N_8244,N_9377);
xnor UO_554 (O_554,N_9884,N_9944);
nor UO_555 (O_555,N_7892,N_9787);
xor UO_556 (O_556,N_7784,N_9416);
nand UO_557 (O_557,N_9760,N_9885);
xor UO_558 (O_558,N_9554,N_8584);
or UO_559 (O_559,N_9818,N_8086);
and UO_560 (O_560,N_8529,N_8095);
or UO_561 (O_561,N_9033,N_9939);
nand UO_562 (O_562,N_7960,N_8977);
and UO_563 (O_563,N_9233,N_9353);
nand UO_564 (O_564,N_8921,N_8917);
and UO_565 (O_565,N_9687,N_9632);
and UO_566 (O_566,N_9732,N_8805);
and UO_567 (O_567,N_8748,N_9100);
and UO_568 (O_568,N_8594,N_8857);
and UO_569 (O_569,N_8951,N_9768);
xnor UO_570 (O_570,N_8349,N_7742);
and UO_571 (O_571,N_8826,N_8789);
nor UO_572 (O_572,N_8888,N_8455);
xnor UO_573 (O_573,N_7995,N_9329);
or UO_574 (O_574,N_9079,N_9750);
xor UO_575 (O_575,N_9269,N_9937);
or UO_576 (O_576,N_8041,N_9478);
or UO_577 (O_577,N_9889,N_7934);
xnor UO_578 (O_578,N_7514,N_9950);
or UO_579 (O_579,N_7716,N_8758);
nand UO_580 (O_580,N_7925,N_9999);
and UO_581 (O_581,N_9958,N_8711);
and UO_582 (O_582,N_9255,N_9977);
nor UO_583 (O_583,N_9736,N_8090);
and UO_584 (O_584,N_8717,N_9102);
nor UO_585 (O_585,N_8658,N_7522);
and UO_586 (O_586,N_9753,N_8313);
nor UO_587 (O_587,N_8024,N_9989);
and UO_588 (O_588,N_9354,N_8176);
nor UO_589 (O_589,N_7546,N_8169);
nor UO_590 (O_590,N_8093,N_7788);
xnor UO_591 (O_591,N_7866,N_7555);
or UO_592 (O_592,N_9222,N_8559);
and UO_593 (O_593,N_8960,N_9647);
nand UO_594 (O_594,N_8869,N_8092);
and UO_595 (O_595,N_9271,N_9158);
and UO_596 (O_596,N_9134,N_7994);
xor UO_597 (O_597,N_8604,N_9908);
and UO_598 (O_598,N_8959,N_8155);
and UO_599 (O_599,N_9763,N_8259);
nor UO_600 (O_600,N_9247,N_8543);
xor UO_601 (O_601,N_9014,N_8393);
and UO_602 (O_602,N_8164,N_9701);
xor UO_603 (O_603,N_9145,N_8392);
xnor UO_604 (O_604,N_9471,N_7542);
xnor UO_605 (O_605,N_9439,N_9492);
nor UO_606 (O_606,N_8301,N_8878);
and UO_607 (O_607,N_9659,N_9926);
nand UO_608 (O_608,N_8776,N_7988);
or UO_609 (O_609,N_9321,N_8179);
and UO_610 (O_610,N_8417,N_9515);
nand UO_611 (O_611,N_8534,N_7990);
nor UO_612 (O_612,N_7951,N_9463);
and UO_613 (O_613,N_9835,N_9386);
xnor UO_614 (O_614,N_9919,N_9902);
nor UO_615 (O_615,N_9570,N_8823);
or UO_616 (O_616,N_9397,N_9448);
nor UO_617 (O_617,N_8007,N_9974);
xnor UO_618 (O_618,N_9039,N_9703);
xnor UO_619 (O_619,N_8223,N_7748);
nand UO_620 (O_620,N_7831,N_8486);
nor UO_621 (O_621,N_8560,N_7843);
xnor UO_622 (O_622,N_8521,N_9500);
xor UO_623 (O_623,N_9093,N_8948);
or UO_624 (O_624,N_9270,N_7883);
or UO_625 (O_625,N_8596,N_8566);
nand UO_626 (O_626,N_8525,N_8269);
nand UO_627 (O_627,N_8729,N_7769);
xnor UO_628 (O_628,N_9117,N_8858);
or UO_629 (O_629,N_8564,N_8297);
and UO_630 (O_630,N_7701,N_8364);
nand UO_631 (O_631,N_8701,N_8104);
nand UO_632 (O_632,N_9096,N_9235);
or UO_633 (O_633,N_7955,N_8931);
nor UO_634 (O_634,N_7765,N_9652);
nand UO_635 (O_635,N_9784,N_7754);
and UO_636 (O_636,N_9444,N_8895);
or UO_637 (O_637,N_9210,N_8714);
nor UO_638 (O_638,N_9059,N_7570);
nand UO_639 (O_639,N_9192,N_9456);
nand UO_640 (O_640,N_9026,N_8745);
nor UO_641 (O_641,N_7986,N_8950);
or UO_642 (O_642,N_9543,N_7594);
and UO_643 (O_643,N_8519,N_7777);
nor UO_644 (O_644,N_9636,N_8405);
and UO_645 (O_645,N_9474,N_9923);
nand UO_646 (O_646,N_9291,N_8884);
and UO_647 (O_647,N_8029,N_9344);
nor UO_648 (O_648,N_8845,N_9244);
xnor UO_649 (O_649,N_8268,N_9490);
nand UO_650 (O_650,N_7753,N_8109);
and UO_651 (O_651,N_9563,N_9533);
nand UO_652 (O_652,N_7929,N_8469);
or UO_653 (O_653,N_9385,N_9451);
and UO_654 (O_654,N_9022,N_9836);
or UO_655 (O_655,N_9304,N_8936);
or UO_656 (O_656,N_8010,N_9169);
nand UO_657 (O_657,N_8603,N_8781);
or UO_658 (O_658,N_9952,N_9755);
xnor UO_659 (O_659,N_8949,N_8757);
nand UO_660 (O_660,N_9367,N_8920);
nor UO_661 (O_661,N_7885,N_9230);
or UO_662 (O_662,N_8198,N_8180);
nor UO_663 (O_663,N_9104,N_9862);
or UO_664 (O_664,N_9366,N_9984);
and UO_665 (O_665,N_7936,N_8299);
nand UO_666 (O_666,N_7657,N_9581);
nor UO_667 (O_667,N_7683,N_8722);
nand UO_668 (O_668,N_7975,N_9272);
xor UO_669 (O_669,N_8460,N_8407);
xnor UO_670 (O_670,N_9018,N_9346);
or UO_671 (O_671,N_9858,N_8479);
nand UO_672 (O_672,N_7721,N_8883);
and UO_673 (O_673,N_8436,N_8044);
or UO_674 (O_674,N_9011,N_9137);
nand UO_675 (O_675,N_9183,N_7635);
xnor UO_676 (O_676,N_9853,N_8157);
or UO_677 (O_677,N_8663,N_7758);
and UO_678 (O_678,N_8125,N_8636);
nor UO_679 (O_679,N_7857,N_8014);
and UO_680 (O_680,N_8033,N_8839);
or UO_681 (O_681,N_9815,N_7973);
xor UO_682 (O_682,N_8767,N_9538);
and UO_683 (O_683,N_9128,N_7876);
nor UO_684 (O_684,N_8262,N_8300);
nand UO_685 (O_685,N_8930,N_7545);
nor UO_686 (O_686,N_8910,N_9980);
nand UO_687 (O_687,N_7987,N_8730);
xor UO_688 (O_688,N_8689,N_8498);
nand UO_689 (O_689,N_8675,N_7824);
and UO_690 (O_690,N_7965,N_7560);
nor UO_691 (O_691,N_7723,N_8457);
or UO_692 (O_692,N_7535,N_9560);
and UO_693 (O_693,N_8279,N_8724);
or UO_694 (O_694,N_7580,N_8232);
xnor UO_695 (O_695,N_7530,N_7915);
or UO_696 (O_696,N_9252,N_8492);
and UO_697 (O_697,N_8769,N_8048);
xnor UO_698 (O_698,N_9053,N_9502);
xor UO_699 (O_699,N_8697,N_9516);
nand UO_700 (O_700,N_7898,N_8051);
xor UO_701 (O_701,N_7515,N_7772);
xnor UO_702 (O_702,N_7566,N_7927);
nor UO_703 (O_703,N_7551,N_7858);
nand UO_704 (O_704,N_8384,N_8449);
and UO_705 (O_705,N_8330,N_9035);
or UO_706 (O_706,N_7540,N_9851);
nand UO_707 (O_707,N_8015,N_9390);
nor UO_708 (O_708,N_7648,N_9081);
nand UO_709 (O_709,N_9348,N_9811);
or UO_710 (O_710,N_8388,N_8914);
and UO_711 (O_711,N_9030,N_8432);
and UO_712 (O_712,N_7905,N_9121);
nor UO_713 (O_713,N_7623,N_9118);
or UO_714 (O_714,N_7985,N_8522);
xnor UO_715 (O_715,N_9951,N_8819);
nand UO_716 (O_716,N_9901,N_8900);
nand UO_717 (O_717,N_8002,N_7893);
nand UO_718 (O_718,N_8067,N_7599);
xnor UO_719 (O_719,N_8337,N_8726);
and UO_720 (O_720,N_9467,N_8333);
nand UO_721 (O_721,N_8768,N_8527);
nand UO_722 (O_722,N_9948,N_9551);
nor UO_723 (O_723,N_8343,N_7640);
or UO_724 (O_724,N_8204,N_9374);
or UO_725 (O_725,N_9063,N_9147);
nor UO_726 (O_726,N_7682,N_7652);
xnor UO_727 (O_727,N_9779,N_7531);
and UO_728 (O_728,N_9473,N_9166);
nor UO_729 (O_729,N_9119,N_9029);
and UO_730 (O_730,N_8991,N_8556);
nor UO_731 (O_731,N_8832,N_7600);
nor UO_732 (O_732,N_9834,N_8829);
and UO_733 (O_733,N_8329,N_8727);
or UO_734 (O_734,N_9949,N_9203);
or UO_735 (O_735,N_9105,N_8988);
or UO_736 (O_736,N_8008,N_8611);
and UO_737 (O_737,N_8670,N_8676);
and UO_738 (O_738,N_7593,N_8267);
xnor UO_739 (O_739,N_7981,N_9323);
or UO_740 (O_740,N_7962,N_9501);
nand UO_741 (O_741,N_8325,N_9707);
and UO_742 (O_742,N_8061,N_7579);
and UO_743 (O_743,N_9556,N_9719);
nor UO_744 (O_744,N_9577,N_8468);
xnor UO_745 (O_745,N_7647,N_9879);
xnor UO_746 (O_746,N_8409,N_8756);
nor UO_747 (O_747,N_8631,N_9667);
and UO_748 (O_748,N_9909,N_9016);
nor UO_749 (O_749,N_8212,N_9899);
or UO_750 (O_750,N_8280,N_7872);
xor UO_751 (O_751,N_7720,N_8552);
and UO_752 (O_752,N_8160,N_9905);
nor UO_753 (O_753,N_9820,N_9653);
nor UO_754 (O_754,N_7548,N_9106);
nand UO_755 (O_755,N_9175,N_9002);
nor UO_756 (O_756,N_7692,N_9572);
xnor UO_757 (O_757,N_8625,N_8815);
nand UO_758 (O_758,N_9669,N_7861);
or UO_759 (O_759,N_8050,N_8371);
or UO_760 (O_760,N_8352,N_9418);
nor UO_761 (O_761,N_9979,N_8302);
and UO_762 (O_762,N_7688,N_9328);
xnor UO_763 (O_763,N_8647,N_9472);
nor UO_764 (O_764,N_8289,N_9256);
or UO_765 (O_765,N_7792,N_9610);
nand UO_766 (O_766,N_9049,N_8932);
nand UO_767 (O_767,N_8696,N_9173);
and UO_768 (O_768,N_8142,N_9398);
or UO_769 (O_769,N_7826,N_7592);
and UO_770 (O_770,N_9698,N_9124);
or UO_771 (O_771,N_8115,N_9677);
nor UO_772 (O_772,N_9725,N_9828);
xnor UO_773 (O_773,N_9437,N_9810);
xor UO_774 (O_774,N_9232,N_8191);
nor UO_775 (O_775,N_8013,N_8063);
or UO_776 (O_776,N_8341,N_8835);
nor UO_777 (O_777,N_9722,N_8402);
nor UO_778 (O_778,N_9619,N_7737);
nor UO_779 (O_779,N_8502,N_8463);
nor UO_780 (O_780,N_8507,N_8747);
and UO_781 (O_781,N_8985,N_8332);
or UO_782 (O_782,N_7739,N_8963);
or UO_783 (O_783,N_7747,N_8181);
nor UO_784 (O_784,N_7694,N_7601);
and UO_785 (O_785,N_8217,N_9819);
and UO_786 (O_786,N_7733,N_8851);
xnor UO_787 (O_787,N_8524,N_8303);
nand UO_788 (O_788,N_9411,N_8445);
nor UO_789 (O_789,N_8022,N_9914);
or UO_790 (O_790,N_8188,N_8898);
or UO_791 (O_791,N_8547,N_9746);
or UO_792 (O_792,N_9213,N_9891);
or UO_793 (O_793,N_7817,N_9308);
or UO_794 (O_794,N_8565,N_9369);
and UO_795 (O_795,N_7774,N_9665);
or UO_796 (O_796,N_8374,N_9696);
nor UO_797 (O_797,N_7660,N_9655);
nor UO_798 (O_798,N_7991,N_9876);
xnor UO_799 (O_799,N_9388,N_9396);
and UO_800 (O_800,N_8593,N_9161);
nand UO_801 (O_801,N_7846,N_9475);
xor UO_802 (O_802,N_7714,N_9536);
nand UO_803 (O_803,N_8146,N_8570);
nand UO_804 (O_804,N_9679,N_7899);
nand UO_805 (O_805,N_9916,N_7553);
xor UO_806 (O_806,N_8075,N_8307);
or UO_807 (O_807,N_7634,N_9873);
nand UO_808 (O_808,N_8957,N_7952);
nor UO_809 (O_809,N_8208,N_8966);
nand UO_810 (O_810,N_8218,N_8579);
nand UO_811 (O_811,N_7572,N_9962);
nand UO_812 (O_812,N_8906,N_9897);
and UO_813 (O_813,N_9400,N_9723);
nand UO_814 (O_814,N_8123,N_7796);
xor UO_815 (O_815,N_8156,N_9296);
nand UO_816 (O_816,N_8915,N_9870);
and UO_817 (O_817,N_9383,N_9508);
or UO_818 (O_818,N_7849,N_9587);
and UO_819 (O_819,N_8540,N_7556);
and UO_820 (O_820,N_9931,N_8091);
nor UO_821 (O_821,N_9277,N_8017);
or UO_822 (O_822,N_9594,N_8975);
xnor UO_823 (O_823,N_7644,N_7752);
xnor UO_824 (O_824,N_9796,N_7618);
nand UO_825 (O_825,N_7853,N_9480);
nand UO_826 (O_826,N_7897,N_9313);
or UO_827 (O_827,N_9115,N_7845);
and UO_828 (O_828,N_7906,N_8257);
or UO_829 (O_829,N_7939,N_8621);
nor UO_830 (O_830,N_9207,N_7937);
nand UO_831 (O_831,N_8563,N_8335);
and UO_832 (O_832,N_9684,N_9345);
or UO_833 (O_833,N_8386,N_8554);
nor UO_834 (O_834,N_9550,N_8590);
and UO_835 (O_835,N_7856,N_9027);
or UO_836 (O_836,N_9322,N_9985);
nor UO_837 (O_837,N_8342,N_9114);
xor UO_838 (O_838,N_8134,N_8544);
or UO_839 (O_839,N_9420,N_9637);
or UO_840 (O_840,N_9956,N_8694);
and UO_841 (O_841,N_7681,N_8166);
and UO_842 (O_842,N_9678,N_8934);
xnor UO_843 (O_843,N_7646,N_8113);
and UO_844 (O_844,N_9704,N_9274);
or UO_845 (O_845,N_7519,N_7779);
and UO_846 (O_846,N_8425,N_9591);
xor UO_847 (O_847,N_8377,N_9064);
xor UO_848 (O_848,N_9483,N_9141);
xor UO_849 (O_849,N_7972,N_9431);
xnor UO_850 (O_850,N_9013,N_8615);
nand UO_851 (O_851,N_8533,N_8348);
xnor UO_852 (O_852,N_9564,N_9198);
and UO_853 (O_853,N_8253,N_7554);
nand UO_854 (O_854,N_8843,N_8643);
or UO_855 (O_855,N_7901,N_8999);
or UO_856 (O_856,N_9424,N_8997);
and UO_857 (O_857,N_7677,N_7617);
nand UO_858 (O_858,N_9545,N_8426);
nor UO_859 (O_859,N_7528,N_8372);
or UO_860 (O_860,N_8808,N_9263);
xnor UO_861 (O_861,N_8264,N_9888);
nor UO_862 (O_862,N_8824,N_9415);
nor UO_863 (O_863,N_7808,N_9527);
nand UO_864 (O_864,N_8446,N_8792);
and UO_865 (O_865,N_9910,N_8116);
and UO_866 (O_866,N_7643,N_8992);
xor UO_867 (O_867,N_7942,N_8222);
nand UO_868 (O_868,N_9082,N_8710);
xnor UO_869 (O_869,N_9360,N_8353);
xor UO_870 (O_870,N_7526,N_8698);
and UO_871 (O_871,N_8746,N_9848);
and UO_872 (O_872,N_8167,N_8881);
or UO_873 (O_873,N_9600,N_9176);
nand UO_874 (O_874,N_9975,N_7717);
and UO_875 (O_875,N_8679,N_9185);
and UO_876 (O_876,N_8794,N_7571);
nor UO_877 (O_877,N_9896,N_9103);
or UO_878 (O_878,N_9743,N_8318);
or UO_879 (O_879,N_8230,N_8183);
nor UO_880 (O_880,N_7517,N_7668);
and UO_881 (O_881,N_8023,N_8820);
xnor UO_882 (O_882,N_9842,N_9756);
and UO_883 (O_883,N_7963,N_9314);
nand UO_884 (O_884,N_9645,N_8503);
and UO_885 (O_885,N_9765,N_9237);
and UO_886 (O_886,N_7559,N_9657);
nor UO_887 (O_887,N_7770,N_9738);
or UO_888 (O_888,N_8891,N_7912);
nand UO_889 (O_889,N_7670,N_8072);
xor UO_890 (O_890,N_9206,N_7932);
xnor UO_891 (O_891,N_8876,N_8344);
xnor UO_892 (O_892,N_9132,N_9793);
nand UO_893 (O_893,N_9762,N_8415);
nand UO_894 (O_894,N_9990,N_8310);
or UO_895 (O_895,N_8172,N_8954);
and UO_896 (O_896,N_8630,N_8152);
nor UO_897 (O_897,N_8523,N_7665);
nand UO_898 (O_898,N_8404,N_8812);
nor UO_899 (O_899,N_9805,N_9180);
xor UO_900 (O_900,N_9299,N_9218);
xnor UO_901 (O_901,N_9708,N_7550);
or UO_902 (O_902,N_9605,N_7802);
or UO_903 (O_903,N_8355,N_7649);
nand UO_904 (O_904,N_9214,N_8387);
or UO_905 (O_905,N_8973,N_8716);
nand UO_906 (O_906,N_9292,N_8944);
nor UO_907 (O_907,N_9076,N_9976);
and UO_908 (O_908,N_7574,N_7686);
or UO_909 (O_909,N_9055,N_8713);
nand UO_910 (O_910,N_8807,N_8001);
nand UO_911 (O_911,N_8668,N_7862);
nand UO_912 (O_912,N_9426,N_7620);
nor UO_913 (O_913,N_9539,N_8700);
and UO_914 (O_914,N_9487,N_7760);
or UO_915 (O_915,N_8274,N_9892);
nand UO_916 (O_916,N_8403,N_8391);
or UO_917 (O_917,N_9379,N_7807);
or UO_918 (O_918,N_7584,N_9017);
xnor UO_919 (O_919,N_9863,N_9157);
xnor UO_920 (O_920,N_7819,N_8965);
nand UO_921 (O_921,N_7710,N_8495);
or UO_922 (O_922,N_9932,N_8509);
nand UO_923 (O_923,N_9280,N_8504);
nand UO_924 (O_924,N_8410,N_8601);
xor UO_925 (O_925,N_7775,N_8577);
or UO_926 (O_926,N_8189,N_7576);
nor UO_927 (O_927,N_8511,N_9394);
and UO_928 (O_928,N_9799,N_9730);
and UO_929 (O_929,N_9643,N_7759);
and UO_930 (O_930,N_9814,N_7855);
xnor UO_931 (O_931,N_8510,N_7533);
and UO_932 (O_932,N_9285,N_8158);
xnor UO_933 (O_933,N_8373,N_7890);
nor UO_934 (O_934,N_9282,N_7608);
nand UO_935 (O_935,N_8712,N_8201);
nand UO_936 (O_936,N_8863,N_7527);
nor UO_937 (O_937,N_9251,N_9193);
xor UO_938 (O_938,N_9052,N_8935);
or UO_939 (O_939,N_8706,N_9534);
and UO_940 (O_940,N_9150,N_9243);
or UO_941 (O_941,N_7565,N_9179);
and UO_942 (O_942,N_8234,N_8309);
xor UO_943 (O_943,N_9546,N_8583);
and UO_944 (O_944,N_8439,N_8219);
and UO_945 (O_945,N_8467,N_9152);
and UO_946 (O_946,N_8531,N_9571);
xor UO_947 (O_947,N_8569,N_8945);
nor UO_948 (O_948,N_9223,N_8699);
or UO_949 (O_949,N_9646,N_9123);
nor UO_950 (O_950,N_8036,N_9859);
or UO_951 (O_951,N_9380,N_7859);
nor UO_952 (O_952,N_7904,N_7800);
and UO_953 (O_953,N_9074,N_9867);
and UO_954 (O_954,N_8648,N_8277);
and UO_955 (O_955,N_8825,N_9125);
or UO_956 (O_956,N_8296,N_8802);
and UO_957 (O_957,N_9089,N_9528);
nand UO_958 (O_958,N_9469,N_7616);
nor UO_959 (O_959,N_9654,N_9776);
xor UO_960 (O_960,N_9001,N_8810);
xor UO_961 (O_961,N_7884,N_8771);
or UO_962 (O_962,N_8031,N_8894);
or UO_963 (O_963,N_9491,N_8173);
nand UO_964 (O_964,N_9993,N_8549);
or UO_965 (O_965,N_9942,N_7518);
or UO_966 (O_966,N_9061,N_9110);
xnor UO_967 (O_967,N_7693,N_8635);
or UO_968 (O_968,N_7709,N_9749);
and UO_969 (O_969,N_9464,N_8434);
and UO_970 (O_970,N_9757,N_8759);
and UO_971 (O_971,N_9204,N_7935);
and UO_972 (O_972,N_9146,N_8326);
or UO_973 (O_973,N_9742,N_8582);
or UO_974 (O_974,N_7516,N_8667);
xnor UO_975 (O_975,N_7719,N_8605);
xnor UO_976 (O_976,N_8578,N_8270);
nor UO_977 (O_977,N_8130,N_7655);
and UO_978 (O_978,N_9559,N_8456);
xnor UO_979 (O_979,N_9585,N_7782);
xor UO_980 (O_980,N_8128,N_8471);
or UO_981 (O_981,N_9405,N_9693);
and UO_982 (O_982,N_9310,N_9804);
xnor UO_983 (O_983,N_8862,N_9302);
xnor UO_984 (O_984,N_8197,N_9988);
nand UO_985 (O_985,N_9880,N_9486);
nor UO_986 (O_986,N_7839,N_8121);
xor UO_987 (O_987,N_9336,N_8213);
and UO_988 (O_988,N_8874,N_9005);
xor UO_989 (O_989,N_8990,N_8339);
nand UO_990 (O_990,N_7907,N_9253);
xor UO_991 (O_991,N_8363,N_8000);
nand UO_992 (O_992,N_8924,N_8245);
xor UO_993 (O_993,N_7794,N_9261);
xnor UO_994 (O_994,N_8983,N_7744);
nand UO_995 (O_995,N_8443,N_9307);
or UO_996 (O_996,N_9126,N_8346);
and UO_997 (O_997,N_9935,N_7953);
and UO_998 (O_998,N_9375,N_9479);
nor UO_999 (O_999,N_8702,N_8225);
and UO_1000 (O_1000,N_8796,N_7663);
and UO_1001 (O_1001,N_8942,N_9670);
and UO_1002 (O_1002,N_8065,N_9260);
nor UO_1003 (O_1003,N_8674,N_9540);
xor UO_1004 (O_1004,N_9455,N_8899);
or UO_1005 (O_1005,N_8610,N_8703);
or UO_1006 (O_1006,N_7666,N_8071);
or UO_1007 (O_1007,N_8860,N_8258);
xnor UO_1008 (O_1008,N_8465,N_8174);
and UO_1009 (O_1009,N_9767,N_7825);
or UO_1010 (O_1010,N_8249,N_9461);
and UO_1011 (O_1011,N_8376,N_8736);
xnor UO_1012 (O_1012,N_8887,N_8657);
nand UO_1013 (O_1013,N_7722,N_8351);
nor UO_1014 (O_1014,N_9918,N_9327);
nand UO_1015 (O_1015,N_8974,N_9403);
nor UO_1016 (O_1016,N_8872,N_8020);
nor UO_1017 (O_1017,N_7948,N_9582);
or UO_1018 (O_1018,N_7656,N_9599);
or UO_1019 (O_1019,N_9007,N_8731);
or UO_1020 (O_1020,N_8919,N_9098);
and UO_1021 (O_1021,N_8416,N_7642);
or UO_1022 (O_1022,N_8962,N_9972);
or UO_1023 (O_1023,N_8107,N_9031);
nand UO_1024 (O_1024,N_7889,N_9727);
and UO_1025 (O_1025,N_9877,N_8680);
or UO_1026 (O_1026,N_8634,N_7536);
xor UO_1027 (O_1027,N_9497,N_9347);
or UO_1028 (O_1028,N_9000,N_7735);
or UO_1029 (O_1029,N_9047,N_8545);
xnor UO_1030 (O_1030,N_8624,N_7728);
nor UO_1031 (O_1031,N_9350,N_8846);
and UO_1032 (O_1032,N_9827,N_8617);
and UO_1033 (O_1033,N_8442,N_9574);
or UO_1034 (O_1034,N_8752,N_8447);
and UO_1035 (O_1035,N_8284,N_9668);
and UO_1036 (O_1036,N_7558,N_8553);
and UO_1037 (O_1037,N_8896,N_8038);
or UO_1038 (O_1038,N_9392,N_8119);
or UO_1039 (O_1039,N_8800,N_9202);
or UO_1040 (O_1040,N_9886,N_9276);
and UO_1041 (O_1041,N_7511,N_7778);
nand UO_1042 (O_1042,N_9925,N_7680);
xnor UO_1043 (O_1043,N_8021,N_7900);
or UO_1044 (O_1044,N_9967,N_8848);
and UO_1045 (O_1045,N_8705,N_8028);
nor UO_1046 (O_1046,N_8046,N_8367);
nand UO_1047 (O_1047,N_7697,N_7575);
or UO_1048 (O_1048,N_9936,N_8732);
nand UO_1049 (O_1049,N_8420,N_9122);
or UO_1050 (O_1050,N_8263,N_8897);
or UO_1051 (O_1051,N_8661,N_7989);
or UO_1052 (O_1052,N_9864,N_9596);
or UO_1053 (O_1053,N_9558,N_9281);
or UO_1054 (O_1054,N_9780,N_9056);
or UO_1055 (O_1055,N_7637,N_8606);
nor UO_1056 (O_1056,N_9043,N_7930);
xnor UO_1057 (O_1057,N_9945,N_8691);
or UO_1058 (O_1058,N_8032,N_7913);
or UO_1059 (O_1059,N_8737,N_8074);
and UO_1060 (O_1060,N_9567,N_7509);
xnor UO_1061 (O_1061,N_8847,N_9991);
nand UO_1062 (O_1062,N_8185,N_9170);
nand UO_1063 (O_1063,N_8518,N_7971);
nor UO_1064 (O_1064,N_9662,N_7614);
xor UO_1065 (O_1065,N_7564,N_8541);
and UO_1066 (O_1066,N_9625,N_8192);
and UO_1067 (O_1067,N_8555,N_8755);
or UO_1068 (O_1068,N_9075,N_8485);
nand UO_1069 (O_1069,N_8688,N_9453);
or UO_1070 (O_1070,N_7674,N_9801);
nand UO_1071 (O_1071,N_8052,N_9664);
nor UO_1072 (O_1072,N_9060,N_8273);
xor UO_1073 (O_1073,N_8317,N_8871);
nor UO_1074 (O_1074,N_8163,N_8641);
or UO_1075 (O_1075,N_8678,N_8118);
or UO_1076 (O_1076,N_8911,N_7732);
nor UO_1077 (O_1077,N_9584,N_7886);
nor UO_1078 (O_1078,N_8039,N_9162);
nor UO_1079 (O_1079,N_8613,N_9520);
xnor UO_1080 (O_1080,N_8754,N_9929);
nor UO_1081 (O_1081,N_9156,N_9399);
and UO_1082 (O_1082,N_8822,N_7650);
nor UO_1083 (O_1083,N_8390,N_7755);
nor UO_1084 (O_1084,N_9217,N_8666);
and UO_1085 (O_1085,N_8271,N_7525);
xnor UO_1086 (O_1086,N_8034,N_9086);
nor UO_1087 (O_1087,N_8323,N_8671);
nand UO_1088 (O_1088,N_8082,N_8690);
nor UO_1089 (O_1089,N_7512,N_9716);
nand UO_1090 (O_1090,N_8475,N_8866);
or UO_1091 (O_1091,N_9633,N_7944);
or UO_1092 (O_1092,N_8831,N_9699);
or UO_1093 (O_1093,N_8939,N_9595);
or UO_1094 (O_1094,N_9268,N_9062);
and UO_1095 (O_1095,N_9326,N_7708);
nor UO_1096 (O_1096,N_8018,N_9715);
and UO_1097 (O_1097,N_8505,N_8627);
nand UO_1098 (O_1098,N_9438,N_7629);
nor UO_1099 (O_1099,N_8662,N_7671);
or UO_1100 (O_1100,N_9603,N_9733);
nand UO_1101 (O_1101,N_8070,N_7895);
or UO_1102 (O_1102,N_8777,N_8005);
nor UO_1103 (O_1103,N_7621,N_9168);
xnor UO_1104 (O_1104,N_9352,N_9015);
xnor UO_1105 (O_1105,N_8608,N_8114);
xor UO_1106 (O_1106,N_7791,N_9737);
nand UO_1107 (O_1107,N_9575,N_8725);
xor UO_1108 (O_1108,N_8623,N_7787);
nor UO_1109 (O_1109,N_9981,N_8190);
nor UO_1110 (O_1110,N_9209,N_8120);
and UO_1111 (O_1111,N_8127,N_8153);
and UO_1112 (O_1112,N_7718,N_9996);
nand UO_1113 (O_1113,N_7978,N_7830);
and UO_1114 (O_1114,N_7673,N_7966);
and UO_1115 (O_1115,N_9215,N_7628);
xor UO_1116 (O_1116,N_9057,N_9745);
or UO_1117 (O_1117,N_8685,N_8193);
xor UO_1118 (O_1118,N_9712,N_9613);
or UO_1119 (O_1119,N_7806,N_7604);
or UO_1120 (O_1120,N_8281,N_7803);
nand UO_1121 (O_1121,N_7882,N_8971);
nor UO_1122 (O_1122,N_8787,N_9212);
and UO_1123 (O_1123,N_9883,N_9181);
or UO_1124 (O_1124,N_7746,N_8818);
nor UO_1125 (O_1125,N_7724,N_9832);
and UO_1126 (O_1126,N_7757,N_8241);
nor UO_1127 (O_1127,N_8224,N_9021);
nor UO_1128 (O_1128,N_9881,N_9159);
xnor UO_1129 (O_1129,N_7627,N_9036);
or UO_1130 (O_1130,N_8025,N_8418);
nor UO_1131 (O_1131,N_9933,N_8354);
xor UO_1132 (O_1132,N_8828,N_9466);
nor UO_1133 (O_1133,N_9216,N_8801);
nand UO_1134 (O_1134,N_8750,N_7745);
nand UO_1135 (O_1135,N_7894,N_8536);
nor UO_1136 (O_1136,N_8684,N_8850);
and UO_1137 (O_1137,N_7598,N_9535);
nand UO_1138 (O_1138,N_7586,N_9153);
xnor UO_1139 (O_1139,N_8370,N_7547);
or UO_1140 (O_1140,N_8473,N_7943);
nor UO_1141 (O_1141,N_7513,N_8571);
nand UO_1142 (O_1142,N_7848,N_7828);
xor UO_1143 (O_1143,N_8489,N_7875);
nand UO_1144 (O_1144,N_9465,N_8202);
nand UO_1145 (O_1145,N_9068,N_9822);
xor UO_1146 (O_1146,N_7505,N_9771);
nand UO_1147 (O_1147,N_8304,N_9837);
xnor UO_1148 (O_1148,N_8145,N_9893);
and UO_1149 (O_1149,N_9856,N_9542);
nor UO_1150 (O_1150,N_7881,N_8150);
and UO_1151 (O_1151,N_8433,N_7938);
nand UO_1152 (O_1152,N_9250,N_8561);
or UO_1153 (O_1153,N_7977,N_9387);
or UO_1154 (O_1154,N_8186,N_8772);
nor UO_1155 (O_1155,N_7715,N_9739);
nand UO_1156 (O_1156,N_9430,N_7713);
nand UO_1157 (O_1157,N_9608,N_9111);
xnor UO_1158 (O_1158,N_8248,N_8762);
or UO_1159 (O_1159,N_9298,N_7850);
and UO_1160 (O_1160,N_7705,N_7567);
nand UO_1161 (O_1161,N_9120,N_8487);
nand UO_1162 (O_1162,N_9953,N_9194);
xnor UO_1163 (O_1163,N_7983,N_9095);
xnor UO_1164 (O_1164,N_8692,N_8986);
xnor UO_1165 (O_1165,N_9381,N_8775);
nand UO_1166 (O_1166,N_7672,N_7730);
nand UO_1167 (O_1167,N_8006,N_9025);
and UO_1168 (O_1168,N_8673,N_8629);
nor UO_1169 (O_1169,N_9190,N_8246);
nor UO_1170 (O_1170,N_9671,N_8078);
nor UO_1171 (O_1171,N_8660,N_9630);
or UO_1172 (O_1172,N_9598,N_7924);
and UO_1173 (O_1173,N_9278,N_9364);
or UO_1174 (O_1174,N_8382,N_9681);
xor UO_1175 (O_1175,N_9429,N_9961);
xor UO_1176 (O_1176,N_9648,N_9199);
or UO_1177 (O_1177,N_9066,N_9447);
and UO_1178 (O_1178,N_9821,N_9713);
nand UO_1179 (O_1179,N_7700,N_9136);
and UO_1180 (O_1180,N_8283,N_8139);
nor UO_1181 (O_1181,N_9408,N_9236);
or UO_1182 (O_1182,N_9624,N_8499);
nand UO_1183 (O_1183,N_9109,N_9735);
nand UO_1184 (O_1184,N_9404,N_8976);
nand UO_1185 (O_1185,N_8586,N_8733);
and UO_1186 (O_1186,N_8528,N_9219);
nor UO_1187 (O_1187,N_9934,N_8609);
nand UO_1188 (O_1188,N_7860,N_8011);
nand UO_1189 (O_1189,N_9425,N_9004);
and UO_1190 (O_1190,N_9312,N_8126);
xor UO_1191 (O_1191,N_8140,N_7829);
xor UO_1192 (O_1192,N_9825,N_9907);
nand UO_1193 (O_1193,N_8840,N_9127);
xor UO_1194 (O_1194,N_8047,N_7702);
or UO_1195 (O_1195,N_8413,N_9108);
and UO_1196 (O_1196,N_7639,N_7731);
nor UO_1197 (O_1197,N_7874,N_9714);
or UO_1198 (O_1198,N_8004,N_7789);
and UO_1199 (O_1199,N_8622,N_8937);
and UO_1200 (O_1200,N_9376,N_8821);
nand UO_1201 (O_1201,N_9855,N_8749);
and UO_1202 (O_1202,N_8867,N_8989);
nand UO_1203 (O_1203,N_9495,N_8646);
and UO_1204 (O_1204,N_7506,N_9854);
and UO_1205 (O_1205,N_9666,N_9549);
nand UO_1206 (O_1206,N_8799,N_7736);
and UO_1207 (O_1207,N_8833,N_7805);
or UO_1208 (O_1208,N_8350,N_9442);
xnor UO_1209 (O_1209,N_8497,N_8797);
and UO_1210 (O_1210,N_9144,N_7588);
or UO_1211 (O_1211,N_9616,N_8589);
nand UO_1212 (O_1212,N_8440,N_8842);
and UO_1213 (O_1213,N_9882,N_7841);
nand UO_1214 (O_1214,N_8054,N_8854);
xnor UO_1215 (O_1215,N_7837,N_8542);
or UO_1216 (O_1216,N_7537,N_9830);
or UO_1217 (O_1217,N_8834,N_8784);
and UO_1218 (O_1218,N_8880,N_9706);
or UO_1219 (O_1219,N_9786,N_7704);
and UO_1220 (O_1220,N_8970,N_8743);
xnor UO_1221 (O_1221,N_9019,N_9782);
xor UO_1222 (O_1222,N_8400,N_7847);
nand UO_1223 (O_1223,N_8664,N_8059);
nand UO_1224 (O_1224,N_7865,N_9357);
nand UO_1225 (O_1225,N_7581,N_9337);
xor UO_1226 (O_1226,N_9289,N_8686);
nor UO_1227 (O_1227,N_7685,N_8194);
xor UO_1228 (O_1228,N_9943,N_8907);
or UO_1229 (O_1229,N_9257,N_7691);
xor UO_1230 (O_1230,N_9434,N_8043);
nand UO_1231 (O_1231,N_7923,N_8947);
and UO_1232 (O_1232,N_8616,N_7654);
and UO_1233 (O_1233,N_8357,N_8838);
xnor UO_1234 (O_1234,N_7633,N_9046);
xnor UO_1235 (O_1235,N_8055,N_9741);
and UO_1236 (O_1236,N_9524,N_9894);
and UO_1237 (O_1237,N_9189,N_8105);
or UO_1238 (O_1238,N_8260,N_9371);
nand UO_1239 (O_1239,N_7902,N_7638);
nor UO_1240 (O_1240,N_9258,N_7822);
nor UO_1241 (O_1241,N_9488,N_8462);
and UO_1242 (O_1242,N_7541,N_8905);
nor UO_1243 (O_1243,N_7529,N_9050);
nor UO_1244 (O_1244,N_8060,N_7669);
and UO_1245 (O_1245,N_9838,N_8841);
nand UO_1246 (O_1246,N_8369,N_9443);
xor UO_1247 (O_1247,N_7793,N_8592);
or UO_1248 (O_1248,N_7993,N_8735);
and UO_1249 (O_1249,N_9149,N_7970);
and UO_1250 (O_1250,N_9304,N_9213);
nand UO_1251 (O_1251,N_8814,N_9197);
or UO_1252 (O_1252,N_8396,N_8132);
and UO_1253 (O_1253,N_9286,N_9554);
or UO_1254 (O_1254,N_7579,N_9804);
xnor UO_1255 (O_1255,N_8061,N_9143);
xnor UO_1256 (O_1256,N_7835,N_9002);
xnor UO_1257 (O_1257,N_9239,N_8605);
or UO_1258 (O_1258,N_8059,N_9132);
xnor UO_1259 (O_1259,N_8645,N_8853);
nand UO_1260 (O_1260,N_8684,N_8132);
nor UO_1261 (O_1261,N_8261,N_9852);
and UO_1262 (O_1262,N_9637,N_8086);
xnor UO_1263 (O_1263,N_9490,N_7500);
or UO_1264 (O_1264,N_9388,N_8727);
nand UO_1265 (O_1265,N_8276,N_9082);
or UO_1266 (O_1266,N_7721,N_8720);
nand UO_1267 (O_1267,N_9988,N_9412);
and UO_1268 (O_1268,N_9300,N_9515);
or UO_1269 (O_1269,N_7699,N_8193);
or UO_1270 (O_1270,N_9886,N_7535);
xor UO_1271 (O_1271,N_9660,N_7811);
xor UO_1272 (O_1272,N_9037,N_8083);
or UO_1273 (O_1273,N_8843,N_8737);
or UO_1274 (O_1274,N_8149,N_8788);
xnor UO_1275 (O_1275,N_8252,N_9840);
or UO_1276 (O_1276,N_7544,N_9696);
xor UO_1277 (O_1277,N_8632,N_7811);
xnor UO_1278 (O_1278,N_8349,N_8399);
and UO_1279 (O_1279,N_9755,N_9770);
xor UO_1280 (O_1280,N_9052,N_8949);
or UO_1281 (O_1281,N_9815,N_9501);
or UO_1282 (O_1282,N_7723,N_8417);
nand UO_1283 (O_1283,N_8938,N_7859);
or UO_1284 (O_1284,N_9476,N_9110);
or UO_1285 (O_1285,N_8582,N_8651);
nor UO_1286 (O_1286,N_8531,N_9907);
nor UO_1287 (O_1287,N_8337,N_8764);
nand UO_1288 (O_1288,N_8949,N_9605);
nand UO_1289 (O_1289,N_8118,N_8903);
nor UO_1290 (O_1290,N_9930,N_8891);
or UO_1291 (O_1291,N_8329,N_8127);
nand UO_1292 (O_1292,N_8732,N_7621);
and UO_1293 (O_1293,N_9157,N_9621);
xnor UO_1294 (O_1294,N_8223,N_9863);
or UO_1295 (O_1295,N_7587,N_9193);
nand UO_1296 (O_1296,N_8865,N_9845);
nor UO_1297 (O_1297,N_7820,N_8830);
nand UO_1298 (O_1298,N_9739,N_8862);
nor UO_1299 (O_1299,N_9447,N_8076);
nand UO_1300 (O_1300,N_8978,N_8036);
nor UO_1301 (O_1301,N_8157,N_9117);
or UO_1302 (O_1302,N_8373,N_8413);
and UO_1303 (O_1303,N_9754,N_9738);
nor UO_1304 (O_1304,N_8806,N_9028);
or UO_1305 (O_1305,N_9839,N_8653);
xor UO_1306 (O_1306,N_8258,N_9220);
xnor UO_1307 (O_1307,N_8254,N_8471);
or UO_1308 (O_1308,N_7575,N_7800);
nor UO_1309 (O_1309,N_9996,N_7592);
nand UO_1310 (O_1310,N_9599,N_8392);
xor UO_1311 (O_1311,N_9819,N_9685);
and UO_1312 (O_1312,N_8023,N_8205);
nor UO_1313 (O_1313,N_7540,N_7830);
and UO_1314 (O_1314,N_7969,N_8756);
and UO_1315 (O_1315,N_7890,N_9159);
or UO_1316 (O_1316,N_9288,N_9510);
nand UO_1317 (O_1317,N_9454,N_8178);
xnor UO_1318 (O_1318,N_8657,N_9941);
or UO_1319 (O_1319,N_8590,N_9369);
and UO_1320 (O_1320,N_8533,N_8646);
nor UO_1321 (O_1321,N_8428,N_9186);
nand UO_1322 (O_1322,N_8933,N_8284);
xnor UO_1323 (O_1323,N_9845,N_7911);
and UO_1324 (O_1324,N_8321,N_7767);
nor UO_1325 (O_1325,N_9256,N_9701);
nand UO_1326 (O_1326,N_8336,N_9930);
or UO_1327 (O_1327,N_8619,N_8666);
nand UO_1328 (O_1328,N_8331,N_9443);
xor UO_1329 (O_1329,N_9777,N_7870);
nand UO_1330 (O_1330,N_9737,N_8620);
and UO_1331 (O_1331,N_9329,N_9242);
and UO_1332 (O_1332,N_7561,N_8955);
nand UO_1333 (O_1333,N_9676,N_7817);
or UO_1334 (O_1334,N_8533,N_8545);
and UO_1335 (O_1335,N_9370,N_8663);
and UO_1336 (O_1336,N_8227,N_8963);
or UO_1337 (O_1337,N_8101,N_9388);
nor UO_1338 (O_1338,N_9171,N_8668);
nand UO_1339 (O_1339,N_7538,N_9737);
nand UO_1340 (O_1340,N_9050,N_8332);
and UO_1341 (O_1341,N_7545,N_8026);
and UO_1342 (O_1342,N_9179,N_9711);
nor UO_1343 (O_1343,N_8033,N_8061);
nor UO_1344 (O_1344,N_8220,N_8998);
nor UO_1345 (O_1345,N_7704,N_8247);
nand UO_1346 (O_1346,N_8206,N_8923);
xnor UO_1347 (O_1347,N_8072,N_8320);
or UO_1348 (O_1348,N_9520,N_8077);
or UO_1349 (O_1349,N_9249,N_7672);
or UO_1350 (O_1350,N_9586,N_9900);
nor UO_1351 (O_1351,N_9967,N_7530);
or UO_1352 (O_1352,N_9281,N_9146);
nand UO_1353 (O_1353,N_8638,N_9150);
nor UO_1354 (O_1354,N_9130,N_9641);
nand UO_1355 (O_1355,N_9291,N_9814);
or UO_1356 (O_1356,N_8929,N_9992);
xor UO_1357 (O_1357,N_9384,N_7969);
nand UO_1358 (O_1358,N_9549,N_7528);
and UO_1359 (O_1359,N_8326,N_9870);
or UO_1360 (O_1360,N_9187,N_8334);
or UO_1361 (O_1361,N_8845,N_8126);
xor UO_1362 (O_1362,N_7814,N_9219);
nor UO_1363 (O_1363,N_9297,N_8951);
nor UO_1364 (O_1364,N_9147,N_9127);
nor UO_1365 (O_1365,N_8228,N_8858);
xor UO_1366 (O_1366,N_8628,N_8313);
nor UO_1367 (O_1367,N_9561,N_7576);
and UO_1368 (O_1368,N_9734,N_8175);
and UO_1369 (O_1369,N_9970,N_9232);
nor UO_1370 (O_1370,N_8191,N_7816);
nand UO_1371 (O_1371,N_9226,N_8730);
or UO_1372 (O_1372,N_8641,N_8690);
nand UO_1373 (O_1373,N_7674,N_7790);
or UO_1374 (O_1374,N_7757,N_7906);
or UO_1375 (O_1375,N_8162,N_8307);
xnor UO_1376 (O_1376,N_8079,N_9543);
nand UO_1377 (O_1377,N_9383,N_8270);
nor UO_1378 (O_1378,N_8016,N_7769);
xor UO_1379 (O_1379,N_9987,N_8279);
and UO_1380 (O_1380,N_8874,N_9636);
and UO_1381 (O_1381,N_8413,N_7767);
xnor UO_1382 (O_1382,N_8012,N_7935);
nand UO_1383 (O_1383,N_9702,N_8262);
nor UO_1384 (O_1384,N_8053,N_8336);
and UO_1385 (O_1385,N_9221,N_9734);
nand UO_1386 (O_1386,N_8886,N_9315);
or UO_1387 (O_1387,N_9511,N_9294);
and UO_1388 (O_1388,N_7683,N_8337);
nor UO_1389 (O_1389,N_8508,N_8111);
and UO_1390 (O_1390,N_9235,N_8991);
nor UO_1391 (O_1391,N_9280,N_8024);
and UO_1392 (O_1392,N_9812,N_9185);
and UO_1393 (O_1393,N_7792,N_9211);
and UO_1394 (O_1394,N_9904,N_8654);
or UO_1395 (O_1395,N_9157,N_9735);
nor UO_1396 (O_1396,N_9863,N_8757);
nand UO_1397 (O_1397,N_7627,N_8924);
xor UO_1398 (O_1398,N_7845,N_9364);
or UO_1399 (O_1399,N_7928,N_9753);
nor UO_1400 (O_1400,N_8811,N_8067);
and UO_1401 (O_1401,N_9474,N_9310);
nand UO_1402 (O_1402,N_8533,N_9462);
or UO_1403 (O_1403,N_9333,N_8080);
xor UO_1404 (O_1404,N_9801,N_7582);
nand UO_1405 (O_1405,N_8783,N_9839);
or UO_1406 (O_1406,N_9790,N_8713);
or UO_1407 (O_1407,N_7693,N_8941);
nor UO_1408 (O_1408,N_8571,N_9635);
nor UO_1409 (O_1409,N_8747,N_7548);
and UO_1410 (O_1410,N_8391,N_9715);
xnor UO_1411 (O_1411,N_9420,N_9012);
and UO_1412 (O_1412,N_8655,N_9516);
nor UO_1413 (O_1413,N_9070,N_9211);
xnor UO_1414 (O_1414,N_8289,N_8793);
or UO_1415 (O_1415,N_7666,N_8931);
and UO_1416 (O_1416,N_7700,N_9244);
nor UO_1417 (O_1417,N_9339,N_7753);
and UO_1418 (O_1418,N_8413,N_8001);
xor UO_1419 (O_1419,N_7804,N_9478);
nor UO_1420 (O_1420,N_7808,N_9811);
nor UO_1421 (O_1421,N_9451,N_9164);
or UO_1422 (O_1422,N_9239,N_7740);
nor UO_1423 (O_1423,N_9708,N_9517);
nand UO_1424 (O_1424,N_7823,N_8819);
and UO_1425 (O_1425,N_7571,N_8247);
nor UO_1426 (O_1426,N_9153,N_8145);
nand UO_1427 (O_1427,N_9105,N_9223);
nand UO_1428 (O_1428,N_9611,N_8822);
and UO_1429 (O_1429,N_9492,N_8179);
or UO_1430 (O_1430,N_9178,N_9938);
xnor UO_1431 (O_1431,N_8634,N_8759);
nand UO_1432 (O_1432,N_8221,N_8084);
or UO_1433 (O_1433,N_7874,N_8743);
and UO_1434 (O_1434,N_8886,N_7599);
nand UO_1435 (O_1435,N_8083,N_8924);
xor UO_1436 (O_1436,N_7981,N_8706);
and UO_1437 (O_1437,N_9271,N_8663);
and UO_1438 (O_1438,N_9802,N_8898);
and UO_1439 (O_1439,N_8340,N_7856);
xnor UO_1440 (O_1440,N_7843,N_9969);
nor UO_1441 (O_1441,N_8620,N_8390);
and UO_1442 (O_1442,N_9018,N_7941);
nand UO_1443 (O_1443,N_9955,N_8536);
xnor UO_1444 (O_1444,N_8455,N_9098);
or UO_1445 (O_1445,N_8704,N_7851);
or UO_1446 (O_1446,N_8641,N_7734);
nor UO_1447 (O_1447,N_9259,N_7650);
or UO_1448 (O_1448,N_8474,N_9179);
or UO_1449 (O_1449,N_8680,N_9364);
nand UO_1450 (O_1450,N_9730,N_9162);
and UO_1451 (O_1451,N_9412,N_9331);
nor UO_1452 (O_1452,N_7916,N_7664);
and UO_1453 (O_1453,N_9935,N_8397);
and UO_1454 (O_1454,N_8768,N_7851);
or UO_1455 (O_1455,N_8106,N_9072);
xor UO_1456 (O_1456,N_8805,N_8016);
nand UO_1457 (O_1457,N_8903,N_8647);
xor UO_1458 (O_1458,N_9807,N_9780);
nor UO_1459 (O_1459,N_9419,N_9201);
nor UO_1460 (O_1460,N_8796,N_7554);
and UO_1461 (O_1461,N_9662,N_9295);
xor UO_1462 (O_1462,N_8118,N_9567);
xor UO_1463 (O_1463,N_7550,N_9565);
xnor UO_1464 (O_1464,N_9178,N_9752);
nand UO_1465 (O_1465,N_7595,N_8241);
xnor UO_1466 (O_1466,N_8239,N_8370);
and UO_1467 (O_1467,N_7675,N_8158);
xnor UO_1468 (O_1468,N_8131,N_7542);
or UO_1469 (O_1469,N_8287,N_8998);
or UO_1470 (O_1470,N_8650,N_9205);
nor UO_1471 (O_1471,N_8168,N_8755);
nor UO_1472 (O_1472,N_9519,N_8927);
and UO_1473 (O_1473,N_8322,N_9896);
xor UO_1474 (O_1474,N_8167,N_9950);
nor UO_1475 (O_1475,N_8809,N_8131);
or UO_1476 (O_1476,N_7588,N_8390);
and UO_1477 (O_1477,N_9858,N_9165);
nand UO_1478 (O_1478,N_9110,N_8813);
and UO_1479 (O_1479,N_7840,N_9773);
nor UO_1480 (O_1480,N_9595,N_9202);
nand UO_1481 (O_1481,N_9475,N_7698);
xor UO_1482 (O_1482,N_9218,N_8040);
or UO_1483 (O_1483,N_7604,N_7941);
or UO_1484 (O_1484,N_7506,N_8557);
or UO_1485 (O_1485,N_8988,N_7694);
or UO_1486 (O_1486,N_8137,N_7640);
xor UO_1487 (O_1487,N_9832,N_9046);
and UO_1488 (O_1488,N_8373,N_9068);
or UO_1489 (O_1489,N_9812,N_8278);
nand UO_1490 (O_1490,N_7831,N_9347);
and UO_1491 (O_1491,N_9377,N_9000);
nand UO_1492 (O_1492,N_7615,N_9223);
nand UO_1493 (O_1493,N_8093,N_9440);
or UO_1494 (O_1494,N_9824,N_8662);
and UO_1495 (O_1495,N_8184,N_7824);
nand UO_1496 (O_1496,N_9145,N_8957);
or UO_1497 (O_1497,N_8628,N_8666);
and UO_1498 (O_1498,N_9429,N_9171);
xor UO_1499 (O_1499,N_8877,N_9439);
endmodule