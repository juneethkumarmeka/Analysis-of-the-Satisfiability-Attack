module basic_500_3000_500_6_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_262,In_250);
xnor U1 (N_1,In_198,In_466);
or U2 (N_2,In_6,In_149);
xor U3 (N_3,In_209,In_84);
nor U4 (N_4,In_307,In_311);
nor U5 (N_5,In_168,In_202);
or U6 (N_6,In_496,In_458);
nand U7 (N_7,In_179,In_86);
nand U8 (N_8,In_288,In_54);
nor U9 (N_9,In_428,In_349);
xor U10 (N_10,In_482,In_328);
and U11 (N_11,In_479,In_368);
nand U12 (N_12,In_219,In_48);
xnor U13 (N_13,In_254,In_358);
or U14 (N_14,In_227,In_5);
and U15 (N_15,In_108,In_419);
nand U16 (N_16,In_85,In_277);
xor U17 (N_17,In_304,In_295);
nor U18 (N_18,In_140,In_370);
nand U19 (N_19,In_470,In_398);
and U20 (N_20,In_119,In_240);
nor U21 (N_21,In_389,In_352);
nor U22 (N_22,In_210,In_266);
nor U23 (N_23,In_20,In_498);
nand U24 (N_24,In_180,In_95);
nor U25 (N_25,In_445,In_226);
nor U26 (N_26,In_111,In_245);
xnor U27 (N_27,In_252,In_120);
nor U28 (N_28,In_382,In_36);
nand U29 (N_29,In_193,In_185);
xor U30 (N_30,In_484,In_153);
xnor U31 (N_31,In_132,In_53);
nor U32 (N_32,In_112,In_261);
nor U33 (N_33,In_271,In_115);
nand U34 (N_34,In_380,In_93);
or U35 (N_35,In_281,In_124);
nand U36 (N_36,In_497,In_127);
nor U37 (N_37,In_15,In_222);
or U38 (N_38,In_367,In_372);
xnor U39 (N_39,In_291,In_18);
xor U40 (N_40,In_74,In_265);
or U41 (N_41,In_89,In_206);
or U42 (N_42,In_467,In_437);
nand U43 (N_43,In_57,In_29);
and U44 (N_44,In_465,In_139);
nand U45 (N_45,In_489,In_280);
and U46 (N_46,In_199,In_224);
xor U47 (N_47,In_107,In_19);
or U48 (N_48,In_73,In_371);
nand U49 (N_49,In_378,In_141);
or U50 (N_50,In_71,In_96);
or U51 (N_51,In_303,In_109);
or U52 (N_52,In_456,In_259);
nor U53 (N_53,In_285,In_369);
xnor U54 (N_54,In_460,In_208);
nor U55 (N_55,In_101,In_172);
xor U56 (N_56,In_409,In_282);
xor U57 (N_57,In_312,In_420);
and U58 (N_58,In_381,In_346);
xnor U59 (N_59,In_8,In_454);
nand U60 (N_60,In_39,In_411);
and U61 (N_61,In_0,In_205);
xnor U62 (N_62,In_402,In_329);
or U63 (N_63,In_194,In_313);
nand U64 (N_64,In_204,In_330);
and U65 (N_65,In_87,In_302);
and U66 (N_66,In_322,In_9);
or U67 (N_67,In_401,In_175);
nand U68 (N_68,In_491,In_196);
xnor U69 (N_69,In_231,In_97);
nand U70 (N_70,In_394,In_464);
nand U71 (N_71,In_481,In_293);
nor U72 (N_72,In_338,In_326);
or U73 (N_73,In_455,In_238);
and U74 (N_74,In_365,In_417);
nand U75 (N_75,In_121,In_52);
nor U76 (N_76,In_397,In_413);
xor U77 (N_77,In_333,In_123);
xor U78 (N_78,In_493,In_220);
nand U79 (N_79,In_343,In_263);
nor U80 (N_80,In_116,In_396);
xnor U81 (N_81,In_13,In_450);
or U82 (N_82,In_64,In_348);
nor U83 (N_83,In_106,In_197);
or U84 (N_84,In_237,In_294);
nand U85 (N_85,In_340,In_427);
nor U86 (N_86,In_395,In_192);
nand U87 (N_87,In_190,In_225);
or U88 (N_88,In_327,In_159);
xor U89 (N_89,In_158,In_213);
and U90 (N_90,In_228,In_289);
nor U91 (N_91,In_157,In_81);
nor U92 (N_92,In_21,In_212);
xor U93 (N_93,In_270,In_154);
and U94 (N_94,In_130,In_353);
or U95 (N_95,In_135,In_477);
nor U96 (N_96,In_336,In_59);
nor U97 (N_97,In_490,In_286);
xnor U98 (N_98,In_436,In_278);
or U99 (N_99,In_386,In_473);
and U100 (N_100,In_246,In_173);
nand U101 (N_101,In_177,In_267);
xor U102 (N_102,In_306,In_251);
nor U103 (N_103,In_430,In_218);
nand U104 (N_104,In_347,In_244);
xnor U105 (N_105,In_102,In_248);
nand U106 (N_106,In_374,In_70);
and U107 (N_107,In_42,In_283);
nand U108 (N_108,In_230,In_174);
xnor U109 (N_109,In_27,In_191);
nand U110 (N_110,In_40,In_345);
nand U111 (N_111,In_442,In_82);
or U112 (N_112,In_148,In_12);
nor U113 (N_113,In_58,In_90);
nor U114 (N_114,In_26,In_236);
xnor U115 (N_115,In_463,In_184);
or U116 (N_116,In_393,In_217);
nor U117 (N_117,In_492,In_399);
xnor U118 (N_118,In_145,In_79);
xnor U119 (N_119,In_214,In_475);
or U120 (N_120,In_453,In_471);
xnor U121 (N_121,In_488,In_301);
and U122 (N_122,In_23,In_361);
nand U123 (N_123,In_187,In_150);
and U124 (N_124,In_418,In_356);
and U125 (N_125,In_404,In_163);
and U126 (N_126,In_67,In_221);
nor U127 (N_127,In_166,In_406);
or U128 (N_128,In_451,In_320);
and U129 (N_129,In_152,In_485);
xor U130 (N_130,In_438,In_444);
xor U131 (N_131,In_324,In_46);
nor U132 (N_132,In_416,In_415);
nand U133 (N_133,In_383,In_56);
or U134 (N_134,In_379,In_354);
and U135 (N_135,In_47,In_405);
nor U136 (N_136,In_376,In_77);
or U137 (N_137,In_117,In_300);
nor U138 (N_138,In_441,In_242);
and U139 (N_139,In_51,In_167);
nor U140 (N_140,In_373,In_448);
or U141 (N_141,In_169,In_486);
nor U142 (N_142,In_434,In_215);
nor U143 (N_143,In_400,In_176);
nand U144 (N_144,In_476,In_443);
and U145 (N_145,In_499,In_131);
and U146 (N_146,In_128,In_412);
nand U147 (N_147,In_258,In_207);
xnor U148 (N_148,In_195,In_17);
or U149 (N_149,In_321,In_494);
and U150 (N_150,In_203,In_105);
nor U151 (N_151,In_414,In_146);
xnor U152 (N_152,In_305,In_474);
nand U153 (N_153,In_314,In_273);
xnor U154 (N_154,In_92,In_24);
and U155 (N_155,In_78,In_249);
nand U156 (N_156,In_144,In_182);
xor U157 (N_157,In_104,In_432);
xor U158 (N_158,In_377,In_452);
and U159 (N_159,In_318,In_151);
or U160 (N_160,In_7,In_459);
or U161 (N_161,In_255,In_309);
or U162 (N_162,In_384,In_260);
or U163 (N_163,In_61,In_435);
and U164 (N_164,In_3,In_125);
xor U165 (N_165,In_355,In_10);
and U166 (N_166,In_200,In_425);
xor U167 (N_167,In_316,In_216);
and U168 (N_168,In_129,In_99);
or U169 (N_169,In_49,In_14);
xor U170 (N_170,In_387,In_103);
xor U171 (N_171,In_143,In_480);
xor U172 (N_172,In_360,In_60);
xnor U173 (N_173,In_41,In_433);
nor U174 (N_174,In_31,In_337);
nor U175 (N_175,In_165,In_331);
and U176 (N_176,In_233,In_133);
nor U177 (N_177,In_34,In_66);
or U178 (N_178,In_38,In_325);
nor U179 (N_179,In_332,In_298);
and U180 (N_180,In_161,In_366);
nand U181 (N_181,In_317,In_446);
and U182 (N_182,In_410,In_80);
nor U183 (N_183,In_335,In_342);
xnor U184 (N_184,In_339,In_341);
or U185 (N_185,In_274,In_275);
nor U186 (N_186,In_28,In_170);
xnor U187 (N_187,In_241,In_279);
nand U188 (N_188,In_391,In_268);
nor U189 (N_189,In_392,In_136);
nand U190 (N_190,In_239,In_315);
xor U191 (N_191,In_4,In_100);
and U192 (N_192,In_43,In_308);
nor U193 (N_193,In_211,In_247);
and U194 (N_194,In_138,In_257);
and U195 (N_195,In_122,In_287);
nand U196 (N_196,In_344,In_147);
or U197 (N_197,In_264,In_375);
xor U198 (N_198,In_284,In_468);
xnor U199 (N_199,In_75,In_234);
nand U200 (N_200,In_439,In_68);
nor U201 (N_201,In_183,In_33);
nor U202 (N_202,In_426,In_357);
and U203 (N_203,In_160,In_440);
nand U204 (N_204,In_171,In_359);
nor U205 (N_205,In_126,In_483);
or U206 (N_206,In_76,In_88);
or U207 (N_207,In_296,In_408);
and U208 (N_208,In_423,In_110);
nor U209 (N_209,In_32,In_292);
and U210 (N_210,In_98,In_256);
and U211 (N_211,In_114,In_319);
nand U212 (N_212,In_1,In_30);
nor U213 (N_213,In_25,In_310);
and U214 (N_214,In_478,In_155);
or U215 (N_215,In_290,In_156);
and U216 (N_216,In_299,In_403);
xor U217 (N_217,In_35,In_422);
and U218 (N_218,In_385,In_323);
or U219 (N_219,In_447,In_45);
xor U220 (N_220,In_334,In_457);
and U221 (N_221,In_487,In_11);
and U222 (N_222,In_37,In_421);
xor U223 (N_223,In_223,In_462);
nor U224 (N_224,In_235,In_16);
or U225 (N_225,In_276,In_162);
nand U226 (N_226,In_2,In_178);
nor U227 (N_227,In_118,In_472);
nand U228 (N_228,In_364,In_243);
nand U229 (N_229,In_69,In_188);
nand U230 (N_230,In_495,In_449);
nand U231 (N_231,In_407,In_362);
or U232 (N_232,In_253,In_50);
and U233 (N_233,In_186,In_390);
or U234 (N_234,In_469,In_388);
or U235 (N_235,In_232,In_269);
nor U236 (N_236,In_137,In_297);
xnor U237 (N_237,In_44,In_91);
and U238 (N_238,In_55,In_431);
and U239 (N_239,In_351,In_229);
and U240 (N_240,In_164,In_272);
nor U241 (N_241,In_65,In_181);
nand U242 (N_242,In_363,In_22);
nor U243 (N_243,In_63,In_94);
nor U244 (N_244,In_350,In_429);
xor U245 (N_245,In_189,In_83);
and U246 (N_246,In_72,In_424);
nand U247 (N_247,In_201,In_62);
nand U248 (N_248,In_134,In_142);
nor U249 (N_249,In_461,In_113);
nor U250 (N_250,In_349,In_375);
xnor U251 (N_251,In_131,In_239);
or U252 (N_252,In_124,In_487);
and U253 (N_253,In_330,In_262);
nand U254 (N_254,In_50,In_46);
xnor U255 (N_255,In_443,In_389);
nor U256 (N_256,In_424,In_147);
and U257 (N_257,In_229,In_438);
and U258 (N_258,In_3,In_370);
or U259 (N_259,In_94,In_123);
or U260 (N_260,In_235,In_198);
xnor U261 (N_261,In_42,In_64);
nand U262 (N_262,In_477,In_199);
and U263 (N_263,In_87,In_219);
and U264 (N_264,In_347,In_341);
nor U265 (N_265,In_464,In_125);
nor U266 (N_266,In_434,In_53);
and U267 (N_267,In_17,In_182);
nand U268 (N_268,In_206,In_183);
and U269 (N_269,In_480,In_261);
xor U270 (N_270,In_237,In_426);
xnor U271 (N_271,In_176,In_335);
xor U272 (N_272,In_314,In_423);
and U273 (N_273,In_139,In_84);
xnor U274 (N_274,In_379,In_135);
and U275 (N_275,In_218,In_131);
nor U276 (N_276,In_375,In_206);
and U277 (N_277,In_271,In_53);
nand U278 (N_278,In_221,In_193);
or U279 (N_279,In_459,In_35);
and U280 (N_280,In_37,In_326);
or U281 (N_281,In_152,In_359);
and U282 (N_282,In_42,In_319);
nand U283 (N_283,In_74,In_38);
or U284 (N_284,In_304,In_52);
or U285 (N_285,In_218,In_21);
xnor U286 (N_286,In_213,In_445);
nand U287 (N_287,In_414,In_496);
nand U288 (N_288,In_173,In_151);
and U289 (N_289,In_466,In_260);
nor U290 (N_290,In_1,In_31);
nor U291 (N_291,In_154,In_293);
or U292 (N_292,In_393,In_282);
xnor U293 (N_293,In_220,In_196);
and U294 (N_294,In_207,In_74);
xnor U295 (N_295,In_327,In_119);
xnor U296 (N_296,In_131,In_382);
nand U297 (N_297,In_455,In_465);
xnor U298 (N_298,In_231,In_403);
or U299 (N_299,In_219,In_105);
nand U300 (N_300,In_364,In_60);
and U301 (N_301,In_230,In_133);
nor U302 (N_302,In_252,In_403);
xnor U303 (N_303,In_367,In_446);
xnor U304 (N_304,In_192,In_75);
and U305 (N_305,In_198,In_112);
and U306 (N_306,In_99,In_182);
nor U307 (N_307,In_456,In_359);
or U308 (N_308,In_273,In_55);
nand U309 (N_309,In_446,In_330);
nor U310 (N_310,In_96,In_148);
nor U311 (N_311,In_421,In_203);
and U312 (N_312,In_443,In_434);
nand U313 (N_313,In_110,In_251);
and U314 (N_314,In_247,In_354);
or U315 (N_315,In_267,In_434);
nor U316 (N_316,In_377,In_145);
nor U317 (N_317,In_68,In_482);
nor U318 (N_318,In_462,In_274);
or U319 (N_319,In_282,In_91);
or U320 (N_320,In_259,In_320);
or U321 (N_321,In_225,In_182);
or U322 (N_322,In_282,In_20);
or U323 (N_323,In_68,In_231);
nand U324 (N_324,In_53,In_221);
and U325 (N_325,In_118,In_109);
and U326 (N_326,In_178,In_24);
nand U327 (N_327,In_389,In_187);
xor U328 (N_328,In_290,In_119);
nor U329 (N_329,In_419,In_94);
nor U330 (N_330,In_400,In_339);
nor U331 (N_331,In_298,In_421);
xor U332 (N_332,In_171,In_370);
and U333 (N_333,In_444,In_185);
nor U334 (N_334,In_1,In_152);
xor U335 (N_335,In_300,In_325);
or U336 (N_336,In_209,In_88);
nor U337 (N_337,In_319,In_191);
xnor U338 (N_338,In_81,In_37);
and U339 (N_339,In_364,In_207);
nor U340 (N_340,In_274,In_76);
or U341 (N_341,In_342,In_16);
and U342 (N_342,In_169,In_429);
and U343 (N_343,In_348,In_289);
nand U344 (N_344,In_42,In_363);
nor U345 (N_345,In_218,In_327);
or U346 (N_346,In_456,In_310);
and U347 (N_347,In_385,In_334);
nand U348 (N_348,In_498,In_195);
nor U349 (N_349,In_222,In_145);
and U350 (N_350,In_247,In_440);
nand U351 (N_351,In_302,In_304);
nor U352 (N_352,In_263,In_162);
or U353 (N_353,In_86,In_285);
nand U354 (N_354,In_139,In_433);
nand U355 (N_355,In_8,In_254);
or U356 (N_356,In_351,In_275);
nand U357 (N_357,In_107,In_328);
nand U358 (N_358,In_374,In_163);
or U359 (N_359,In_18,In_143);
nor U360 (N_360,In_346,In_325);
and U361 (N_361,In_334,In_141);
nor U362 (N_362,In_131,In_384);
nor U363 (N_363,In_149,In_197);
xnor U364 (N_364,In_443,In_433);
or U365 (N_365,In_203,In_349);
or U366 (N_366,In_488,In_250);
xnor U367 (N_367,In_140,In_190);
xnor U368 (N_368,In_263,In_237);
nor U369 (N_369,In_178,In_262);
nand U370 (N_370,In_314,In_107);
nand U371 (N_371,In_11,In_245);
nor U372 (N_372,In_344,In_282);
or U373 (N_373,In_441,In_455);
or U374 (N_374,In_32,In_348);
nor U375 (N_375,In_284,In_155);
or U376 (N_376,In_158,In_358);
and U377 (N_377,In_365,In_499);
nor U378 (N_378,In_243,In_209);
nor U379 (N_379,In_183,In_70);
nand U380 (N_380,In_390,In_189);
nand U381 (N_381,In_58,In_437);
nand U382 (N_382,In_108,In_158);
nor U383 (N_383,In_193,In_300);
nor U384 (N_384,In_4,In_83);
xnor U385 (N_385,In_408,In_33);
nand U386 (N_386,In_310,In_204);
nand U387 (N_387,In_466,In_277);
xnor U388 (N_388,In_97,In_2);
and U389 (N_389,In_442,In_423);
nand U390 (N_390,In_330,In_377);
nand U391 (N_391,In_301,In_257);
nand U392 (N_392,In_337,In_294);
nor U393 (N_393,In_288,In_45);
xnor U394 (N_394,In_335,In_187);
or U395 (N_395,In_494,In_335);
or U396 (N_396,In_365,In_254);
and U397 (N_397,In_420,In_411);
or U398 (N_398,In_221,In_327);
or U399 (N_399,In_245,In_279);
nor U400 (N_400,In_180,In_475);
or U401 (N_401,In_337,In_367);
or U402 (N_402,In_34,In_232);
nand U403 (N_403,In_492,In_345);
and U404 (N_404,In_218,In_388);
xnor U405 (N_405,In_17,In_215);
or U406 (N_406,In_178,In_112);
nand U407 (N_407,In_153,In_488);
and U408 (N_408,In_150,In_209);
xnor U409 (N_409,In_6,In_219);
nor U410 (N_410,In_6,In_208);
nand U411 (N_411,In_132,In_162);
or U412 (N_412,In_167,In_173);
xnor U413 (N_413,In_112,In_413);
nor U414 (N_414,In_306,In_87);
and U415 (N_415,In_349,In_450);
xnor U416 (N_416,In_492,In_180);
nor U417 (N_417,In_483,In_275);
xor U418 (N_418,In_126,In_16);
nand U419 (N_419,In_493,In_429);
or U420 (N_420,In_374,In_5);
and U421 (N_421,In_381,In_482);
nand U422 (N_422,In_352,In_308);
nand U423 (N_423,In_10,In_55);
and U424 (N_424,In_459,In_27);
and U425 (N_425,In_48,In_228);
or U426 (N_426,In_335,In_228);
or U427 (N_427,In_5,In_399);
or U428 (N_428,In_112,In_449);
nor U429 (N_429,In_23,In_144);
or U430 (N_430,In_352,In_79);
and U431 (N_431,In_193,In_470);
nand U432 (N_432,In_361,In_258);
nor U433 (N_433,In_475,In_102);
and U434 (N_434,In_319,In_442);
and U435 (N_435,In_141,In_175);
and U436 (N_436,In_160,In_81);
nor U437 (N_437,In_152,In_233);
or U438 (N_438,In_14,In_47);
nor U439 (N_439,In_158,In_329);
nand U440 (N_440,In_309,In_67);
nand U441 (N_441,In_177,In_492);
xnor U442 (N_442,In_339,In_194);
and U443 (N_443,In_322,In_413);
xor U444 (N_444,In_231,In_340);
or U445 (N_445,In_236,In_432);
nand U446 (N_446,In_422,In_240);
xor U447 (N_447,In_350,In_294);
nand U448 (N_448,In_363,In_404);
and U449 (N_449,In_154,In_445);
or U450 (N_450,In_45,In_244);
xnor U451 (N_451,In_333,In_90);
and U452 (N_452,In_195,In_477);
or U453 (N_453,In_216,In_469);
nand U454 (N_454,In_245,In_299);
or U455 (N_455,In_41,In_306);
nor U456 (N_456,In_141,In_178);
or U457 (N_457,In_472,In_334);
or U458 (N_458,In_326,In_67);
and U459 (N_459,In_364,In_424);
nor U460 (N_460,In_121,In_450);
nor U461 (N_461,In_175,In_233);
and U462 (N_462,In_127,In_484);
xor U463 (N_463,In_291,In_428);
nand U464 (N_464,In_117,In_69);
and U465 (N_465,In_253,In_336);
nand U466 (N_466,In_421,In_307);
xor U467 (N_467,In_372,In_462);
nand U468 (N_468,In_313,In_285);
xor U469 (N_469,In_72,In_450);
nand U470 (N_470,In_214,In_394);
nand U471 (N_471,In_11,In_285);
or U472 (N_472,In_369,In_287);
nor U473 (N_473,In_223,In_403);
xor U474 (N_474,In_455,In_14);
nor U475 (N_475,In_287,In_456);
nand U476 (N_476,In_276,In_90);
nor U477 (N_477,In_4,In_251);
and U478 (N_478,In_267,In_85);
nand U479 (N_479,In_67,In_268);
nand U480 (N_480,In_42,In_137);
xnor U481 (N_481,In_362,In_237);
or U482 (N_482,In_13,In_277);
or U483 (N_483,In_321,In_81);
nor U484 (N_484,In_179,In_218);
nand U485 (N_485,In_301,In_347);
nor U486 (N_486,In_24,In_71);
or U487 (N_487,In_56,In_211);
xor U488 (N_488,In_341,In_342);
and U489 (N_489,In_230,In_4);
nand U490 (N_490,In_286,In_46);
and U491 (N_491,In_172,In_364);
nor U492 (N_492,In_46,In_465);
nor U493 (N_493,In_94,In_264);
nor U494 (N_494,In_33,In_231);
nand U495 (N_495,In_197,In_120);
and U496 (N_496,In_94,In_451);
nand U497 (N_497,In_107,In_339);
nor U498 (N_498,In_258,In_188);
nor U499 (N_499,In_105,In_50);
xnor U500 (N_500,N_78,N_192);
or U501 (N_501,N_462,N_283);
nor U502 (N_502,N_405,N_252);
or U503 (N_503,N_122,N_362);
nand U504 (N_504,N_479,N_125);
and U505 (N_505,N_367,N_288);
and U506 (N_506,N_411,N_349);
and U507 (N_507,N_476,N_147);
nor U508 (N_508,N_57,N_270);
or U509 (N_509,N_35,N_265);
and U510 (N_510,N_272,N_148);
nor U511 (N_511,N_285,N_41);
nand U512 (N_512,N_281,N_130);
nand U513 (N_513,N_317,N_186);
nor U514 (N_514,N_467,N_99);
nor U515 (N_515,N_79,N_451);
or U516 (N_516,N_71,N_216);
or U517 (N_517,N_188,N_158);
xor U518 (N_518,N_46,N_131);
or U519 (N_519,N_497,N_402);
xnor U520 (N_520,N_396,N_103);
xnor U521 (N_521,N_316,N_269);
nand U522 (N_522,N_32,N_218);
nor U523 (N_523,N_350,N_143);
xnor U524 (N_524,N_76,N_355);
nor U525 (N_525,N_408,N_110);
or U526 (N_526,N_498,N_257);
and U527 (N_527,N_149,N_441);
and U528 (N_528,N_50,N_23);
and U529 (N_529,N_132,N_453);
and U530 (N_530,N_455,N_219);
nor U531 (N_531,N_39,N_189);
nor U532 (N_532,N_201,N_211);
nor U533 (N_533,N_3,N_304);
nor U534 (N_534,N_138,N_404);
xor U535 (N_535,N_255,N_488);
nand U536 (N_536,N_440,N_484);
nand U537 (N_537,N_429,N_207);
or U538 (N_538,N_121,N_302);
nor U539 (N_539,N_458,N_221);
nor U540 (N_540,N_259,N_452);
or U541 (N_541,N_204,N_301);
and U542 (N_542,N_150,N_61);
or U543 (N_543,N_213,N_51);
xor U544 (N_544,N_210,N_347);
xnor U545 (N_545,N_318,N_313);
and U546 (N_546,N_67,N_494);
nand U547 (N_547,N_415,N_80);
nor U548 (N_548,N_181,N_49);
or U549 (N_549,N_63,N_351);
xnor U550 (N_550,N_320,N_397);
and U551 (N_551,N_209,N_28);
xnor U552 (N_552,N_424,N_433);
or U553 (N_553,N_275,N_258);
nor U554 (N_554,N_124,N_492);
or U555 (N_555,N_354,N_229);
or U556 (N_556,N_442,N_469);
or U557 (N_557,N_450,N_296);
and U558 (N_558,N_152,N_12);
and U559 (N_559,N_200,N_416);
and U560 (N_560,N_115,N_162);
xnor U561 (N_561,N_375,N_254);
xor U562 (N_562,N_206,N_203);
or U563 (N_563,N_273,N_14);
xor U564 (N_564,N_250,N_438);
nand U565 (N_565,N_92,N_168);
and U566 (N_566,N_136,N_86);
nand U567 (N_567,N_456,N_482);
xnor U568 (N_568,N_289,N_15);
or U569 (N_569,N_297,N_65);
and U570 (N_570,N_231,N_113);
or U571 (N_571,N_217,N_21);
nor U572 (N_572,N_238,N_214);
xor U573 (N_573,N_154,N_374);
and U574 (N_574,N_34,N_98);
nand U575 (N_575,N_454,N_324);
or U576 (N_576,N_127,N_197);
or U577 (N_577,N_268,N_277);
nand U578 (N_578,N_242,N_391);
and U579 (N_579,N_325,N_341);
nor U580 (N_580,N_220,N_377);
or U581 (N_581,N_36,N_73);
or U582 (N_582,N_180,N_245);
xor U583 (N_583,N_4,N_319);
and U584 (N_584,N_223,N_437);
xnor U585 (N_585,N_48,N_295);
xnor U586 (N_586,N_348,N_118);
and U587 (N_587,N_309,N_382);
xnor U588 (N_588,N_222,N_202);
and U589 (N_589,N_195,N_190);
nor U590 (N_590,N_13,N_261);
nor U591 (N_591,N_499,N_226);
and U592 (N_592,N_159,N_100);
nor U593 (N_593,N_398,N_308);
and U594 (N_594,N_81,N_55);
nand U595 (N_595,N_17,N_228);
or U596 (N_596,N_191,N_133);
xor U597 (N_597,N_77,N_385);
nor U598 (N_598,N_365,N_326);
or U599 (N_599,N_88,N_106);
nor U600 (N_600,N_42,N_380);
xor U601 (N_601,N_475,N_300);
and U602 (N_602,N_193,N_291);
xnor U603 (N_603,N_178,N_495);
nand U604 (N_604,N_493,N_298);
and U605 (N_605,N_431,N_353);
nor U606 (N_606,N_37,N_135);
xor U607 (N_607,N_109,N_134);
and U608 (N_608,N_9,N_290);
xnor U609 (N_609,N_435,N_463);
nand U610 (N_610,N_471,N_339);
nor U611 (N_611,N_129,N_423);
and U612 (N_612,N_434,N_262);
nand U613 (N_613,N_327,N_102);
nand U614 (N_614,N_457,N_436);
nand U615 (N_615,N_389,N_107);
nor U616 (N_616,N_409,N_306);
nand U617 (N_617,N_62,N_95);
and U618 (N_618,N_116,N_139);
xnor U619 (N_619,N_315,N_432);
xor U620 (N_620,N_399,N_141);
xor U621 (N_621,N_430,N_108);
nand U622 (N_622,N_368,N_418);
nor U623 (N_623,N_140,N_464);
nor U624 (N_624,N_312,N_422);
nand U625 (N_625,N_68,N_322);
or U626 (N_626,N_310,N_445);
nand U627 (N_627,N_428,N_271);
nand U628 (N_628,N_421,N_280);
xnor U629 (N_629,N_94,N_256);
or U630 (N_630,N_241,N_90);
and U631 (N_631,N_331,N_263);
xor U632 (N_632,N_439,N_164);
and U633 (N_633,N_343,N_372);
and U634 (N_634,N_406,N_387);
and U635 (N_635,N_232,N_246);
and U636 (N_636,N_194,N_87);
nand U637 (N_637,N_307,N_444);
nand U638 (N_638,N_356,N_184);
xor U639 (N_639,N_419,N_364);
nand U640 (N_640,N_26,N_1);
nand U641 (N_641,N_234,N_395);
nand U642 (N_642,N_279,N_111);
xnor U643 (N_643,N_361,N_366);
and U644 (N_644,N_260,N_371);
or U645 (N_645,N_91,N_239);
or U646 (N_646,N_276,N_359);
and U647 (N_647,N_10,N_69);
or U648 (N_648,N_25,N_403);
and U649 (N_649,N_244,N_491);
xor U650 (N_650,N_470,N_6);
nand U651 (N_651,N_170,N_425);
and U652 (N_652,N_27,N_82);
nor U653 (N_653,N_384,N_227);
nand U654 (N_654,N_248,N_43);
xnor U655 (N_655,N_144,N_346);
nand U656 (N_656,N_237,N_52);
and U657 (N_657,N_337,N_179);
nor U658 (N_658,N_60,N_357);
or U659 (N_659,N_173,N_328);
xor U660 (N_660,N_461,N_412);
nor U661 (N_661,N_414,N_177);
or U662 (N_662,N_460,N_16);
xnor U663 (N_663,N_160,N_224);
or U664 (N_664,N_225,N_335);
nor U665 (N_665,N_240,N_292);
or U666 (N_666,N_74,N_420);
and U667 (N_667,N_215,N_24);
nand U668 (N_668,N_369,N_30);
and U669 (N_669,N_314,N_58);
nand U670 (N_670,N_167,N_282);
xnor U671 (N_671,N_104,N_373);
and U672 (N_672,N_392,N_174);
nand U673 (N_673,N_198,N_294);
nor U674 (N_674,N_137,N_11);
or U675 (N_675,N_468,N_443);
or U676 (N_676,N_31,N_7);
nand U677 (N_677,N_235,N_447);
nor U678 (N_678,N_299,N_72);
and U679 (N_679,N_119,N_333);
xnor U680 (N_680,N_112,N_474);
and U681 (N_681,N_40,N_172);
nor U682 (N_682,N_249,N_97);
nand U683 (N_683,N_96,N_410);
nor U684 (N_684,N_407,N_155);
xnor U685 (N_685,N_33,N_305);
or U686 (N_686,N_334,N_381);
nor U687 (N_687,N_253,N_267);
and U688 (N_688,N_5,N_287);
and U689 (N_689,N_176,N_182);
xnor U690 (N_690,N_340,N_93);
nand U691 (N_691,N_236,N_101);
nand U692 (N_692,N_323,N_199);
xnor U693 (N_693,N_394,N_483);
xor U694 (N_694,N_449,N_114);
and U695 (N_695,N_22,N_45);
nor U696 (N_696,N_59,N_196);
nand U697 (N_697,N_338,N_89);
and U698 (N_698,N_336,N_54);
xor U699 (N_699,N_400,N_293);
xnor U700 (N_700,N_332,N_487);
nand U701 (N_701,N_417,N_477);
or U702 (N_702,N_448,N_163);
or U703 (N_703,N_126,N_426);
nand U704 (N_704,N_360,N_187);
or U705 (N_705,N_459,N_146);
and U706 (N_706,N_481,N_496);
xor U707 (N_707,N_183,N_251);
xor U708 (N_708,N_44,N_66);
xnor U709 (N_709,N_378,N_166);
nand U710 (N_710,N_84,N_70);
nor U711 (N_711,N_205,N_370);
nand U712 (N_712,N_413,N_478);
or U713 (N_713,N_278,N_329);
and U714 (N_714,N_379,N_185);
or U715 (N_715,N_303,N_473);
and U716 (N_716,N_401,N_208);
nand U717 (N_717,N_156,N_490);
nor U718 (N_718,N_151,N_117);
nand U719 (N_719,N_274,N_393);
nand U720 (N_720,N_284,N_390);
nor U721 (N_721,N_157,N_175);
nor U722 (N_722,N_345,N_20);
or U723 (N_723,N_0,N_2);
or U724 (N_724,N_153,N_427);
and U725 (N_725,N_29,N_358);
nor U726 (N_726,N_165,N_480);
or U727 (N_727,N_388,N_230);
nand U728 (N_728,N_145,N_489);
nand U729 (N_729,N_266,N_344);
or U730 (N_730,N_465,N_18);
nand U731 (N_731,N_171,N_120);
nor U732 (N_732,N_47,N_19);
xor U733 (N_733,N_56,N_311);
nand U734 (N_734,N_330,N_38);
nand U735 (N_735,N_83,N_85);
nand U736 (N_736,N_75,N_8);
or U737 (N_737,N_142,N_105);
nand U738 (N_738,N_233,N_466);
nor U739 (N_739,N_128,N_383);
xnor U740 (N_740,N_486,N_386);
nand U741 (N_741,N_123,N_485);
and U742 (N_742,N_243,N_212);
nand U743 (N_743,N_53,N_472);
nand U744 (N_744,N_446,N_342);
or U745 (N_745,N_247,N_169);
nor U746 (N_746,N_161,N_352);
and U747 (N_747,N_321,N_286);
xor U748 (N_748,N_376,N_64);
or U749 (N_749,N_363,N_264);
xor U750 (N_750,N_428,N_267);
nand U751 (N_751,N_441,N_161);
xor U752 (N_752,N_213,N_25);
nand U753 (N_753,N_487,N_440);
or U754 (N_754,N_128,N_52);
nand U755 (N_755,N_425,N_248);
or U756 (N_756,N_228,N_194);
xnor U757 (N_757,N_124,N_367);
and U758 (N_758,N_476,N_105);
nand U759 (N_759,N_346,N_338);
and U760 (N_760,N_79,N_199);
and U761 (N_761,N_68,N_431);
xor U762 (N_762,N_313,N_373);
or U763 (N_763,N_153,N_387);
nand U764 (N_764,N_63,N_348);
nor U765 (N_765,N_123,N_342);
and U766 (N_766,N_224,N_373);
xnor U767 (N_767,N_81,N_158);
xnor U768 (N_768,N_52,N_74);
or U769 (N_769,N_211,N_380);
nor U770 (N_770,N_430,N_389);
xnor U771 (N_771,N_266,N_117);
nor U772 (N_772,N_398,N_366);
xor U773 (N_773,N_319,N_375);
nor U774 (N_774,N_367,N_241);
and U775 (N_775,N_452,N_11);
nor U776 (N_776,N_159,N_58);
nand U777 (N_777,N_355,N_437);
nor U778 (N_778,N_200,N_259);
and U779 (N_779,N_86,N_477);
and U780 (N_780,N_183,N_388);
and U781 (N_781,N_111,N_109);
xor U782 (N_782,N_33,N_205);
xor U783 (N_783,N_220,N_105);
nand U784 (N_784,N_483,N_7);
nor U785 (N_785,N_194,N_405);
nand U786 (N_786,N_263,N_367);
or U787 (N_787,N_389,N_304);
nand U788 (N_788,N_408,N_106);
or U789 (N_789,N_252,N_442);
and U790 (N_790,N_266,N_186);
nor U791 (N_791,N_297,N_15);
and U792 (N_792,N_40,N_65);
nand U793 (N_793,N_416,N_208);
nor U794 (N_794,N_6,N_195);
or U795 (N_795,N_402,N_461);
nand U796 (N_796,N_112,N_321);
xor U797 (N_797,N_28,N_207);
nor U798 (N_798,N_59,N_397);
nand U799 (N_799,N_362,N_386);
and U800 (N_800,N_462,N_292);
nor U801 (N_801,N_14,N_113);
nor U802 (N_802,N_202,N_396);
or U803 (N_803,N_273,N_113);
or U804 (N_804,N_448,N_69);
nand U805 (N_805,N_348,N_9);
xnor U806 (N_806,N_246,N_217);
and U807 (N_807,N_350,N_497);
xnor U808 (N_808,N_233,N_384);
or U809 (N_809,N_28,N_56);
and U810 (N_810,N_110,N_316);
and U811 (N_811,N_300,N_13);
nor U812 (N_812,N_384,N_480);
nand U813 (N_813,N_71,N_314);
nand U814 (N_814,N_327,N_155);
xor U815 (N_815,N_226,N_108);
nor U816 (N_816,N_206,N_304);
nor U817 (N_817,N_484,N_8);
nor U818 (N_818,N_445,N_23);
or U819 (N_819,N_282,N_482);
or U820 (N_820,N_243,N_471);
xnor U821 (N_821,N_451,N_363);
nand U822 (N_822,N_398,N_38);
or U823 (N_823,N_133,N_489);
nor U824 (N_824,N_197,N_292);
xnor U825 (N_825,N_412,N_199);
or U826 (N_826,N_130,N_49);
nand U827 (N_827,N_390,N_167);
and U828 (N_828,N_309,N_291);
nand U829 (N_829,N_285,N_431);
xor U830 (N_830,N_494,N_355);
nand U831 (N_831,N_149,N_351);
nor U832 (N_832,N_349,N_290);
nand U833 (N_833,N_421,N_228);
and U834 (N_834,N_461,N_454);
xor U835 (N_835,N_382,N_85);
nor U836 (N_836,N_374,N_180);
and U837 (N_837,N_366,N_41);
or U838 (N_838,N_254,N_100);
nand U839 (N_839,N_293,N_183);
nor U840 (N_840,N_487,N_236);
or U841 (N_841,N_170,N_347);
and U842 (N_842,N_22,N_453);
xor U843 (N_843,N_468,N_205);
or U844 (N_844,N_345,N_234);
and U845 (N_845,N_333,N_413);
xor U846 (N_846,N_441,N_484);
and U847 (N_847,N_453,N_377);
nand U848 (N_848,N_180,N_28);
xor U849 (N_849,N_204,N_229);
nor U850 (N_850,N_56,N_109);
and U851 (N_851,N_164,N_483);
or U852 (N_852,N_470,N_257);
or U853 (N_853,N_315,N_108);
or U854 (N_854,N_13,N_456);
nor U855 (N_855,N_470,N_290);
and U856 (N_856,N_11,N_107);
nor U857 (N_857,N_203,N_320);
or U858 (N_858,N_414,N_62);
or U859 (N_859,N_157,N_259);
xnor U860 (N_860,N_274,N_81);
or U861 (N_861,N_372,N_151);
or U862 (N_862,N_115,N_460);
xor U863 (N_863,N_322,N_487);
nand U864 (N_864,N_233,N_183);
or U865 (N_865,N_322,N_491);
xor U866 (N_866,N_133,N_104);
nand U867 (N_867,N_349,N_87);
and U868 (N_868,N_460,N_183);
or U869 (N_869,N_86,N_377);
nor U870 (N_870,N_138,N_422);
nand U871 (N_871,N_258,N_70);
nor U872 (N_872,N_101,N_71);
or U873 (N_873,N_158,N_127);
nand U874 (N_874,N_164,N_63);
and U875 (N_875,N_163,N_50);
xnor U876 (N_876,N_187,N_40);
and U877 (N_877,N_190,N_483);
xnor U878 (N_878,N_197,N_146);
nor U879 (N_879,N_485,N_495);
or U880 (N_880,N_101,N_338);
xnor U881 (N_881,N_377,N_214);
nor U882 (N_882,N_117,N_165);
and U883 (N_883,N_294,N_469);
and U884 (N_884,N_353,N_343);
and U885 (N_885,N_11,N_196);
or U886 (N_886,N_412,N_364);
nor U887 (N_887,N_450,N_12);
or U888 (N_888,N_86,N_112);
and U889 (N_889,N_464,N_119);
nand U890 (N_890,N_492,N_440);
and U891 (N_891,N_438,N_22);
xor U892 (N_892,N_74,N_306);
nor U893 (N_893,N_335,N_446);
or U894 (N_894,N_176,N_151);
and U895 (N_895,N_110,N_294);
nor U896 (N_896,N_48,N_156);
and U897 (N_897,N_63,N_10);
and U898 (N_898,N_253,N_459);
nand U899 (N_899,N_204,N_78);
nor U900 (N_900,N_394,N_399);
nand U901 (N_901,N_447,N_180);
xnor U902 (N_902,N_433,N_244);
and U903 (N_903,N_57,N_190);
or U904 (N_904,N_204,N_86);
nand U905 (N_905,N_130,N_16);
nand U906 (N_906,N_160,N_427);
or U907 (N_907,N_229,N_26);
or U908 (N_908,N_5,N_421);
nand U909 (N_909,N_223,N_85);
xnor U910 (N_910,N_54,N_220);
nand U911 (N_911,N_219,N_204);
xnor U912 (N_912,N_20,N_305);
nor U913 (N_913,N_13,N_222);
and U914 (N_914,N_90,N_58);
and U915 (N_915,N_106,N_38);
and U916 (N_916,N_284,N_93);
nor U917 (N_917,N_314,N_37);
or U918 (N_918,N_189,N_173);
and U919 (N_919,N_37,N_491);
and U920 (N_920,N_322,N_452);
and U921 (N_921,N_116,N_416);
and U922 (N_922,N_231,N_329);
xor U923 (N_923,N_231,N_286);
nor U924 (N_924,N_329,N_146);
xnor U925 (N_925,N_281,N_336);
nand U926 (N_926,N_67,N_43);
xor U927 (N_927,N_292,N_128);
nor U928 (N_928,N_283,N_146);
and U929 (N_929,N_8,N_480);
nor U930 (N_930,N_498,N_348);
nand U931 (N_931,N_424,N_119);
nor U932 (N_932,N_130,N_238);
nand U933 (N_933,N_292,N_50);
or U934 (N_934,N_318,N_262);
xor U935 (N_935,N_448,N_153);
or U936 (N_936,N_403,N_122);
or U937 (N_937,N_210,N_109);
or U938 (N_938,N_426,N_165);
nor U939 (N_939,N_272,N_216);
nor U940 (N_940,N_375,N_0);
nor U941 (N_941,N_338,N_441);
nand U942 (N_942,N_307,N_408);
nor U943 (N_943,N_276,N_364);
nor U944 (N_944,N_153,N_173);
or U945 (N_945,N_358,N_166);
nand U946 (N_946,N_165,N_392);
nand U947 (N_947,N_51,N_65);
xor U948 (N_948,N_243,N_445);
xor U949 (N_949,N_255,N_471);
xnor U950 (N_950,N_23,N_143);
nor U951 (N_951,N_404,N_234);
or U952 (N_952,N_67,N_266);
nand U953 (N_953,N_114,N_244);
and U954 (N_954,N_375,N_233);
nand U955 (N_955,N_1,N_372);
and U956 (N_956,N_362,N_107);
nand U957 (N_957,N_230,N_442);
and U958 (N_958,N_496,N_411);
nor U959 (N_959,N_384,N_264);
nor U960 (N_960,N_227,N_80);
nor U961 (N_961,N_70,N_85);
nand U962 (N_962,N_462,N_469);
nand U963 (N_963,N_477,N_480);
nand U964 (N_964,N_163,N_173);
nor U965 (N_965,N_418,N_356);
xnor U966 (N_966,N_314,N_347);
xor U967 (N_967,N_317,N_87);
or U968 (N_968,N_437,N_360);
nor U969 (N_969,N_318,N_44);
and U970 (N_970,N_195,N_199);
or U971 (N_971,N_420,N_215);
nand U972 (N_972,N_207,N_79);
nand U973 (N_973,N_431,N_236);
nand U974 (N_974,N_237,N_300);
or U975 (N_975,N_133,N_178);
nor U976 (N_976,N_201,N_90);
nand U977 (N_977,N_54,N_158);
xor U978 (N_978,N_126,N_487);
nand U979 (N_979,N_175,N_381);
nor U980 (N_980,N_391,N_146);
nand U981 (N_981,N_67,N_430);
xnor U982 (N_982,N_410,N_290);
and U983 (N_983,N_236,N_493);
xor U984 (N_984,N_17,N_407);
and U985 (N_985,N_355,N_127);
nor U986 (N_986,N_374,N_118);
or U987 (N_987,N_146,N_90);
or U988 (N_988,N_182,N_309);
nor U989 (N_989,N_112,N_91);
xor U990 (N_990,N_325,N_428);
xnor U991 (N_991,N_291,N_86);
and U992 (N_992,N_193,N_362);
nand U993 (N_993,N_57,N_61);
nand U994 (N_994,N_423,N_426);
nand U995 (N_995,N_226,N_58);
nand U996 (N_996,N_216,N_226);
nor U997 (N_997,N_379,N_4);
xnor U998 (N_998,N_351,N_64);
and U999 (N_999,N_486,N_53);
xnor U1000 (N_1000,N_552,N_989);
nor U1001 (N_1001,N_822,N_941);
nor U1002 (N_1002,N_951,N_804);
and U1003 (N_1003,N_782,N_665);
xor U1004 (N_1004,N_667,N_717);
nor U1005 (N_1005,N_960,N_506);
nor U1006 (N_1006,N_980,N_728);
and U1007 (N_1007,N_678,N_981);
or U1008 (N_1008,N_501,N_952);
or U1009 (N_1009,N_684,N_550);
and U1010 (N_1010,N_685,N_636);
xor U1011 (N_1011,N_521,N_771);
and U1012 (N_1012,N_809,N_695);
nor U1013 (N_1013,N_624,N_876);
nor U1014 (N_1014,N_762,N_650);
or U1015 (N_1015,N_997,N_851);
xnor U1016 (N_1016,N_713,N_765);
nor U1017 (N_1017,N_926,N_587);
or U1018 (N_1018,N_969,N_743);
nand U1019 (N_1019,N_567,N_617);
and U1020 (N_1020,N_548,N_640);
xnor U1021 (N_1021,N_930,N_718);
and U1022 (N_1022,N_884,N_693);
nor U1023 (N_1023,N_527,N_612);
and U1024 (N_1024,N_858,N_599);
xor U1025 (N_1025,N_634,N_996);
or U1026 (N_1026,N_918,N_803);
nand U1027 (N_1027,N_616,N_572);
and U1028 (N_1028,N_838,N_615);
nand U1029 (N_1029,N_559,N_625);
nand U1030 (N_1030,N_998,N_748);
nand U1031 (N_1031,N_915,N_878);
nand U1032 (N_1032,N_919,N_710);
nand U1033 (N_1033,N_985,N_833);
and U1034 (N_1034,N_794,N_917);
and U1035 (N_1035,N_757,N_979);
xnor U1036 (N_1036,N_842,N_764);
nor U1037 (N_1037,N_775,N_909);
nand U1038 (N_1038,N_977,N_744);
nor U1039 (N_1039,N_712,N_912);
nand U1040 (N_1040,N_541,N_651);
nand U1041 (N_1041,N_646,N_538);
or U1042 (N_1042,N_921,N_654);
and U1043 (N_1043,N_702,N_807);
nand U1044 (N_1044,N_533,N_633);
nand U1045 (N_1045,N_701,N_729);
xor U1046 (N_1046,N_781,N_545);
nand U1047 (N_1047,N_620,N_813);
or U1048 (N_1048,N_895,N_938);
and U1049 (N_1049,N_819,N_609);
or U1050 (N_1050,N_711,N_671);
or U1051 (N_1051,N_860,N_818);
nand U1052 (N_1052,N_940,N_539);
nor U1053 (N_1053,N_956,N_867);
and U1054 (N_1054,N_534,N_834);
xor U1055 (N_1055,N_735,N_734);
xnor U1056 (N_1056,N_546,N_768);
or U1057 (N_1057,N_741,N_516);
and U1058 (N_1058,N_773,N_797);
and U1059 (N_1059,N_655,N_935);
or U1060 (N_1060,N_508,N_856);
xnor U1061 (N_1061,N_510,N_690);
nand U1062 (N_1062,N_847,N_815);
or U1063 (N_1063,N_716,N_628);
or U1064 (N_1064,N_512,N_673);
xor U1065 (N_1065,N_845,N_772);
nand U1066 (N_1066,N_631,N_879);
or U1067 (N_1067,N_857,N_836);
or U1068 (N_1068,N_754,N_630);
and U1069 (N_1069,N_814,N_928);
xnor U1070 (N_1070,N_611,N_528);
nand U1071 (N_1071,N_732,N_529);
and U1072 (N_1072,N_519,N_944);
nor U1073 (N_1073,N_937,N_544);
or U1074 (N_1074,N_780,N_635);
nor U1075 (N_1075,N_747,N_707);
nor U1076 (N_1076,N_874,N_827);
xnor U1077 (N_1077,N_578,N_598);
nand U1078 (N_1078,N_719,N_756);
or U1079 (N_1079,N_812,N_666);
xor U1080 (N_1080,N_664,N_639);
xor U1081 (N_1081,N_504,N_513);
nor U1082 (N_1082,N_901,N_869);
xor U1083 (N_1083,N_904,N_890);
nor U1084 (N_1084,N_709,N_626);
and U1085 (N_1085,N_829,N_948);
nor U1086 (N_1086,N_505,N_680);
and U1087 (N_1087,N_811,N_575);
xor U1088 (N_1088,N_686,N_608);
and U1089 (N_1089,N_900,N_726);
nand U1090 (N_1090,N_720,N_698);
and U1091 (N_1091,N_677,N_826);
nor U1092 (N_1092,N_532,N_742);
or U1093 (N_1093,N_848,N_689);
nand U1094 (N_1094,N_779,N_555);
nor U1095 (N_1095,N_540,N_849);
or U1096 (N_1096,N_841,N_911);
nand U1097 (N_1097,N_975,N_658);
or U1098 (N_1098,N_502,N_576);
nand U1099 (N_1099,N_872,N_793);
nand U1100 (N_1100,N_563,N_562);
nor U1101 (N_1101,N_753,N_854);
xnor U1102 (N_1102,N_913,N_557);
or U1103 (N_1103,N_882,N_873);
xor U1104 (N_1104,N_916,N_517);
xnor U1105 (N_1105,N_843,N_991);
nor U1106 (N_1106,N_607,N_929);
xor U1107 (N_1107,N_755,N_888);
or U1108 (N_1108,N_520,N_579);
or U1109 (N_1109,N_887,N_638);
or U1110 (N_1110,N_524,N_697);
and U1111 (N_1111,N_933,N_610);
nor U1112 (N_1112,N_687,N_652);
xor U1113 (N_1113,N_808,N_586);
nand U1114 (N_1114,N_902,N_580);
xnor U1115 (N_1115,N_589,N_958);
and U1116 (N_1116,N_964,N_721);
or U1117 (N_1117,N_623,N_880);
and U1118 (N_1118,N_522,N_606);
nand U1119 (N_1119,N_730,N_681);
nand U1120 (N_1120,N_973,N_643);
nor U1121 (N_1121,N_866,N_708);
and U1122 (N_1122,N_507,N_704);
and U1123 (N_1123,N_832,N_789);
nor U1124 (N_1124,N_592,N_798);
nand U1125 (N_1125,N_657,N_692);
or U1126 (N_1126,N_825,N_927);
and U1127 (N_1127,N_959,N_770);
or U1128 (N_1128,N_817,N_569);
nor U1129 (N_1129,N_968,N_503);
and U1130 (N_1130,N_805,N_865);
nand U1131 (N_1131,N_543,N_792);
nor U1132 (N_1132,N_554,N_723);
and U1133 (N_1133,N_733,N_816);
nand U1134 (N_1134,N_637,N_514);
xor U1135 (N_1135,N_844,N_703);
nor U1136 (N_1136,N_893,N_602);
or U1137 (N_1137,N_897,N_571);
nor U1138 (N_1138,N_566,N_992);
nand U1139 (N_1139,N_542,N_936);
or U1140 (N_1140,N_668,N_549);
nand U1141 (N_1141,N_953,N_896);
and U1142 (N_1142,N_604,N_961);
or U1143 (N_1143,N_763,N_932);
nand U1144 (N_1144,N_594,N_661);
xor U1145 (N_1145,N_669,N_537);
nand U1146 (N_1146,N_972,N_988);
or U1147 (N_1147,N_785,N_995);
nor U1148 (N_1148,N_839,N_820);
or U1149 (N_1149,N_778,N_791);
and U1150 (N_1150,N_931,N_801);
nand U1151 (N_1151,N_894,N_568);
nand U1152 (N_1152,N_601,N_802);
nand U1153 (N_1153,N_600,N_760);
or U1154 (N_1154,N_864,N_889);
nor U1155 (N_1155,N_954,N_853);
xor U1156 (N_1156,N_910,N_526);
nand U1157 (N_1157,N_993,N_824);
and U1158 (N_1158,N_863,N_535);
or U1159 (N_1159,N_786,N_581);
and U1160 (N_1160,N_725,N_565);
or U1161 (N_1161,N_536,N_957);
or U1162 (N_1162,N_783,N_746);
and U1163 (N_1163,N_588,N_663);
nand U1164 (N_1164,N_577,N_583);
and U1165 (N_1165,N_831,N_971);
nand U1166 (N_1166,N_727,N_976);
xor U1167 (N_1167,N_675,N_947);
or U1168 (N_1168,N_547,N_596);
xor U1169 (N_1169,N_672,N_525);
nor U1170 (N_1170,N_945,N_974);
nand U1171 (N_1171,N_642,N_593);
nor U1172 (N_1172,N_553,N_777);
or U1173 (N_1173,N_881,N_759);
or U1174 (N_1174,N_556,N_800);
nand U1175 (N_1175,N_850,N_705);
xnor U1176 (N_1176,N_696,N_823);
nor U1177 (N_1177,N_871,N_920);
or U1178 (N_1178,N_564,N_821);
or U1179 (N_1179,N_560,N_752);
nand U1180 (N_1180,N_605,N_699);
and U1181 (N_1181,N_715,N_530);
and U1182 (N_1182,N_670,N_694);
xor U1183 (N_1183,N_906,N_899);
and U1184 (N_1184,N_774,N_674);
xnor U1185 (N_1185,N_982,N_810);
and U1186 (N_1186,N_885,N_922);
and U1187 (N_1187,N_840,N_776);
xor U1188 (N_1188,N_787,N_619);
xor U1189 (N_1189,N_799,N_603);
nor U1190 (N_1190,N_835,N_622);
nand U1191 (N_1191,N_632,N_644);
nand U1192 (N_1192,N_962,N_722);
or U1193 (N_1193,N_738,N_648);
nor U1194 (N_1194,N_629,N_987);
nor U1195 (N_1195,N_994,N_846);
or U1196 (N_1196,N_551,N_597);
and U1197 (N_1197,N_641,N_855);
or U1198 (N_1198,N_868,N_828);
xnor U1199 (N_1199,N_795,N_923);
xor U1200 (N_1200,N_518,N_946);
nand U1201 (N_1201,N_939,N_903);
nor U1202 (N_1202,N_892,N_558);
xor U1203 (N_1203,N_925,N_761);
or U1204 (N_1204,N_758,N_570);
and U1205 (N_1205,N_749,N_796);
xor U1206 (N_1206,N_990,N_618);
and U1207 (N_1207,N_739,N_837);
and U1208 (N_1208,N_595,N_891);
xor U1209 (N_1209,N_613,N_965);
and U1210 (N_1210,N_591,N_688);
or U1211 (N_1211,N_676,N_905);
or U1212 (N_1212,N_766,N_509);
nand U1213 (N_1213,N_963,N_590);
xnor U1214 (N_1214,N_875,N_830);
and U1215 (N_1215,N_614,N_500);
and U1216 (N_1216,N_806,N_706);
and U1217 (N_1217,N_714,N_767);
nand U1218 (N_1218,N_573,N_967);
or U1219 (N_1219,N_970,N_914);
xnor U1220 (N_1220,N_561,N_898);
or U1221 (N_1221,N_942,N_966);
nand U1222 (N_1222,N_523,N_907);
nand U1223 (N_1223,N_784,N_955);
and U1224 (N_1224,N_740,N_790);
xnor U1225 (N_1225,N_737,N_852);
nor U1226 (N_1226,N_621,N_751);
and U1227 (N_1227,N_886,N_531);
or U1228 (N_1228,N_682,N_584);
or U1229 (N_1229,N_585,N_862);
xnor U1230 (N_1230,N_662,N_649);
and U1231 (N_1231,N_950,N_574);
xnor U1232 (N_1232,N_883,N_691);
nand U1233 (N_1233,N_660,N_515);
or U1234 (N_1234,N_679,N_769);
nor U1235 (N_1235,N_999,N_627);
and U1236 (N_1236,N_986,N_647);
and U1237 (N_1237,N_750,N_731);
nor U1238 (N_1238,N_511,N_877);
nor U1239 (N_1239,N_659,N_924);
and U1240 (N_1240,N_683,N_653);
or U1241 (N_1241,N_984,N_788);
or U1242 (N_1242,N_859,N_934);
and U1243 (N_1243,N_908,N_870);
xor U1244 (N_1244,N_736,N_745);
and U1245 (N_1245,N_656,N_700);
or U1246 (N_1246,N_645,N_978);
or U1247 (N_1247,N_983,N_943);
or U1248 (N_1248,N_861,N_949);
nand U1249 (N_1249,N_724,N_582);
or U1250 (N_1250,N_795,N_664);
nor U1251 (N_1251,N_529,N_577);
and U1252 (N_1252,N_747,N_977);
xor U1253 (N_1253,N_660,N_566);
nand U1254 (N_1254,N_945,N_541);
nand U1255 (N_1255,N_640,N_816);
nor U1256 (N_1256,N_824,N_730);
nor U1257 (N_1257,N_890,N_644);
nand U1258 (N_1258,N_628,N_510);
and U1259 (N_1259,N_549,N_991);
nand U1260 (N_1260,N_932,N_914);
xnor U1261 (N_1261,N_981,N_840);
and U1262 (N_1262,N_982,N_647);
or U1263 (N_1263,N_975,N_802);
and U1264 (N_1264,N_974,N_933);
or U1265 (N_1265,N_695,N_995);
and U1266 (N_1266,N_845,N_507);
and U1267 (N_1267,N_823,N_615);
nor U1268 (N_1268,N_995,N_946);
or U1269 (N_1269,N_967,N_948);
nand U1270 (N_1270,N_561,N_751);
xor U1271 (N_1271,N_618,N_617);
or U1272 (N_1272,N_521,N_873);
or U1273 (N_1273,N_789,N_997);
or U1274 (N_1274,N_512,N_596);
or U1275 (N_1275,N_521,N_921);
nor U1276 (N_1276,N_804,N_762);
nand U1277 (N_1277,N_761,N_948);
nand U1278 (N_1278,N_539,N_881);
xor U1279 (N_1279,N_963,N_790);
or U1280 (N_1280,N_894,N_729);
xnor U1281 (N_1281,N_960,N_686);
xnor U1282 (N_1282,N_612,N_923);
nor U1283 (N_1283,N_799,N_536);
nand U1284 (N_1284,N_726,N_888);
or U1285 (N_1285,N_683,N_859);
xor U1286 (N_1286,N_976,N_833);
nor U1287 (N_1287,N_965,N_591);
nor U1288 (N_1288,N_707,N_678);
nor U1289 (N_1289,N_760,N_666);
nor U1290 (N_1290,N_936,N_906);
nor U1291 (N_1291,N_825,N_841);
or U1292 (N_1292,N_815,N_894);
or U1293 (N_1293,N_990,N_551);
nor U1294 (N_1294,N_511,N_572);
and U1295 (N_1295,N_785,N_816);
and U1296 (N_1296,N_879,N_809);
nor U1297 (N_1297,N_712,N_998);
nor U1298 (N_1298,N_903,N_960);
nor U1299 (N_1299,N_685,N_533);
and U1300 (N_1300,N_958,N_997);
xor U1301 (N_1301,N_837,N_616);
xor U1302 (N_1302,N_856,N_854);
nand U1303 (N_1303,N_824,N_832);
xnor U1304 (N_1304,N_921,N_910);
and U1305 (N_1305,N_971,N_631);
nand U1306 (N_1306,N_937,N_839);
and U1307 (N_1307,N_977,N_516);
nor U1308 (N_1308,N_710,N_977);
nor U1309 (N_1309,N_822,N_833);
or U1310 (N_1310,N_662,N_973);
xor U1311 (N_1311,N_974,N_904);
xor U1312 (N_1312,N_880,N_625);
or U1313 (N_1313,N_612,N_993);
nand U1314 (N_1314,N_723,N_777);
xnor U1315 (N_1315,N_669,N_686);
xor U1316 (N_1316,N_899,N_879);
or U1317 (N_1317,N_956,N_592);
xnor U1318 (N_1318,N_768,N_942);
xnor U1319 (N_1319,N_572,N_917);
nand U1320 (N_1320,N_713,N_910);
nor U1321 (N_1321,N_924,N_603);
nor U1322 (N_1322,N_573,N_783);
and U1323 (N_1323,N_675,N_928);
or U1324 (N_1324,N_535,N_962);
xor U1325 (N_1325,N_671,N_761);
nand U1326 (N_1326,N_806,N_714);
nand U1327 (N_1327,N_840,N_615);
xor U1328 (N_1328,N_593,N_608);
xnor U1329 (N_1329,N_676,N_550);
nor U1330 (N_1330,N_604,N_903);
nor U1331 (N_1331,N_551,N_862);
and U1332 (N_1332,N_591,N_913);
and U1333 (N_1333,N_719,N_694);
xor U1334 (N_1334,N_875,N_966);
and U1335 (N_1335,N_804,N_888);
and U1336 (N_1336,N_541,N_782);
xor U1337 (N_1337,N_595,N_904);
nand U1338 (N_1338,N_513,N_859);
nand U1339 (N_1339,N_662,N_550);
xnor U1340 (N_1340,N_717,N_672);
or U1341 (N_1341,N_507,N_726);
and U1342 (N_1342,N_586,N_548);
and U1343 (N_1343,N_637,N_735);
or U1344 (N_1344,N_622,N_968);
nand U1345 (N_1345,N_699,N_712);
or U1346 (N_1346,N_699,N_952);
and U1347 (N_1347,N_719,N_697);
or U1348 (N_1348,N_872,N_697);
nor U1349 (N_1349,N_651,N_857);
nor U1350 (N_1350,N_627,N_706);
xnor U1351 (N_1351,N_940,N_740);
and U1352 (N_1352,N_980,N_775);
nor U1353 (N_1353,N_859,N_660);
or U1354 (N_1354,N_887,N_752);
nor U1355 (N_1355,N_520,N_928);
and U1356 (N_1356,N_806,N_598);
or U1357 (N_1357,N_709,N_751);
nor U1358 (N_1358,N_828,N_507);
xnor U1359 (N_1359,N_929,N_951);
nand U1360 (N_1360,N_980,N_755);
nor U1361 (N_1361,N_815,N_502);
xnor U1362 (N_1362,N_828,N_941);
xnor U1363 (N_1363,N_716,N_623);
and U1364 (N_1364,N_731,N_614);
nand U1365 (N_1365,N_787,N_996);
nand U1366 (N_1366,N_572,N_891);
and U1367 (N_1367,N_629,N_810);
or U1368 (N_1368,N_693,N_974);
nand U1369 (N_1369,N_598,N_943);
or U1370 (N_1370,N_675,N_713);
nand U1371 (N_1371,N_567,N_794);
or U1372 (N_1372,N_718,N_937);
and U1373 (N_1373,N_834,N_948);
xor U1374 (N_1374,N_926,N_556);
xor U1375 (N_1375,N_788,N_803);
nor U1376 (N_1376,N_976,N_938);
or U1377 (N_1377,N_824,N_937);
nor U1378 (N_1378,N_835,N_716);
nand U1379 (N_1379,N_782,N_660);
or U1380 (N_1380,N_914,N_535);
and U1381 (N_1381,N_747,N_729);
nand U1382 (N_1382,N_984,N_900);
and U1383 (N_1383,N_550,N_763);
nor U1384 (N_1384,N_595,N_991);
or U1385 (N_1385,N_855,N_897);
xor U1386 (N_1386,N_608,N_729);
nor U1387 (N_1387,N_802,N_762);
nor U1388 (N_1388,N_715,N_632);
nor U1389 (N_1389,N_710,N_737);
and U1390 (N_1390,N_611,N_992);
and U1391 (N_1391,N_506,N_638);
xor U1392 (N_1392,N_612,N_545);
xnor U1393 (N_1393,N_855,N_570);
xnor U1394 (N_1394,N_525,N_773);
nor U1395 (N_1395,N_516,N_727);
or U1396 (N_1396,N_666,N_800);
nand U1397 (N_1397,N_913,N_519);
nand U1398 (N_1398,N_556,N_589);
or U1399 (N_1399,N_689,N_906);
or U1400 (N_1400,N_671,N_690);
and U1401 (N_1401,N_802,N_921);
and U1402 (N_1402,N_653,N_634);
nor U1403 (N_1403,N_544,N_707);
or U1404 (N_1404,N_984,N_688);
and U1405 (N_1405,N_839,N_994);
or U1406 (N_1406,N_569,N_911);
nand U1407 (N_1407,N_590,N_983);
nand U1408 (N_1408,N_625,N_983);
xnor U1409 (N_1409,N_834,N_740);
nand U1410 (N_1410,N_629,N_926);
nand U1411 (N_1411,N_642,N_615);
or U1412 (N_1412,N_512,N_923);
or U1413 (N_1413,N_701,N_794);
xnor U1414 (N_1414,N_756,N_949);
or U1415 (N_1415,N_952,N_616);
and U1416 (N_1416,N_529,N_959);
or U1417 (N_1417,N_737,N_627);
xnor U1418 (N_1418,N_597,N_515);
nor U1419 (N_1419,N_746,N_709);
nor U1420 (N_1420,N_784,N_695);
or U1421 (N_1421,N_661,N_765);
and U1422 (N_1422,N_584,N_583);
xnor U1423 (N_1423,N_761,N_975);
nand U1424 (N_1424,N_541,N_743);
nor U1425 (N_1425,N_510,N_838);
nand U1426 (N_1426,N_806,N_775);
xor U1427 (N_1427,N_688,N_927);
nand U1428 (N_1428,N_555,N_530);
nand U1429 (N_1429,N_638,N_701);
xor U1430 (N_1430,N_826,N_864);
nor U1431 (N_1431,N_543,N_509);
or U1432 (N_1432,N_573,N_597);
or U1433 (N_1433,N_893,N_813);
nor U1434 (N_1434,N_607,N_789);
or U1435 (N_1435,N_978,N_560);
xor U1436 (N_1436,N_807,N_776);
xor U1437 (N_1437,N_798,N_988);
or U1438 (N_1438,N_617,N_725);
nand U1439 (N_1439,N_714,N_907);
nand U1440 (N_1440,N_962,N_748);
nand U1441 (N_1441,N_669,N_706);
nand U1442 (N_1442,N_709,N_752);
xor U1443 (N_1443,N_763,N_720);
nor U1444 (N_1444,N_609,N_908);
and U1445 (N_1445,N_969,N_923);
and U1446 (N_1446,N_886,N_969);
or U1447 (N_1447,N_792,N_691);
or U1448 (N_1448,N_781,N_825);
nand U1449 (N_1449,N_985,N_710);
nand U1450 (N_1450,N_899,N_991);
nor U1451 (N_1451,N_793,N_916);
and U1452 (N_1452,N_669,N_915);
nor U1453 (N_1453,N_765,N_769);
nand U1454 (N_1454,N_823,N_757);
nor U1455 (N_1455,N_514,N_882);
and U1456 (N_1456,N_672,N_814);
or U1457 (N_1457,N_561,N_620);
nor U1458 (N_1458,N_509,N_617);
or U1459 (N_1459,N_725,N_863);
or U1460 (N_1460,N_918,N_556);
nor U1461 (N_1461,N_932,N_535);
xor U1462 (N_1462,N_711,N_923);
xnor U1463 (N_1463,N_523,N_515);
nor U1464 (N_1464,N_900,N_590);
nand U1465 (N_1465,N_786,N_891);
nor U1466 (N_1466,N_585,N_736);
or U1467 (N_1467,N_717,N_766);
nor U1468 (N_1468,N_757,N_728);
xor U1469 (N_1469,N_996,N_762);
xnor U1470 (N_1470,N_564,N_895);
or U1471 (N_1471,N_544,N_748);
nor U1472 (N_1472,N_683,N_741);
nor U1473 (N_1473,N_610,N_717);
nor U1474 (N_1474,N_671,N_984);
or U1475 (N_1475,N_895,N_555);
nor U1476 (N_1476,N_538,N_888);
nand U1477 (N_1477,N_788,N_995);
or U1478 (N_1478,N_956,N_799);
or U1479 (N_1479,N_968,N_809);
xor U1480 (N_1480,N_961,N_537);
nand U1481 (N_1481,N_896,N_724);
nor U1482 (N_1482,N_528,N_684);
or U1483 (N_1483,N_655,N_842);
or U1484 (N_1484,N_966,N_726);
nor U1485 (N_1485,N_881,N_540);
or U1486 (N_1486,N_528,N_778);
xnor U1487 (N_1487,N_808,N_996);
nand U1488 (N_1488,N_882,N_919);
nor U1489 (N_1489,N_554,N_609);
xnor U1490 (N_1490,N_965,N_748);
or U1491 (N_1491,N_638,N_578);
nor U1492 (N_1492,N_936,N_615);
nor U1493 (N_1493,N_680,N_851);
nand U1494 (N_1494,N_679,N_584);
nand U1495 (N_1495,N_943,N_641);
and U1496 (N_1496,N_983,N_904);
nand U1497 (N_1497,N_722,N_500);
nor U1498 (N_1498,N_792,N_621);
or U1499 (N_1499,N_700,N_695);
or U1500 (N_1500,N_1472,N_1128);
xor U1501 (N_1501,N_1457,N_1251);
and U1502 (N_1502,N_1487,N_1443);
and U1503 (N_1503,N_1162,N_1151);
and U1504 (N_1504,N_1489,N_1070);
and U1505 (N_1505,N_1034,N_1125);
or U1506 (N_1506,N_1382,N_1355);
or U1507 (N_1507,N_1079,N_1248);
xor U1508 (N_1508,N_1337,N_1340);
xor U1509 (N_1509,N_1243,N_1395);
xnor U1510 (N_1510,N_1245,N_1038);
and U1511 (N_1511,N_1013,N_1447);
and U1512 (N_1512,N_1496,N_1313);
or U1513 (N_1513,N_1372,N_1390);
nand U1514 (N_1514,N_1271,N_1482);
nor U1515 (N_1515,N_1131,N_1366);
nor U1516 (N_1516,N_1189,N_1119);
nand U1517 (N_1517,N_1221,N_1270);
and U1518 (N_1518,N_1422,N_1357);
nor U1519 (N_1519,N_1264,N_1413);
nor U1520 (N_1520,N_1166,N_1027);
xnor U1521 (N_1521,N_1268,N_1102);
nor U1522 (N_1522,N_1406,N_1399);
and U1523 (N_1523,N_1330,N_1396);
nor U1524 (N_1524,N_1228,N_1242);
nor U1525 (N_1525,N_1109,N_1209);
or U1526 (N_1526,N_1187,N_1481);
nand U1527 (N_1527,N_1025,N_1118);
and U1528 (N_1528,N_1419,N_1218);
nand U1529 (N_1529,N_1149,N_1167);
and U1530 (N_1530,N_1344,N_1492);
or U1531 (N_1531,N_1081,N_1222);
nor U1532 (N_1532,N_1193,N_1021);
nand U1533 (N_1533,N_1283,N_1460);
xnor U1534 (N_1534,N_1009,N_1152);
xnor U1535 (N_1535,N_1381,N_1068);
xnor U1536 (N_1536,N_1310,N_1153);
or U1537 (N_1537,N_1425,N_1073);
nor U1538 (N_1538,N_1062,N_1142);
and U1539 (N_1539,N_1106,N_1232);
xor U1540 (N_1540,N_1329,N_1060);
or U1541 (N_1541,N_1072,N_1332);
or U1542 (N_1542,N_1449,N_1143);
or U1543 (N_1543,N_1050,N_1345);
nor U1544 (N_1544,N_1176,N_1173);
and U1545 (N_1545,N_1373,N_1227);
xnor U1546 (N_1546,N_1088,N_1260);
or U1547 (N_1547,N_1250,N_1308);
xor U1548 (N_1548,N_1266,N_1309);
nor U1549 (N_1549,N_1444,N_1331);
or U1550 (N_1550,N_1130,N_1219);
and U1551 (N_1551,N_1114,N_1277);
nand U1552 (N_1552,N_1267,N_1414);
nor U1553 (N_1553,N_1044,N_1324);
and U1554 (N_1554,N_1285,N_1158);
or U1555 (N_1555,N_1058,N_1233);
nand U1556 (N_1556,N_1354,N_1346);
nor U1557 (N_1557,N_1442,N_1408);
xnor U1558 (N_1558,N_1299,N_1090);
or U1559 (N_1559,N_1302,N_1418);
or U1560 (N_1560,N_1446,N_1435);
or U1561 (N_1561,N_1012,N_1104);
and U1562 (N_1562,N_1431,N_1107);
and U1563 (N_1563,N_1317,N_1005);
and U1564 (N_1564,N_1319,N_1279);
and U1565 (N_1565,N_1210,N_1469);
or U1566 (N_1566,N_1015,N_1334);
nor U1567 (N_1567,N_1259,N_1067);
or U1568 (N_1568,N_1437,N_1429);
and U1569 (N_1569,N_1365,N_1342);
nand U1570 (N_1570,N_1298,N_1179);
xor U1571 (N_1571,N_1402,N_1237);
nand U1572 (N_1572,N_1117,N_1417);
nand U1573 (N_1573,N_1111,N_1287);
and U1574 (N_1574,N_1147,N_1059);
or U1575 (N_1575,N_1076,N_1180);
nor U1576 (N_1576,N_1471,N_1273);
nand U1577 (N_1577,N_1224,N_1284);
nor U1578 (N_1578,N_1410,N_1083);
or U1579 (N_1579,N_1473,N_1168);
and U1580 (N_1580,N_1236,N_1007);
nand U1581 (N_1581,N_1363,N_1339);
nor U1582 (N_1582,N_1276,N_1169);
nand U1583 (N_1583,N_1433,N_1023);
nor U1584 (N_1584,N_1291,N_1199);
nor U1585 (N_1585,N_1369,N_1338);
xnor U1586 (N_1586,N_1001,N_1064);
nor U1587 (N_1587,N_1175,N_1392);
or U1588 (N_1588,N_1490,N_1141);
and U1589 (N_1589,N_1003,N_1416);
xnor U1590 (N_1590,N_1371,N_1010);
or U1591 (N_1591,N_1052,N_1434);
xnor U1592 (N_1592,N_1211,N_1108);
and U1593 (N_1593,N_1486,N_1470);
or U1594 (N_1594,N_1056,N_1194);
or U1595 (N_1595,N_1049,N_1134);
xor U1596 (N_1596,N_1451,N_1077);
or U1597 (N_1597,N_1439,N_1074);
or U1598 (N_1598,N_1499,N_1039);
nor U1599 (N_1599,N_1315,N_1206);
nand U1600 (N_1600,N_1322,N_1148);
xnor U1601 (N_1601,N_1184,N_1051);
and U1602 (N_1602,N_1293,N_1154);
xnor U1603 (N_1603,N_1030,N_1040);
nor U1604 (N_1604,N_1341,N_1286);
and U1605 (N_1605,N_1085,N_1105);
xor U1606 (N_1606,N_1181,N_1491);
nor U1607 (N_1607,N_1116,N_1412);
and U1608 (N_1608,N_1031,N_1476);
nand U1609 (N_1609,N_1378,N_1212);
or U1610 (N_1610,N_1427,N_1198);
or U1611 (N_1611,N_1343,N_1426);
or U1612 (N_1612,N_1132,N_1225);
nor U1613 (N_1613,N_1328,N_1098);
xor U1614 (N_1614,N_1112,N_1127);
nand U1615 (N_1615,N_1008,N_1288);
and U1616 (N_1616,N_1360,N_1367);
nor U1617 (N_1617,N_1475,N_1139);
and U1618 (N_1618,N_1186,N_1216);
or U1619 (N_1619,N_1424,N_1170);
and U1620 (N_1620,N_1163,N_1280);
or U1621 (N_1621,N_1485,N_1458);
and U1622 (N_1622,N_1226,N_1205);
xnor U1623 (N_1623,N_1230,N_1325);
xor U1624 (N_1624,N_1203,N_1483);
nor U1625 (N_1625,N_1089,N_1269);
or U1626 (N_1626,N_1071,N_1135);
or U1627 (N_1627,N_1235,N_1215);
and U1628 (N_1628,N_1093,N_1022);
nor U1629 (N_1629,N_1488,N_1327);
nor U1630 (N_1630,N_1004,N_1459);
xnor U1631 (N_1631,N_1465,N_1409);
nor U1632 (N_1632,N_1349,N_1249);
nor U1633 (N_1633,N_1165,N_1407);
nor U1634 (N_1634,N_1385,N_1454);
nor U1635 (N_1635,N_1244,N_1467);
nand U1636 (N_1636,N_1144,N_1024);
xor U1637 (N_1637,N_1188,N_1061);
nand U1638 (N_1638,N_1078,N_1045);
nand U1639 (N_1639,N_1404,N_1026);
and U1640 (N_1640,N_1428,N_1217);
nor U1641 (N_1641,N_1397,N_1042);
nor U1642 (N_1642,N_1137,N_1350);
or U1643 (N_1643,N_1182,N_1479);
or U1644 (N_1644,N_1359,N_1468);
nand U1645 (N_1645,N_1377,N_1477);
or U1646 (N_1646,N_1238,N_1438);
xnor U1647 (N_1647,N_1423,N_1202);
nor U1648 (N_1648,N_1497,N_1110);
or U1649 (N_1649,N_1281,N_1080);
xor U1650 (N_1650,N_1311,N_1348);
nand U1651 (N_1651,N_1290,N_1415);
xnor U1652 (N_1652,N_1095,N_1361);
nor U1653 (N_1653,N_1054,N_1140);
xnor U1654 (N_1654,N_1303,N_1389);
or U1655 (N_1655,N_1474,N_1032);
or U1656 (N_1656,N_1380,N_1306);
xnor U1657 (N_1657,N_1272,N_1033);
nor U1658 (N_1658,N_1092,N_1208);
and U1659 (N_1659,N_1261,N_1041);
nand U1660 (N_1660,N_1394,N_1048);
nor U1661 (N_1661,N_1164,N_1278);
xnor U1662 (N_1662,N_1159,N_1006);
and U1663 (N_1663,N_1126,N_1196);
xnor U1664 (N_1664,N_1150,N_1115);
or U1665 (N_1665,N_1157,N_1136);
or U1666 (N_1666,N_1352,N_1387);
xnor U1667 (N_1667,N_1047,N_1133);
nand U1668 (N_1668,N_1011,N_1453);
nand U1669 (N_1669,N_1065,N_1351);
nor U1670 (N_1670,N_1197,N_1314);
xor U1671 (N_1671,N_1356,N_1411);
nor U1672 (N_1672,N_1436,N_1375);
and U1673 (N_1673,N_1124,N_1300);
and U1674 (N_1674,N_1234,N_1020);
and U1675 (N_1675,N_1019,N_1318);
and U1676 (N_1676,N_1043,N_1246);
or U1677 (N_1677,N_1190,N_1174);
nand U1678 (N_1678,N_1214,N_1000);
and U1679 (N_1679,N_1305,N_1384);
xnor U1680 (N_1680,N_1069,N_1441);
xor U1681 (N_1681,N_1201,N_1253);
nand U1682 (N_1682,N_1240,N_1075);
and U1683 (N_1683,N_1057,N_1129);
or U1684 (N_1684,N_1018,N_1084);
and U1685 (N_1685,N_1398,N_1231);
or U1686 (N_1686,N_1401,N_1445);
xnor U1687 (N_1687,N_1494,N_1358);
nor U1688 (N_1688,N_1239,N_1316);
nor U1689 (N_1689,N_1220,N_1274);
xor U1690 (N_1690,N_1430,N_1323);
nand U1691 (N_1691,N_1333,N_1046);
nand U1692 (N_1692,N_1452,N_1321);
or U1693 (N_1693,N_1145,N_1263);
nand U1694 (N_1694,N_1368,N_1053);
nor U1695 (N_1695,N_1403,N_1002);
nand U1696 (N_1696,N_1461,N_1029);
nand U1697 (N_1697,N_1066,N_1466);
and U1698 (N_1698,N_1086,N_1087);
nor U1699 (N_1699,N_1036,N_1335);
nor U1700 (N_1700,N_1379,N_1495);
and U1701 (N_1701,N_1282,N_1037);
xor U1702 (N_1702,N_1462,N_1364);
and U1703 (N_1703,N_1195,N_1493);
nor U1704 (N_1704,N_1456,N_1320);
and U1705 (N_1705,N_1450,N_1391);
xor U1706 (N_1706,N_1156,N_1297);
nor U1707 (N_1707,N_1097,N_1405);
or U1708 (N_1708,N_1480,N_1160);
or U1709 (N_1709,N_1185,N_1241);
and U1710 (N_1710,N_1304,N_1183);
and U1711 (N_1711,N_1014,N_1207);
and U1712 (N_1712,N_1099,N_1296);
xnor U1713 (N_1713,N_1101,N_1258);
or U1714 (N_1714,N_1254,N_1312);
or U1715 (N_1715,N_1420,N_1123);
or U1716 (N_1716,N_1347,N_1055);
xor U1717 (N_1717,N_1388,N_1171);
nor U1718 (N_1718,N_1229,N_1155);
or U1719 (N_1719,N_1113,N_1200);
nor U1720 (N_1720,N_1301,N_1376);
and U1721 (N_1721,N_1256,N_1386);
or U1722 (N_1722,N_1172,N_1255);
or U1723 (N_1723,N_1063,N_1146);
nand U1724 (N_1724,N_1262,N_1383);
nor U1725 (N_1725,N_1478,N_1103);
nor U1726 (N_1726,N_1307,N_1275);
or U1727 (N_1727,N_1370,N_1138);
nor U1728 (N_1728,N_1265,N_1091);
and U1729 (N_1729,N_1464,N_1096);
nand U1730 (N_1730,N_1498,N_1161);
xor U1731 (N_1731,N_1421,N_1178);
xnor U1732 (N_1732,N_1035,N_1100);
nor U1733 (N_1733,N_1353,N_1393);
nand U1734 (N_1734,N_1294,N_1336);
xor U1735 (N_1735,N_1295,N_1463);
and U1736 (N_1736,N_1028,N_1121);
or U1737 (N_1737,N_1362,N_1292);
or U1738 (N_1738,N_1247,N_1400);
xnor U1739 (N_1739,N_1177,N_1440);
and U1740 (N_1740,N_1448,N_1374);
or U1741 (N_1741,N_1326,N_1016);
xnor U1742 (N_1742,N_1252,N_1432);
xor U1743 (N_1743,N_1082,N_1289);
nand U1744 (N_1744,N_1213,N_1455);
xor U1745 (N_1745,N_1191,N_1192);
xnor U1746 (N_1746,N_1257,N_1017);
or U1747 (N_1747,N_1204,N_1120);
and U1748 (N_1748,N_1122,N_1223);
nand U1749 (N_1749,N_1094,N_1484);
nor U1750 (N_1750,N_1132,N_1209);
or U1751 (N_1751,N_1437,N_1482);
nor U1752 (N_1752,N_1236,N_1402);
nor U1753 (N_1753,N_1035,N_1128);
and U1754 (N_1754,N_1078,N_1155);
and U1755 (N_1755,N_1070,N_1412);
nand U1756 (N_1756,N_1289,N_1086);
or U1757 (N_1757,N_1474,N_1197);
and U1758 (N_1758,N_1197,N_1342);
nand U1759 (N_1759,N_1018,N_1273);
nor U1760 (N_1760,N_1377,N_1106);
nand U1761 (N_1761,N_1000,N_1418);
xor U1762 (N_1762,N_1049,N_1276);
nand U1763 (N_1763,N_1137,N_1271);
xnor U1764 (N_1764,N_1292,N_1179);
or U1765 (N_1765,N_1393,N_1408);
nor U1766 (N_1766,N_1018,N_1198);
or U1767 (N_1767,N_1126,N_1127);
and U1768 (N_1768,N_1068,N_1127);
and U1769 (N_1769,N_1178,N_1470);
xor U1770 (N_1770,N_1338,N_1474);
and U1771 (N_1771,N_1113,N_1098);
xnor U1772 (N_1772,N_1251,N_1177);
xnor U1773 (N_1773,N_1390,N_1368);
or U1774 (N_1774,N_1213,N_1449);
or U1775 (N_1775,N_1327,N_1445);
xor U1776 (N_1776,N_1395,N_1354);
nand U1777 (N_1777,N_1174,N_1055);
nor U1778 (N_1778,N_1392,N_1447);
nor U1779 (N_1779,N_1066,N_1311);
xor U1780 (N_1780,N_1374,N_1227);
nand U1781 (N_1781,N_1466,N_1030);
nor U1782 (N_1782,N_1490,N_1497);
nor U1783 (N_1783,N_1166,N_1387);
or U1784 (N_1784,N_1349,N_1287);
nor U1785 (N_1785,N_1203,N_1256);
and U1786 (N_1786,N_1046,N_1212);
xor U1787 (N_1787,N_1396,N_1466);
nor U1788 (N_1788,N_1120,N_1229);
nand U1789 (N_1789,N_1357,N_1428);
and U1790 (N_1790,N_1488,N_1394);
xor U1791 (N_1791,N_1103,N_1012);
xnor U1792 (N_1792,N_1383,N_1399);
and U1793 (N_1793,N_1303,N_1346);
nand U1794 (N_1794,N_1206,N_1033);
or U1795 (N_1795,N_1126,N_1035);
nand U1796 (N_1796,N_1310,N_1279);
nor U1797 (N_1797,N_1177,N_1312);
or U1798 (N_1798,N_1022,N_1434);
xor U1799 (N_1799,N_1452,N_1448);
nand U1800 (N_1800,N_1478,N_1462);
nor U1801 (N_1801,N_1382,N_1428);
nand U1802 (N_1802,N_1412,N_1228);
and U1803 (N_1803,N_1441,N_1395);
nand U1804 (N_1804,N_1081,N_1475);
xor U1805 (N_1805,N_1469,N_1296);
and U1806 (N_1806,N_1215,N_1294);
or U1807 (N_1807,N_1376,N_1185);
or U1808 (N_1808,N_1211,N_1496);
xnor U1809 (N_1809,N_1382,N_1239);
nor U1810 (N_1810,N_1398,N_1484);
nor U1811 (N_1811,N_1113,N_1032);
or U1812 (N_1812,N_1168,N_1397);
nand U1813 (N_1813,N_1107,N_1220);
nor U1814 (N_1814,N_1218,N_1097);
or U1815 (N_1815,N_1325,N_1438);
xor U1816 (N_1816,N_1499,N_1323);
and U1817 (N_1817,N_1072,N_1184);
nor U1818 (N_1818,N_1281,N_1126);
or U1819 (N_1819,N_1318,N_1013);
nand U1820 (N_1820,N_1098,N_1114);
or U1821 (N_1821,N_1308,N_1433);
xnor U1822 (N_1822,N_1448,N_1139);
xnor U1823 (N_1823,N_1328,N_1006);
or U1824 (N_1824,N_1193,N_1113);
nor U1825 (N_1825,N_1017,N_1143);
and U1826 (N_1826,N_1023,N_1425);
or U1827 (N_1827,N_1120,N_1371);
nor U1828 (N_1828,N_1327,N_1395);
xnor U1829 (N_1829,N_1475,N_1025);
or U1830 (N_1830,N_1273,N_1096);
nor U1831 (N_1831,N_1084,N_1024);
nand U1832 (N_1832,N_1265,N_1155);
or U1833 (N_1833,N_1189,N_1192);
nand U1834 (N_1834,N_1432,N_1206);
and U1835 (N_1835,N_1239,N_1486);
or U1836 (N_1836,N_1165,N_1183);
nor U1837 (N_1837,N_1443,N_1284);
or U1838 (N_1838,N_1210,N_1402);
nor U1839 (N_1839,N_1415,N_1365);
nor U1840 (N_1840,N_1469,N_1223);
or U1841 (N_1841,N_1007,N_1439);
nand U1842 (N_1842,N_1077,N_1439);
or U1843 (N_1843,N_1364,N_1013);
and U1844 (N_1844,N_1451,N_1122);
and U1845 (N_1845,N_1413,N_1225);
xnor U1846 (N_1846,N_1332,N_1079);
nand U1847 (N_1847,N_1472,N_1273);
or U1848 (N_1848,N_1453,N_1358);
and U1849 (N_1849,N_1157,N_1087);
nor U1850 (N_1850,N_1180,N_1168);
or U1851 (N_1851,N_1013,N_1235);
xnor U1852 (N_1852,N_1480,N_1344);
and U1853 (N_1853,N_1088,N_1157);
xnor U1854 (N_1854,N_1232,N_1065);
xor U1855 (N_1855,N_1241,N_1298);
or U1856 (N_1856,N_1067,N_1499);
nor U1857 (N_1857,N_1303,N_1290);
or U1858 (N_1858,N_1248,N_1449);
xor U1859 (N_1859,N_1216,N_1490);
nand U1860 (N_1860,N_1287,N_1402);
or U1861 (N_1861,N_1091,N_1273);
xor U1862 (N_1862,N_1004,N_1467);
nor U1863 (N_1863,N_1084,N_1205);
and U1864 (N_1864,N_1359,N_1175);
or U1865 (N_1865,N_1224,N_1142);
and U1866 (N_1866,N_1386,N_1128);
or U1867 (N_1867,N_1446,N_1136);
nand U1868 (N_1868,N_1029,N_1448);
or U1869 (N_1869,N_1030,N_1108);
and U1870 (N_1870,N_1334,N_1345);
nand U1871 (N_1871,N_1456,N_1195);
and U1872 (N_1872,N_1012,N_1092);
nor U1873 (N_1873,N_1200,N_1039);
or U1874 (N_1874,N_1416,N_1196);
nand U1875 (N_1875,N_1030,N_1412);
or U1876 (N_1876,N_1228,N_1257);
nand U1877 (N_1877,N_1121,N_1313);
and U1878 (N_1878,N_1360,N_1300);
nand U1879 (N_1879,N_1296,N_1404);
and U1880 (N_1880,N_1362,N_1080);
nor U1881 (N_1881,N_1393,N_1172);
xor U1882 (N_1882,N_1306,N_1387);
xor U1883 (N_1883,N_1070,N_1430);
xnor U1884 (N_1884,N_1444,N_1314);
or U1885 (N_1885,N_1448,N_1379);
xor U1886 (N_1886,N_1343,N_1498);
nor U1887 (N_1887,N_1487,N_1281);
or U1888 (N_1888,N_1330,N_1135);
and U1889 (N_1889,N_1048,N_1184);
or U1890 (N_1890,N_1108,N_1359);
or U1891 (N_1891,N_1355,N_1419);
or U1892 (N_1892,N_1023,N_1049);
xor U1893 (N_1893,N_1417,N_1311);
and U1894 (N_1894,N_1186,N_1148);
nor U1895 (N_1895,N_1142,N_1287);
and U1896 (N_1896,N_1288,N_1284);
xnor U1897 (N_1897,N_1279,N_1400);
nand U1898 (N_1898,N_1054,N_1348);
or U1899 (N_1899,N_1087,N_1016);
nand U1900 (N_1900,N_1421,N_1176);
nand U1901 (N_1901,N_1315,N_1124);
nand U1902 (N_1902,N_1482,N_1246);
nand U1903 (N_1903,N_1132,N_1001);
and U1904 (N_1904,N_1030,N_1413);
or U1905 (N_1905,N_1128,N_1222);
or U1906 (N_1906,N_1102,N_1338);
nor U1907 (N_1907,N_1141,N_1261);
or U1908 (N_1908,N_1027,N_1321);
nor U1909 (N_1909,N_1143,N_1178);
nand U1910 (N_1910,N_1364,N_1041);
nor U1911 (N_1911,N_1431,N_1233);
and U1912 (N_1912,N_1431,N_1101);
nor U1913 (N_1913,N_1356,N_1453);
nand U1914 (N_1914,N_1431,N_1244);
nand U1915 (N_1915,N_1161,N_1484);
nand U1916 (N_1916,N_1051,N_1016);
or U1917 (N_1917,N_1243,N_1295);
nor U1918 (N_1918,N_1194,N_1123);
and U1919 (N_1919,N_1125,N_1035);
and U1920 (N_1920,N_1209,N_1281);
xnor U1921 (N_1921,N_1323,N_1159);
or U1922 (N_1922,N_1078,N_1261);
xnor U1923 (N_1923,N_1128,N_1366);
nor U1924 (N_1924,N_1446,N_1402);
xnor U1925 (N_1925,N_1056,N_1030);
nand U1926 (N_1926,N_1067,N_1111);
nor U1927 (N_1927,N_1090,N_1274);
xnor U1928 (N_1928,N_1208,N_1197);
nand U1929 (N_1929,N_1317,N_1212);
xor U1930 (N_1930,N_1375,N_1061);
nor U1931 (N_1931,N_1446,N_1422);
nand U1932 (N_1932,N_1411,N_1424);
xnor U1933 (N_1933,N_1264,N_1421);
nand U1934 (N_1934,N_1424,N_1225);
nand U1935 (N_1935,N_1354,N_1147);
nor U1936 (N_1936,N_1131,N_1077);
and U1937 (N_1937,N_1124,N_1100);
nand U1938 (N_1938,N_1268,N_1269);
nor U1939 (N_1939,N_1341,N_1316);
nand U1940 (N_1940,N_1183,N_1414);
or U1941 (N_1941,N_1211,N_1170);
or U1942 (N_1942,N_1468,N_1270);
xnor U1943 (N_1943,N_1442,N_1190);
or U1944 (N_1944,N_1456,N_1353);
and U1945 (N_1945,N_1302,N_1031);
and U1946 (N_1946,N_1372,N_1135);
nor U1947 (N_1947,N_1023,N_1202);
nor U1948 (N_1948,N_1345,N_1482);
xnor U1949 (N_1949,N_1470,N_1346);
nand U1950 (N_1950,N_1043,N_1378);
xnor U1951 (N_1951,N_1411,N_1324);
and U1952 (N_1952,N_1474,N_1350);
nor U1953 (N_1953,N_1479,N_1197);
nand U1954 (N_1954,N_1146,N_1223);
or U1955 (N_1955,N_1011,N_1043);
nand U1956 (N_1956,N_1159,N_1195);
xnor U1957 (N_1957,N_1440,N_1081);
and U1958 (N_1958,N_1359,N_1205);
or U1959 (N_1959,N_1187,N_1266);
and U1960 (N_1960,N_1215,N_1063);
nand U1961 (N_1961,N_1003,N_1367);
nor U1962 (N_1962,N_1058,N_1308);
and U1963 (N_1963,N_1141,N_1396);
and U1964 (N_1964,N_1138,N_1111);
or U1965 (N_1965,N_1150,N_1455);
or U1966 (N_1966,N_1326,N_1242);
or U1967 (N_1967,N_1107,N_1127);
nor U1968 (N_1968,N_1266,N_1359);
or U1969 (N_1969,N_1260,N_1480);
nand U1970 (N_1970,N_1156,N_1375);
or U1971 (N_1971,N_1275,N_1116);
or U1972 (N_1972,N_1450,N_1203);
nor U1973 (N_1973,N_1460,N_1288);
nand U1974 (N_1974,N_1346,N_1180);
and U1975 (N_1975,N_1373,N_1034);
or U1976 (N_1976,N_1210,N_1006);
and U1977 (N_1977,N_1416,N_1480);
or U1978 (N_1978,N_1320,N_1413);
and U1979 (N_1979,N_1413,N_1441);
or U1980 (N_1980,N_1494,N_1288);
and U1981 (N_1981,N_1442,N_1062);
and U1982 (N_1982,N_1439,N_1258);
or U1983 (N_1983,N_1286,N_1129);
nand U1984 (N_1984,N_1115,N_1341);
and U1985 (N_1985,N_1278,N_1049);
xnor U1986 (N_1986,N_1009,N_1425);
and U1987 (N_1987,N_1075,N_1353);
or U1988 (N_1988,N_1374,N_1189);
and U1989 (N_1989,N_1378,N_1240);
or U1990 (N_1990,N_1488,N_1345);
or U1991 (N_1991,N_1123,N_1362);
nor U1992 (N_1992,N_1355,N_1397);
nand U1993 (N_1993,N_1390,N_1495);
or U1994 (N_1994,N_1217,N_1385);
nand U1995 (N_1995,N_1232,N_1133);
nor U1996 (N_1996,N_1172,N_1141);
xnor U1997 (N_1997,N_1349,N_1124);
xnor U1998 (N_1998,N_1370,N_1308);
xnor U1999 (N_1999,N_1316,N_1479);
nand U2000 (N_2000,N_1791,N_1793);
or U2001 (N_2001,N_1821,N_1705);
xor U2002 (N_2002,N_1538,N_1586);
xor U2003 (N_2003,N_1978,N_1870);
nand U2004 (N_2004,N_1945,N_1703);
xor U2005 (N_2005,N_1588,N_1755);
xor U2006 (N_2006,N_1545,N_1908);
or U2007 (N_2007,N_1925,N_1949);
or U2008 (N_2008,N_1604,N_1515);
xor U2009 (N_2009,N_1943,N_1894);
nor U2010 (N_2010,N_1546,N_1881);
nor U2011 (N_2011,N_1552,N_1666);
xor U2012 (N_2012,N_1979,N_1628);
nand U2013 (N_2013,N_1873,N_1960);
xor U2014 (N_2014,N_1686,N_1562);
nand U2015 (N_2015,N_1851,N_1688);
nand U2016 (N_2016,N_1748,N_1639);
or U2017 (N_2017,N_1939,N_1869);
and U2018 (N_2018,N_1579,N_1745);
nor U2019 (N_2019,N_1836,N_1554);
nor U2020 (N_2020,N_1665,N_1685);
nand U2021 (N_2021,N_1569,N_1811);
and U2022 (N_2022,N_1504,N_1996);
or U2023 (N_2023,N_1754,N_1935);
xor U2024 (N_2024,N_1541,N_1779);
nor U2025 (N_2025,N_1721,N_1601);
nand U2026 (N_2026,N_1809,N_1897);
nor U2027 (N_2027,N_1929,N_1618);
nand U2028 (N_2028,N_1527,N_1884);
xor U2029 (N_2029,N_1875,N_1871);
nor U2030 (N_2030,N_1623,N_1673);
nor U2031 (N_2031,N_1531,N_1612);
and U2032 (N_2032,N_1707,N_1728);
and U2033 (N_2033,N_1550,N_1994);
xnor U2034 (N_2034,N_1933,N_1658);
xnor U2035 (N_2035,N_1764,N_1828);
and U2036 (N_2036,N_1891,N_1782);
nor U2037 (N_2037,N_1906,N_1563);
xor U2038 (N_2038,N_1578,N_1787);
nand U2039 (N_2039,N_1689,N_1656);
or U2040 (N_2040,N_1711,N_1564);
nor U2041 (N_2041,N_1700,N_1566);
nand U2042 (N_2042,N_1766,N_1786);
nor U2043 (N_2043,N_1885,N_1937);
nand U2044 (N_2044,N_1626,N_1972);
nand U2045 (N_2045,N_1681,N_1931);
nor U2046 (N_2046,N_1610,N_1888);
nor U2047 (N_2047,N_1968,N_1783);
and U2048 (N_2048,N_1505,N_1962);
nand U2049 (N_2049,N_1825,N_1558);
xnor U2050 (N_2050,N_1990,N_1989);
and U2051 (N_2051,N_1657,N_1668);
and U2052 (N_2052,N_1544,N_1606);
nand U2053 (N_2053,N_1892,N_1854);
xor U2054 (N_2054,N_1723,N_1502);
nor U2055 (N_2055,N_1820,N_1918);
nor U2056 (N_2056,N_1777,N_1883);
nor U2057 (N_2057,N_1549,N_1812);
xor U2058 (N_2058,N_1636,N_1722);
nor U2059 (N_2059,N_1853,N_1773);
nor U2060 (N_2060,N_1838,N_1655);
nor U2061 (N_2061,N_1907,N_1739);
and U2062 (N_2062,N_1613,N_1852);
and U2063 (N_2063,N_1916,N_1924);
nor U2064 (N_2064,N_1800,N_1726);
and U2065 (N_2065,N_1518,N_1631);
nor U2066 (N_2066,N_1983,N_1622);
and U2067 (N_2067,N_1860,N_1798);
nand U2068 (N_2068,N_1704,N_1583);
nand U2069 (N_2069,N_1827,N_1734);
and U2070 (N_2070,N_1915,N_1625);
nand U2071 (N_2071,N_1950,N_1605);
nor U2072 (N_2072,N_1671,N_1822);
or U2073 (N_2073,N_1732,N_1946);
nand U2074 (N_2074,N_1620,N_1682);
and U2075 (N_2075,N_1697,N_1910);
xor U2076 (N_2076,N_1667,N_1751);
nor U2077 (N_2077,N_1699,N_1857);
and U2078 (N_2078,N_1867,N_1815);
xnor U2079 (N_2079,N_1953,N_1535);
and U2080 (N_2080,N_1593,N_1634);
and U2081 (N_2081,N_1547,N_1517);
or U2082 (N_2082,N_1847,N_1765);
xor U2083 (N_2083,N_1619,N_1647);
nand U2084 (N_2084,N_1584,N_1621);
xor U2085 (N_2085,N_1653,N_1927);
or U2086 (N_2086,N_1904,N_1698);
nor U2087 (N_2087,N_1823,N_1900);
nand U2088 (N_2088,N_1651,N_1780);
xnor U2089 (N_2089,N_1982,N_1794);
and U2090 (N_2090,N_1887,N_1540);
nor U2091 (N_2091,N_1942,N_1627);
and U2092 (N_2092,N_1767,N_1865);
or U2093 (N_2093,N_1992,N_1679);
xnor U2094 (N_2094,N_1642,N_1874);
or U2095 (N_2095,N_1597,N_1724);
nand U2096 (N_2096,N_1720,N_1781);
nor U2097 (N_2097,N_1889,N_1746);
nand U2098 (N_2098,N_1824,N_1980);
xor U2099 (N_2099,N_1633,N_1839);
xnor U2100 (N_2100,N_1876,N_1961);
nand U2101 (N_2101,N_1710,N_1810);
nor U2102 (N_2102,N_1877,N_1941);
nand U2103 (N_2103,N_1737,N_1932);
and U2104 (N_2104,N_1696,N_1760);
nand U2105 (N_2105,N_1947,N_1714);
or U2106 (N_2106,N_1801,N_1757);
and U2107 (N_2107,N_1512,N_1784);
nor U2108 (N_2108,N_1832,N_1997);
or U2109 (N_2109,N_1845,N_1572);
nand U2110 (N_2110,N_1725,N_1763);
nor U2111 (N_2111,N_1969,N_1591);
or U2112 (N_2112,N_1774,N_1635);
or U2113 (N_2113,N_1955,N_1503);
nor U2114 (N_2114,N_1829,N_1596);
and U2115 (N_2115,N_1802,N_1848);
and U2116 (N_2116,N_1902,N_1532);
xnor U2117 (N_2117,N_1690,N_1988);
nor U2118 (N_2118,N_1501,N_1510);
xnor U2119 (N_2119,N_1589,N_1818);
nand U2120 (N_2120,N_1788,N_1921);
xor U2121 (N_2121,N_1677,N_1716);
or U2122 (N_2122,N_1542,N_1903);
xor U2123 (N_2123,N_1617,N_1598);
or U2124 (N_2124,N_1956,N_1567);
or U2125 (N_2125,N_1595,N_1736);
xnor U2126 (N_2126,N_1500,N_1599);
and U2127 (N_2127,N_1831,N_1930);
nand U2128 (N_2128,N_1514,N_1638);
nand U2129 (N_2129,N_1749,N_1813);
and U2130 (N_2130,N_1652,N_1523);
nand U2131 (N_2131,N_1521,N_1806);
nand U2132 (N_2132,N_1646,N_1528);
xnor U2133 (N_2133,N_1731,N_1624);
or U2134 (N_2134,N_1967,N_1868);
and U2135 (N_2135,N_1923,N_1835);
xor U2136 (N_2136,N_1592,N_1577);
nand U2137 (N_2137,N_1938,N_1778);
or U2138 (N_2138,N_1678,N_1609);
nand U2139 (N_2139,N_1744,N_1849);
or U2140 (N_2140,N_1742,N_1758);
or U2141 (N_2141,N_1603,N_1664);
or U2142 (N_2142,N_1808,N_1743);
or U2143 (N_2143,N_1899,N_1555);
nor U2144 (N_2144,N_1833,N_1675);
nor U2145 (N_2145,N_1785,N_1771);
nand U2146 (N_2146,N_1807,N_1981);
nand U2147 (N_2147,N_1987,N_1843);
nor U2148 (N_2148,N_1525,N_1740);
nor U2149 (N_2149,N_1896,N_1600);
or U2150 (N_2150,N_1975,N_1973);
nor U2151 (N_2151,N_1886,N_1509);
and U2152 (N_2152,N_1640,N_1846);
xor U2153 (N_2153,N_1676,N_1669);
and U2154 (N_2154,N_1615,N_1752);
and U2155 (N_2155,N_1717,N_1893);
and U2156 (N_2156,N_1861,N_1805);
nand U2157 (N_2157,N_1692,N_1934);
nor U2158 (N_2158,N_1702,N_1912);
xor U2159 (N_2159,N_1769,N_1650);
and U2160 (N_2160,N_1993,N_1574);
nand U2161 (N_2161,N_1630,N_1855);
nand U2162 (N_2162,N_1970,N_1995);
nor U2163 (N_2163,N_1866,N_1901);
or U2164 (N_2164,N_1837,N_1695);
nand U2165 (N_2165,N_1898,N_1984);
nand U2166 (N_2166,N_1706,N_1506);
and U2167 (N_2167,N_1952,N_1772);
or U2168 (N_2168,N_1738,N_1519);
or U2169 (N_2169,N_1804,N_1974);
and U2170 (N_2170,N_1641,N_1797);
or U2171 (N_2171,N_1928,N_1733);
or U2172 (N_2172,N_1520,N_1850);
nand U2173 (N_2173,N_1998,N_1911);
nand U2174 (N_2174,N_1880,N_1963);
xnor U2175 (N_2175,N_1792,N_1580);
and U2176 (N_2176,N_1718,N_1663);
or U2177 (N_2177,N_1844,N_1922);
nand U2178 (N_2178,N_1560,N_1856);
nand U2179 (N_2179,N_1735,N_1576);
or U2180 (N_2180,N_1795,N_1776);
xor U2181 (N_2181,N_1712,N_1645);
xnor U2182 (N_2182,N_1661,N_1878);
or U2183 (N_2183,N_1819,N_1954);
and U2184 (N_2184,N_1557,N_1608);
xor U2185 (N_2185,N_1508,N_1834);
and U2186 (N_2186,N_1602,N_1693);
and U2187 (N_2187,N_1709,N_1660);
or U2188 (N_2188,N_1985,N_1756);
nor U2189 (N_2189,N_1768,N_1533);
nand U2190 (N_2190,N_1529,N_1530);
nand U2191 (N_2191,N_1537,N_1775);
or U2192 (N_2192,N_1715,N_1582);
and U2193 (N_2193,N_1573,N_1522);
or U2194 (N_2194,N_1799,N_1536);
or U2195 (N_2195,N_1687,N_1770);
nor U2196 (N_2196,N_1614,N_1971);
nor U2197 (N_2197,N_1571,N_1581);
nor U2198 (N_2198,N_1905,N_1548);
and U2199 (N_2199,N_1914,N_1882);
and U2200 (N_2200,N_1513,N_1729);
nand U2201 (N_2201,N_1659,N_1859);
nand U2202 (N_2202,N_1830,N_1649);
xor U2203 (N_2203,N_1858,N_1919);
or U2204 (N_2204,N_1568,N_1790);
xor U2205 (N_2205,N_1727,N_1803);
nand U2206 (N_2206,N_1879,N_1585);
and U2207 (N_2207,N_1570,N_1977);
or U2208 (N_2208,N_1670,N_1926);
or U2209 (N_2209,N_1594,N_1951);
or U2210 (N_2210,N_1936,N_1730);
xnor U2211 (N_2211,N_1637,N_1959);
or U2212 (N_2212,N_1511,N_1565);
and U2213 (N_2213,N_1920,N_1999);
nand U2214 (N_2214,N_1862,N_1826);
or U2215 (N_2215,N_1587,N_1762);
or U2216 (N_2216,N_1632,N_1539);
and U2217 (N_2217,N_1691,N_1607);
nand U2218 (N_2218,N_1648,N_1543);
or U2219 (N_2219,N_1913,N_1611);
or U2220 (N_2220,N_1551,N_1948);
xor U2221 (N_2221,N_1629,N_1840);
nor U2222 (N_2222,N_1556,N_1864);
or U2223 (N_2223,N_1741,N_1701);
or U2224 (N_2224,N_1672,N_1817);
nand U2225 (N_2225,N_1507,N_1863);
xor U2226 (N_2226,N_1753,N_1680);
nand U2227 (N_2227,N_1986,N_1814);
or U2228 (N_2228,N_1684,N_1524);
and U2229 (N_2229,N_1654,N_1516);
or U2230 (N_2230,N_1872,N_1957);
nand U2231 (N_2231,N_1958,N_1674);
or U2232 (N_2232,N_1761,N_1976);
or U2233 (N_2233,N_1944,N_1917);
nand U2234 (N_2234,N_1940,N_1842);
and U2235 (N_2235,N_1747,N_1816);
or U2236 (N_2236,N_1719,N_1694);
nand U2237 (N_2237,N_1964,N_1683);
or U2238 (N_2238,N_1750,N_1708);
or U2239 (N_2239,N_1662,N_1561);
or U2240 (N_2240,N_1643,N_1616);
or U2241 (N_2241,N_1526,N_1759);
xnor U2242 (N_2242,N_1991,N_1575);
or U2243 (N_2243,N_1644,N_1965);
nor U2244 (N_2244,N_1909,N_1796);
or U2245 (N_2245,N_1713,N_1966);
nand U2246 (N_2246,N_1559,N_1590);
and U2247 (N_2247,N_1841,N_1789);
xor U2248 (N_2248,N_1553,N_1895);
and U2249 (N_2249,N_1534,N_1890);
xnor U2250 (N_2250,N_1881,N_1918);
or U2251 (N_2251,N_1730,N_1848);
and U2252 (N_2252,N_1761,N_1794);
nand U2253 (N_2253,N_1867,N_1633);
or U2254 (N_2254,N_1620,N_1986);
or U2255 (N_2255,N_1889,N_1766);
or U2256 (N_2256,N_1816,N_1905);
or U2257 (N_2257,N_1889,N_1747);
and U2258 (N_2258,N_1910,N_1892);
nor U2259 (N_2259,N_1663,N_1788);
nand U2260 (N_2260,N_1733,N_1625);
or U2261 (N_2261,N_1652,N_1870);
xnor U2262 (N_2262,N_1708,N_1584);
nand U2263 (N_2263,N_1848,N_1617);
and U2264 (N_2264,N_1806,N_1944);
xor U2265 (N_2265,N_1846,N_1801);
nand U2266 (N_2266,N_1963,N_1780);
or U2267 (N_2267,N_1966,N_1564);
and U2268 (N_2268,N_1901,N_1653);
xor U2269 (N_2269,N_1616,N_1606);
xor U2270 (N_2270,N_1692,N_1608);
nor U2271 (N_2271,N_1626,N_1888);
or U2272 (N_2272,N_1864,N_1841);
xor U2273 (N_2273,N_1718,N_1792);
nor U2274 (N_2274,N_1521,N_1979);
nand U2275 (N_2275,N_1750,N_1600);
xor U2276 (N_2276,N_1959,N_1604);
nand U2277 (N_2277,N_1659,N_1614);
xor U2278 (N_2278,N_1941,N_1989);
xnor U2279 (N_2279,N_1961,N_1850);
and U2280 (N_2280,N_1962,N_1595);
xor U2281 (N_2281,N_1825,N_1514);
or U2282 (N_2282,N_1668,N_1862);
nor U2283 (N_2283,N_1945,N_1883);
or U2284 (N_2284,N_1984,N_1654);
nor U2285 (N_2285,N_1751,N_1669);
xnor U2286 (N_2286,N_1616,N_1842);
and U2287 (N_2287,N_1513,N_1622);
xor U2288 (N_2288,N_1528,N_1754);
and U2289 (N_2289,N_1774,N_1507);
nor U2290 (N_2290,N_1979,N_1549);
nor U2291 (N_2291,N_1620,N_1696);
or U2292 (N_2292,N_1706,N_1618);
or U2293 (N_2293,N_1688,N_1574);
and U2294 (N_2294,N_1840,N_1816);
nand U2295 (N_2295,N_1500,N_1720);
or U2296 (N_2296,N_1726,N_1799);
xnor U2297 (N_2297,N_1680,N_1708);
and U2298 (N_2298,N_1546,N_1582);
and U2299 (N_2299,N_1930,N_1858);
or U2300 (N_2300,N_1850,N_1741);
and U2301 (N_2301,N_1671,N_1813);
xnor U2302 (N_2302,N_1612,N_1953);
nand U2303 (N_2303,N_1760,N_1572);
or U2304 (N_2304,N_1748,N_1545);
nor U2305 (N_2305,N_1504,N_1979);
and U2306 (N_2306,N_1624,N_1786);
nor U2307 (N_2307,N_1516,N_1699);
and U2308 (N_2308,N_1943,N_1680);
nand U2309 (N_2309,N_1535,N_1735);
nand U2310 (N_2310,N_1715,N_1759);
xor U2311 (N_2311,N_1896,N_1760);
nand U2312 (N_2312,N_1952,N_1823);
nor U2313 (N_2313,N_1653,N_1536);
nor U2314 (N_2314,N_1927,N_1513);
or U2315 (N_2315,N_1920,N_1842);
nor U2316 (N_2316,N_1555,N_1666);
and U2317 (N_2317,N_1512,N_1697);
or U2318 (N_2318,N_1811,N_1686);
nor U2319 (N_2319,N_1887,N_1706);
xor U2320 (N_2320,N_1711,N_1861);
xnor U2321 (N_2321,N_1529,N_1719);
xor U2322 (N_2322,N_1943,N_1582);
xnor U2323 (N_2323,N_1909,N_1801);
xor U2324 (N_2324,N_1660,N_1539);
xnor U2325 (N_2325,N_1708,N_1843);
nand U2326 (N_2326,N_1619,N_1622);
xor U2327 (N_2327,N_1575,N_1769);
xor U2328 (N_2328,N_1603,N_1940);
nor U2329 (N_2329,N_1717,N_1828);
and U2330 (N_2330,N_1624,N_1752);
or U2331 (N_2331,N_1714,N_1899);
and U2332 (N_2332,N_1907,N_1569);
and U2333 (N_2333,N_1672,N_1846);
or U2334 (N_2334,N_1675,N_1929);
and U2335 (N_2335,N_1908,N_1503);
nand U2336 (N_2336,N_1821,N_1735);
xnor U2337 (N_2337,N_1864,N_1684);
nor U2338 (N_2338,N_1706,N_1885);
nand U2339 (N_2339,N_1687,N_1608);
and U2340 (N_2340,N_1947,N_1929);
or U2341 (N_2341,N_1967,N_1991);
or U2342 (N_2342,N_1874,N_1772);
nor U2343 (N_2343,N_1928,N_1831);
nor U2344 (N_2344,N_1926,N_1727);
xor U2345 (N_2345,N_1810,N_1576);
nor U2346 (N_2346,N_1702,N_1960);
or U2347 (N_2347,N_1819,N_1516);
and U2348 (N_2348,N_1924,N_1757);
or U2349 (N_2349,N_1993,N_1698);
and U2350 (N_2350,N_1821,N_1520);
xnor U2351 (N_2351,N_1504,N_1845);
nand U2352 (N_2352,N_1622,N_1675);
or U2353 (N_2353,N_1561,N_1635);
xnor U2354 (N_2354,N_1901,N_1887);
or U2355 (N_2355,N_1754,N_1948);
nor U2356 (N_2356,N_1996,N_1516);
nor U2357 (N_2357,N_1637,N_1872);
and U2358 (N_2358,N_1735,N_1508);
and U2359 (N_2359,N_1989,N_1872);
and U2360 (N_2360,N_1852,N_1997);
nand U2361 (N_2361,N_1726,N_1607);
and U2362 (N_2362,N_1971,N_1647);
or U2363 (N_2363,N_1785,N_1743);
nor U2364 (N_2364,N_1793,N_1869);
or U2365 (N_2365,N_1645,N_1698);
or U2366 (N_2366,N_1675,N_1505);
nor U2367 (N_2367,N_1715,N_1885);
nand U2368 (N_2368,N_1590,N_1738);
nor U2369 (N_2369,N_1966,N_1707);
xor U2370 (N_2370,N_1799,N_1822);
and U2371 (N_2371,N_1615,N_1654);
or U2372 (N_2372,N_1984,N_1688);
and U2373 (N_2373,N_1718,N_1969);
and U2374 (N_2374,N_1607,N_1787);
and U2375 (N_2375,N_1591,N_1811);
xnor U2376 (N_2376,N_1653,N_1986);
or U2377 (N_2377,N_1744,N_1640);
and U2378 (N_2378,N_1867,N_1989);
xor U2379 (N_2379,N_1621,N_1931);
or U2380 (N_2380,N_1659,N_1662);
nor U2381 (N_2381,N_1923,N_1561);
nand U2382 (N_2382,N_1827,N_1890);
nor U2383 (N_2383,N_1722,N_1529);
nand U2384 (N_2384,N_1653,N_1512);
xor U2385 (N_2385,N_1527,N_1824);
nand U2386 (N_2386,N_1922,N_1562);
and U2387 (N_2387,N_1823,N_1951);
or U2388 (N_2388,N_1669,N_1944);
and U2389 (N_2389,N_1917,N_1503);
or U2390 (N_2390,N_1833,N_1618);
and U2391 (N_2391,N_1851,N_1542);
or U2392 (N_2392,N_1860,N_1931);
or U2393 (N_2393,N_1950,N_1683);
nand U2394 (N_2394,N_1841,N_1576);
or U2395 (N_2395,N_1657,N_1957);
xor U2396 (N_2396,N_1929,N_1536);
and U2397 (N_2397,N_1552,N_1894);
nor U2398 (N_2398,N_1884,N_1902);
or U2399 (N_2399,N_1609,N_1602);
or U2400 (N_2400,N_1562,N_1648);
or U2401 (N_2401,N_1942,N_1767);
nand U2402 (N_2402,N_1655,N_1821);
and U2403 (N_2403,N_1565,N_1876);
and U2404 (N_2404,N_1791,N_1948);
and U2405 (N_2405,N_1871,N_1782);
or U2406 (N_2406,N_1636,N_1609);
nor U2407 (N_2407,N_1602,N_1526);
nand U2408 (N_2408,N_1732,N_1758);
nor U2409 (N_2409,N_1867,N_1826);
xnor U2410 (N_2410,N_1971,N_1994);
nand U2411 (N_2411,N_1764,N_1891);
nand U2412 (N_2412,N_1716,N_1523);
or U2413 (N_2413,N_1817,N_1587);
and U2414 (N_2414,N_1800,N_1692);
nand U2415 (N_2415,N_1941,N_1824);
xnor U2416 (N_2416,N_1963,N_1987);
and U2417 (N_2417,N_1857,N_1723);
nor U2418 (N_2418,N_1602,N_1538);
and U2419 (N_2419,N_1699,N_1838);
nand U2420 (N_2420,N_1588,N_1917);
xnor U2421 (N_2421,N_1726,N_1951);
nor U2422 (N_2422,N_1939,N_1516);
xnor U2423 (N_2423,N_1626,N_1727);
nand U2424 (N_2424,N_1946,N_1594);
xnor U2425 (N_2425,N_1795,N_1726);
and U2426 (N_2426,N_1792,N_1541);
or U2427 (N_2427,N_1738,N_1960);
and U2428 (N_2428,N_1793,N_1618);
nand U2429 (N_2429,N_1787,N_1844);
nor U2430 (N_2430,N_1660,N_1673);
xor U2431 (N_2431,N_1810,N_1566);
nor U2432 (N_2432,N_1699,N_1711);
or U2433 (N_2433,N_1883,N_1900);
nand U2434 (N_2434,N_1809,N_1847);
nor U2435 (N_2435,N_1921,N_1505);
and U2436 (N_2436,N_1653,N_1668);
xnor U2437 (N_2437,N_1632,N_1721);
xor U2438 (N_2438,N_1659,N_1952);
nand U2439 (N_2439,N_1558,N_1926);
and U2440 (N_2440,N_1568,N_1507);
nand U2441 (N_2441,N_1821,N_1512);
and U2442 (N_2442,N_1603,N_1767);
nor U2443 (N_2443,N_1593,N_1571);
or U2444 (N_2444,N_1765,N_1655);
or U2445 (N_2445,N_1553,N_1551);
or U2446 (N_2446,N_1634,N_1961);
and U2447 (N_2447,N_1698,N_1644);
nand U2448 (N_2448,N_1585,N_1682);
xnor U2449 (N_2449,N_1926,N_1536);
or U2450 (N_2450,N_1800,N_1558);
xnor U2451 (N_2451,N_1976,N_1603);
xnor U2452 (N_2452,N_1634,N_1660);
nor U2453 (N_2453,N_1717,N_1732);
nor U2454 (N_2454,N_1583,N_1891);
nand U2455 (N_2455,N_1836,N_1888);
xnor U2456 (N_2456,N_1797,N_1632);
and U2457 (N_2457,N_1727,N_1814);
xnor U2458 (N_2458,N_1853,N_1723);
and U2459 (N_2459,N_1680,N_1904);
nor U2460 (N_2460,N_1601,N_1505);
nand U2461 (N_2461,N_1826,N_1538);
or U2462 (N_2462,N_1695,N_1601);
and U2463 (N_2463,N_1693,N_1622);
xor U2464 (N_2464,N_1830,N_1697);
xor U2465 (N_2465,N_1880,N_1997);
or U2466 (N_2466,N_1712,N_1970);
nand U2467 (N_2467,N_1539,N_1530);
and U2468 (N_2468,N_1508,N_1793);
nand U2469 (N_2469,N_1917,N_1828);
and U2470 (N_2470,N_1859,N_1680);
and U2471 (N_2471,N_1922,N_1734);
nor U2472 (N_2472,N_1806,N_1526);
xor U2473 (N_2473,N_1981,N_1727);
and U2474 (N_2474,N_1735,N_1924);
and U2475 (N_2475,N_1929,N_1767);
nand U2476 (N_2476,N_1685,N_1671);
nand U2477 (N_2477,N_1815,N_1907);
xor U2478 (N_2478,N_1704,N_1875);
nand U2479 (N_2479,N_1746,N_1996);
nor U2480 (N_2480,N_1659,N_1549);
and U2481 (N_2481,N_1909,N_1919);
xor U2482 (N_2482,N_1682,N_1837);
and U2483 (N_2483,N_1665,N_1905);
nand U2484 (N_2484,N_1665,N_1628);
nor U2485 (N_2485,N_1615,N_1694);
xnor U2486 (N_2486,N_1839,N_1735);
nand U2487 (N_2487,N_1711,N_1741);
nand U2488 (N_2488,N_1786,N_1719);
xor U2489 (N_2489,N_1504,N_1959);
or U2490 (N_2490,N_1800,N_1898);
nor U2491 (N_2491,N_1965,N_1533);
or U2492 (N_2492,N_1549,N_1597);
and U2493 (N_2493,N_1680,N_1812);
nor U2494 (N_2494,N_1567,N_1716);
nor U2495 (N_2495,N_1869,N_1721);
nor U2496 (N_2496,N_1895,N_1587);
and U2497 (N_2497,N_1992,N_1529);
xnor U2498 (N_2498,N_1655,N_1608);
and U2499 (N_2499,N_1546,N_1677);
or U2500 (N_2500,N_2433,N_2386);
and U2501 (N_2501,N_2369,N_2481);
nand U2502 (N_2502,N_2385,N_2151);
or U2503 (N_2503,N_2488,N_2462);
xnor U2504 (N_2504,N_2147,N_2222);
nand U2505 (N_2505,N_2145,N_2317);
and U2506 (N_2506,N_2059,N_2336);
nand U2507 (N_2507,N_2326,N_2171);
and U2508 (N_2508,N_2069,N_2475);
or U2509 (N_2509,N_2003,N_2377);
xnor U2510 (N_2510,N_2306,N_2409);
and U2511 (N_2511,N_2008,N_2213);
xnor U2512 (N_2512,N_2159,N_2262);
and U2513 (N_2513,N_2299,N_2286);
nand U2514 (N_2514,N_2248,N_2174);
nor U2515 (N_2515,N_2494,N_2391);
or U2516 (N_2516,N_2132,N_2044);
xor U2517 (N_2517,N_2428,N_2035);
xnor U2518 (N_2518,N_2071,N_2247);
nand U2519 (N_2519,N_2404,N_2118);
or U2520 (N_2520,N_2129,N_2175);
xnor U2521 (N_2521,N_2162,N_2339);
nor U2522 (N_2522,N_2446,N_2289);
xnor U2523 (N_2523,N_2472,N_2471);
nand U2524 (N_2524,N_2414,N_2215);
nor U2525 (N_2525,N_2293,N_2020);
nand U2526 (N_2526,N_2070,N_2013);
or U2527 (N_2527,N_2460,N_2359);
and U2528 (N_2528,N_2148,N_2100);
nand U2529 (N_2529,N_2393,N_2420);
nand U2530 (N_2530,N_2028,N_2250);
or U2531 (N_2531,N_2268,N_2373);
nor U2532 (N_2532,N_2130,N_2455);
and U2533 (N_2533,N_2240,N_2001);
xor U2534 (N_2534,N_2410,N_2018);
xnor U2535 (N_2535,N_2218,N_2110);
and U2536 (N_2536,N_2038,N_2115);
and U2537 (N_2537,N_2355,N_2083);
and U2538 (N_2538,N_2439,N_2228);
or U2539 (N_2539,N_2040,N_2170);
nor U2540 (N_2540,N_2492,N_2114);
nand U2541 (N_2541,N_2036,N_2230);
nand U2542 (N_2542,N_2353,N_2382);
nand U2543 (N_2543,N_2352,N_2113);
or U2544 (N_2544,N_2011,N_2208);
nor U2545 (N_2545,N_2107,N_2039);
nor U2546 (N_2546,N_2201,N_2067);
xnor U2547 (N_2547,N_2229,N_2027);
and U2548 (N_2548,N_2227,N_2241);
or U2549 (N_2549,N_2243,N_2088);
or U2550 (N_2550,N_2368,N_2180);
nor U2551 (N_2551,N_2402,N_2161);
and U2552 (N_2552,N_2146,N_2451);
and U2553 (N_2553,N_2477,N_2205);
nor U2554 (N_2554,N_2023,N_2275);
nor U2555 (N_2555,N_2407,N_2032);
and U2556 (N_2556,N_2127,N_2281);
and U2557 (N_2557,N_2330,N_2366);
nor U2558 (N_2558,N_2332,N_2342);
nor U2559 (N_2559,N_2207,N_2497);
xor U2560 (N_2560,N_2046,N_2450);
xnor U2561 (N_2561,N_2438,N_2285);
xnor U2562 (N_2562,N_2469,N_2102);
nor U2563 (N_2563,N_2394,N_2203);
and U2564 (N_2564,N_2349,N_2133);
or U2565 (N_2565,N_2436,N_2081);
nor U2566 (N_2566,N_2406,N_2354);
nand U2567 (N_2567,N_2097,N_2112);
and U2568 (N_2568,N_2474,N_2362);
xnor U2569 (N_2569,N_2415,N_2264);
and U2570 (N_2570,N_2154,N_2026);
xnor U2571 (N_2571,N_2290,N_2282);
or U2572 (N_2572,N_2374,N_2186);
xor U2573 (N_2573,N_2403,N_2172);
nand U2574 (N_2574,N_2379,N_2153);
or U2575 (N_2575,N_2210,N_2358);
or U2576 (N_2576,N_2395,N_2237);
nor U2577 (N_2577,N_2457,N_2164);
nor U2578 (N_2578,N_2074,N_2337);
nand U2579 (N_2579,N_2126,N_2273);
nand U2580 (N_2580,N_2284,N_2263);
and U2581 (N_2581,N_2425,N_2421);
xor U2582 (N_2582,N_2177,N_2458);
or U2583 (N_2583,N_2217,N_2104);
or U2584 (N_2584,N_2198,N_2030);
nor U2585 (N_2585,N_2328,N_2052);
or U2586 (N_2586,N_2291,N_2183);
or U2587 (N_2587,N_2463,N_2086);
nand U2588 (N_2588,N_2305,N_2370);
and U2589 (N_2589,N_2345,N_2189);
nor U2590 (N_2590,N_2312,N_2223);
nor U2591 (N_2591,N_2434,N_2489);
nand U2592 (N_2592,N_2004,N_2109);
or U2593 (N_2593,N_2271,N_2192);
nor U2594 (N_2594,N_2065,N_2498);
and U2595 (N_2595,N_2002,N_2194);
xnor U2596 (N_2596,N_2412,N_2288);
nor U2597 (N_2597,N_2350,N_2343);
and U2598 (N_2598,N_2371,N_2009);
nor U2599 (N_2599,N_2378,N_2453);
and U2600 (N_2600,N_2231,N_2466);
and U2601 (N_2601,N_2125,N_2401);
nand U2602 (N_2602,N_2033,N_2073);
nor U2603 (N_2603,N_2155,N_2441);
or U2604 (N_2604,N_2259,N_2445);
nand U2605 (N_2605,N_2120,N_2266);
and U2606 (N_2606,N_2051,N_2260);
and U2607 (N_2607,N_2322,N_2456);
nor U2608 (N_2608,N_2238,N_2309);
or U2609 (N_2609,N_2021,N_2209);
and U2610 (N_2610,N_2485,N_2478);
nor U2611 (N_2611,N_2212,N_2117);
nor U2612 (N_2612,N_2029,N_2276);
xnor U2613 (N_2613,N_2136,N_2448);
and U2614 (N_2614,N_2311,N_2007);
or U2615 (N_2615,N_2016,N_2157);
nand U2616 (N_2616,N_2211,N_2224);
and U2617 (N_2617,N_2464,N_2307);
xnor U2618 (N_2618,N_2341,N_2367);
xor U2619 (N_2619,N_2054,N_2300);
and U2620 (N_2620,N_2200,N_2142);
or U2621 (N_2621,N_2356,N_2252);
and U2622 (N_2622,N_2078,N_2495);
or U2623 (N_2623,N_2010,N_2169);
or U2624 (N_2624,N_2048,N_2121);
xnor U2625 (N_2625,N_2150,N_2184);
xor U2626 (N_2626,N_2105,N_2167);
or U2627 (N_2627,N_2221,N_2465);
and U2628 (N_2628,N_2216,N_2031);
nand U2629 (N_2629,N_2427,N_2388);
xnor U2630 (N_2630,N_2302,N_2050);
nand U2631 (N_2631,N_2075,N_2443);
xnor U2632 (N_2632,N_2123,N_2079);
xnor U2633 (N_2633,N_2043,N_2015);
or U2634 (N_2634,N_2012,N_2098);
nand U2635 (N_2635,N_2139,N_2468);
nor U2636 (N_2636,N_2258,N_2249);
nand U2637 (N_2637,N_2197,N_2178);
or U2638 (N_2638,N_2041,N_2274);
xor U2639 (N_2639,N_2442,N_2017);
nand U2640 (N_2640,N_2049,N_2236);
or U2641 (N_2641,N_2255,N_2280);
nand U2642 (N_2642,N_2483,N_2437);
nand U2643 (N_2643,N_2314,N_2246);
nand U2644 (N_2644,N_2072,N_2278);
nand U2645 (N_2645,N_2400,N_2480);
xnor U2646 (N_2646,N_2424,N_2068);
nand U2647 (N_2647,N_2430,N_2411);
and U2648 (N_2648,N_2242,N_2256);
nor U2649 (N_2649,N_2364,N_2496);
nand U2650 (N_2650,N_2426,N_2484);
or U2651 (N_2651,N_2296,N_2416);
or U2652 (N_2652,N_2333,N_2270);
and U2653 (N_2653,N_2389,N_2063);
or U2654 (N_2654,N_2392,N_2251);
xnor U2655 (N_2655,N_2181,N_2323);
and U2656 (N_2656,N_2327,N_2479);
xnor U2657 (N_2657,N_2244,N_2057);
nand U2658 (N_2658,N_2094,N_2091);
and U2659 (N_2659,N_2099,N_2316);
or U2660 (N_2660,N_2160,N_2396);
or U2661 (N_2661,N_2245,N_2076);
or U2662 (N_2662,N_2253,N_2319);
xnor U2663 (N_2663,N_2085,N_2152);
and U2664 (N_2664,N_2380,N_2297);
or U2665 (N_2665,N_2025,N_2053);
xor U2666 (N_2666,N_2493,N_2196);
xor U2667 (N_2667,N_2476,N_2254);
xnor U2668 (N_2668,N_2348,N_2277);
and U2669 (N_2669,N_2234,N_2419);
nand U2670 (N_2670,N_2335,N_2166);
nand U2671 (N_2671,N_2357,N_2173);
and U2672 (N_2672,N_2176,N_2056);
or U2673 (N_2673,N_2320,N_2321);
nand U2674 (N_2674,N_2179,N_2141);
or U2675 (N_2675,N_2116,N_2313);
nor U2676 (N_2676,N_2294,N_2204);
nor U2677 (N_2677,N_2324,N_2301);
and U2678 (N_2678,N_2344,N_2449);
nand U2679 (N_2679,N_2137,N_2444);
nand U2680 (N_2680,N_2233,N_2135);
nor U2681 (N_2681,N_2206,N_2019);
and U2682 (N_2682,N_2066,N_2077);
xnor U2683 (N_2683,N_2239,N_2232);
or U2684 (N_2684,N_2287,N_2214);
xnor U2685 (N_2685,N_2134,N_2191);
nand U2686 (N_2686,N_2383,N_2226);
nand U2687 (N_2687,N_2408,N_2140);
xor U2688 (N_2688,N_2417,N_2338);
xor U2689 (N_2689,N_2062,N_2340);
xnor U2690 (N_2690,N_2045,N_2461);
xor U2691 (N_2691,N_2034,N_2398);
nor U2692 (N_2692,N_2363,N_2298);
nor U2693 (N_2693,N_2482,N_2101);
and U2694 (N_2694,N_2225,N_2182);
or U2695 (N_2695,N_2304,N_2199);
or U2696 (N_2696,N_2149,N_2156);
or U2697 (N_2697,N_2390,N_2108);
or U2698 (N_2698,N_2470,N_2318);
xor U2699 (N_2699,N_2459,N_2202);
xor U2700 (N_2700,N_2060,N_2376);
xor U2701 (N_2701,N_2190,N_2165);
nor U2702 (N_2702,N_2005,N_2124);
nand U2703 (N_2703,N_2257,N_2014);
xor U2704 (N_2704,N_2486,N_2490);
and U2705 (N_2705,N_2095,N_2128);
xnor U2706 (N_2706,N_2106,N_2087);
nand U2707 (N_2707,N_2384,N_2447);
nand U2708 (N_2708,N_2315,N_2295);
nand U2709 (N_2709,N_2047,N_2283);
nor U2710 (N_2710,N_2090,N_2413);
or U2711 (N_2711,N_2055,N_2487);
and U2712 (N_2712,N_2185,N_2397);
nand U2713 (N_2713,N_2022,N_2122);
nand U2714 (N_2714,N_2452,N_2000);
nand U2715 (N_2715,N_2308,N_2096);
xor U2716 (N_2716,N_2279,N_2499);
and U2717 (N_2717,N_2361,N_2405);
xnor U2718 (N_2718,N_2360,N_2372);
nand U2719 (N_2719,N_2331,N_2491);
xnor U2720 (N_2720,N_2061,N_2292);
or U2721 (N_2721,N_2435,N_2473);
nor U2722 (N_2722,N_2265,N_2163);
xor U2723 (N_2723,N_2058,N_2423);
and U2724 (N_2724,N_2387,N_2334);
nor U2725 (N_2725,N_2235,N_2467);
nand U2726 (N_2726,N_2347,N_2024);
or U2727 (N_2727,N_2351,N_2440);
nor U2728 (N_2728,N_2219,N_2381);
nor U2729 (N_2729,N_2365,N_2158);
or U2730 (N_2730,N_2143,N_2272);
or U2731 (N_2731,N_2111,N_2310);
and U2732 (N_2732,N_2267,N_2064);
nand U2733 (N_2733,N_2269,N_2080);
nor U2734 (N_2734,N_2187,N_2093);
xnor U2735 (N_2735,N_2422,N_2084);
and U2736 (N_2736,N_2193,N_2375);
and U2737 (N_2737,N_2454,N_2399);
nor U2738 (N_2738,N_2325,N_2082);
or U2739 (N_2739,N_2119,N_2188);
and U2740 (N_2740,N_2089,N_2037);
xor U2741 (N_2741,N_2092,N_2429);
xnor U2742 (N_2742,N_2168,N_2138);
xnor U2743 (N_2743,N_2220,N_2131);
nand U2744 (N_2744,N_2431,N_2418);
or U2745 (N_2745,N_2329,N_2042);
or U2746 (N_2746,N_2006,N_2261);
nor U2747 (N_2747,N_2432,N_2103);
nor U2748 (N_2748,N_2346,N_2144);
or U2749 (N_2749,N_2195,N_2303);
or U2750 (N_2750,N_2164,N_2089);
nand U2751 (N_2751,N_2235,N_2454);
nand U2752 (N_2752,N_2123,N_2087);
xnor U2753 (N_2753,N_2332,N_2387);
and U2754 (N_2754,N_2402,N_2289);
or U2755 (N_2755,N_2294,N_2039);
nor U2756 (N_2756,N_2289,N_2386);
or U2757 (N_2757,N_2331,N_2482);
or U2758 (N_2758,N_2182,N_2106);
xnor U2759 (N_2759,N_2350,N_2083);
or U2760 (N_2760,N_2367,N_2134);
and U2761 (N_2761,N_2386,N_2442);
and U2762 (N_2762,N_2426,N_2435);
xor U2763 (N_2763,N_2338,N_2458);
or U2764 (N_2764,N_2371,N_2166);
or U2765 (N_2765,N_2150,N_2361);
and U2766 (N_2766,N_2300,N_2469);
or U2767 (N_2767,N_2485,N_2448);
or U2768 (N_2768,N_2147,N_2157);
xnor U2769 (N_2769,N_2281,N_2286);
or U2770 (N_2770,N_2075,N_2199);
nand U2771 (N_2771,N_2159,N_2104);
and U2772 (N_2772,N_2390,N_2492);
nor U2773 (N_2773,N_2148,N_2154);
nor U2774 (N_2774,N_2369,N_2021);
or U2775 (N_2775,N_2205,N_2450);
nor U2776 (N_2776,N_2042,N_2116);
xnor U2777 (N_2777,N_2229,N_2269);
xor U2778 (N_2778,N_2034,N_2428);
xor U2779 (N_2779,N_2049,N_2235);
xnor U2780 (N_2780,N_2034,N_2449);
xor U2781 (N_2781,N_2016,N_2293);
xor U2782 (N_2782,N_2242,N_2198);
or U2783 (N_2783,N_2160,N_2037);
and U2784 (N_2784,N_2111,N_2005);
and U2785 (N_2785,N_2014,N_2304);
nor U2786 (N_2786,N_2176,N_2304);
xor U2787 (N_2787,N_2390,N_2064);
nor U2788 (N_2788,N_2043,N_2063);
nand U2789 (N_2789,N_2003,N_2211);
nand U2790 (N_2790,N_2112,N_2429);
xor U2791 (N_2791,N_2350,N_2458);
or U2792 (N_2792,N_2038,N_2102);
nand U2793 (N_2793,N_2363,N_2456);
and U2794 (N_2794,N_2423,N_2025);
or U2795 (N_2795,N_2021,N_2441);
xor U2796 (N_2796,N_2149,N_2444);
or U2797 (N_2797,N_2298,N_2140);
and U2798 (N_2798,N_2332,N_2038);
and U2799 (N_2799,N_2342,N_2093);
nand U2800 (N_2800,N_2167,N_2268);
and U2801 (N_2801,N_2164,N_2088);
xor U2802 (N_2802,N_2354,N_2116);
and U2803 (N_2803,N_2351,N_2157);
or U2804 (N_2804,N_2014,N_2174);
and U2805 (N_2805,N_2179,N_2394);
and U2806 (N_2806,N_2395,N_2218);
xnor U2807 (N_2807,N_2378,N_2158);
xnor U2808 (N_2808,N_2387,N_2024);
xnor U2809 (N_2809,N_2410,N_2217);
nand U2810 (N_2810,N_2015,N_2341);
and U2811 (N_2811,N_2068,N_2293);
or U2812 (N_2812,N_2283,N_2458);
nor U2813 (N_2813,N_2011,N_2311);
and U2814 (N_2814,N_2131,N_2349);
nor U2815 (N_2815,N_2312,N_2207);
xor U2816 (N_2816,N_2099,N_2255);
nand U2817 (N_2817,N_2113,N_2118);
or U2818 (N_2818,N_2337,N_2272);
or U2819 (N_2819,N_2163,N_2418);
nand U2820 (N_2820,N_2037,N_2151);
nand U2821 (N_2821,N_2296,N_2221);
nor U2822 (N_2822,N_2111,N_2212);
nand U2823 (N_2823,N_2082,N_2066);
nor U2824 (N_2824,N_2133,N_2132);
xor U2825 (N_2825,N_2048,N_2054);
and U2826 (N_2826,N_2443,N_2042);
nand U2827 (N_2827,N_2349,N_2088);
and U2828 (N_2828,N_2133,N_2437);
xnor U2829 (N_2829,N_2238,N_2083);
or U2830 (N_2830,N_2368,N_2039);
nand U2831 (N_2831,N_2220,N_2355);
and U2832 (N_2832,N_2125,N_2094);
xor U2833 (N_2833,N_2102,N_2359);
nand U2834 (N_2834,N_2090,N_2068);
nand U2835 (N_2835,N_2307,N_2198);
nand U2836 (N_2836,N_2223,N_2044);
and U2837 (N_2837,N_2155,N_2382);
xor U2838 (N_2838,N_2218,N_2012);
xor U2839 (N_2839,N_2173,N_2432);
and U2840 (N_2840,N_2156,N_2391);
and U2841 (N_2841,N_2351,N_2066);
nand U2842 (N_2842,N_2229,N_2366);
nand U2843 (N_2843,N_2283,N_2300);
nor U2844 (N_2844,N_2383,N_2079);
nor U2845 (N_2845,N_2071,N_2005);
nand U2846 (N_2846,N_2102,N_2393);
nand U2847 (N_2847,N_2487,N_2048);
or U2848 (N_2848,N_2198,N_2393);
xnor U2849 (N_2849,N_2358,N_2396);
nand U2850 (N_2850,N_2411,N_2424);
nand U2851 (N_2851,N_2316,N_2388);
and U2852 (N_2852,N_2428,N_2455);
xor U2853 (N_2853,N_2015,N_2158);
and U2854 (N_2854,N_2460,N_2467);
xor U2855 (N_2855,N_2332,N_2205);
nand U2856 (N_2856,N_2300,N_2251);
and U2857 (N_2857,N_2458,N_2152);
nor U2858 (N_2858,N_2301,N_2087);
xor U2859 (N_2859,N_2417,N_2468);
and U2860 (N_2860,N_2110,N_2347);
and U2861 (N_2861,N_2332,N_2408);
xor U2862 (N_2862,N_2062,N_2153);
nor U2863 (N_2863,N_2343,N_2298);
nand U2864 (N_2864,N_2040,N_2256);
and U2865 (N_2865,N_2424,N_2105);
or U2866 (N_2866,N_2017,N_2361);
and U2867 (N_2867,N_2341,N_2014);
and U2868 (N_2868,N_2016,N_2310);
nor U2869 (N_2869,N_2365,N_2243);
or U2870 (N_2870,N_2097,N_2294);
and U2871 (N_2871,N_2464,N_2390);
and U2872 (N_2872,N_2433,N_2106);
nor U2873 (N_2873,N_2232,N_2021);
nand U2874 (N_2874,N_2498,N_2073);
and U2875 (N_2875,N_2452,N_2306);
and U2876 (N_2876,N_2373,N_2393);
nand U2877 (N_2877,N_2440,N_2338);
or U2878 (N_2878,N_2379,N_2371);
and U2879 (N_2879,N_2290,N_2112);
xnor U2880 (N_2880,N_2068,N_2197);
nand U2881 (N_2881,N_2144,N_2361);
nand U2882 (N_2882,N_2444,N_2190);
or U2883 (N_2883,N_2420,N_2321);
xor U2884 (N_2884,N_2190,N_2219);
nor U2885 (N_2885,N_2143,N_2253);
xnor U2886 (N_2886,N_2266,N_2476);
or U2887 (N_2887,N_2205,N_2129);
and U2888 (N_2888,N_2057,N_2490);
xor U2889 (N_2889,N_2260,N_2359);
nor U2890 (N_2890,N_2161,N_2469);
nor U2891 (N_2891,N_2092,N_2280);
xor U2892 (N_2892,N_2027,N_2315);
xnor U2893 (N_2893,N_2427,N_2221);
nand U2894 (N_2894,N_2338,N_2339);
xnor U2895 (N_2895,N_2235,N_2017);
nand U2896 (N_2896,N_2017,N_2419);
xnor U2897 (N_2897,N_2230,N_2084);
nand U2898 (N_2898,N_2373,N_2213);
xor U2899 (N_2899,N_2224,N_2415);
nor U2900 (N_2900,N_2285,N_2353);
or U2901 (N_2901,N_2330,N_2425);
and U2902 (N_2902,N_2191,N_2064);
and U2903 (N_2903,N_2001,N_2035);
xnor U2904 (N_2904,N_2302,N_2147);
or U2905 (N_2905,N_2001,N_2034);
nor U2906 (N_2906,N_2151,N_2033);
and U2907 (N_2907,N_2490,N_2436);
and U2908 (N_2908,N_2043,N_2241);
nand U2909 (N_2909,N_2082,N_2210);
xor U2910 (N_2910,N_2179,N_2305);
nor U2911 (N_2911,N_2489,N_2136);
and U2912 (N_2912,N_2046,N_2261);
nand U2913 (N_2913,N_2299,N_2450);
nor U2914 (N_2914,N_2454,N_2432);
nand U2915 (N_2915,N_2090,N_2114);
nand U2916 (N_2916,N_2418,N_2351);
nand U2917 (N_2917,N_2462,N_2295);
and U2918 (N_2918,N_2355,N_2244);
nand U2919 (N_2919,N_2094,N_2313);
and U2920 (N_2920,N_2342,N_2462);
nor U2921 (N_2921,N_2328,N_2043);
xor U2922 (N_2922,N_2329,N_2050);
or U2923 (N_2923,N_2334,N_2073);
or U2924 (N_2924,N_2366,N_2034);
or U2925 (N_2925,N_2424,N_2072);
nor U2926 (N_2926,N_2044,N_2443);
nor U2927 (N_2927,N_2012,N_2128);
or U2928 (N_2928,N_2451,N_2314);
xnor U2929 (N_2929,N_2141,N_2185);
nand U2930 (N_2930,N_2297,N_2121);
nand U2931 (N_2931,N_2009,N_2175);
nor U2932 (N_2932,N_2101,N_2058);
xnor U2933 (N_2933,N_2447,N_2084);
nand U2934 (N_2934,N_2156,N_2108);
nor U2935 (N_2935,N_2180,N_2470);
nand U2936 (N_2936,N_2463,N_2102);
xor U2937 (N_2937,N_2343,N_2281);
nor U2938 (N_2938,N_2336,N_2268);
or U2939 (N_2939,N_2180,N_2284);
or U2940 (N_2940,N_2150,N_2274);
or U2941 (N_2941,N_2459,N_2233);
or U2942 (N_2942,N_2109,N_2053);
or U2943 (N_2943,N_2244,N_2121);
or U2944 (N_2944,N_2042,N_2251);
nor U2945 (N_2945,N_2230,N_2426);
nand U2946 (N_2946,N_2221,N_2327);
and U2947 (N_2947,N_2361,N_2383);
and U2948 (N_2948,N_2235,N_2461);
nand U2949 (N_2949,N_2005,N_2416);
or U2950 (N_2950,N_2199,N_2423);
and U2951 (N_2951,N_2470,N_2186);
and U2952 (N_2952,N_2432,N_2433);
nor U2953 (N_2953,N_2090,N_2340);
nor U2954 (N_2954,N_2379,N_2150);
xor U2955 (N_2955,N_2334,N_2466);
or U2956 (N_2956,N_2455,N_2075);
and U2957 (N_2957,N_2240,N_2266);
xnor U2958 (N_2958,N_2105,N_2440);
nor U2959 (N_2959,N_2077,N_2065);
and U2960 (N_2960,N_2265,N_2110);
nand U2961 (N_2961,N_2233,N_2495);
nor U2962 (N_2962,N_2264,N_2341);
nand U2963 (N_2963,N_2352,N_2311);
nand U2964 (N_2964,N_2450,N_2487);
nand U2965 (N_2965,N_2218,N_2254);
nor U2966 (N_2966,N_2497,N_2327);
nor U2967 (N_2967,N_2220,N_2488);
xnor U2968 (N_2968,N_2312,N_2083);
or U2969 (N_2969,N_2254,N_2284);
or U2970 (N_2970,N_2494,N_2217);
nand U2971 (N_2971,N_2001,N_2467);
xor U2972 (N_2972,N_2103,N_2328);
and U2973 (N_2973,N_2382,N_2436);
or U2974 (N_2974,N_2186,N_2440);
xnor U2975 (N_2975,N_2476,N_2223);
nor U2976 (N_2976,N_2179,N_2199);
nand U2977 (N_2977,N_2413,N_2111);
nor U2978 (N_2978,N_2056,N_2354);
nand U2979 (N_2979,N_2496,N_2214);
xor U2980 (N_2980,N_2438,N_2333);
nor U2981 (N_2981,N_2210,N_2112);
nand U2982 (N_2982,N_2016,N_2324);
nand U2983 (N_2983,N_2002,N_2120);
xnor U2984 (N_2984,N_2178,N_2005);
xnor U2985 (N_2985,N_2190,N_2157);
xnor U2986 (N_2986,N_2037,N_2485);
or U2987 (N_2987,N_2474,N_2042);
nand U2988 (N_2988,N_2048,N_2284);
xnor U2989 (N_2989,N_2449,N_2498);
nand U2990 (N_2990,N_2410,N_2174);
nor U2991 (N_2991,N_2208,N_2251);
or U2992 (N_2992,N_2196,N_2107);
xnor U2993 (N_2993,N_2255,N_2366);
xor U2994 (N_2994,N_2060,N_2036);
or U2995 (N_2995,N_2405,N_2040);
nand U2996 (N_2996,N_2149,N_2203);
xor U2997 (N_2997,N_2402,N_2050);
xnor U2998 (N_2998,N_2446,N_2052);
or U2999 (N_2999,N_2032,N_2112);
xnor UO_0 (O_0,N_2571,N_2941);
nand UO_1 (O_1,N_2808,N_2956);
nand UO_2 (O_2,N_2987,N_2848);
or UO_3 (O_3,N_2612,N_2781);
or UO_4 (O_4,N_2677,N_2880);
or UO_5 (O_5,N_2702,N_2641);
xnor UO_6 (O_6,N_2748,N_2503);
and UO_7 (O_7,N_2632,N_2603);
nand UO_8 (O_8,N_2629,N_2901);
or UO_9 (O_9,N_2528,N_2943);
and UO_10 (O_10,N_2950,N_2546);
nor UO_11 (O_11,N_2580,N_2538);
or UO_12 (O_12,N_2593,N_2878);
nand UO_13 (O_13,N_2715,N_2533);
or UO_14 (O_14,N_2542,N_2611);
and UO_15 (O_15,N_2960,N_2930);
xnor UO_16 (O_16,N_2852,N_2825);
nor UO_17 (O_17,N_2635,N_2574);
nor UO_18 (O_18,N_2886,N_2917);
and UO_19 (O_19,N_2615,N_2722);
nand UO_20 (O_20,N_2934,N_2621);
nor UO_21 (O_21,N_2681,N_2671);
or UO_22 (O_22,N_2773,N_2753);
or UO_23 (O_23,N_2689,N_2623);
xnor UO_24 (O_24,N_2973,N_2797);
nand UO_25 (O_25,N_2839,N_2863);
and UO_26 (O_26,N_2714,N_2798);
nand UO_27 (O_27,N_2522,N_2962);
nor UO_28 (O_28,N_2888,N_2706);
xnor UO_29 (O_29,N_2816,N_2974);
nor UO_30 (O_30,N_2596,N_2764);
xnor UO_31 (O_31,N_2556,N_2657);
nor UO_32 (O_32,N_2918,N_2819);
and UO_33 (O_33,N_2573,N_2576);
or UO_34 (O_34,N_2840,N_2992);
xnor UO_35 (O_35,N_2949,N_2766);
nand UO_36 (O_36,N_2645,N_2659);
nand UO_37 (O_37,N_2982,N_2674);
nor UO_38 (O_38,N_2860,N_2907);
nor UO_39 (O_39,N_2958,N_2724);
and UO_40 (O_40,N_2953,N_2920);
xnor UO_41 (O_41,N_2905,N_2730);
or UO_42 (O_42,N_2544,N_2991);
nor UO_43 (O_43,N_2999,N_2820);
or UO_44 (O_44,N_2509,N_2775);
and UO_45 (O_45,N_2640,N_2590);
xor UO_46 (O_46,N_2661,N_2535);
and UO_47 (O_47,N_2900,N_2877);
and UO_48 (O_48,N_2527,N_2817);
nand UO_49 (O_49,N_2595,N_2912);
or UO_50 (O_50,N_2919,N_2647);
nand UO_51 (O_51,N_2608,N_2678);
nor UO_52 (O_52,N_2872,N_2989);
or UO_53 (O_53,N_2968,N_2957);
or UO_54 (O_54,N_2586,N_2606);
nor UO_55 (O_55,N_2772,N_2742);
xor UO_56 (O_56,N_2804,N_2909);
xnor UO_57 (O_57,N_2807,N_2857);
and UO_58 (O_58,N_2884,N_2510);
nor UO_59 (O_59,N_2827,N_2793);
nor UO_60 (O_60,N_2876,N_2910);
and UO_61 (O_61,N_2747,N_2837);
nand UO_62 (O_62,N_2897,N_2990);
or UO_63 (O_63,N_2966,N_2521);
nor UO_64 (O_64,N_2687,N_2662);
xnor UO_65 (O_65,N_2942,N_2630);
nand UO_66 (O_66,N_2740,N_2996);
and UO_67 (O_67,N_2902,N_2805);
nor UO_68 (O_68,N_2898,N_2847);
nor UO_69 (O_69,N_2868,N_2899);
and UO_70 (O_70,N_2708,N_2993);
nor UO_71 (O_71,N_2667,N_2988);
or UO_72 (O_72,N_2642,N_2757);
nand UO_73 (O_73,N_2655,N_2836);
and UO_74 (O_74,N_2695,N_2931);
or UO_75 (O_75,N_2646,N_2507);
or UO_76 (O_76,N_2944,N_2849);
xor UO_77 (O_77,N_2639,N_2703);
nand UO_78 (O_78,N_2532,N_2961);
xnor UO_79 (O_79,N_2833,N_2653);
xnor UO_80 (O_80,N_2799,N_2887);
or UO_81 (O_81,N_2965,N_2745);
nand UO_82 (O_82,N_2997,N_2758);
nor UO_83 (O_83,N_2566,N_2664);
nand UO_84 (O_84,N_2728,N_2822);
xor UO_85 (O_85,N_2505,N_2511);
or UO_86 (O_86,N_2523,N_2927);
or UO_87 (O_87,N_2624,N_2995);
nand UO_88 (O_88,N_2506,N_2756);
or UO_89 (O_89,N_2828,N_2769);
xnor UO_90 (O_90,N_2759,N_2738);
xor UO_91 (O_91,N_2540,N_2866);
and UO_92 (O_92,N_2952,N_2946);
nor UO_93 (O_93,N_2913,N_2776);
and UO_94 (O_94,N_2578,N_2679);
nand UO_95 (O_95,N_2971,N_2734);
and UO_96 (O_96,N_2795,N_2829);
nand UO_97 (O_97,N_2796,N_2543);
and UO_98 (O_98,N_2903,N_2508);
and UO_99 (O_99,N_2696,N_2592);
nor UO_100 (O_100,N_2788,N_2801);
nand UO_101 (O_101,N_2939,N_2552);
or UO_102 (O_102,N_2732,N_2550);
xnor UO_103 (O_103,N_2959,N_2626);
nand UO_104 (O_104,N_2534,N_2697);
nor UO_105 (O_105,N_2713,N_2587);
xnor UO_106 (O_106,N_2978,N_2834);
nand UO_107 (O_107,N_2693,N_2867);
nand UO_108 (O_108,N_2690,N_2760);
nand UO_109 (O_109,N_2806,N_2660);
nor UO_110 (O_110,N_2869,N_2892);
or UO_111 (O_111,N_2735,N_2707);
or UO_112 (O_112,N_2744,N_2894);
xnor UO_113 (O_113,N_2832,N_2783);
and UO_114 (O_114,N_2582,N_2864);
or UO_115 (O_115,N_2846,N_2743);
nand UO_116 (O_116,N_2810,N_2648);
xor UO_117 (O_117,N_2895,N_2780);
and UO_118 (O_118,N_2545,N_2779);
nor UO_119 (O_119,N_2812,N_2599);
and UO_120 (O_120,N_2739,N_2802);
nor UO_121 (O_121,N_2890,N_2865);
nand UO_122 (O_122,N_2964,N_2983);
xnor UO_123 (O_123,N_2975,N_2838);
nand UO_124 (O_124,N_2625,N_2613);
or UO_125 (O_125,N_2610,N_2637);
nand UO_126 (O_126,N_2710,N_2557);
xor UO_127 (O_127,N_2699,N_2826);
nand UO_128 (O_128,N_2994,N_2924);
or UO_129 (O_129,N_2518,N_2502);
nor UO_130 (O_130,N_2844,N_2786);
nor UO_131 (O_131,N_2565,N_2584);
nor UO_132 (O_132,N_2948,N_2685);
xor UO_133 (O_133,N_2906,N_2673);
and UO_134 (O_134,N_2561,N_2515);
nand UO_135 (O_135,N_2688,N_2570);
nand UO_136 (O_136,N_2784,N_2602);
and UO_137 (O_137,N_2785,N_2733);
or UO_138 (O_138,N_2512,N_2951);
or UO_139 (O_139,N_2843,N_2815);
nand UO_140 (O_140,N_2516,N_2851);
and UO_141 (O_141,N_2908,N_2789);
or UO_142 (O_142,N_2955,N_2666);
xnor UO_143 (O_143,N_2985,N_2691);
or UO_144 (O_144,N_2600,N_2861);
and UO_145 (O_145,N_2870,N_2601);
or UO_146 (O_146,N_2554,N_2762);
nor UO_147 (O_147,N_2519,N_2536);
nand UO_148 (O_148,N_2588,N_2854);
xor UO_149 (O_149,N_2676,N_2520);
nand UO_150 (O_150,N_2617,N_2682);
nor UO_151 (O_151,N_2850,N_2741);
or UO_152 (O_152,N_2716,N_2607);
and UO_153 (O_153,N_2879,N_2636);
nand UO_154 (O_154,N_2569,N_2976);
nand UO_155 (O_155,N_2628,N_2800);
nor UO_156 (O_156,N_2813,N_2932);
nand UO_157 (O_157,N_2853,N_2874);
and UO_158 (O_158,N_2729,N_2889);
and UO_159 (O_159,N_2531,N_2782);
nor UO_160 (O_160,N_2700,N_2774);
xor UO_161 (O_161,N_2814,N_2928);
or UO_162 (O_162,N_2591,N_2881);
nand UO_163 (O_163,N_2577,N_2616);
nor UO_164 (O_164,N_2692,N_2792);
xor UO_165 (O_165,N_2597,N_2891);
and UO_166 (O_166,N_2929,N_2559);
or UO_167 (O_167,N_2842,N_2787);
nor UO_168 (O_168,N_2720,N_2925);
nand UO_169 (O_169,N_2675,N_2719);
nand UO_170 (O_170,N_2529,N_2539);
nand UO_171 (O_171,N_2914,N_2513);
or UO_172 (O_172,N_2972,N_2922);
nand UO_173 (O_173,N_2604,N_2589);
and UO_174 (O_174,N_2885,N_2936);
nand UO_175 (O_175,N_2663,N_2524);
or UO_176 (O_176,N_2768,N_2575);
nand UO_177 (O_177,N_2649,N_2609);
or UO_178 (O_178,N_2711,N_2916);
nor UO_179 (O_179,N_2767,N_2670);
or UO_180 (O_180,N_2551,N_2858);
or UO_181 (O_181,N_2638,N_2594);
xor UO_182 (O_182,N_2709,N_2835);
or UO_183 (O_183,N_2755,N_2749);
nand UO_184 (O_184,N_2500,N_2771);
nand UO_185 (O_185,N_2618,N_2633);
nor UO_186 (O_186,N_2643,N_2859);
xor UO_187 (O_187,N_2530,N_2751);
nor UO_188 (O_188,N_2970,N_2684);
and UO_189 (O_189,N_2627,N_2548);
or UO_190 (O_190,N_2809,N_2778);
or UO_191 (O_191,N_2504,N_2514);
nand UO_192 (O_192,N_2911,N_2963);
xor UO_193 (O_193,N_2614,N_2721);
nand UO_194 (O_194,N_2672,N_2979);
nor UO_195 (O_195,N_2821,N_2526);
xor UO_196 (O_196,N_2765,N_2754);
xnor UO_197 (O_197,N_2652,N_2893);
and UO_198 (O_198,N_2537,N_2830);
nor UO_199 (O_199,N_2777,N_2977);
or UO_200 (O_200,N_2701,N_2723);
xor UO_201 (O_201,N_2935,N_2954);
nor UO_202 (O_202,N_2680,N_2605);
or UO_203 (O_203,N_2572,N_2882);
or UO_204 (O_204,N_2694,N_2704);
and UO_205 (O_205,N_2705,N_2558);
xnor UO_206 (O_206,N_2717,N_2945);
and UO_207 (O_207,N_2585,N_2669);
nand UO_208 (O_208,N_2871,N_2501);
nor UO_209 (O_209,N_2750,N_2541);
or UO_210 (O_210,N_2581,N_2598);
xor UO_211 (O_211,N_2547,N_2818);
or UO_212 (O_212,N_2725,N_2790);
nand UO_213 (O_213,N_2856,N_2658);
xor UO_214 (O_214,N_2650,N_2824);
xnor UO_215 (O_215,N_2583,N_2763);
nor UO_216 (O_216,N_2634,N_2980);
nor UO_217 (O_217,N_2947,N_2967);
xor UO_218 (O_218,N_2875,N_2926);
xnor UO_219 (O_219,N_2746,N_2940);
xor UO_220 (O_220,N_2712,N_2620);
nor UO_221 (O_221,N_2563,N_2644);
xnor UO_222 (O_222,N_2718,N_2794);
and UO_223 (O_223,N_2915,N_2845);
or UO_224 (O_224,N_2862,N_2567);
nor UO_225 (O_225,N_2654,N_2752);
or UO_226 (O_226,N_2568,N_2938);
nor UO_227 (O_227,N_2562,N_2668);
or UO_228 (O_228,N_2726,N_2549);
or UO_229 (O_229,N_2727,N_2698);
or UO_230 (O_230,N_2656,N_2761);
nand UO_231 (O_231,N_2933,N_2896);
and UO_232 (O_232,N_2553,N_2921);
and UO_233 (O_233,N_2683,N_2731);
nor UO_234 (O_234,N_2736,N_2811);
or UO_235 (O_235,N_2803,N_2998);
xnor UO_236 (O_236,N_2791,N_2841);
and UO_237 (O_237,N_2665,N_2823);
xnor UO_238 (O_238,N_2686,N_2981);
and UO_239 (O_239,N_2923,N_2560);
xnor UO_240 (O_240,N_2579,N_2969);
xnor UO_241 (O_241,N_2855,N_2622);
or UO_242 (O_242,N_2619,N_2651);
and UO_243 (O_243,N_2770,N_2883);
nand UO_244 (O_244,N_2631,N_2517);
nand UO_245 (O_245,N_2984,N_2831);
nand UO_246 (O_246,N_2525,N_2737);
and UO_247 (O_247,N_2555,N_2873);
nand UO_248 (O_248,N_2986,N_2904);
or UO_249 (O_249,N_2564,N_2937);
or UO_250 (O_250,N_2651,N_2895);
xnor UO_251 (O_251,N_2788,N_2668);
nor UO_252 (O_252,N_2907,N_2715);
xor UO_253 (O_253,N_2516,N_2899);
xnor UO_254 (O_254,N_2837,N_2771);
nand UO_255 (O_255,N_2951,N_2996);
or UO_256 (O_256,N_2883,N_2986);
and UO_257 (O_257,N_2740,N_2655);
nand UO_258 (O_258,N_2610,N_2530);
and UO_259 (O_259,N_2706,N_2581);
or UO_260 (O_260,N_2760,N_2695);
and UO_261 (O_261,N_2777,N_2623);
and UO_262 (O_262,N_2860,N_2975);
and UO_263 (O_263,N_2896,N_2978);
xor UO_264 (O_264,N_2853,N_2532);
nand UO_265 (O_265,N_2814,N_2958);
xor UO_266 (O_266,N_2664,N_2676);
nand UO_267 (O_267,N_2949,N_2993);
nand UO_268 (O_268,N_2875,N_2902);
nand UO_269 (O_269,N_2941,N_2778);
nand UO_270 (O_270,N_2598,N_2509);
nand UO_271 (O_271,N_2971,N_2832);
xnor UO_272 (O_272,N_2713,N_2622);
and UO_273 (O_273,N_2599,N_2677);
nor UO_274 (O_274,N_2668,N_2589);
and UO_275 (O_275,N_2915,N_2636);
and UO_276 (O_276,N_2914,N_2531);
or UO_277 (O_277,N_2841,N_2667);
or UO_278 (O_278,N_2547,N_2659);
xor UO_279 (O_279,N_2585,N_2985);
nor UO_280 (O_280,N_2556,N_2529);
or UO_281 (O_281,N_2667,N_2932);
nor UO_282 (O_282,N_2911,N_2679);
xor UO_283 (O_283,N_2746,N_2749);
nor UO_284 (O_284,N_2797,N_2977);
nor UO_285 (O_285,N_2755,N_2502);
xnor UO_286 (O_286,N_2580,N_2998);
xnor UO_287 (O_287,N_2884,N_2772);
nand UO_288 (O_288,N_2769,N_2714);
nor UO_289 (O_289,N_2864,N_2777);
xor UO_290 (O_290,N_2779,N_2625);
and UO_291 (O_291,N_2983,N_2535);
and UO_292 (O_292,N_2980,N_2646);
or UO_293 (O_293,N_2779,N_2596);
nor UO_294 (O_294,N_2916,N_2990);
or UO_295 (O_295,N_2547,N_2570);
and UO_296 (O_296,N_2550,N_2697);
nor UO_297 (O_297,N_2990,N_2996);
nand UO_298 (O_298,N_2528,N_2969);
and UO_299 (O_299,N_2771,N_2990);
or UO_300 (O_300,N_2641,N_2865);
and UO_301 (O_301,N_2894,N_2520);
or UO_302 (O_302,N_2775,N_2899);
xnor UO_303 (O_303,N_2502,N_2686);
nand UO_304 (O_304,N_2714,N_2607);
xor UO_305 (O_305,N_2816,N_2500);
xnor UO_306 (O_306,N_2556,N_2786);
nand UO_307 (O_307,N_2964,N_2515);
nand UO_308 (O_308,N_2760,N_2858);
nand UO_309 (O_309,N_2734,N_2892);
xnor UO_310 (O_310,N_2712,N_2682);
and UO_311 (O_311,N_2706,N_2950);
or UO_312 (O_312,N_2712,N_2995);
nor UO_313 (O_313,N_2864,N_2595);
and UO_314 (O_314,N_2627,N_2936);
xor UO_315 (O_315,N_2947,N_2507);
nor UO_316 (O_316,N_2764,N_2802);
xnor UO_317 (O_317,N_2555,N_2532);
xor UO_318 (O_318,N_2812,N_2661);
nor UO_319 (O_319,N_2613,N_2745);
xnor UO_320 (O_320,N_2931,N_2807);
and UO_321 (O_321,N_2636,N_2965);
or UO_322 (O_322,N_2660,N_2666);
or UO_323 (O_323,N_2505,N_2812);
or UO_324 (O_324,N_2851,N_2928);
or UO_325 (O_325,N_2949,N_2733);
nor UO_326 (O_326,N_2591,N_2965);
or UO_327 (O_327,N_2930,N_2730);
xor UO_328 (O_328,N_2592,N_2587);
and UO_329 (O_329,N_2802,N_2533);
and UO_330 (O_330,N_2994,N_2669);
nor UO_331 (O_331,N_2622,N_2536);
nand UO_332 (O_332,N_2657,N_2817);
or UO_333 (O_333,N_2563,N_2846);
nor UO_334 (O_334,N_2765,N_2724);
and UO_335 (O_335,N_2834,N_2790);
and UO_336 (O_336,N_2768,N_2523);
nand UO_337 (O_337,N_2569,N_2793);
xnor UO_338 (O_338,N_2603,N_2961);
nor UO_339 (O_339,N_2684,N_2515);
nor UO_340 (O_340,N_2503,N_2707);
and UO_341 (O_341,N_2883,N_2697);
nand UO_342 (O_342,N_2891,N_2561);
or UO_343 (O_343,N_2892,N_2911);
nand UO_344 (O_344,N_2585,N_2889);
and UO_345 (O_345,N_2830,N_2687);
xnor UO_346 (O_346,N_2508,N_2651);
or UO_347 (O_347,N_2864,N_2928);
nor UO_348 (O_348,N_2915,N_2750);
or UO_349 (O_349,N_2691,N_2800);
nand UO_350 (O_350,N_2678,N_2799);
xnor UO_351 (O_351,N_2617,N_2616);
xnor UO_352 (O_352,N_2832,N_2919);
xor UO_353 (O_353,N_2843,N_2747);
nand UO_354 (O_354,N_2977,N_2612);
or UO_355 (O_355,N_2560,N_2808);
and UO_356 (O_356,N_2656,N_2774);
xnor UO_357 (O_357,N_2546,N_2918);
xor UO_358 (O_358,N_2888,N_2609);
nand UO_359 (O_359,N_2669,N_2817);
nand UO_360 (O_360,N_2518,N_2565);
nand UO_361 (O_361,N_2745,N_2807);
and UO_362 (O_362,N_2917,N_2820);
nand UO_363 (O_363,N_2640,N_2618);
nand UO_364 (O_364,N_2673,N_2799);
xnor UO_365 (O_365,N_2728,N_2560);
nand UO_366 (O_366,N_2545,N_2564);
and UO_367 (O_367,N_2648,N_2884);
xnor UO_368 (O_368,N_2501,N_2993);
nor UO_369 (O_369,N_2806,N_2690);
nand UO_370 (O_370,N_2966,N_2601);
and UO_371 (O_371,N_2809,N_2661);
and UO_372 (O_372,N_2887,N_2871);
nor UO_373 (O_373,N_2603,N_2709);
xor UO_374 (O_374,N_2936,N_2584);
xnor UO_375 (O_375,N_2715,N_2564);
and UO_376 (O_376,N_2691,N_2892);
nor UO_377 (O_377,N_2901,N_2772);
nor UO_378 (O_378,N_2912,N_2702);
nand UO_379 (O_379,N_2580,N_2791);
nand UO_380 (O_380,N_2568,N_2571);
nor UO_381 (O_381,N_2937,N_2630);
or UO_382 (O_382,N_2818,N_2670);
and UO_383 (O_383,N_2885,N_2703);
xor UO_384 (O_384,N_2732,N_2710);
nand UO_385 (O_385,N_2980,N_2693);
nand UO_386 (O_386,N_2516,N_2636);
and UO_387 (O_387,N_2653,N_2575);
nor UO_388 (O_388,N_2506,N_2902);
xor UO_389 (O_389,N_2685,N_2619);
nor UO_390 (O_390,N_2936,N_2769);
nand UO_391 (O_391,N_2508,N_2691);
and UO_392 (O_392,N_2990,N_2674);
and UO_393 (O_393,N_2696,N_2731);
and UO_394 (O_394,N_2546,N_2851);
nor UO_395 (O_395,N_2987,N_2916);
and UO_396 (O_396,N_2701,N_2761);
nor UO_397 (O_397,N_2726,N_2637);
nand UO_398 (O_398,N_2660,N_2781);
nor UO_399 (O_399,N_2942,N_2673);
and UO_400 (O_400,N_2650,N_2955);
and UO_401 (O_401,N_2684,N_2619);
or UO_402 (O_402,N_2841,N_2952);
or UO_403 (O_403,N_2799,N_2841);
nand UO_404 (O_404,N_2778,N_2885);
and UO_405 (O_405,N_2641,N_2577);
xor UO_406 (O_406,N_2511,N_2622);
or UO_407 (O_407,N_2737,N_2676);
or UO_408 (O_408,N_2719,N_2603);
xor UO_409 (O_409,N_2695,N_2852);
nand UO_410 (O_410,N_2687,N_2916);
nand UO_411 (O_411,N_2759,N_2925);
or UO_412 (O_412,N_2850,N_2631);
or UO_413 (O_413,N_2989,N_2564);
xnor UO_414 (O_414,N_2753,N_2504);
nand UO_415 (O_415,N_2832,N_2809);
nor UO_416 (O_416,N_2923,N_2604);
or UO_417 (O_417,N_2505,N_2926);
or UO_418 (O_418,N_2506,N_2719);
nand UO_419 (O_419,N_2877,N_2871);
and UO_420 (O_420,N_2634,N_2760);
or UO_421 (O_421,N_2814,N_2675);
nor UO_422 (O_422,N_2768,N_2678);
and UO_423 (O_423,N_2924,N_2755);
nor UO_424 (O_424,N_2664,N_2887);
or UO_425 (O_425,N_2756,N_2791);
nor UO_426 (O_426,N_2521,N_2964);
nand UO_427 (O_427,N_2816,N_2758);
or UO_428 (O_428,N_2897,N_2579);
nand UO_429 (O_429,N_2897,N_2831);
xnor UO_430 (O_430,N_2739,N_2765);
nand UO_431 (O_431,N_2948,N_2951);
nand UO_432 (O_432,N_2931,N_2512);
or UO_433 (O_433,N_2646,N_2880);
nor UO_434 (O_434,N_2966,N_2649);
xnor UO_435 (O_435,N_2755,N_2568);
or UO_436 (O_436,N_2783,N_2668);
nand UO_437 (O_437,N_2610,N_2841);
and UO_438 (O_438,N_2586,N_2663);
xnor UO_439 (O_439,N_2540,N_2801);
or UO_440 (O_440,N_2801,N_2933);
nor UO_441 (O_441,N_2823,N_2931);
nand UO_442 (O_442,N_2710,N_2636);
nand UO_443 (O_443,N_2621,N_2874);
or UO_444 (O_444,N_2676,N_2701);
and UO_445 (O_445,N_2870,N_2903);
nor UO_446 (O_446,N_2580,N_2872);
xor UO_447 (O_447,N_2797,N_2867);
or UO_448 (O_448,N_2962,N_2910);
nor UO_449 (O_449,N_2850,N_2810);
xor UO_450 (O_450,N_2525,N_2540);
or UO_451 (O_451,N_2859,N_2852);
or UO_452 (O_452,N_2864,N_2753);
nand UO_453 (O_453,N_2997,N_2692);
and UO_454 (O_454,N_2542,N_2664);
and UO_455 (O_455,N_2657,N_2875);
or UO_456 (O_456,N_2595,N_2814);
xnor UO_457 (O_457,N_2503,N_2829);
nand UO_458 (O_458,N_2531,N_2862);
xnor UO_459 (O_459,N_2970,N_2539);
or UO_460 (O_460,N_2677,N_2979);
xor UO_461 (O_461,N_2771,N_2972);
or UO_462 (O_462,N_2921,N_2606);
nand UO_463 (O_463,N_2700,N_2910);
nand UO_464 (O_464,N_2927,N_2519);
xnor UO_465 (O_465,N_2761,N_2990);
or UO_466 (O_466,N_2911,N_2974);
nand UO_467 (O_467,N_2535,N_2749);
nand UO_468 (O_468,N_2554,N_2520);
nand UO_469 (O_469,N_2988,N_2897);
xor UO_470 (O_470,N_2793,N_2849);
or UO_471 (O_471,N_2987,N_2998);
nor UO_472 (O_472,N_2561,N_2974);
nor UO_473 (O_473,N_2545,N_2855);
nor UO_474 (O_474,N_2512,N_2694);
nor UO_475 (O_475,N_2757,N_2796);
nor UO_476 (O_476,N_2914,N_2959);
or UO_477 (O_477,N_2500,N_2729);
and UO_478 (O_478,N_2905,N_2832);
and UO_479 (O_479,N_2906,N_2694);
or UO_480 (O_480,N_2831,N_2739);
and UO_481 (O_481,N_2874,N_2842);
xnor UO_482 (O_482,N_2516,N_2874);
and UO_483 (O_483,N_2522,N_2604);
nor UO_484 (O_484,N_2521,N_2806);
nand UO_485 (O_485,N_2739,N_2572);
xnor UO_486 (O_486,N_2821,N_2802);
nand UO_487 (O_487,N_2765,N_2945);
and UO_488 (O_488,N_2602,N_2978);
and UO_489 (O_489,N_2801,N_2893);
and UO_490 (O_490,N_2549,N_2782);
nand UO_491 (O_491,N_2887,N_2897);
xor UO_492 (O_492,N_2996,N_2947);
and UO_493 (O_493,N_2819,N_2782);
xor UO_494 (O_494,N_2704,N_2862);
xnor UO_495 (O_495,N_2791,N_2721);
nand UO_496 (O_496,N_2761,N_2535);
or UO_497 (O_497,N_2950,N_2812);
nand UO_498 (O_498,N_2807,N_2645);
or UO_499 (O_499,N_2962,N_2977);
endmodule