module basic_1500_15000_2000_10_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_576,In_1155);
nor U1 (N_1,In_1371,In_45);
or U2 (N_2,In_784,In_1356);
or U3 (N_3,In_435,In_719);
and U4 (N_4,In_13,In_197);
and U5 (N_5,In_668,In_1361);
and U6 (N_6,In_1306,In_375);
nand U7 (N_7,In_1319,In_786);
or U8 (N_8,In_564,In_1307);
nand U9 (N_9,In_123,In_693);
xnor U10 (N_10,In_762,In_1421);
nand U11 (N_11,In_571,In_5);
and U12 (N_12,In_1200,In_236);
and U13 (N_13,In_1106,In_569);
or U14 (N_14,In_900,In_678);
or U15 (N_15,In_366,In_956);
nor U16 (N_16,In_912,In_163);
nor U17 (N_17,In_526,In_121);
or U18 (N_18,In_1495,In_1491);
nor U19 (N_19,In_766,In_1157);
or U20 (N_20,In_1303,In_771);
or U21 (N_21,In_239,In_403);
or U22 (N_22,In_559,In_1402);
and U23 (N_23,In_1261,In_889);
xor U24 (N_24,In_1073,In_640);
nand U25 (N_25,In_1055,In_1005);
and U26 (N_26,In_846,In_83);
or U27 (N_27,In_814,In_1426);
and U28 (N_28,In_294,In_1052);
nand U29 (N_29,In_189,In_824);
and U30 (N_30,In_1084,In_918);
or U31 (N_31,In_481,In_544);
nand U32 (N_32,In_15,In_679);
nand U33 (N_33,In_1116,In_922);
nor U34 (N_34,In_1412,In_1375);
or U35 (N_35,In_1445,In_408);
and U36 (N_36,In_517,In_1080);
and U37 (N_37,In_1478,In_1203);
or U38 (N_38,In_734,In_175);
nor U39 (N_39,In_82,In_399);
nand U40 (N_40,In_348,In_1082);
and U41 (N_41,In_880,In_166);
nand U42 (N_42,In_835,In_1069);
and U43 (N_43,In_165,In_192);
nor U44 (N_44,In_367,In_1204);
nand U45 (N_45,In_258,In_606);
nor U46 (N_46,In_184,In_518);
nor U47 (N_47,In_568,In_1345);
nand U48 (N_48,In_352,In_478);
and U49 (N_49,In_952,In_1031);
nor U50 (N_50,In_924,In_154);
nor U51 (N_51,In_174,In_864);
and U52 (N_52,In_675,In_479);
nor U53 (N_53,In_574,In_1413);
or U54 (N_54,In_217,In_190);
or U55 (N_55,In_622,In_1420);
or U56 (N_56,In_1459,In_556);
nand U57 (N_57,In_1035,In_1085);
and U58 (N_58,In_809,In_428);
and U59 (N_59,In_510,In_904);
nor U60 (N_60,In_291,In_1047);
nor U61 (N_61,In_1440,In_595);
nand U62 (N_62,In_508,In_681);
and U63 (N_63,In_1399,In_1387);
nand U64 (N_64,In_703,In_859);
or U65 (N_65,In_1074,In_832);
or U66 (N_66,In_1453,In_725);
or U67 (N_67,In_292,In_474);
or U68 (N_68,In_583,In_851);
and U69 (N_69,In_277,In_872);
and U70 (N_70,In_630,In_1062);
nand U71 (N_71,In_1451,In_42);
nand U72 (N_72,In_1024,In_1271);
nand U73 (N_73,In_460,In_818);
or U74 (N_74,In_1262,In_759);
nor U75 (N_75,In_1151,In_1000);
nor U76 (N_76,In_999,In_127);
nor U77 (N_77,In_1170,In_1314);
or U78 (N_78,In_393,In_747);
nor U79 (N_79,In_1336,In_834);
or U80 (N_80,In_370,In_271);
and U81 (N_81,In_505,In_930);
nand U82 (N_82,In_99,In_682);
or U83 (N_83,In_967,In_1334);
and U84 (N_84,In_577,In_372);
nand U85 (N_85,In_785,In_749);
nor U86 (N_86,In_635,In_187);
or U87 (N_87,In_157,In_1229);
and U88 (N_88,In_1343,In_492);
or U89 (N_89,In_1161,In_37);
nor U90 (N_90,In_1175,In_712);
or U91 (N_91,In_1312,In_171);
and U92 (N_92,In_1480,In_513);
or U93 (N_93,In_1075,In_17);
nor U94 (N_94,In_1471,In_426);
xnor U95 (N_95,In_642,In_1446);
or U96 (N_96,In_242,In_1246);
and U97 (N_97,In_1169,In_246);
nand U98 (N_98,In_204,In_928);
xor U99 (N_99,In_425,In_404);
nor U100 (N_100,In_1077,In_585);
or U101 (N_101,In_73,In_301);
nor U102 (N_102,In_1444,In_400);
and U103 (N_103,In_887,In_1023);
and U104 (N_104,In_3,In_50);
nor U105 (N_105,In_799,In_688);
and U106 (N_106,In_983,In_262);
nand U107 (N_107,In_782,In_1452);
nand U108 (N_108,In_112,In_368);
and U109 (N_109,In_386,In_883);
nor U110 (N_110,In_516,In_1027);
or U111 (N_111,In_917,In_103);
nand U112 (N_112,In_676,In_627);
or U113 (N_113,In_1164,In_772);
nor U114 (N_114,In_1273,In_1252);
nand U115 (N_115,In_414,In_1342);
and U116 (N_116,In_283,In_274);
and U117 (N_117,In_1003,In_950);
and U118 (N_118,In_1096,In_421);
and U119 (N_119,In_495,In_915);
or U120 (N_120,In_153,In_760);
nand U121 (N_121,In_134,In_1283);
nor U122 (N_122,In_427,In_298);
nor U123 (N_123,In_836,In_1379);
nor U124 (N_124,In_80,In_1294);
nor U125 (N_125,In_24,In_971);
and U126 (N_126,In_1267,In_973);
or U127 (N_127,In_162,In_390);
xnor U128 (N_128,In_1322,In_245);
nor U129 (N_129,In_664,In_1469);
nand U130 (N_130,In_145,In_355);
nor U131 (N_131,In_1441,In_490);
and U132 (N_132,In_588,In_1220);
and U133 (N_133,In_139,In_51);
nand U134 (N_134,In_763,In_1070);
or U135 (N_135,In_483,In_1184);
nor U136 (N_136,In_1234,In_43);
or U137 (N_137,In_1275,In_238);
or U138 (N_138,In_838,In_1227);
nand U139 (N_139,In_954,In_700);
nand U140 (N_140,In_927,In_106);
nand U141 (N_141,In_1217,In_921);
nor U142 (N_142,In_152,In_1428);
and U143 (N_143,In_605,In_618);
or U144 (N_144,In_506,In_385);
xor U145 (N_145,In_394,In_970);
nor U146 (N_146,In_1274,In_519);
and U147 (N_147,In_614,In_228);
or U148 (N_148,In_1192,In_58);
nand U149 (N_149,In_199,In_79);
nand U150 (N_150,In_198,In_111);
nand U151 (N_151,In_1408,In_338);
nand U152 (N_152,In_995,In_940);
nor U153 (N_153,In_1373,In_302);
and U154 (N_154,In_631,In_966);
nand U155 (N_155,In_1468,In_1245);
and U156 (N_156,In_667,In_336);
and U157 (N_157,In_767,In_1207);
nor U158 (N_158,In_164,In_1160);
nand U159 (N_159,In_11,In_133);
nor U160 (N_160,In_801,In_235);
nand U161 (N_161,In_487,In_329);
or U162 (N_162,In_1310,In_739);
nor U163 (N_163,In_1357,In_934);
nor U164 (N_164,In_1429,In_469);
or U165 (N_165,In_176,In_829);
nor U166 (N_166,In_1110,In_105);
and U167 (N_167,In_444,In_641);
and U168 (N_168,In_376,In_1393);
or U169 (N_169,In_412,In_1410);
nor U170 (N_170,In_436,In_1038);
nor U171 (N_171,In_1060,In_828);
nand U172 (N_172,In_1390,In_695);
nor U173 (N_173,In_268,In_991);
nand U174 (N_174,In_1012,In_669);
and U175 (N_175,In_533,In_363);
nor U176 (N_176,In_318,In_473);
nand U177 (N_177,In_1297,In_1434);
nor U178 (N_178,In_852,In_1368);
or U179 (N_179,In_1071,In_1409);
and U180 (N_180,In_1079,In_503);
or U181 (N_181,In_951,In_567);
xor U182 (N_182,In_706,In_259);
and U183 (N_183,In_827,In_1406);
or U184 (N_184,In_735,In_196);
and U185 (N_185,In_587,In_126);
nor U186 (N_186,In_1340,In_1465);
nor U187 (N_187,In_1320,In_59);
nand U188 (N_188,In_1285,In_430);
nand U189 (N_189,In_645,In_148);
nand U190 (N_190,In_989,In_1225);
and U191 (N_191,In_781,In_415);
xnor U192 (N_192,In_1094,In_774);
xor U193 (N_193,In_990,In_18);
nor U194 (N_194,In_1033,In_497);
nand U195 (N_195,In_876,In_1330);
nor U196 (N_196,In_1332,In_1432);
nand U197 (N_197,In_694,In_1442);
nor U198 (N_198,In_1001,In_109);
or U199 (N_199,In_457,In_334);
nor U200 (N_200,In_69,In_216);
or U201 (N_201,In_1091,In_434);
and U202 (N_202,In_488,In_1448);
nand U203 (N_203,In_1455,In_705);
nand U204 (N_204,In_750,In_1111);
nand U205 (N_205,In_1467,In_888);
or U206 (N_206,In_1221,In_874);
and U207 (N_207,In_1017,In_1014);
nor U208 (N_208,In_1250,In_396);
and U209 (N_209,In_29,In_795);
nor U210 (N_210,In_1190,In_773);
nand U211 (N_211,In_1403,In_644);
and U212 (N_212,In_293,In_683);
nor U213 (N_213,In_100,In_916);
nand U214 (N_214,In_466,In_72);
and U215 (N_215,In_458,In_448);
nor U216 (N_216,In_233,In_1232);
nand U217 (N_217,In_1078,In_674);
or U218 (N_218,In_1366,In_344);
nor U219 (N_219,In_498,In_961);
and U220 (N_220,In_551,In_57);
and U221 (N_221,In_450,In_637);
nand U222 (N_222,In_440,In_114);
nor U223 (N_223,In_264,In_282);
or U224 (N_224,In_1456,In_628);
or U225 (N_225,In_493,In_1264);
and U226 (N_226,In_267,In_21);
nand U227 (N_227,In_737,In_462);
nor U228 (N_228,In_169,In_1066);
nand U229 (N_229,In_191,In_288);
xnor U230 (N_230,In_1235,In_1427);
or U231 (N_231,In_295,In_306);
and U232 (N_232,In_1166,In_33);
nand U233 (N_233,In_793,In_512);
nand U234 (N_234,In_1417,In_905);
or U235 (N_235,In_1329,In_1394);
or U236 (N_236,In_252,In_132);
nand U237 (N_237,In_477,In_756);
nand U238 (N_238,In_1479,In_1327);
nand U239 (N_239,In_721,In_636);
and U240 (N_240,In_1051,In_1211);
and U241 (N_241,In_63,In_1386);
and U242 (N_242,In_1112,In_1381);
and U243 (N_243,In_1049,In_580);
nor U244 (N_244,In_619,In_54);
nor U245 (N_245,In_261,In_1253);
and U246 (N_246,In_1133,In_974);
nor U247 (N_247,In_672,In_729);
nand U248 (N_248,In_1022,In_979);
xnor U249 (N_249,In_1212,In_557);
and U250 (N_250,In_1109,In_770);
nor U251 (N_251,In_514,In_34);
and U252 (N_252,In_545,In_1020);
nand U253 (N_253,In_279,In_1202);
nor U254 (N_254,In_1376,In_323);
nor U255 (N_255,In_964,In_208);
and U256 (N_256,In_155,In_1400);
nor U257 (N_257,In_877,In_1067);
nor U258 (N_258,In_920,In_1256);
nand U259 (N_259,In_933,In_555);
and U260 (N_260,In_243,In_1362);
nand U261 (N_261,In_1280,In_908);
nor U262 (N_262,In_1475,In_798);
and U263 (N_263,In_1325,In_167);
and U264 (N_264,In_406,In_603);
or U265 (N_265,In_1099,In_1279);
or U266 (N_266,In_647,In_303);
and U267 (N_267,In_407,In_1162);
nand U268 (N_268,In_733,In_161);
or U269 (N_269,In_496,In_596);
nor U270 (N_270,In_1378,In_875);
and U271 (N_271,In_1257,In_1107);
or U272 (N_272,In_23,In_232);
nand U273 (N_273,In_840,In_313);
nor U274 (N_274,In_981,In_881);
and U275 (N_275,In_945,In_178);
nor U276 (N_276,In_351,In_590);
and U277 (N_277,In_953,In_270);
or U278 (N_278,In_468,In_1411);
and U279 (N_279,In_982,In_1087);
nand U280 (N_280,In_311,In_125);
and U281 (N_281,In_692,In_1143);
nor U282 (N_282,In_998,In_276);
nand U283 (N_283,In_1176,In_1258);
nor U284 (N_284,In_224,In_857);
nor U285 (N_285,In_1130,In_620);
nand U286 (N_286,In_796,In_377);
nor U287 (N_287,In_753,In_312);
or U288 (N_288,In_1344,In_1337);
or U289 (N_289,In_854,In_955);
or U290 (N_290,In_1072,In_752);
and U291 (N_291,In_1487,In_858);
or U292 (N_292,In_8,In_1183);
and U293 (N_293,In_269,In_459);
or U294 (N_294,In_776,In_1187);
and U295 (N_295,In_214,In_49);
nor U296 (N_296,In_790,In_783);
nor U297 (N_297,In_1260,In_609);
or U298 (N_298,In_87,In_661);
or U299 (N_299,In_994,In_53);
and U300 (N_300,In_823,In_1147);
or U301 (N_301,In_443,In_1058);
nor U302 (N_302,In_1097,In_1119);
or U303 (N_303,In_1450,In_968);
or U304 (N_304,In_621,In_1174);
and U305 (N_305,In_1150,In_527);
nor U306 (N_306,In_1168,In_398);
and U307 (N_307,In_855,In_128);
or U308 (N_308,In_464,In_543);
or U309 (N_309,In_816,In_1124);
or U310 (N_310,In_1497,In_599);
or U311 (N_311,In_1259,In_831);
xor U312 (N_312,In_986,In_213);
nor U313 (N_313,In_1457,In_227);
and U314 (N_314,In_379,In_1438);
and U315 (N_315,In_101,In_1237);
and U316 (N_316,In_1064,In_1392);
nand U317 (N_317,In_751,In_1136);
or U318 (N_318,In_1142,In_931);
nand U319 (N_319,In_454,In_135);
or U320 (N_320,In_575,In_93);
nand U321 (N_321,In_1238,In_249);
nor U322 (N_322,In_563,In_476);
nor U323 (N_323,In_108,In_1300);
or U324 (N_324,In_1348,In_720);
and U325 (N_325,In_1145,In_1333);
nand U326 (N_326,In_489,In_1193);
or U327 (N_327,In_780,In_320);
or U328 (N_328,In_594,In_1132);
nor U329 (N_329,In_328,In_14);
nor U330 (N_330,In_1236,In_451);
nand U331 (N_331,In_122,In_309);
or U332 (N_332,In_1419,In_652);
or U333 (N_333,In_251,In_470);
nand U334 (N_334,In_707,In_1430);
and U335 (N_335,In_46,In_708);
and U336 (N_336,In_442,In_1036);
or U337 (N_337,In_1401,In_12);
or U338 (N_338,In_405,In_1199);
and U339 (N_339,In_422,In_119);
nor U340 (N_340,In_511,In_1443);
nor U341 (N_341,In_388,In_1324);
nor U342 (N_342,In_485,In_715);
nor U343 (N_343,In_237,In_947);
and U344 (N_344,In_537,In_826);
nor U345 (N_345,In_849,In_680);
or U346 (N_346,In_1268,In_345);
nand U347 (N_347,In_1377,In_260);
nand U348 (N_348,In_491,In_949);
nand U349 (N_349,In_1290,In_718);
and U350 (N_350,In_391,In_1040);
nand U351 (N_351,In_1063,In_1269);
nor U352 (N_352,In_1293,In_1189);
and U353 (N_353,In_1156,In_20);
nand U354 (N_354,In_361,In_1359);
nand U355 (N_355,In_102,In_322);
or U356 (N_356,In_1102,In_1369);
nor U357 (N_357,In_978,In_44);
nor U358 (N_358,In_1315,In_1182);
or U359 (N_359,In_528,In_1414);
or U360 (N_360,In_1382,In_717);
nand U361 (N_361,In_1194,In_1418);
and U362 (N_362,In_183,In_253);
nor U363 (N_363,In_446,In_653);
or U364 (N_364,In_140,In_1205);
and U365 (N_365,In_327,In_1115);
or U366 (N_366,In_1154,In_633);
nor U367 (N_367,In_130,In_1464);
and U368 (N_368,In_47,In_634);
nor U369 (N_369,In_297,In_35);
and U370 (N_370,In_1365,In_467);
nand U371 (N_371,In_75,In_755);
nor U372 (N_372,In_1372,In_1435);
nor U373 (N_373,In_92,In_1311);
and U374 (N_374,In_55,In_873);
nor U375 (N_375,In_359,In_1278);
nand U376 (N_376,In_156,In_602);
or U377 (N_377,In_1149,In_1);
or U378 (N_378,In_330,In_263);
nand U379 (N_379,In_1172,In_48);
and U380 (N_380,In_378,In_1191);
nand U381 (N_381,In_1088,In_1331);
nor U382 (N_382,In_1181,In_980);
and U383 (N_383,In_1163,In_494);
nand U384 (N_384,In_1493,In_4);
and U385 (N_385,In_608,In_910);
and U386 (N_386,In_757,In_819);
nand U387 (N_387,In_1423,In_461);
xnor U388 (N_388,In_315,In_64);
nand U389 (N_389,In_1231,In_244);
or U390 (N_390,In_1249,In_1032);
and U391 (N_391,In_1349,In_202);
nand U392 (N_392,In_1186,In_808);
or U393 (N_393,In_9,In_870);
or U394 (N_394,In_429,In_646);
nand U395 (N_395,In_66,In_151);
or U396 (N_396,In_656,In_825);
nor U397 (N_397,In_552,In_898);
nand U398 (N_398,In_222,In_671);
nor U399 (N_399,In_1265,In_229);
nand U400 (N_400,In_539,In_833);
nor U401 (N_401,In_565,In_1422);
or U402 (N_402,In_206,In_914);
and U403 (N_403,In_1206,In_1059);
nand U404 (N_404,In_16,In_195);
nand U405 (N_405,In_331,In_340);
nor U406 (N_406,In_534,In_413);
nand U407 (N_407,In_901,In_365);
nand U408 (N_408,In_1137,In_182);
xnor U409 (N_409,In_765,In_472);
or U410 (N_410,In_515,In_943);
or U411 (N_411,In_1057,In_579);
and U412 (N_412,In_884,In_598);
xor U413 (N_413,In_1042,In_52);
nor U414 (N_414,In_778,In_1025);
and U415 (N_415,In_1083,In_1018);
nand U416 (N_416,In_1405,In_741);
nand U417 (N_417,In_1460,In_821);
nor U418 (N_418,In_1044,In_1385);
nor U419 (N_419,In_113,In_1043);
or U420 (N_420,In_856,In_1086);
and U421 (N_421,In_389,In_1360);
nor U422 (N_422,In_97,In_744);
nand U423 (N_423,In_1011,In_502);
and U424 (N_424,In_938,In_584);
xnor U425 (N_425,In_179,In_696);
nor U426 (N_426,In_639,In_1284);
or U427 (N_427,In_853,In_1351);
and U428 (N_428,In_186,In_1167);
and U429 (N_429,In_848,In_617);
nand U430 (N_430,In_1065,In_1198);
or U431 (N_431,In_1416,In_959);
nand U432 (N_432,In_146,In_1050);
and U433 (N_433,In_432,In_1251);
nand U434 (N_434,In_136,In_659);
or U435 (N_435,In_1355,In_319);
nor U436 (N_436,In_1123,In_241);
and U437 (N_437,In_354,In_592);
nand U438 (N_438,In_850,In_310);
and U439 (N_439,In_1118,In_300);
nand U440 (N_440,In_919,In_221);
nand U441 (N_441,In_702,In_965);
and U442 (N_442,In_1431,In_266);
nand U443 (N_443,In_1439,In_578);
nand U444 (N_444,In_1139,In_572);
and U445 (N_445,In_168,In_1296);
nor U446 (N_446,In_307,In_988);
nand U447 (N_447,In_343,In_1498);
and U448 (N_448,In_19,In_305);
and U449 (N_449,In_1436,In_147);
xnor U450 (N_450,In_1489,In_1289);
or U451 (N_451,In_730,In_560);
nand U452 (N_452,In_392,In_1254);
nand U453 (N_453,In_638,In_1210);
and U454 (N_454,In_463,In_1358);
nand U455 (N_455,In_969,In_1095);
nand U456 (N_456,In_445,In_895);
and U457 (N_457,In_159,In_1054);
nand U458 (N_458,In_709,In_548);
or U459 (N_459,In_1391,In_1173);
and U460 (N_460,In_768,In_532);
nand U461 (N_461,In_475,In_1383);
and U462 (N_462,In_86,In_81);
nand U463 (N_463,In_1178,In_424);
nor U464 (N_464,In_177,In_697);
and U465 (N_465,In_1287,In_417);
or U466 (N_466,In_643,In_797);
nor U467 (N_467,In_369,In_815);
and U468 (N_468,In_731,In_843);
nand U469 (N_469,In_381,In_1007);
and U470 (N_470,In_1415,In_885);
and U471 (N_471,In_1449,In_240);
and U472 (N_472,In_1335,In_1352);
or U473 (N_473,In_1128,In_350);
or U474 (N_474,In_754,In_586);
nor U475 (N_475,In_380,In_686);
nand U476 (N_476,In_992,In_504);
and U477 (N_477,In_1046,In_939);
nand U478 (N_478,In_1101,In_742);
or U479 (N_479,In_562,In_962);
nand U480 (N_480,In_632,In_1216);
nor U481 (N_481,In_597,In_649);
or U482 (N_482,In_1270,In_936);
and U483 (N_483,In_1240,In_822);
and U484 (N_484,In_234,In_1197);
or U485 (N_485,In_736,In_1053);
nor U486 (N_486,In_225,In_150);
nor U487 (N_487,In_1370,In_250);
and U488 (N_488,In_871,In_1218);
and U489 (N_489,In_1288,In_1494);
nor U490 (N_490,In_272,In_1482);
and U491 (N_491,In_1474,In_629);
nor U492 (N_492,In_673,In_1447);
and U493 (N_493,In_1425,In_1148);
or U494 (N_494,In_847,In_677);
nor U495 (N_495,In_521,In_70);
nand U496 (N_496,In_441,In_1126);
and U497 (N_497,In_316,In_658);
and U498 (N_498,In_813,In_626);
nand U499 (N_499,In_255,In_1013);
or U500 (N_500,In_1223,In_1048);
nand U501 (N_501,In_203,In_1129);
xnor U502 (N_502,In_1028,In_85);
and U503 (N_503,In_358,In_817);
and U504 (N_504,In_1466,In_779);
or U505 (N_505,In_56,In_612);
nor U506 (N_506,In_520,In_1222);
and U507 (N_507,In_623,In_713);
nor U508 (N_508,In_1321,In_173);
and U509 (N_509,In_447,In_941);
and U510 (N_510,In_732,In_41);
or U511 (N_511,In_339,In_1291);
or U512 (N_512,In_1228,In_879);
nor U513 (N_513,In_1034,In_104);
or U514 (N_514,In_863,In_610);
or U515 (N_515,In_890,In_714);
or U516 (N_516,In_304,In_972);
or U517 (N_517,In_1188,In_286);
nor U518 (N_518,In_185,In_1477);
nand U519 (N_519,In_554,In_1304);
nand U520 (N_520,In_1363,In_761);
or U521 (N_521,In_699,In_746);
nand U522 (N_522,In_611,In_841);
or U523 (N_523,In_275,In_704);
or U524 (N_524,In_438,In_573);
nand U525 (N_525,In_27,In_28);
or U526 (N_526,In_61,In_529);
nand U527 (N_527,In_791,In_531);
nor U528 (N_528,In_1233,In_226);
and U529 (N_529,In_830,In_1219);
or U530 (N_530,In_1180,In_287);
nand U531 (N_531,In_1045,In_1093);
nand U532 (N_532,In_482,In_869);
or U533 (N_533,In_738,In_1243);
and U534 (N_534,In_395,In_94);
and U535 (N_535,In_589,In_1248);
nand U536 (N_536,In_625,In_1339);
or U537 (N_537,In_1266,In_284);
nand U538 (N_538,In_180,In_769);
nor U539 (N_539,In_1002,In_1483);
nand U540 (N_540,In_465,In_74);
nand U541 (N_541,In_71,In_1242);
nand U542 (N_542,In_317,In_1021);
and U543 (N_543,In_726,In_1346);
nand U544 (N_544,In_98,In_792);
nor U545 (N_545,In_280,In_342);
or U546 (N_546,In_373,In_1215);
and U547 (N_547,In_1029,In_698);
and U548 (N_548,In_1282,In_581);
nor U549 (N_549,In_77,In_899);
and U550 (N_550,In_975,In_1039);
nand U551 (N_551,In_902,In_158);
or U552 (N_552,In_321,In_326);
xnor U553 (N_553,In_996,In_6);
or U554 (N_554,In_120,In_1488);
nor U555 (N_555,In_807,In_1138);
and U556 (N_556,In_1277,In_837);
or U557 (N_557,In_957,In_600);
nor U558 (N_558,In_570,In_654);
or U559 (N_559,In_346,In_1286);
nor U560 (N_560,In_231,In_1121);
and U561 (N_561,In_411,In_341);
and U562 (N_562,In_278,In_397);
and U563 (N_563,In_745,In_862);
or U564 (N_564,In_131,In_1276);
nand U565 (N_565,In_1458,In_1120);
nor U566 (N_566,In_1473,In_897);
and U567 (N_567,In_691,In_1424);
or U568 (N_568,In_1470,In_728);
or U569 (N_569,In_7,In_290);
nand U570 (N_570,In_892,In_281);
nor U571 (N_571,In_1076,In_170);
and U572 (N_572,In_1131,In_1195);
and U573 (N_573,In_1239,In_88);
nand U574 (N_574,In_1263,In_1328);
and U575 (N_575,In_894,In_1317);
or U576 (N_576,In_181,In_558);
or U577 (N_577,In_687,In_923);
and U578 (N_578,In_256,In_78);
or U579 (N_579,In_802,In_68);
nor U580 (N_580,In_215,In_985);
nor U581 (N_581,In_716,In_1006);
or U582 (N_582,In_1404,In_803);
nor U583 (N_583,In_507,In_1354);
nor U584 (N_584,In_794,In_1454);
or U585 (N_585,In_1030,In_789);
nand U586 (N_586,In_723,In_499);
or U587 (N_587,In_689,In_743);
nand U588 (N_588,In_1397,In_690);
and U589 (N_589,In_1165,In_1159);
or U590 (N_590,In_878,In_1127);
nor U591 (N_591,In_1272,In_218);
or U592 (N_592,In_811,In_207);
nand U593 (N_593,In_775,In_1241);
and U594 (N_594,In_893,In_1484);
xor U595 (N_595,In_1171,In_804);
and U596 (N_596,In_1103,In_546);
or U597 (N_597,In_1015,In_958);
and U598 (N_598,In_500,In_1326);
xor U599 (N_599,In_220,In_613);
or U600 (N_600,In_431,In_1114);
nor U601 (N_601,In_1490,In_1308);
nand U602 (N_602,In_1305,In_948);
nor U603 (N_603,In_62,In_925);
nand U604 (N_604,In_536,In_1125);
nor U605 (N_605,In_913,In_387);
nor U606 (N_606,In_655,In_116);
nor U607 (N_607,In_374,In_561);
nand U608 (N_608,In_371,In_337);
or U609 (N_609,In_418,In_553);
and U610 (N_610,In_455,In_650);
nor U611 (N_611,In_882,In_296);
nor U612 (N_612,In_866,In_701);
nor U613 (N_613,In_660,In_844);
nor U614 (N_614,In_205,In_138);
nor U615 (N_615,In_1299,In_91);
nor U616 (N_616,In_1224,In_25);
nor U617 (N_617,In_509,In_541);
nor U618 (N_618,In_727,In_710);
or U619 (N_619,In_219,In_1108);
or U620 (N_620,In_740,In_997);
nor U621 (N_621,In_1398,In_201);
nand U622 (N_622,In_384,In_247);
or U623 (N_623,In_210,In_960);
or U624 (N_624,In_360,In_1230);
and U625 (N_625,In_524,In_1098);
or U626 (N_626,In_987,In_484);
nand U627 (N_627,In_95,In_437);
nand U628 (N_628,In_842,In_1226);
or U629 (N_629,In_907,In_1309);
xor U630 (N_630,In_1341,In_1208);
nor U631 (N_631,In_1213,In_117);
nor U632 (N_632,In_903,In_1367);
and U633 (N_633,In_160,In_685);
nand U634 (N_634,In_648,In_1353);
and U635 (N_635,In_926,In_805);
nor U636 (N_636,In_416,In_230);
or U637 (N_637,In_525,In_36);
or U638 (N_638,In_449,In_984);
and U639 (N_639,In_142,In_891);
nor U640 (N_640,In_1476,In_722);
xnor U641 (N_641,In_1008,In_149);
or U642 (N_642,In_911,In_38);
nor U643 (N_643,In_273,In_1201);
or U644 (N_644,In_624,In_1026);
and U645 (N_645,In_538,In_942);
and U646 (N_646,In_200,In_223);
xnor U647 (N_647,In_1179,In_349);
nor U648 (N_648,In_1122,In_1019);
or U649 (N_649,In_129,In_1350);
nand U650 (N_650,In_1462,In_820);
nor U651 (N_651,In_549,In_1037);
and U652 (N_652,In_1100,In_929);
or U653 (N_653,In_550,In_1009);
and U654 (N_654,In_666,In_1004);
and U655 (N_655,In_84,In_410);
nor U656 (N_656,In_593,In_860);
and U657 (N_657,In_401,In_110);
and U658 (N_658,In_777,In_684);
nand U659 (N_659,In_800,In_353);
nor U660 (N_660,In_896,In_1152);
or U661 (N_661,In_906,In_591);
nor U662 (N_662,In_90,In_868);
nand U663 (N_663,In_1041,In_1113);
nand U664 (N_664,In_1255,In_1496);
nor U665 (N_665,In_946,In_886);
and U666 (N_666,In_285,In_530);
nand U667 (N_667,In_1185,In_1395);
nor U668 (N_668,In_616,In_107);
or U669 (N_669,In_522,In_663);
or U670 (N_670,In_937,In_1153);
and U671 (N_671,In_362,In_1244);
nand U672 (N_672,In_748,In_1089);
xor U673 (N_673,In_453,In_433);
nand U674 (N_674,In_423,In_1485);
and U675 (N_675,In_409,In_299);
and U676 (N_676,In_935,In_1177);
nand U677 (N_677,In_944,In_1104);
and U678 (N_678,In_364,In_582);
and U679 (N_679,In_188,In_67);
nand U680 (N_680,In_60,In_788);
nor U681 (N_681,In_96,In_2);
or U682 (N_682,In_1364,In_1081);
nand U683 (N_683,In_314,In_542);
nor U684 (N_684,In_209,In_1214);
nor U685 (N_685,In_993,In_535);
nand U686 (N_686,In_420,In_471);
nor U687 (N_687,In_1384,In_724);
nor U688 (N_688,In_547,In_711);
or U689 (N_689,In_1492,In_1298);
and U690 (N_690,In_787,In_1146);
nor U691 (N_691,In_265,In_1141);
nand U692 (N_692,In_601,In_1313);
and U693 (N_693,In_615,In_194);
and U694 (N_694,In_39,In_26);
nor U695 (N_695,In_118,In_480);
nand U696 (N_696,In_607,In_383);
nor U697 (N_697,In_1140,In_566);
nand U698 (N_698,In_172,In_812);
and U699 (N_699,In_662,In_10);
nand U700 (N_700,In_861,In_248);
and U701 (N_701,In_419,In_137);
and U702 (N_702,In_1323,In_402);
xnor U703 (N_703,In_932,In_115);
nor U704 (N_704,In_1134,In_1090);
nor U705 (N_705,In_356,In_124);
or U706 (N_706,In_143,In_335);
xnor U707 (N_707,In_845,In_501);
and U708 (N_708,In_651,In_977);
nand U709 (N_709,In_1388,In_439);
and U710 (N_710,In_212,In_1486);
nor U711 (N_711,In_1316,In_865);
or U712 (N_712,In_22,In_1016);
nor U713 (N_713,In_1407,In_963);
nand U714 (N_714,In_1380,In_308);
nor U715 (N_715,In_1301,In_764);
and U716 (N_716,In_211,In_32);
and U717 (N_717,In_289,In_1144);
and U718 (N_718,In_76,In_382);
or U719 (N_719,In_1481,In_333);
and U720 (N_720,In_65,In_806);
or U721 (N_721,In_1117,In_1092);
and U722 (N_722,In_1463,In_325);
nor U723 (N_723,In_1247,In_486);
and U724 (N_724,In_0,In_1068);
nor U725 (N_725,In_1338,In_1158);
or U726 (N_726,In_324,In_1105);
and U727 (N_727,In_1389,In_31);
nand U728 (N_728,In_193,In_1347);
nand U729 (N_729,In_332,In_758);
and U730 (N_730,In_604,In_976);
nand U731 (N_731,In_540,In_89);
nand U732 (N_732,In_1318,In_839);
nor U733 (N_733,In_141,In_657);
and U734 (N_734,In_1461,In_1281);
or U735 (N_735,In_867,In_1437);
nand U736 (N_736,In_665,In_810);
or U737 (N_737,In_456,In_254);
nor U738 (N_738,In_1295,In_1061);
or U739 (N_739,In_1302,In_452);
or U740 (N_740,In_357,In_257);
or U741 (N_741,In_1056,In_1472);
or U742 (N_742,In_1374,In_1499);
and U743 (N_743,In_40,In_1209);
or U744 (N_744,In_30,In_1010);
nor U745 (N_745,In_347,In_1135);
and U746 (N_746,In_1292,In_1433);
nor U747 (N_747,In_909,In_144);
nand U748 (N_748,In_670,In_523);
or U749 (N_749,In_1196,In_1396);
nand U750 (N_750,In_1411,In_394);
and U751 (N_751,In_1494,In_401);
or U752 (N_752,In_1334,In_347);
or U753 (N_753,In_1062,In_159);
and U754 (N_754,In_1169,In_1397);
nor U755 (N_755,In_863,In_0);
nand U756 (N_756,In_1261,In_1371);
or U757 (N_757,In_627,In_426);
nor U758 (N_758,In_1342,In_660);
nand U759 (N_759,In_1269,In_573);
nor U760 (N_760,In_1312,In_924);
nand U761 (N_761,In_484,In_447);
or U762 (N_762,In_1174,In_480);
nand U763 (N_763,In_776,In_439);
and U764 (N_764,In_286,In_497);
or U765 (N_765,In_1480,In_1279);
or U766 (N_766,In_201,In_182);
nor U767 (N_767,In_327,In_222);
and U768 (N_768,In_1295,In_592);
or U769 (N_769,In_317,In_513);
nor U770 (N_770,In_527,In_1441);
and U771 (N_771,In_1082,In_1489);
nor U772 (N_772,In_290,In_208);
xor U773 (N_773,In_1177,In_42);
and U774 (N_774,In_612,In_707);
nand U775 (N_775,In_444,In_91);
nand U776 (N_776,In_1323,In_1372);
nand U777 (N_777,In_797,In_864);
or U778 (N_778,In_1171,In_622);
xor U779 (N_779,In_564,In_1155);
and U780 (N_780,In_586,In_352);
nor U781 (N_781,In_44,In_106);
xnor U782 (N_782,In_1219,In_684);
nor U783 (N_783,In_1371,In_881);
or U784 (N_784,In_198,In_802);
nand U785 (N_785,In_905,In_1426);
and U786 (N_786,In_700,In_1067);
and U787 (N_787,In_1172,In_770);
nor U788 (N_788,In_365,In_880);
nand U789 (N_789,In_1365,In_211);
nor U790 (N_790,In_1487,In_233);
nor U791 (N_791,In_1021,In_794);
nor U792 (N_792,In_395,In_422);
and U793 (N_793,In_108,In_1339);
and U794 (N_794,In_396,In_448);
nor U795 (N_795,In_1389,In_554);
nor U796 (N_796,In_1440,In_763);
nor U797 (N_797,In_1322,In_615);
nand U798 (N_798,In_995,In_483);
and U799 (N_799,In_1301,In_116);
nand U800 (N_800,In_1369,In_283);
nor U801 (N_801,In_819,In_1482);
and U802 (N_802,In_1146,In_637);
nand U803 (N_803,In_1408,In_4);
nor U804 (N_804,In_547,In_486);
or U805 (N_805,In_135,In_1305);
nor U806 (N_806,In_683,In_633);
and U807 (N_807,In_633,In_897);
nand U808 (N_808,In_104,In_170);
or U809 (N_809,In_845,In_1291);
and U810 (N_810,In_43,In_314);
nor U811 (N_811,In_1287,In_537);
nor U812 (N_812,In_778,In_766);
nand U813 (N_813,In_943,In_1177);
xnor U814 (N_814,In_948,In_821);
nor U815 (N_815,In_1312,In_606);
and U816 (N_816,In_1396,In_493);
nand U817 (N_817,In_1258,In_68);
nor U818 (N_818,In_175,In_958);
nand U819 (N_819,In_90,In_689);
nor U820 (N_820,In_1271,In_907);
and U821 (N_821,In_10,In_491);
and U822 (N_822,In_1079,In_1249);
or U823 (N_823,In_642,In_281);
nand U824 (N_824,In_901,In_1073);
xnor U825 (N_825,In_1057,In_1178);
or U826 (N_826,In_865,In_332);
or U827 (N_827,In_419,In_514);
or U828 (N_828,In_965,In_398);
nor U829 (N_829,In_396,In_651);
and U830 (N_830,In_1314,In_1127);
nor U831 (N_831,In_537,In_993);
or U832 (N_832,In_330,In_1023);
xnor U833 (N_833,In_326,In_833);
nor U834 (N_834,In_393,In_989);
nor U835 (N_835,In_1160,In_1220);
nand U836 (N_836,In_765,In_514);
or U837 (N_837,In_517,In_585);
and U838 (N_838,In_1161,In_1328);
nand U839 (N_839,In_523,In_230);
nor U840 (N_840,In_1460,In_625);
nand U841 (N_841,In_350,In_95);
or U842 (N_842,In_277,In_1075);
and U843 (N_843,In_449,In_868);
xnor U844 (N_844,In_783,In_183);
or U845 (N_845,In_1265,In_759);
and U846 (N_846,In_40,In_410);
nor U847 (N_847,In_1425,In_1163);
and U848 (N_848,In_1318,In_389);
nand U849 (N_849,In_1406,In_1291);
and U850 (N_850,In_229,In_359);
and U851 (N_851,In_542,In_1344);
nor U852 (N_852,In_511,In_364);
nand U853 (N_853,In_370,In_1482);
and U854 (N_854,In_350,In_1112);
nor U855 (N_855,In_1194,In_996);
nor U856 (N_856,In_142,In_315);
and U857 (N_857,In_732,In_226);
nand U858 (N_858,In_838,In_121);
nand U859 (N_859,In_367,In_180);
and U860 (N_860,In_253,In_671);
xor U861 (N_861,In_1366,In_757);
and U862 (N_862,In_1374,In_594);
nand U863 (N_863,In_732,In_393);
xnor U864 (N_864,In_708,In_1346);
and U865 (N_865,In_1165,In_982);
nor U866 (N_866,In_1418,In_1064);
or U867 (N_867,In_413,In_1177);
and U868 (N_868,In_1098,In_35);
or U869 (N_869,In_268,In_1285);
nand U870 (N_870,In_793,In_784);
or U871 (N_871,In_809,In_565);
nand U872 (N_872,In_1137,In_881);
nand U873 (N_873,In_1359,In_1163);
xor U874 (N_874,In_374,In_1128);
or U875 (N_875,In_239,In_1068);
nand U876 (N_876,In_823,In_293);
or U877 (N_877,In_735,In_1103);
nand U878 (N_878,In_653,In_808);
or U879 (N_879,In_1056,In_314);
or U880 (N_880,In_1014,In_1360);
and U881 (N_881,In_169,In_1374);
nand U882 (N_882,In_511,In_577);
nand U883 (N_883,In_1001,In_311);
or U884 (N_884,In_1055,In_1112);
or U885 (N_885,In_374,In_86);
nand U886 (N_886,In_301,In_1154);
nand U887 (N_887,In_60,In_155);
and U888 (N_888,In_1064,In_1311);
or U889 (N_889,In_108,In_735);
or U890 (N_890,In_1388,In_256);
nor U891 (N_891,In_250,In_258);
nand U892 (N_892,In_982,In_517);
or U893 (N_893,In_1029,In_1349);
or U894 (N_894,In_72,In_731);
nor U895 (N_895,In_218,In_2);
nand U896 (N_896,In_997,In_9);
nor U897 (N_897,In_892,In_153);
nor U898 (N_898,In_159,In_1070);
and U899 (N_899,In_1198,In_207);
or U900 (N_900,In_719,In_254);
nor U901 (N_901,In_1301,In_679);
nand U902 (N_902,In_603,In_375);
nand U903 (N_903,In_899,In_61);
and U904 (N_904,In_167,In_1063);
nand U905 (N_905,In_227,In_1133);
xnor U906 (N_906,In_789,In_111);
and U907 (N_907,In_1296,In_87);
and U908 (N_908,In_983,In_788);
nor U909 (N_909,In_333,In_1031);
and U910 (N_910,In_423,In_321);
nand U911 (N_911,In_1280,In_405);
nor U912 (N_912,In_346,In_1253);
or U913 (N_913,In_62,In_525);
or U914 (N_914,In_360,In_291);
or U915 (N_915,In_1202,In_1124);
nor U916 (N_916,In_1264,In_1405);
or U917 (N_917,In_592,In_579);
nor U918 (N_918,In_996,In_982);
nor U919 (N_919,In_738,In_998);
or U920 (N_920,In_928,In_352);
and U921 (N_921,In_1038,In_783);
nand U922 (N_922,In_1066,In_445);
nor U923 (N_923,In_316,In_678);
and U924 (N_924,In_1079,In_287);
nor U925 (N_925,In_127,In_1254);
nor U926 (N_926,In_529,In_331);
and U927 (N_927,In_1443,In_710);
nand U928 (N_928,In_79,In_72);
nor U929 (N_929,In_777,In_1191);
nor U930 (N_930,In_124,In_297);
or U931 (N_931,In_127,In_1286);
nor U932 (N_932,In_1417,In_1062);
and U933 (N_933,In_940,In_671);
and U934 (N_934,In_987,In_55);
or U935 (N_935,In_1263,In_212);
nand U936 (N_936,In_522,In_991);
nand U937 (N_937,In_1286,In_868);
nor U938 (N_938,In_19,In_879);
nor U939 (N_939,In_5,In_519);
or U940 (N_940,In_1012,In_674);
nor U941 (N_941,In_963,In_1215);
or U942 (N_942,In_694,In_627);
nand U943 (N_943,In_78,In_307);
xor U944 (N_944,In_1275,In_1410);
nand U945 (N_945,In_291,In_1357);
nor U946 (N_946,In_957,In_1054);
nand U947 (N_947,In_280,In_1343);
or U948 (N_948,In_1258,In_524);
nor U949 (N_949,In_1296,In_199);
or U950 (N_950,In_198,In_499);
nand U951 (N_951,In_826,In_1476);
and U952 (N_952,In_382,In_44);
nor U953 (N_953,In_1430,In_796);
or U954 (N_954,In_1368,In_1076);
nand U955 (N_955,In_482,In_250);
or U956 (N_956,In_247,In_897);
nand U957 (N_957,In_176,In_534);
nand U958 (N_958,In_1261,In_674);
or U959 (N_959,In_517,In_557);
and U960 (N_960,In_886,In_1129);
or U961 (N_961,In_1372,In_548);
or U962 (N_962,In_150,In_305);
nand U963 (N_963,In_1447,In_1036);
or U964 (N_964,In_257,In_641);
or U965 (N_965,In_1266,In_1491);
nand U966 (N_966,In_2,In_676);
and U967 (N_967,In_596,In_1045);
nor U968 (N_968,In_186,In_757);
and U969 (N_969,In_251,In_901);
or U970 (N_970,In_470,In_404);
and U971 (N_971,In_361,In_693);
nand U972 (N_972,In_1270,In_1007);
nand U973 (N_973,In_528,In_432);
and U974 (N_974,In_874,In_958);
xnor U975 (N_975,In_593,In_414);
or U976 (N_976,In_444,In_462);
nand U977 (N_977,In_1434,In_719);
and U978 (N_978,In_563,In_378);
and U979 (N_979,In_16,In_908);
or U980 (N_980,In_226,In_111);
and U981 (N_981,In_343,In_472);
and U982 (N_982,In_1,In_471);
or U983 (N_983,In_1091,In_284);
or U984 (N_984,In_625,In_735);
nand U985 (N_985,In_1020,In_1210);
nor U986 (N_986,In_814,In_658);
nor U987 (N_987,In_796,In_270);
or U988 (N_988,In_148,In_1090);
and U989 (N_989,In_452,In_281);
nand U990 (N_990,In_1309,In_594);
and U991 (N_991,In_945,In_1487);
nand U992 (N_992,In_871,In_988);
and U993 (N_993,In_1187,In_580);
and U994 (N_994,In_890,In_944);
nor U995 (N_995,In_1249,In_357);
or U996 (N_996,In_732,In_784);
and U997 (N_997,In_397,In_647);
and U998 (N_998,In_221,In_1118);
or U999 (N_999,In_1487,In_1326);
nand U1000 (N_1000,In_567,In_910);
nand U1001 (N_1001,In_39,In_1323);
nor U1002 (N_1002,In_1028,In_364);
or U1003 (N_1003,In_625,In_1349);
or U1004 (N_1004,In_303,In_1490);
or U1005 (N_1005,In_837,In_1137);
or U1006 (N_1006,In_1498,In_249);
and U1007 (N_1007,In_577,In_1006);
nor U1008 (N_1008,In_1348,In_823);
and U1009 (N_1009,In_385,In_481);
or U1010 (N_1010,In_96,In_308);
or U1011 (N_1011,In_1401,In_325);
nand U1012 (N_1012,In_1115,In_30);
and U1013 (N_1013,In_773,In_535);
nand U1014 (N_1014,In_1480,In_694);
or U1015 (N_1015,In_213,In_906);
nor U1016 (N_1016,In_1402,In_1171);
or U1017 (N_1017,In_772,In_1371);
and U1018 (N_1018,In_1289,In_887);
and U1019 (N_1019,In_690,In_580);
nand U1020 (N_1020,In_1220,In_584);
and U1021 (N_1021,In_756,In_700);
nand U1022 (N_1022,In_39,In_1197);
nand U1023 (N_1023,In_141,In_831);
nor U1024 (N_1024,In_864,In_280);
nor U1025 (N_1025,In_543,In_248);
and U1026 (N_1026,In_293,In_814);
and U1027 (N_1027,In_1304,In_637);
nor U1028 (N_1028,In_145,In_583);
and U1029 (N_1029,In_761,In_457);
and U1030 (N_1030,In_1020,In_1235);
or U1031 (N_1031,In_9,In_1250);
or U1032 (N_1032,In_267,In_1379);
nor U1033 (N_1033,In_1411,In_62);
and U1034 (N_1034,In_14,In_1190);
nor U1035 (N_1035,In_555,In_585);
xnor U1036 (N_1036,In_1274,In_1231);
or U1037 (N_1037,In_665,In_656);
and U1038 (N_1038,In_1473,In_288);
nor U1039 (N_1039,In_484,In_1179);
nor U1040 (N_1040,In_1333,In_583);
and U1041 (N_1041,In_1055,In_524);
or U1042 (N_1042,In_847,In_1256);
nor U1043 (N_1043,In_330,In_1490);
nand U1044 (N_1044,In_660,In_641);
or U1045 (N_1045,In_277,In_534);
nor U1046 (N_1046,In_1022,In_1130);
nor U1047 (N_1047,In_985,In_1088);
or U1048 (N_1048,In_1304,In_505);
nand U1049 (N_1049,In_1052,In_1077);
and U1050 (N_1050,In_933,In_869);
nor U1051 (N_1051,In_1172,In_1327);
nor U1052 (N_1052,In_325,In_1056);
nand U1053 (N_1053,In_968,In_741);
xor U1054 (N_1054,In_1036,In_770);
nand U1055 (N_1055,In_1291,In_303);
nand U1056 (N_1056,In_233,In_169);
or U1057 (N_1057,In_1263,In_824);
nand U1058 (N_1058,In_764,In_885);
nor U1059 (N_1059,In_1432,In_675);
xor U1060 (N_1060,In_633,In_649);
or U1061 (N_1061,In_807,In_683);
and U1062 (N_1062,In_22,In_445);
and U1063 (N_1063,In_1058,In_1445);
and U1064 (N_1064,In_611,In_494);
and U1065 (N_1065,In_266,In_185);
nand U1066 (N_1066,In_1022,In_26);
nand U1067 (N_1067,In_779,In_405);
or U1068 (N_1068,In_1484,In_151);
nand U1069 (N_1069,In_121,In_771);
and U1070 (N_1070,In_346,In_317);
and U1071 (N_1071,In_1083,In_792);
and U1072 (N_1072,In_426,In_353);
nor U1073 (N_1073,In_664,In_486);
or U1074 (N_1074,In_868,In_695);
or U1075 (N_1075,In_248,In_196);
nand U1076 (N_1076,In_160,In_1486);
or U1077 (N_1077,In_1445,In_100);
nor U1078 (N_1078,In_906,In_708);
nand U1079 (N_1079,In_45,In_1386);
nor U1080 (N_1080,In_32,In_1199);
nand U1081 (N_1081,In_878,In_170);
nor U1082 (N_1082,In_731,In_303);
nor U1083 (N_1083,In_1253,In_465);
nand U1084 (N_1084,In_679,In_754);
or U1085 (N_1085,In_550,In_830);
or U1086 (N_1086,In_560,In_168);
nor U1087 (N_1087,In_1069,In_672);
nor U1088 (N_1088,In_107,In_1080);
or U1089 (N_1089,In_677,In_1117);
and U1090 (N_1090,In_1004,In_134);
and U1091 (N_1091,In_690,In_435);
or U1092 (N_1092,In_412,In_500);
and U1093 (N_1093,In_1219,In_1272);
nand U1094 (N_1094,In_777,In_379);
nand U1095 (N_1095,In_360,In_94);
or U1096 (N_1096,In_1229,In_1030);
nor U1097 (N_1097,In_796,In_352);
nor U1098 (N_1098,In_276,In_1475);
or U1099 (N_1099,In_1215,In_223);
nand U1100 (N_1100,In_795,In_947);
or U1101 (N_1101,In_1161,In_917);
and U1102 (N_1102,In_274,In_1336);
nor U1103 (N_1103,In_901,In_1033);
nand U1104 (N_1104,In_824,In_125);
and U1105 (N_1105,In_1217,In_1370);
nor U1106 (N_1106,In_1097,In_1341);
nand U1107 (N_1107,In_762,In_935);
or U1108 (N_1108,In_317,In_1382);
nand U1109 (N_1109,In_625,In_502);
nor U1110 (N_1110,In_58,In_1479);
nor U1111 (N_1111,In_1162,In_1387);
and U1112 (N_1112,In_211,In_1311);
or U1113 (N_1113,In_413,In_645);
nor U1114 (N_1114,In_577,In_738);
or U1115 (N_1115,In_387,In_246);
and U1116 (N_1116,In_1167,In_846);
nor U1117 (N_1117,In_698,In_1209);
nor U1118 (N_1118,In_473,In_257);
and U1119 (N_1119,In_1179,In_661);
nor U1120 (N_1120,In_1387,In_675);
or U1121 (N_1121,In_598,In_1018);
or U1122 (N_1122,In_724,In_1336);
and U1123 (N_1123,In_140,In_308);
and U1124 (N_1124,In_537,In_1468);
nand U1125 (N_1125,In_970,In_1142);
nor U1126 (N_1126,In_1464,In_834);
or U1127 (N_1127,In_1422,In_951);
nor U1128 (N_1128,In_1407,In_1359);
nand U1129 (N_1129,In_1488,In_816);
or U1130 (N_1130,In_1017,In_737);
or U1131 (N_1131,In_1251,In_1250);
and U1132 (N_1132,In_811,In_373);
nand U1133 (N_1133,In_1439,In_935);
nor U1134 (N_1134,In_903,In_812);
and U1135 (N_1135,In_1279,In_1164);
nor U1136 (N_1136,In_1145,In_416);
nand U1137 (N_1137,In_89,In_497);
nand U1138 (N_1138,In_178,In_1130);
nand U1139 (N_1139,In_856,In_460);
nand U1140 (N_1140,In_105,In_191);
or U1141 (N_1141,In_616,In_830);
xor U1142 (N_1142,In_1438,In_867);
and U1143 (N_1143,In_1055,In_785);
xnor U1144 (N_1144,In_1081,In_264);
nand U1145 (N_1145,In_586,In_683);
or U1146 (N_1146,In_726,In_1122);
and U1147 (N_1147,In_647,In_1341);
xor U1148 (N_1148,In_775,In_85);
nor U1149 (N_1149,In_113,In_1386);
or U1150 (N_1150,In_541,In_929);
or U1151 (N_1151,In_767,In_90);
nor U1152 (N_1152,In_246,In_723);
or U1153 (N_1153,In_544,In_1079);
or U1154 (N_1154,In_638,In_418);
and U1155 (N_1155,In_282,In_239);
or U1156 (N_1156,In_1281,In_609);
and U1157 (N_1157,In_1281,In_1394);
or U1158 (N_1158,In_868,In_552);
and U1159 (N_1159,In_682,In_871);
nor U1160 (N_1160,In_173,In_49);
or U1161 (N_1161,In_1309,In_589);
nand U1162 (N_1162,In_850,In_778);
xnor U1163 (N_1163,In_247,In_1282);
nand U1164 (N_1164,In_1142,In_497);
nor U1165 (N_1165,In_1228,In_454);
nand U1166 (N_1166,In_25,In_1328);
nor U1167 (N_1167,In_1482,In_343);
or U1168 (N_1168,In_902,In_320);
and U1169 (N_1169,In_204,In_414);
nand U1170 (N_1170,In_646,In_1337);
or U1171 (N_1171,In_1441,In_336);
and U1172 (N_1172,In_1202,In_1382);
or U1173 (N_1173,In_832,In_831);
or U1174 (N_1174,In_769,In_315);
nand U1175 (N_1175,In_475,In_1403);
or U1176 (N_1176,In_1420,In_152);
nand U1177 (N_1177,In_959,In_966);
and U1178 (N_1178,In_1012,In_818);
and U1179 (N_1179,In_1249,In_219);
or U1180 (N_1180,In_1428,In_1325);
nor U1181 (N_1181,In_1017,In_1366);
nor U1182 (N_1182,In_381,In_1107);
or U1183 (N_1183,In_1470,In_1020);
nor U1184 (N_1184,In_1108,In_1184);
xor U1185 (N_1185,In_1361,In_533);
and U1186 (N_1186,In_675,In_1361);
and U1187 (N_1187,In_1238,In_1055);
or U1188 (N_1188,In_1037,In_721);
nor U1189 (N_1189,In_136,In_948);
and U1190 (N_1190,In_725,In_768);
or U1191 (N_1191,In_251,In_1452);
xnor U1192 (N_1192,In_1374,In_542);
nand U1193 (N_1193,In_154,In_580);
nor U1194 (N_1194,In_1396,In_332);
or U1195 (N_1195,In_768,In_1102);
and U1196 (N_1196,In_450,In_379);
xor U1197 (N_1197,In_471,In_683);
or U1198 (N_1198,In_976,In_717);
nor U1199 (N_1199,In_83,In_286);
nand U1200 (N_1200,In_621,In_127);
and U1201 (N_1201,In_302,In_1144);
and U1202 (N_1202,In_855,In_1296);
nand U1203 (N_1203,In_1264,In_1415);
and U1204 (N_1204,In_54,In_766);
nor U1205 (N_1205,In_481,In_511);
nand U1206 (N_1206,In_929,In_93);
or U1207 (N_1207,In_809,In_1375);
nand U1208 (N_1208,In_403,In_1441);
nand U1209 (N_1209,In_870,In_218);
or U1210 (N_1210,In_736,In_282);
or U1211 (N_1211,In_92,In_493);
or U1212 (N_1212,In_797,In_810);
nor U1213 (N_1213,In_312,In_118);
nand U1214 (N_1214,In_166,In_277);
and U1215 (N_1215,In_817,In_171);
and U1216 (N_1216,In_1351,In_1013);
xnor U1217 (N_1217,In_593,In_208);
or U1218 (N_1218,In_1392,In_608);
nor U1219 (N_1219,In_1238,In_37);
or U1220 (N_1220,In_1034,In_263);
or U1221 (N_1221,In_1035,In_398);
and U1222 (N_1222,In_1026,In_362);
nor U1223 (N_1223,In_1373,In_950);
nand U1224 (N_1224,In_1168,In_317);
nand U1225 (N_1225,In_302,In_1097);
nand U1226 (N_1226,In_350,In_45);
and U1227 (N_1227,In_1136,In_811);
and U1228 (N_1228,In_539,In_294);
and U1229 (N_1229,In_1368,In_809);
nand U1230 (N_1230,In_269,In_855);
or U1231 (N_1231,In_275,In_44);
and U1232 (N_1232,In_634,In_1135);
and U1233 (N_1233,In_52,In_88);
nor U1234 (N_1234,In_130,In_758);
or U1235 (N_1235,In_12,In_14);
and U1236 (N_1236,In_1049,In_1199);
and U1237 (N_1237,In_187,In_1054);
nand U1238 (N_1238,In_1111,In_31);
or U1239 (N_1239,In_352,In_415);
xnor U1240 (N_1240,In_445,In_773);
nand U1241 (N_1241,In_1346,In_1148);
nor U1242 (N_1242,In_1317,In_590);
and U1243 (N_1243,In_1203,In_105);
and U1244 (N_1244,In_787,In_604);
and U1245 (N_1245,In_1371,In_489);
or U1246 (N_1246,In_162,In_1354);
nor U1247 (N_1247,In_1308,In_776);
and U1248 (N_1248,In_151,In_1019);
nor U1249 (N_1249,In_315,In_519);
nor U1250 (N_1250,In_613,In_519);
and U1251 (N_1251,In_265,In_670);
and U1252 (N_1252,In_1370,In_1044);
or U1253 (N_1253,In_1360,In_954);
nand U1254 (N_1254,In_1072,In_1487);
or U1255 (N_1255,In_1091,In_424);
nand U1256 (N_1256,In_434,In_1372);
and U1257 (N_1257,In_1394,In_413);
nand U1258 (N_1258,In_1498,In_1407);
nand U1259 (N_1259,In_245,In_1190);
and U1260 (N_1260,In_915,In_1019);
or U1261 (N_1261,In_97,In_768);
nor U1262 (N_1262,In_1499,In_1389);
or U1263 (N_1263,In_1278,In_350);
nand U1264 (N_1264,In_595,In_1221);
nor U1265 (N_1265,In_515,In_1332);
or U1266 (N_1266,In_259,In_1152);
or U1267 (N_1267,In_569,In_1298);
or U1268 (N_1268,In_523,In_1428);
nor U1269 (N_1269,In_977,In_766);
or U1270 (N_1270,In_1020,In_1032);
nand U1271 (N_1271,In_779,In_383);
or U1272 (N_1272,In_1038,In_36);
and U1273 (N_1273,In_116,In_1048);
xor U1274 (N_1274,In_223,In_513);
and U1275 (N_1275,In_554,In_582);
and U1276 (N_1276,In_133,In_137);
nor U1277 (N_1277,In_843,In_421);
or U1278 (N_1278,In_381,In_77);
nor U1279 (N_1279,In_2,In_88);
xor U1280 (N_1280,In_1073,In_1010);
nor U1281 (N_1281,In_952,In_254);
or U1282 (N_1282,In_589,In_444);
and U1283 (N_1283,In_1432,In_236);
nor U1284 (N_1284,In_645,In_1339);
nand U1285 (N_1285,In_1366,In_1277);
nor U1286 (N_1286,In_1141,In_970);
and U1287 (N_1287,In_1096,In_243);
nor U1288 (N_1288,In_658,In_785);
and U1289 (N_1289,In_725,In_419);
nand U1290 (N_1290,In_404,In_688);
nor U1291 (N_1291,In_479,In_1213);
and U1292 (N_1292,In_1333,In_114);
nor U1293 (N_1293,In_1401,In_879);
and U1294 (N_1294,In_367,In_558);
nor U1295 (N_1295,In_51,In_1227);
nor U1296 (N_1296,In_868,In_1310);
nor U1297 (N_1297,In_1389,In_1044);
or U1298 (N_1298,In_965,In_59);
and U1299 (N_1299,In_684,In_917);
or U1300 (N_1300,In_766,In_1430);
nor U1301 (N_1301,In_1045,In_1388);
or U1302 (N_1302,In_75,In_1181);
and U1303 (N_1303,In_327,In_844);
or U1304 (N_1304,In_132,In_1220);
nor U1305 (N_1305,In_749,In_217);
nand U1306 (N_1306,In_1258,In_1380);
or U1307 (N_1307,In_1311,In_911);
nand U1308 (N_1308,In_302,In_592);
nand U1309 (N_1309,In_819,In_1329);
nor U1310 (N_1310,In_832,In_714);
nand U1311 (N_1311,In_702,In_619);
or U1312 (N_1312,In_1471,In_239);
nand U1313 (N_1313,In_1490,In_1085);
nand U1314 (N_1314,In_1011,In_462);
and U1315 (N_1315,In_647,In_745);
xor U1316 (N_1316,In_1459,In_26);
nor U1317 (N_1317,In_1020,In_991);
nand U1318 (N_1318,In_1032,In_300);
and U1319 (N_1319,In_581,In_633);
nor U1320 (N_1320,In_453,In_903);
and U1321 (N_1321,In_689,In_541);
or U1322 (N_1322,In_1412,In_872);
nor U1323 (N_1323,In_248,In_756);
nand U1324 (N_1324,In_177,In_1151);
nand U1325 (N_1325,In_846,In_410);
and U1326 (N_1326,In_404,In_906);
and U1327 (N_1327,In_471,In_995);
and U1328 (N_1328,In_314,In_1033);
nand U1329 (N_1329,In_1116,In_107);
and U1330 (N_1330,In_816,In_504);
nand U1331 (N_1331,In_837,In_886);
nor U1332 (N_1332,In_980,In_1036);
xnor U1333 (N_1333,In_1075,In_663);
nand U1334 (N_1334,In_1240,In_358);
and U1335 (N_1335,In_908,In_1250);
nand U1336 (N_1336,In_501,In_1426);
and U1337 (N_1337,In_101,In_1121);
or U1338 (N_1338,In_222,In_70);
nor U1339 (N_1339,In_674,In_1457);
nand U1340 (N_1340,In_676,In_1078);
nand U1341 (N_1341,In_1459,In_253);
and U1342 (N_1342,In_944,In_169);
nor U1343 (N_1343,In_1330,In_689);
and U1344 (N_1344,In_1270,In_70);
or U1345 (N_1345,In_471,In_1021);
or U1346 (N_1346,In_1036,In_1459);
nor U1347 (N_1347,In_1083,In_1054);
and U1348 (N_1348,In_748,In_887);
nand U1349 (N_1349,In_38,In_826);
nand U1350 (N_1350,In_229,In_1370);
nand U1351 (N_1351,In_937,In_1412);
and U1352 (N_1352,In_371,In_1023);
and U1353 (N_1353,In_1021,In_920);
and U1354 (N_1354,In_1105,In_180);
nor U1355 (N_1355,In_254,In_38);
or U1356 (N_1356,In_31,In_329);
and U1357 (N_1357,In_123,In_1090);
and U1358 (N_1358,In_779,In_460);
nand U1359 (N_1359,In_1371,In_1207);
and U1360 (N_1360,In_576,In_1413);
nand U1361 (N_1361,In_198,In_432);
nand U1362 (N_1362,In_1133,In_420);
and U1363 (N_1363,In_42,In_1379);
nor U1364 (N_1364,In_923,In_1435);
and U1365 (N_1365,In_1416,In_851);
and U1366 (N_1366,In_1136,In_452);
and U1367 (N_1367,In_351,In_1436);
xnor U1368 (N_1368,In_177,In_1185);
xnor U1369 (N_1369,In_632,In_1355);
nand U1370 (N_1370,In_913,In_563);
nor U1371 (N_1371,In_366,In_1017);
and U1372 (N_1372,In_729,In_256);
or U1373 (N_1373,In_1156,In_996);
nor U1374 (N_1374,In_1315,In_699);
nand U1375 (N_1375,In_135,In_1413);
and U1376 (N_1376,In_1346,In_285);
xnor U1377 (N_1377,In_556,In_202);
and U1378 (N_1378,In_809,In_883);
and U1379 (N_1379,In_565,In_936);
nor U1380 (N_1380,In_256,In_1064);
or U1381 (N_1381,In_952,In_1245);
nand U1382 (N_1382,In_702,In_116);
nor U1383 (N_1383,In_1148,In_325);
or U1384 (N_1384,In_650,In_449);
or U1385 (N_1385,In_1112,In_704);
nand U1386 (N_1386,In_112,In_1397);
nor U1387 (N_1387,In_651,In_480);
nand U1388 (N_1388,In_1144,In_33);
nor U1389 (N_1389,In_941,In_197);
or U1390 (N_1390,In_292,In_105);
or U1391 (N_1391,In_1421,In_571);
and U1392 (N_1392,In_1232,In_1223);
or U1393 (N_1393,In_669,In_218);
or U1394 (N_1394,In_1070,In_1083);
nand U1395 (N_1395,In_869,In_587);
nand U1396 (N_1396,In_664,In_320);
or U1397 (N_1397,In_402,In_1171);
or U1398 (N_1398,In_580,In_984);
nor U1399 (N_1399,In_1474,In_1122);
and U1400 (N_1400,In_1086,In_94);
nor U1401 (N_1401,In_27,In_1054);
and U1402 (N_1402,In_159,In_1351);
nand U1403 (N_1403,In_1410,In_858);
and U1404 (N_1404,In_1325,In_741);
or U1405 (N_1405,In_977,In_459);
nor U1406 (N_1406,In_621,In_804);
nor U1407 (N_1407,In_478,In_43);
nand U1408 (N_1408,In_1144,In_710);
nand U1409 (N_1409,In_751,In_1344);
nand U1410 (N_1410,In_126,In_557);
nor U1411 (N_1411,In_235,In_1331);
and U1412 (N_1412,In_985,In_255);
and U1413 (N_1413,In_407,In_1467);
or U1414 (N_1414,In_598,In_360);
and U1415 (N_1415,In_570,In_18);
nor U1416 (N_1416,In_170,In_1342);
nor U1417 (N_1417,In_1186,In_394);
or U1418 (N_1418,In_1055,In_855);
nand U1419 (N_1419,In_825,In_16);
and U1420 (N_1420,In_1225,In_1071);
or U1421 (N_1421,In_1110,In_517);
nor U1422 (N_1422,In_1429,In_72);
nor U1423 (N_1423,In_867,In_1216);
or U1424 (N_1424,In_552,In_453);
nand U1425 (N_1425,In_609,In_1480);
or U1426 (N_1426,In_1282,In_218);
and U1427 (N_1427,In_779,In_473);
nor U1428 (N_1428,In_603,In_1032);
and U1429 (N_1429,In_1491,In_99);
nand U1430 (N_1430,In_204,In_1060);
nor U1431 (N_1431,In_1474,In_1424);
nand U1432 (N_1432,In_1053,In_876);
and U1433 (N_1433,In_1375,In_1055);
nand U1434 (N_1434,In_601,In_747);
nor U1435 (N_1435,In_1384,In_1275);
nor U1436 (N_1436,In_899,In_1222);
and U1437 (N_1437,In_344,In_960);
and U1438 (N_1438,In_1071,In_656);
nand U1439 (N_1439,In_1429,In_80);
or U1440 (N_1440,In_992,In_1252);
nand U1441 (N_1441,In_1446,In_705);
or U1442 (N_1442,In_1064,In_1307);
or U1443 (N_1443,In_587,In_759);
nor U1444 (N_1444,In_1087,In_997);
or U1445 (N_1445,In_304,In_391);
nor U1446 (N_1446,In_633,In_691);
nor U1447 (N_1447,In_733,In_249);
and U1448 (N_1448,In_414,In_1126);
and U1449 (N_1449,In_1059,In_1339);
nand U1450 (N_1450,In_687,In_1204);
nand U1451 (N_1451,In_1178,In_1200);
nor U1452 (N_1452,In_330,In_157);
nand U1453 (N_1453,In_302,In_701);
or U1454 (N_1454,In_494,In_414);
or U1455 (N_1455,In_642,In_530);
nand U1456 (N_1456,In_359,In_701);
nand U1457 (N_1457,In_156,In_1137);
and U1458 (N_1458,In_196,In_1056);
nor U1459 (N_1459,In_900,In_774);
nand U1460 (N_1460,In_164,In_666);
nand U1461 (N_1461,In_913,In_226);
or U1462 (N_1462,In_807,In_1182);
nor U1463 (N_1463,In_425,In_1105);
or U1464 (N_1464,In_1431,In_1372);
nor U1465 (N_1465,In_345,In_165);
and U1466 (N_1466,In_1314,In_378);
nor U1467 (N_1467,In_576,In_11);
and U1468 (N_1468,In_1163,In_189);
nand U1469 (N_1469,In_1129,In_701);
and U1470 (N_1470,In_305,In_224);
and U1471 (N_1471,In_1448,In_924);
nor U1472 (N_1472,In_818,In_8);
nand U1473 (N_1473,In_723,In_306);
nor U1474 (N_1474,In_514,In_669);
nor U1475 (N_1475,In_1391,In_1255);
and U1476 (N_1476,In_738,In_624);
nor U1477 (N_1477,In_1248,In_313);
and U1478 (N_1478,In_24,In_257);
or U1479 (N_1479,In_585,In_818);
nand U1480 (N_1480,In_315,In_52);
and U1481 (N_1481,In_219,In_338);
or U1482 (N_1482,In_545,In_22);
nand U1483 (N_1483,In_283,In_1349);
nor U1484 (N_1484,In_1031,In_932);
nand U1485 (N_1485,In_778,In_280);
or U1486 (N_1486,In_660,In_808);
and U1487 (N_1487,In_24,In_539);
or U1488 (N_1488,In_662,In_747);
or U1489 (N_1489,In_410,In_352);
nand U1490 (N_1490,In_578,In_1358);
or U1491 (N_1491,In_1218,In_1386);
xnor U1492 (N_1492,In_328,In_962);
or U1493 (N_1493,In_1112,In_817);
nor U1494 (N_1494,In_196,In_974);
or U1495 (N_1495,In_1202,In_1339);
nand U1496 (N_1496,In_1450,In_754);
xor U1497 (N_1497,In_1004,In_67);
or U1498 (N_1498,In_570,In_79);
nor U1499 (N_1499,In_1155,In_1399);
or U1500 (N_1500,N_758,N_1119);
xor U1501 (N_1501,N_514,N_513);
or U1502 (N_1502,N_831,N_823);
nor U1503 (N_1503,N_90,N_439);
or U1504 (N_1504,N_176,N_1376);
nor U1505 (N_1505,N_685,N_129);
and U1506 (N_1506,N_1308,N_759);
nor U1507 (N_1507,N_338,N_869);
or U1508 (N_1508,N_207,N_1325);
or U1509 (N_1509,N_952,N_447);
or U1510 (N_1510,N_1421,N_433);
nor U1511 (N_1511,N_1480,N_194);
or U1512 (N_1512,N_1171,N_102);
nor U1513 (N_1513,N_246,N_1476);
and U1514 (N_1514,N_1197,N_897);
or U1515 (N_1515,N_9,N_1299);
and U1516 (N_1516,N_566,N_130);
nor U1517 (N_1517,N_645,N_390);
and U1518 (N_1518,N_879,N_943);
nor U1519 (N_1519,N_419,N_260);
nand U1520 (N_1520,N_35,N_697);
nand U1521 (N_1521,N_158,N_1047);
nor U1522 (N_1522,N_1234,N_522);
and U1523 (N_1523,N_767,N_898);
nor U1524 (N_1524,N_1058,N_383);
and U1525 (N_1525,N_425,N_1442);
or U1526 (N_1526,N_1305,N_1387);
and U1527 (N_1527,N_935,N_393);
or U1528 (N_1528,N_545,N_1464);
nor U1529 (N_1529,N_1160,N_405);
or U1530 (N_1530,N_1366,N_934);
or U1531 (N_1531,N_661,N_1200);
nand U1532 (N_1532,N_1333,N_403);
nand U1533 (N_1533,N_615,N_624);
nand U1534 (N_1534,N_1302,N_786);
and U1535 (N_1535,N_1151,N_820);
and U1536 (N_1536,N_472,N_272);
or U1537 (N_1537,N_1395,N_12);
or U1538 (N_1538,N_1493,N_13);
nand U1539 (N_1539,N_1105,N_917);
and U1540 (N_1540,N_722,N_1056);
nor U1541 (N_1541,N_332,N_822);
and U1542 (N_1542,N_835,N_372);
or U1543 (N_1543,N_836,N_427);
and U1544 (N_1544,N_610,N_254);
or U1545 (N_1545,N_1154,N_66);
or U1546 (N_1546,N_1273,N_313);
and U1547 (N_1547,N_475,N_293);
or U1548 (N_1548,N_280,N_595);
nand U1549 (N_1549,N_154,N_817);
nor U1550 (N_1550,N_891,N_551);
nand U1551 (N_1551,N_388,N_8);
or U1552 (N_1552,N_204,N_1436);
nand U1553 (N_1553,N_798,N_533);
or U1554 (N_1554,N_1009,N_818);
nand U1555 (N_1555,N_213,N_371);
nand U1556 (N_1556,N_357,N_1059);
and U1557 (N_1557,N_308,N_165);
and U1558 (N_1558,N_1069,N_97);
or U1559 (N_1559,N_436,N_1022);
or U1560 (N_1560,N_1332,N_775);
and U1561 (N_1561,N_572,N_1445);
nand U1562 (N_1562,N_537,N_1142);
nor U1563 (N_1563,N_67,N_1145);
nand U1564 (N_1564,N_1351,N_755);
nand U1565 (N_1565,N_670,N_988);
and U1566 (N_1566,N_1092,N_501);
nand U1567 (N_1567,N_3,N_1391);
and U1568 (N_1568,N_875,N_957);
xor U1569 (N_1569,N_1446,N_139);
and U1570 (N_1570,N_909,N_143);
nand U1571 (N_1571,N_657,N_526);
or U1572 (N_1572,N_1244,N_951);
or U1573 (N_1573,N_50,N_1348);
nand U1574 (N_1574,N_1250,N_886);
nand U1575 (N_1575,N_1318,N_834);
and U1576 (N_1576,N_1206,N_655);
or U1577 (N_1577,N_772,N_719);
or U1578 (N_1578,N_922,N_1497);
or U1579 (N_1579,N_453,N_1329);
nand U1580 (N_1580,N_350,N_429);
and U1581 (N_1581,N_1282,N_1124);
nor U1582 (N_1582,N_521,N_733);
or U1583 (N_1583,N_1122,N_1107);
nor U1584 (N_1584,N_737,N_1423);
and U1585 (N_1585,N_166,N_679);
nand U1586 (N_1586,N_531,N_747);
and U1587 (N_1587,N_738,N_980);
nand U1588 (N_1588,N_1357,N_1323);
nand U1589 (N_1589,N_1035,N_1134);
nor U1590 (N_1590,N_1456,N_696);
or U1591 (N_1591,N_333,N_250);
and U1592 (N_1592,N_170,N_445);
or U1593 (N_1593,N_1027,N_1211);
or U1594 (N_1594,N_1071,N_451);
nor U1595 (N_1595,N_349,N_159);
xor U1596 (N_1596,N_358,N_412);
or U1597 (N_1597,N_832,N_860);
nand U1598 (N_1598,N_1355,N_274);
or U1599 (N_1599,N_795,N_884);
or U1600 (N_1600,N_420,N_1088);
nand U1601 (N_1601,N_1147,N_219);
or U1602 (N_1602,N_60,N_1219);
or U1603 (N_1603,N_1496,N_226);
nand U1604 (N_1604,N_268,N_725);
or U1605 (N_1605,N_712,N_689);
nor U1606 (N_1606,N_1188,N_112);
and U1607 (N_1607,N_386,N_1430);
nor U1608 (N_1608,N_1065,N_962);
and U1609 (N_1609,N_637,N_1396);
or U1610 (N_1610,N_450,N_981);
nor U1611 (N_1611,N_629,N_1326);
or U1612 (N_1612,N_597,N_257);
and U1613 (N_1613,N_669,N_931);
nand U1614 (N_1614,N_216,N_906);
and U1615 (N_1615,N_62,N_203);
and U1616 (N_1616,N_651,N_1283);
and U1617 (N_1617,N_295,N_585);
and U1618 (N_1618,N_296,N_476);
nor U1619 (N_1619,N_867,N_125);
or U1620 (N_1620,N_653,N_286);
nor U1621 (N_1621,N_106,N_530);
xnor U1622 (N_1622,N_1010,N_1169);
or U1623 (N_1623,N_664,N_298);
and U1624 (N_1624,N_438,N_1070);
xnor U1625 (N_1625,N_155,N_830);
nor U1626 (N_1626,N_381,N_242);
and U1627 (N_1627,N_821,N_1440);
nor U1628 (N_1628,N_1401,N_631);
nor U1629 (N_1629,N_1094,N_810);
nand U1630 (N_1630,N_1472,N_1485);
nor U1631 (N_1631,N_1291,N_1370);
nor U1632 (N_1632,N_168,N_1157);
nor U1633 (N_1633,N_1279,N_83);
or U1634 (N_1634,N_456,N_676);
or U1635 (N_1635,N_948,N_31);
or U1636 (N_1636,N_1265,N_1461);
nor U1637 (N_1637,N_1,N_471);
nand U1638 (N_1638,N_968,N_1300);
or U1639 (N_1639,N_986,N_1490);
nand U1640 (N_1640,N_64,N_1458);
nand U1641 (N_1641,N_1448,N_1191);
and U1642 (N_1642,N_464,N_1114);
nor U1643 (N_1643,N_1095,N_893);
and U1644 (N_1644,N_605,N_763);
or U1645 (N_1645,N_1139,N_147);
and U1646 (N_1646,N_1252,N_10);
nor U1647 (N_1647,N_1249,N_434);
or U1648 (N_1648,N_138,N_237);
nand U1649 (N_1649,N_145,N_959);
xor U1650 (N_1650,N_728,N_1083);
nor U1651 (N_1651,N_1465,N_870);
and U1652 (N_1652,N_105,N_984);
nor U1653 (N_1653,N_1342,N_69);
or U1654 (N_1654,N_1123,N_735);
nor U1655 (N_1655,N_1315,N_500);
or U1656 (N_1656,N_1264,N_1328);
and U1657 (N_1657,N_1150,N_355);
nand U1658 (N_1658,N_1133,N_424);
and U1659 (N_1659,N_838,N_694);
nand U1660 (N_1660,N_61,N_1061);
nand U1661 (N_1661,N_269,N_1138);
and U1662 (N_1662,N_187,N_1416);
and U1663 (N_1663,N_19,N_826);
or U1664 (N_1664,N_292,N_1052);
nand U1665 (N_1665,N_325,N_520);
and U1666 (N_1666,N_1141,N_1316);
or U1667 (N_1667,N_1180,N_1426);
or U1668 (N_1668,N_290,N_1382);
and U1669 (N_1669,N_271,N_604);
and U1670 (N_1670,N_320,N_947);
and U1671 (N_1671,N_532,N_185);
nor U1672 (N_1672,N_792,N_252);
nand U1673 (N_1673,N_1284,N_1477);
or U1674 (N_1674,N_880,N_770);
or U1675 (N_1675,N_787,N_152);
and U1676 (N_1676,N_76,N_360);
nor U1677 (N_1677,N_58,N_568);
nor U1678 (N_1678,N_496,N_273);
nand U1679 (N_1679,N_1335,N_930);
nand U1680 (N_1680,N_233,N_4);
nor U1681 (N_1681,N_1251,N_977);
or U1682 (N_1682,N_748,N_720);
nor U1683 (N_1683,N_394,N_100);
or U1684 (N_1684,N_814,N_294);
and U1685 (N_1685,N_1106,N_938);
or U1686 (N_1686,N_1002,N_137);
nand U1687 (N_1687,N_169,N_1199);
nand U1688 (N_1688,N_970,N_921);
nand U1689 (N_1689,N_1137,N_1347);
or U1690 (N_1690,N_1384,N_515);
nand U1691 (N_1691,N_599,N_583);
nor U1692 (N_1692,N_723,N_994);
nand U1693 (N_1693,N_443,N_1079);
or U1694 (N_1694,N_779,N_861);
and U1695 (N_1695,N_151,N_1008);
or U1696 (N_1696,N_318,N_417);
and U1697 (N_1697,N_908,N_1155);
nor U1698 (N_1698,N_1406,N_741);
nand U1699 (N_1699,N_77,N_1334);
nor U1700 (N_1700,N_606,N_956);
or U1701 (N_1701,N_511,N_55);
nand U1702 (N_1702,N_781,N_1034);
or U1703 (N_1703,N_641,N_841);
nor U1704 (N_1704,N_1025,N_1038);
nand U1705 (N_1705,N_1098,N_1407);
nor U1706 (N_1706,N_201,N_240);
xor U1707 (N_1707,N_542,N_672);
nor U1708 (N_1708,N_400,N_74);
nand U1709 (N_1709,N_756,N_580);
nor U1710 (N_1710,N_1209,N_1452);
and U1711 (N_1711,N_1467,N_714);
nand U1712 (N_1712,N_239,N_704);
nand U1713 (N_1713,N_1078,N_1310);
nand U1714 (N_1714,N_275,N_391);
xor U1715 (N_1715,N_1181,N_1004);
or U1716 (N_1716,N_430,N_866);
nor U1717 (N_1717,N_684,N_1365);
and U1718 (N_1718,N_745,N_251);
nand U1719 (N_1719,N_656,N_1166);
and U1720 (N_1720,N_1330,N_750);
nor U1721 (N_1721,N_964,N_739);
nor U1722 (N_1722,N_340,N_560);
nand U1723 (N_1723,N_309,N_706);
nand U1724 (N_1724,N_768,N_1450);
nand U1725 (N_1725,N_634,N_113);
and U1726 (N_1726,N_1296,N_1463);
nor U1727 (N_1727,N_474,N_71);
and U1728 (N_1728,N_1232,N_470);
nor U1729 (N_1729,N_985,N_1015);
nor U1730 (N_1730,N_721,N_1451);
nor U1731 (N_1731,N_107,N_161);
xor U1732 (N_1732,N_534,N_1156);
and U1733 (N_1733,N_997,N_173);
or U1734 (N_1734,N_746,N_63);
nand U1735 (N_1735,N_398,N_270);
nor U1736 (N_1736,N_912,N_699);
and U1737 (N_1737,N_1491,N_1297);
nand U1738 (N_1738,N_713,N_375);
nand U1739 (N_1739,N_644,N_1431);
nor U1740 (N_1740,N_322,N_849);
or U1741 (N_1741,N_1163,N_224);
nor U1742 (N_1742,N_794,N_498);
nand U1743 (N_1743,N_128,N_1205);
and U1744 (N_1744,N_1410,N_323);
or U1745 (N_1745,N_1322,N_1483);
nor U1746 (N_1746,N_282,N_801);
nor U1747 (N_1747,N_353,N_602);
or U1748 (N_1748,N_1120,N_705);
or U1749 (N_1749,N_1457,N_1019);
or U1750 (N_1750,N_1220,N_15);
or U1751 (N_1751,N_1267,N_691);
nand U1752 (N_1752,N_1230,N_762);
and U1753 (N_1753,N_1076,N_14);
or U1754 (N_1754,N_111,N_379);
and U1755 (N_1755,N_1146,N_234);
nand U1756 (N_1756,N_68,N_1268);
nor U1757 (N_1757,N_1313,N_199);
or U1758 (N_1758,N_592,N_1104);
or U1759 (N_1759,N_1195,N_1100);
or U1760 (N_1760,N_1112,N_1039);
nor U1761 (N_1761,N_1374,N_843);
or U1762 (N_1762,N_180,N_518);
nor U1763 (N_1763,N_965,N_600);
nand U1764 (N_1764,N_1240,N_579);
and U1765 (N_1765,N_42,N_1287);
nand U1766 (N_1766,N_487,N_20);
nand U1767 (N_1767,N_547,N_612);
or U1768 (N_1768,N_1193,N_1375);
and U1769 (N_1769,N_1215,N_1184);
or U1770 (N_1770,N_1016,N_743);
xnor U1771 (N_1771,N_575,N_958);
nand U1772 (N_1772,N_1275,N_478);
and U1773 (N_1773,N_347,N_1482);
nor U1774 (N_1774,N_718,N_556);
or U1775 (N_1775,N_437,N_700);
nand U1776 (N_1776,N_206,N_1050);
and U1777 (N_1777,N_837,N_1398);
xor U1778 (N_1778,N_1201,N_1454);
and U1779 (N_1779,N_611,N_6);
and U1780 (N_1780,N_567,N_562);
or U1781 (N_1781,N_109,N_517);
nor U1782 (N_1782,N_716,N_57);
and U1783 (N_1783,N_1340,N_244);
nand U1784 (N_1784,N_804,N_172);
or U1785 (N_1785,N_217,N_882);
nand U1786 (N_1786,N_131,N_1425);
and U1787 (N_1787,N_2,N_1102);
and U1788 (N_1788,N_119,N_829);
and U1789 (N_1789,N_466,N_724);
or U1790 (N_1790,N_1143,N_380);
nor U1791 (N_1791,N_785,N_1412);
or U1792 (N_1792,N_460,N_382);
nand U1793 (N_1793,N_569,N_1295);
nand U1794 (N_1794,N_319,N_1379);
nor U1795 (N_1795,N_1372,N_284);
nand U1796 (N_1796,N_305,N_334);
nand U1797 (N_1797,N_1130,N_732);
and U1798 (N_1798,N_1363,N_782);
or U1799 (N_1799,N_1017,N_457);
or U1800 (N_1800,N_499,N_1129);
xor U1801 (N_1801,N_1435,N_1177);
and U1802 (N_1802,N_396,N_734);
or U1803 (N_1803,N_1285,N_1449);
nor U1804 (N_1804,N_626,N_1392);
nand U1805 (N_1805,N_30,N_540);
nor U1806 (N_1806,N_202,N_1337);
nor U1807 (N_1807,N_596,N_1224);
nand U1808 (N_1808,N_1368,N_682);
nor U1809 (N_1809,N_619,N_571);
and U1810 (N_1810,N_459,N_955);
and U1811 (N_1811,N_426,N_374);
and U1812 (N_1812,N_625,N_266);
and U1813 (N_1813,N_1266,N_1236);
and U1814 (N_1814,N_285,N_730);
nand U1815 (N_1815,N_1087,N_1116);
and U1816 (N_1816,N_1272,N_847);
or U1817 (N_1817,N_442,N_223);
nor U1818 (N_1818,N_842,N_942);
and U1819 (N_1819,N_1229,N_840);
or U1820 (N_1820,N_197,N_186);
or U1821 (N_1821,N_1460,N_850);
or U1822 (N_1822,N_1045,N_1255);
or U1823 (N_1823,N_409,N_265);
nand U1824 (N_1824,N_805,N_777);
nand U1825 (N_1825,N_707,N_1064);
nor U1826 (N_1826,N_1301,N_407);
nand U1827 (N_1827,N_1020,N_1073);
and U1828 (N_1828,N_34,N_797);
and U1829 (N_1829,N_321,N_1269);
and U1830 (N_1830,N_554,N_1090);
and U1831 (N_1831,N_1060,N_878);
and U1832 (N_1832,N_636,N_330);
and U1833 (N_1833,N_370,N_281);
nand U1834 (N_1834,N_377,N_608);
and U1835 (N_1835,N_923,N_497);
and U1836 (N_1836,N_780,N_489);
or U1837 (N_1837,N_278,N_961);
xor U1838 (N_1838,N_565,N_1400);
and U1839 (N_1839,N_488,N_1492);
nand U1840 (N_1840,N_505,N_78);
or U1841 (N_1841,N_1207,N_70);
and U1842 (N_1842,N_819,N_259);
and U1843 (N_1843,N_261,N_1063);
or U1844 (N_1844,N_1099,N_757);
and U1845 (N_1845,N_493,N_1210);
nand U1846 (N_1846,N_874,N_877);
or U1847 (N_1847,N_473,N_1128);
and U1848 (N_1848,N_1377,N_1189);
nor U1849 (N_1849,N_1053,N_621);
xor U1850 (N_1850,N_364,N_276);
nor U1851 (N_1851,N_1317,N_399);
or U1852 (N_1852,N_616,N_905);
and U1853 (N_1853,N_88,N_751);
nand U1854 (N_1854,N_133,N_647);
nand U1855 (N_1855,N_94,N_7);
nor U1856 (N_1856,N_245,N_969);
nor U1857 (N_1857,N_648,N_277);
nor U1858 (N_1858,N_315,N_235);
nand U1859 (N_1859,N_29,N_573);
nor U1860 (N_1860,N_38,N_925);
nor U1861 (N_1861,N_75,N_465);
and U1862 (N_1862,N_788,N_121);
xnor U1863 (N_1863,N_279,N_535);
nor U1864 (N_1864,N_1049,N_528);
and U1865 (N_1865,N_431,N_96);
nor U1866 (N_1866,N_1204,N_731);
nand U1867 (N_1867,N_300,N_736);
or U1868 (N_1868,N_1242,N_632);
or U1869 (N_1869,N_123,N_116);
and U1870 (N_1870,N_1218,N_126);
or U1871 (N_1871,N_1289,N_22);
nor U1872 (N_1872,N_1380,N_667);
and U1873 (N_1873,N_978,N_1003);
nor U1874 (N_1874,N_548,N_435);
or U1875 (N_1875,N_304,N_359);
and U1876 (N_1876,N_1031,N_26);
and U1877 (N_1877,N_1489,N_559);
and U1878 (N_1878,N_895,N_901);
nand U1879 (N_1879,N_802,N_53);
nand U1880 (N_1880,N_711,N_449);
or U1881 (N_1881,N_576,N_108);
and U1882 (N_1882,N_854,N_885);
nor U1883 (N_1883,N_492,N_1286);
nor U1884 (N_1884,N_41,N_81);
nand U1885 (N_1885,N_727,N_114);
and U1886 (N_1886,N_24,N_638);
nand U1887 (N_1887,N_52,N_715);
and U1888 (N_1888,N_337,N_85);
nand U1889 (N_1889,N_136,N_791);
nor U1890 (N_1890,N_1277,N_665);
nand U1891 (N_1891,N_1126,N_506);
or U1892 (N_1892,N_509,N_228);
and U1893 (N_1893,N_1466,N_156);
and U1894 (N_1894,N_510,N_1074);
or U1895 (N_1895,N_916,N_1422);
nor U1896 (N_1896,N_1292,N_650);
or U1897 (N_1897,N_120,N_222);
and U1898 (N_1898,N_927,N_1113);
nor U1899 (N_1899,N_37,N_1263);
nor U1900 (N_1900,N_402,N_1388);
and U1901 (N_1901,N_799,N_1051);
nor U1902 (N_1902,N_1280,N_454);
and U1903 (N_1903,N_141,N_5);
nor U1904 (N_1904,N_1077,N_1159);
and U1905 (N_1905,N_163,N_1399);
nor U1906 (N_1906,N_844,N_765);
nor U1907 (N_1907,N_1228,N_541);
xor U1908 (N_1908,N_783,N_144);
nand U1909 (N_1909,N_32,N_1080);
or U1910 (N_1910,N_378,N_1178);
or U1911 (N_1911,N_701,N_243);
or U1912 (N_1912,N_79,N_1418);
nand U1913 (N_1913,N_945,N_477);
nor U1914 (N_1914,N_179,N_1420);
nor U1915 (N_1915,N_1203,N_1468);
or U1916 (N_1916,N_1254,N_502);
and U1917 (N_1917,N_744,N_51);
and U1918 (N_1918,N_343,N_1024);
nor U1919 (N_1919,N_1311,N_729);
nor U1920 (N_1920,N_190,N_418);
nand U1921 (N_1921,N_690,N_848);
nand U1922 (N_1922,N_950,N_348);
nand U1923 (N_1923,N_184,N_803);
or U1924 (N_1924,N_1344,N_949);
nand U1925 (N_1925,N_1135,N_618);
or U1926 (N_1926,N_1241,N_221);
nand U1927 (N_1927,N_494,N_577);
nand U1928 (N_1928,N_341,N_793);
or U1929 (N_1929,N_452,N_1350);
or U1930 (N_1930,N_479,N_1258);
nor U1931 (N_1931,N_1028,N_944);
and U1932 (N_1932,N_709,N_483);
and U1933 (N_1933,N_1167,N_584);
and U1934 (N_1934,N_157,N_188);
xor U1935 (N_1935,N_110,N_181);
nor U1936 (N_1936,N_671,N_1213);
and U1937 (N_1937,N_633,N_262);
or U1938 (N_1938,N_1131,N_996);
or U1939 (N_1939,N_1081,N_303);
or U1940 (N_1940,N_845,N_1136);
or U1941 (N_1941,N_95,N_507);
and U1942 (N_1942,N_1115,N_1041);
nor U1943 (N_1943,N_642,N_73);
xor U1944 (N_1944,N_317,N_1443);
nor U1945 (N_1945,N_1362,N_1474);
nand U1946 (N_1946,N_189,N_1462);
and U1947 (N_1947,N_103,N_1349);
and U1948 (N_1948,N_1110,N_873);
nor U1949 (N_1949,N_1037,N_512);
or U1950 (N_1950,N_966,N_859);
or U1951 (N_1951,N_56,N_1498);
nor U1952 (N_1952,N_1026,N_552);
and U1953 (N_1953,N_856,N_1021);
and U1954 (N_1954,N_1470,N_857);
or U1955 (N_1955,N_198,N_227);
and U1956 (N_1956,N_919,N_1226);
nand U1957 (N_1957,N_570,N_915);
xor U1958 (N_1958,N_824,N_708);
and U1959 (N_1959,N_387,N_212);
nand U1960 (N_1960,N_327,N_852);
and U1961 (N_1961,N_134,N_191);
nand U1962 (N_1962,N_59,N_1320);
and U1963 (N_1963,N_900,N_40);
nand U1964 (N_1964,N_283,N_862);
nand U1965 (N_1965,N_306,N_193);
nand U1966 (N_1966,N_1162,N_808);
nor U1967 (N_1967,N_331,N_1486);
nand U1968 (N_1968,N_140,N_833);
nand U1969 (N_1969,N_1262,N_481);
or U1970 (N_1970,N_432,N_1394);
and U1971 (N_1971,N_609,N_1152);
and U1972 (N_1972,N_1086,N_356);
or U1973 (N_1973,N_630,N_33);
or U1974 (N_1974,N_316,N_503);
nand U1975 (N_1975,N_1455,N_1271);
nand U1976 (N_1976,N_1165,N_1438);
nor U1977 (N_1977,N_1014,N_603);
or U1978 (N_1978,N_858,N_749);
nand U1979 (N_1979,N_816,N_345);
nor U1980 (N_1980,N_1404,N_1075);
nor U1981 (N_1981,N_346,N_1040);
nand U1982 (N_1982,N_1298,N_992);
nor U1983 (N_1983,N_504,N_1192);
nor U1984 (N_1984,N_581,N_192);
nor U1985 (N_1985,N_907,N_18);
and U1986 (N_1986,N_936,N_635);
nand U1987 (N_1987,N_48,N_414);
and U1988 (N_1988,N_1386,N_310);
nand U1989 (N_1989,N_1274,N_1190);
or U1990 (N_1990,N_200,N_1231);
nor U1991 (N_1991,N_622,N_389);
and U1992 (N_1992,N_1371,N_1354);
nor U1993 (N_1993,N_839,N_594);
or U1994 (N_1994,N_241,N_1182);
or U1995 (N_1995,N_1411,N_238);
nand U1996 (N_1996,N_659,N_529);
nand U1997 (N_1997,N_1185,N_983);
or U1998 (N_1998,N_1381,N_1259);
nand U1999 (N_1999,N_1005,N_1304);
nand U2000 (N_2000,N_654,N_918);
nand U2001 (N_2001,N_369,N_1243);
nor U2002 (N_2002,N_446,N_1402);
or U2003 (N_2003,N_307,N_1144);
nor U2004 (N_2004,N_1246,N_267);
nand U2005 (N_2005,N_686,N_778);
and U2006 (N_2006,N_1082,N_1356);
nand U2007 (N_2007,N_46,N_693);
or U2008 (N_2008,N_553,N_1453);
and U2009 (N_2009,N_1108,N_1029);
or U2010 (N_2010,N_1012,N_1390);
nor U2011 (N_2011,N_1186,N_21);
or U2012 (N_2012,N_710,N_827);
nor U2013 (N_2013,N_1288,N_543);
nand U2014 (N_2014,N_43,N_146);
and U2015 (N_2015,N_752,N_361);
or U2016 (N_2016,N_1125,N_45);
and U2017 (N_2017,N_160,N_963);
or U2018 (N_2018,N_695,N_301);
or U2019 (N_2019,N_1208,N_591);
nor U2020 (N_2020,N_467,N_1013);
and U2021 (N_2021,N_544,N_411);
nor U2022 (N_2022,N_491,N_27);
or U2023 (N_2023,N_1358,N_678);
nand U2024 (N_2024,N_1383,N_555);
xor U2025 (N_2025,N_1321,N_336);
nor U2026 (N_2026,N_1089,N_84);
and U2027 (N_2027,N_1360,N_872);
nand U2028 (N_2028,N_1212,N_1281);
nand U2029 (N_2029,N_1495,N_539);
nand U2030 (N_2030,N_1117,N_65);
and U2031 (N_2031,N_1033,N_972);
or U2032 (N_2032,N_1161,N_178);
nand U2033 (N_2033,N_776,N_1444);
or U2034 (N_2034,N_516,N_1196);
or U2035 (N_2035,N_1173,N_463);
nor U2036 (N_2036,N_404,N_1307);
or U2037 (N_2037,N_1023,N_1164);
nor U2038 (N_2038,N_894,N_1433);
nand U2039 (N_2039,N_167,N_1256);
and U2040 (N_2040,N_607,N_883);
nand U2041 (N_2041,N_1109,N_329);
and U2042 (N_2042,N_789,N_851);
or U2043 (N_2043,N_586,N_1097);
nor U2044 (N_2044,N_1378,N_311);
nor U2045 (N_2045,N_589,N_876);
nand U2046 (N_2046,N_366,N_210);
nor U2047 (N_2047,N_99,N_326);
or U2048 (N_2048,N_1221,N_211);
and U2049 (N_2049,N_214,N_1397);
or U2050 (N_2050,N_519,N_726);
nor U2051 (N_2051,N_920,N_1174);
nor U2052 (N_2052,N_790,N_954);
and U2053 (N_2053,N_889,N_288);
and U2054 (N_2054,N_253,N_263);
nand U2055 (N_2055,N_1132,N_1409);
or U2056 (N_2056,N_177,N_601);
nor U2057 (N_2057,N_771,N_127);
and U2058 (N_2058,N_220,N_225);
nor U2059 (N_2059,N_312,N_54);
nand U2060 (N_2060,N_769,N_546);
nand U2061 (N_2061,N_1447,N_205);
nand U2062 (N_2062,N_1046,N_423);
or U2063 (N_2063,N_468,N_1385);
nand U2064 (N_2064,N_1149,N_122);
nor U2065 (N_2065,N_287,N_881);
nor U2066 (N_2066,N_392,N_124);
nand U2067 (N_2067,N_1172,N_564);
nand U2068 (N_2068,N_1168,N_742);
or U2069 (N_2069,N_484,N_1260);
and U2070 (N_2070,N_28,N_1176);
or U2071 (N_2071,N_1158,N_914);
or U2072 (N_2072,N_617,N_926);
nand U2073 (N_2073,N_1237,N_1217);
nand U2074 (N_2074,N_1343,N_865);
and U2075 (N_2075,N_218,N_395);
and U2076 (N_2076,N_1091,N_523);
and U2077 (N_2077,N_36,N_643);
or U2078 (N_2078,N_646,N_1441);
or U2079 (N_2079,N_448,N_373);
and U2080 (N_2080,N_384,N_1413);
nand U2081 (N_2081,N_117,N_673);
or U2082 (N_2082,N_328,N_297);
nor U2083 (N_2083,N_774,N_132);
nor U2084 (N_2084,N_153,N_939);
nand U2085 (N_2085,N_230,N_118);
nor U2086 (N_2086,N_688,N_215);
nand U2087 (N_2087,N_1484,N_461);
nor U2088 (N_2088,N_764,N_1000);
nand U2089 (N_2089,N_1499,N_1479);
and U2090 (N_2090,N_1175,N_365);
or U2091 (N_2091,N_974,N_162);
and U2092 (N_2092,N_1306,N_385);
or U2093 (N_2093,N_335,N_932);
or U2094 (N_2094,N_937,N_1032);
or U2095 (N_2095,N_1290,N_1488);
nand U2096 (N_2096,N_904,N_104);
and U2097 (N_2097,N_993,N_998);
nand U2098 (N_2098,N_164,N_209);
nand U2099 (N_2099,N_462,N_853);
nor U2100 (N_2100,N_975,N_1253);
nor U2101 (N_2101,N_652,N_549);
xor U2102 (N_2102,N_761,N_590);
nor U2103 (N_2103,N_1345,N_482);
nor U2104 (N_2104,N_681,N_1216);
nand U2105 (N_2105,N_613,N_753);
and U2106 (N_2106,N_910,N_1369);
and U2107 (N_2107,N_1294,N_809);
nor U2108 (N_2108,N_1352,N_929);
and U2109 (N_2109,N_960,N_588);
nand U2110 (N_2110,N_911,N_1238);
nor U2111 (N_2111,N_813,N_784);
nand U2112 (N_2112,N_229,N_890);
and U2113 (N_2113,N_1361,N_620);
nand U2114 (N_2114,N_558,N_1202);
or U2115 (N_2115,N_413,N_864);
or U2116 (N_2116,N_871,N_1338);
nor U2117 (N_2117,N_903,N_1153);
nor U2118 (N_2118,N_1270,N_1339);
and U2119 (N_2119,N_362,N_415);
nand U2120 (N_2120,N_1373,N_773);
and U2121 (N_2121,N_444,N_39);
and U2122 (N_2122,N_687,N_1011);
nand U2123 (N_2123,N_410,N_98);
nand U2124 (N_2124,N_89,N_538);
nor U2125 (N_2125,N_289,N_351);
or U2126 (N_2126,N_677,N_563);
and U2127 (N_2127,N_249,N_740);
nor U2128 (N_2128,N_1353,N_93);
nor U2129 (N_2129,N_1324,N_663);
or U2130 (N_2130,N_800,N_662);
and U2131 (N_2131,N_1225,N_339);
nor U2132 (N_2132,N_324,N_1140);
or U2133 (N_2133,N_899,N_1432);
or U2134 (N_2134,N_208,N_11);
and U2135 (N_2135,N_582,N_416);
nand U2136 (N_2136,N_1428,N_698);
xor U2137 (N_2137,N_80,N_1096);
or U2138 (N_2138,N_1183,N_1405);
or U2139 (N_2139,N_928,N_25);
nor U2140 (N_2140,N_490,N_1101);
and U2141 (N_2141,N_1437,N_1314);
nand U2142 (N_2142,N_527,N_23);
and U2143 (N_2143,N_999,N_668);
nand U2144 (N_2144,N_587,N_196);
and U2145 (N_2145,N_264,N_376);
xnor U2146 (N_2146,N_760,N_902);
and U2147 (N_2147,N_593,N_485);
or U2148 (N_2148,N_17,N_195);
nand U2149 (N_2149,N_982,N_486);
nand U2150 (N_2150,N_1415,N_1393);
or U2151 (N_2151,N_754,N_422);
nor U2152 (N_2152,N_258,N_1414);
or U2153 (N_2153,N_1331,N_987);
and U2154 (N_2154,N_674,N_408);
and U2155 (N_2155,N_933,N_967);
or U2156 (N_2156,N_255,N_469);
or U2157 (N_2157,N_888,N_990);
nand U2158 (N_2158,N_232,N_354);
nor U2159 (N_2159,N_807,N_495);
nor U2160 (N_2160,N_1245,N_550);
or U2161 (N_2161,N_913,N_639);
and U2162 (N_2162,N_149,N_680);
and U2163 (N_2163,N_989,N_946);
nor U2164 (N_2164,N_1062,N_973);
nand U2165 (N_2165,N_561,N_623);
and U2166 (N_2166,N_302,N_1118);
and U2167 (N_2167,N_557,N_150);
nand U2168 (N_2168,N_1359,N_455);
nand U2169 (N_2169,N_142,N_1036);
xnor U2170 (N_2170,N_525,N_1067);
or U2171 (N_2171,N_811,N_1233);
and U2172 (N_2172,N_868,N_47);
and U2173 (N_2173,N_1248,N_1473);
or U2174 (N_2174,N_941,N_855);
or U2175 (N_2175,N_896,N_1194);
or U2176 (N_2176,N_815,N_649);
nor U2177 (N_2177,N_508,N_1247);
nor U2178 (N_2178,N_995,N_666);
and U2179 (N_2179,N_766,N_1001);
nor U2180 (N_2180,N_1478,N_1346);
and U2181 (N_2181,N_1068,N_1487);
or U2182 (N_2182,N_1429,N_135);
nor U2183 (N_2183,N_406,N_578);
nand U2184 (N_2184,N_344,N_1481);
nor U2185 (N_2185,N_1475,N_248);
nand U2186 (N_2186,N_627,N_1319);
or U2187 (N_2187,N_1419,N_1309);
nand U2188 (N_2188,N_614,N_536);
or U2189 (N_2189,N_0,N_812);
nor U2190 (N_2190,N_1018,N_660);
or U2191 (N_2191,N_1121,N_1367);
and U2192 (N_2192,N_1471,N_675);
or U2193 (N_2193,N_367,N_1222);
and U2194 (N_2194,N_91,N_806);
or U2195 (N_2195,N_401,N_1148);
and U2196 (N_2196,N_887,N_702);
nand U2197 (N_2197,N_1048,N_1469);
and U2198 (N_2198,N_658,N_16);
nand U2199 (N_2199,N_1111,N_1030);
or U2200 (N_2200,N_828,N_1494);
and U2201 (N_2201,N_171,N_101);
nand U2202 (N_2202,N_825,N_1223);
and U2203 (N_2203,N_1054,N_1427);
nand U2204 (N_2204,N_1179,N_247);
nor U2205 (N_2205,N_1261,N_368);
nor U2206 (N_2206,N_1434,N_1327);
and U2207 (N_2207,N_1170,N_44);
or U2208 (N_2208,N_1439,N_440);
nand U2209 (N_2209,N_1042,N_299);
and U2210 (N_2210,N_148,N_574);
or U2211 (N_2211,N_692,N_1239);
and U2212 (N_2212,N_1127,N_182);
or U2213 (N_2213,N_1187,N_1417);
or U2214 (N_2214,N_397,N_1403);
nand U2215 (N_2215,N_183,N_1293);
nand U2216 (N_2216,N_863,N_86);
nand U2217 (N_2217,N_640,N_1227);
or U2218 (N_2218,N_796,N_1103);
and U2219 (N_2219,N_940,N_1278);
nand U2220 (N_2220,N_174,N_1303);
nand U2221 (N_2221,N_1214,N_1007);
nand U2222 (N_2222,N_1389,N_717);
nand U2223 (N_2223,N_1312,N_598);
nor U2224 (N_2224,N_1424,N_291);
nand U2225 (N_2225,N_87,N_480);
nand U2226 (N_2226,N_1093,N_1057);
and U2227 (N_2227,N_231,N_683);
or U2228 (N_2228,N_1459,N_236);
or U2229 (N_2229,N_976,N_1198);
nand U2230 (N_2230,N_82,N_421);
and U2231 (N_2231,N_1085,N_72);
xnor U2232 (N_2232,N_342,N_1084);
or U2233 (N_2233,N_846,N_175);
and U2234 (N_2234,N_953,N_1257);
and U2235 (N_2235,N_363,N_1055);
nor U2236 (N_2236,N_1235,N_1341);
or U2237 (N_2237,N_971,N_428);
nor U2238 (N_2238,N_49,N_1364);
and U2239 (N_2239,N_524,N_115);
or U2240 (N_2240,N_1408,N_1066);
nand U2241 (N_2241,N_256,N_892);
or U2242 (N_2242,N_1276,N_314);
or U2243 (N_2243,N_352,N_458);
or U2244 (N_2244,N_703,N_441);
and U2245 (N_2245,N_92,N_1043);
nand U2246 (N_2246,N_979,N_1336);
nand U2247 (N_2247,N_991,N_1072);
nand U2248 (N_2248,N_1006,N_628);
and U2249 (N_2249,N_924,N_1044);
nor U2250 (N_2250,N_1298,N_699);
nor U2251 (N_2251,N_148,N_1065);
nand U2252 (N_2252,N_268,N_453);
and U2253 (N_2253,N_1186,N_716);
nor U2254 (N_2254,N_349,N_1063);
and U2255 (N_2255,N_1432,N_683);
nand U2256 (N_2256,N_278,N_911);
and U2257 (N_2257,N_274,N_736);
or U2258 (N_2258,N_1336,N_1131);
nor U2259 (N_2259,N_911,N_1096);
or U2260 (N_2260,N_459,N_629);
nand U2261 (N_2261,N_418,N_1199);
nor U2262 (N_2262,N_1377,N_1083);
xnor U2263 (N_2263,N_90,N_1240);
and U2264 (N_2264,N_416,N_1357);
and U2265 (N_2265,N_112,N_1335);
or U2266 (N_2266,N_461,N_550);
or U2267 (N_2267,N_81,N_1272);
and U2268 (N_2268,N_770,N_82);
nand U2269 (N_2269,N_28,N_1111);
nand U2270 (N_2270,N_1220,N_719);
nor U2271 (N_2271,N_102,N_106);
or U2272 (N_2272,N_1070,N_906);
or U2273 (N_2273,N_430,N_467);
nand U2274 (N_2274,N_1101,N_619);
and U2275 (N_2275,N_914,N_781);
nor U2276 (N_2276,N_649,N_1086);
and U2277 (N_2277,N_718,N_407);
nor U2278 (N_2278,N_909,N_999);
and U2279 (N_2279,N_373,N_301);
and U2280 (N_2280,N_1048,N_766);
nand U2281 (N_2281,N_961,N_139);
nand U2282 (N_2282,N_549,N_788);
and U2283 (N_2283,N_92,N_319);
and U2284 (N_2284,N_574,N_713);
nor U2285 (N_2285,N_724,N_1169);
or U2286 (N_2286,N_808,N_962);
and U2287 (N_2287,N_153,N_1245);
nand U2288 (N_2288,N_959,N_301);
nand U2289 (N_2289,N_580,N_628);
nand U2290 (N_2290,N_455,N_740);
nor U2291 (N_2291,N_1426,N_299);
or U2292 (N_2292,N_614,N_12);
and U2293 (N_2293,N_740,N_599);
nor U2294 (N_2294,N_698,N_892);
or U2295 (N_2295,N_794,N_412);
and U2296 (N_2296,N_1183,N_401);
nor U2297 (N_2297,N_502,N_156);
and U2298 (N_2298,N_762,N_884);
and U2299 (N_2299,N_1076,N_740);
and U2300 (N_2300,N_1028,N_140);
or U2301 (N_2301,N_210,N_316);
nand U2302 (N_2302,N_741,N_931);
or U2303 (N_2303,N_191,N_1251);
xnor U2304 (N_2304,N_223,N_647);
nand U2305 (N_2305,N_752,N_627);
nand U2306 (N_2306,N_666,N_1272);
and U2307 (N_2307,N_665,N_808);
nor U2308 (N_2308,N_309,N_1179);
nor U2309 (N_2309,N_1176,N_1404);
nor U2310 (N_2310,N_359,N_458);
or U2311 (N_2311,N_1209,N_306);
nor U2312 (N_2312,N_444,N_185);
and U2313 (N_2313,N_1006,N_328);
nand U2314 (N_2314,N_800,N_1201);
or U2315 (N_2315,N_325,N_1344);
nand U2316 (N_2316,N_557,N_87);
and U2317 (N_2317,N_308,N_329);
and U2318 (N_2318,N_529,N_171);
and U2319 (N_2319,N_564,N_1316);
nor U2320 (N_2320,N_1466,N_1438);
or U2321 (N_2321,N_716,N_724);
nor U2322 (N_2322,N_563,N_1400);
and U2323 (N_2323,N_797,N_1224);
nor U2324 (N_2324,N_1232,N_1428);
nor U2325 (N_2325,N_949,N_1236);
and U2326 (N_2326,N_599,N_482);
nand U2327 (N_2327,N_1089,N_863);
and U2328 (N_2328,N_73,N_520);
nor U2329 (N_2329,N_421,N_471);
or U2330 (N_2330,N_1236,N_647);
nor U2331 (N_2331,N_409,N_1107);
nand U2332 (N_2332,N_104,N_144);
and U2333 (N_2333,N_1055,N_1038);
or U2334 (N_2334,N_594,N_86);
or U2335 (N_2335,N_902,N_1112);
nand U2336 (N_2336,N_474,N_562);
nor U2337 (N_2337,N_1358,N_422);
or U2338 (N_2338,N_788,N_77);
nand U2339 (N_2339,N_1485,N_10);
and U2340 (N_2340,N_82,N_162);
and U2341 (N_2341,N_1342,N_186);
and U2342 (N_2342,N_343,N_1184);
and U2343 (N_2343,N_1405,N_400);
nand U2344 (N_2344,N_1073,N_924);
nand U2345 (N_2345,N_1272,N_483);
or U2346 (N_2346,N_1206,N_188);
or U2347 (N_2347,N_297,N_380);
or U2348 (N_2348,N_1090,N_568);
nand U2349 (N_2349,N_1460,N_48);
nand U2350 (N_2350,N_1251,N_84);
and U2351 (N_2351,N_525,N_422);
and U2352 (N_2352,N_1042,N_39);
and U2353 (N_2353,N_224,N_1171);
or U2354 (N_2354,N_584,N_892);
nor U2355 (N_2355,N_773,N_1452);
and U2356 (N_2356,N_465,N_1331);
nand U2357 (N_2357,N_1070,N_662);
and U2358 (N_2358,N_224,N_94);
or U2359 (N_2359,N_1078,N_94);
and U2360 (N_2360,N_447,N_1079);
nand U2361 (N_2361,N_416,N_754);
nand U2362 (N_2362,N_605,N_732);
nor U2363 (N_2363,N_905,N_1452);
nand U2364 (N_2364,N_687,N_12);
nor U2365 (N_2365,N_748,N_437);
or U2366 (N_2366,N_88,N_1266);
and U2367 (N_2367,N_333,N_1185);
nand U2368 (N_2368,N_1486,N_790);
nand U2369 (N_2369,N_366,N_770);
nand U2370 (N_2370,N_901,N_1316);
or U2371 (N_2371,N_559,N_495);
nor U2372 (N_2372,N_779,N_229);
and U2373 (N_2373,N_497,N_1426);
nor U2374 (N_2374,N_1020,N_1055);
xnor U2375 (N_2375,N_1203,N_197);
nand U2376 (N_2376,N_27,N_903);
nor U2377 (N_2377,N_1455,N_1193);
nor U2378 (N_2378,N_1329,N_1339);
or U2379 (N_2379,N_609,N_42);
or U2380 (N_2380,N_48,N_1061);
xor U2381 (N_2381,N_187,N_1115);
or U2382 (N_2382,N_897,N_376);
nand U2383 (N_2383,N_1498,N_903);
nor U2384 (N_2384,N_675,N_1458);
nand U2385 (N_2385,N_1190,N_1495);
nor U2386 (N_2386,N_1330,N_1354);
nor U2387 (N_2387,N_1417,N_376);
or U2388 (N_2388,N_551,N_935);
and U2389 (N_2389,N_1338,N_1083);
or U2390 (N_2390,N_274,N_711);
and U2391 (N_2391,N_1304,N_1435);
and U2392 (N_2392,N_1150,N_687);
and U2393 (N_2393,N_561,N_932);
or U2394 (N_2394,N_1170,N_1276);
or U2395 (N_2395,N_1131,N_35);
nand U2396 (N_2396,N_454,N_289);
nand U2397 (N_2397,N_18,N_1301);
nand U2398 (N_2398,N_939,N_303);
and U2399 (N_2399,N_770,N_451);
or U2400 (N_2400,N_415,N_649);
nand U2401 (N_2401,N_538,N_1487);
and U2402 (N_2402,N_1443,N_59);
and U2403 (N_2403,N_240,N_365);
or U2404 (N_2404,N_69,N_697);
or U2405 (N_2405,N_256,N_124);
or U2406 (N_2406,N_644,N_883);
or U2407 (N_2407,N_113,N_1368);
nor U2408 (N_2408,N_1052,N_45);
or U2409 (N_2409,N_956,N_571);
nor U2410 (N_2410,N_233,N_699);
nor U2411 (N_2411,N_369,N_730);
nand U2412 (N_2412,N_1263,N_1326);
nand U2413 (N_2413,N_921,N_492);
or U2414 (N_2414,N_424,N_744);
or U2415 (N_2415,N_953,N_343);
nor U2416 (N_2416,N_1317,N_419);
or U2417 (N_2417,N_175,N_1057);
or U2418 (N_2418,N_640,N_1200);
and U2419 (N_2419,N_971,N_591);
and U2420 (N_2420,N_644,N_64);
nor U2421 (N_2421,N_556,N_618);
nand U2422 (N_2422,N_60,N_1297);
nand U2423 (N_2423,N_580,N_51);
or U2424 (N_2424,N_1287,N_828);
and U2425 (N_2425,N_1205,N_56);
nand U2426 (N_2426,N_881,N_49);
xnor U2427 (N_2427,N_878,N_598);
or U2428 (N_2428,N_327,N_360);
nor U2429 (N_2429,N_1045,N_829);
or U2430 (N_2430,N_459,N_552);
nor U2431 (N_2431,N_1457,N_816);
nand U2432 (N_2432,N_680,N_966);
nor U2433 (N_2433,N_148,N_226);
nor U2434 (N_2434,N_816,N_1278);
nand U2435 (N_2435,N_356,N_959);
or U2436 (N_2436,N_1056,N_186);
nor U2437 (N_2437,N_500,N_3);
nand U2438 (N_2438,N_125,N_1247);
or U2439 (N_2439,N_302,N_947);
or U2440 (N_2440,N_1251,N_1045);
and U2441 (N_2441,N_1058,N_416);
nor U2442 (N_2442,N_614,N_229);
and U2443 (N_2443,N_394,N_484);
xnor U2444 (N_2444,N_1419,N_144);
nand U2445 (N_2445,N_890,N_485);
or U2446 (N_2446,N_9,N_787);
nor U2447 (N_2447,N_949,N_1028);
or U2448 (N_2448,N_987,N_438);
nor U2449 (N_2449,N_16,N_772);
or U2450 (N_2450,N_400,N_315);
and U2451 (N_2451,N_72,N_1387);
nand U2452 (N_2452,N_1458,N_1096);
nor U2453 (N_2453,N_322,N_402);
or U2454 (N_2454,N_495,N_826);
or U2455 (N_2455,N_31,N_688);
and U2456 (N_2456,N_982,N_295);
nand U2457 (N_2457,N_729,N_1494);
or U2458 (N_2458,N_413,N_1450);
nor U2459 (N_2459,N_1390,N_109);
or U2460 (N_2460,N_85,N_674);
or U2461 (N_2461,N_1282,N_355);
or U2462 (N_2462,N_1105,N_1340);
and U2463 (N_2463,N_163,N_258);
nand U2464 (N_2464,N_238,N_1377);
nor U2465 (N_2465,N_306,N_1413);
nand U2466 (N_2466,N_243,N_84);
nand U2467 (N_2467,N_1328,N_121);
or U2468 (N_2468,N_332,N_147);
nand U2469 (N_2469,N_298,N_1087);
nor U2470 (N_2470,N_87,N_1295);
or U2471 (N_2471,N_91,N_333);
and U2472 (N_2472,N_684,N_817);
nand U2473 (N_2473,N_829,N_133);
or U2474 (N_2474,N_812,N_368);
nand U2475 (N_2475,N_1300,N_1329);
xnor U2476 (N_2476,N_926,N_760);
and U2477 (N_2477,N_770,N_1049);
nor U2478 (N_2478,N_1227,N_677);
and U2479 (N_2479,N_1091,N_1479);
nor U2480 (N_2480,N_399,N_91);
and U2481 (N_2481,N_1036,N_287);
and U2482 (N_2482,N_1152,N_981);
nand U2483 (N_2483,N_276,N_892);
or U2484 (N_2484,N_97,N_1266);
nand U2485 (N_2485,N_965,N_150);
nor U2486 (N_2486,N_1374,N_1097);
and U2487 (N_2487,N_214,N_748);
nand U2488 (N_2488,N_1149,N_480);
nand U2489 (N_2489,N_880,N_787);
nand U2490 (N_2490,N_1309,N_483);
and U2491 (N_2491,N_613,N_568);
and U2492 (N_2492,N_536,N_1058);
xor U2493 (N_2493,N_1101,N_676);
nand U2494 (N_2494,N_533,N_980);
or U2495 (N_2495,N_641,N_384);
or U2496 (N_2496,N_163,N_230);
and U2497 (N_2497,N_541,N_637);
and U2498 (N_2498,N_629,N_1491);
or U2499 (N_2499,N_56,N_108);
or U2500 (N_2500,N_931,N_1185);
nor U2501 (N_2501,N_424,N_491);
nor U2502 (N_2502,N_93,N_839);
or U2503 (N_2503,N_666,N_938);
or U2504 (N_2504,N_1402,N_794);
or U2505 (N_2505,N_397,N_543);
nand U2506 (N_2506,N_373,N_420);
nor U2507 (N_2507,N_30,N_1338);
and U2508 (N_2508,N_1087,N_1316);
nor U2509 (N_2509,N_466,N_61);
or U2510 (N_2510,N_1205,N_813);
nor U2511 (N_2511,N_1458,N_709);
nand U2512 (N_2512,N_523,N_1204);
and U2513 (N_2513,N_773,N_25);
nand U2514 (N_2514,N_619,N_889);
nand U2515 (N_2515,N_1076,N_214);
nor U2516 (N_2516,N_466,N_22);
xnor U2517 (N_2517,N_991,N_1281);
and U2518 (N_2518,N_1419,N_1325);
and U2519 (N_2519,N_389,N_303);
and U2520 (N_2520,N_144,N_264);
or U2521 (N_2521,N_1437,N_164);
or U2522 (N_2522,N_611,N_146);
nand U2523 (N_2523,N_236,N_673);
nor U2524 (N_2524,N_1289,N_648);
and U2525 (N_2525,N_94,N_1348);
or U2526 (N_2526,N_273,N_434);
or U2527 (N_2527,N_903,N_1047);
or U2528 (N_2528,N_72,N_566);
and U2529 (N_2529,N_212,N_1338);
nor U2530 (N_2530,N_601,N_935);
and U2531 (N_2531,N_413,N_273);
or U2532 (N_2532,N_266,N_841);
and U2533 (N_2533,N_1185,N_430);
nand U2534 (N_2534,N_426,N_801);
or U2535 (N_2535,N_778,N_1305);
or U2536 (N_2536,N_983,N_1138);
nor U2537 (N_2537,N_811,N_382);
xor U2538 (N_2538,N_586,N_819);
nor U2539 (N_2539,N_232,N_464);
or U2540 (N_2540,N_1108,N_260);
and U2541 (N_2541,N_966,N_1429);
nand U2542 (N_2542,N_730,N_1200);
or U2543 (N_2543,N_1126,N_883);
or U2544 (N_2544,N_399,N_1012);
nand U2545 (N_2545,N_656,N_968);
nand U2546 (N_2546,N_1260,N_591);
nor U2547 (N_2547,N_1340,N_591);
nand U2548 (N_2548,N_439,N_935);
nand U2549 (N_2549,N_1053,N_860);
nor U2550 (N_2550,N_871,N_815);
or U2551 (N_2551,N_526,N_913);
or U2552 (N_2552,N_707,N_1273);
and U2553 (N_2553,N_1075,N_1366);
and U2554 (N_2554,N_321,N_263);
nand U2555 (N_2555,N_267,N_1054);
nand U2556 (N_2556,N_1158,N_283);
nor U2557 (N_2557,N_1053,N_858);
nand U2558 (N_2558,N_1009,N_1496);
or U2559 (N_2559,N_1360,N_197);
or U2560 (N_2560,N_40,N_323);
and U2561 (N_2561,N_759,N_466);
or U2562 (N_2562,N_304,N_484);
or U2563 (N_2563,N_1069,N_953);
or U2564 (N_2564,N_398,N_362);
nand U2565 (N_2565,N_749,N_308);
nor U2566 (N_2566,N_123,N_1165);
nand U2567 (N_2567,N_379,N_1397);
or U2568 (N_2568,N_416,N_625);
nand U2569 (N_2569,N_818,N_85);
or U2570 (N_2570,N_381,N_1281);
nor U2571 (N_2571,N_1114,N_1314);
nor U2572 (N_2572,N_358,N_250);
or U2573 (N_2573,N_1138,N_1475);
nor U2574 (N_2574,N_936,N_14);
and U2575 (N_2575,N_1343,N_729);
or U2576 (N_2576,N_1094,N_563);
and U2577 (N_2577,N_1440,N_1130);
nand U2578 (N_2578,N_1239,N_919);
nand U2579 (N_2579,N_22,N_488);
nand U2580 (N_2580,N_6,N_833);
nand U2581 (N_2581,N_1187,N_471);
nand U2582 (N_2582,N_966,N_210);
nand U2583 (N_2583,N_183,N_599);
nor U2584 (N_2584,N_1093,N_846);
and U2585 (N_2585,N_408,N_842);
and U2586 (N_2586,N_1214,N_1349);
nor U2587 (N_2587,N_724,N_969);
nor U2588 (N_2588,N_139,N_180);
and U2589 (N_2589,N_12,N_1054);
nand U2590 (N_2590,N_901,N_1025);
nand U2591 (N_2591,N_1172,N_1014);
or U2592 (N_2592,N_1026,N_600);
or U2593 (N_2593,N_676,N_1410);
nand U2594 (N_2594,N_750,N_1276);
or U2595 (N_2595,N_660,N_1321);
nand U2596 (N_2596,N_605,N_425);
and U2597 (N_2597,N_1168,N_1113);
nor U2598 (N_2598,N_1228,N_1203);
or U2599 (N_2599,N_251,N_983);
nand U2600 (N_2600,N_634,N_473);
and U2601 (N_2601,N_230,N_426);
and U2602 (N_2602,N_226,N_1340);
nand U2603 (N_2603,N_281,N_27);
nor U2604 (N_2604,N_880,N_773);
and U2605 (N_2605,N_778,N_443);
nand U2606 (N_2606,N_1053,N_601);
nand U2607 (N_2607,N_1261,N_514);
and U2608 (N_2608,N_1169,N_1493);
and U2609 (N_2609,N_754,N_295);
nand U2610 (N_2610,N_766,N_130);
nor U2611 (N_2611,N_1369,N_1153);
nor U2612 (N_2612,N_949,N_444);
or U2613 (N_2613,N_275,N_1493);
nand U2614 (N_2614,N_63,N_1322);
and U2615 (N_2615,N_147,N_885);
and U2616 (N_2616,N_1087,N_450);
and U2617 (N_2617,N_1037,N_785);
nand U2618 (N_2618,N_319,N_502);
or U2619 (N_2619,N_1342,N_473);
nor U2620 (N_2620,N_574,N_14);
nand U2621 (N_2621,N_149,N_655);
and U2622 (N_2622,N_303,N_1362);
nand U2623 (N_2623,N_9,N_349);
and U2624 (N_2624,N_921,N_739);
nand U2625 (N_2625,N_618,N_561);
nand U2626 (N_2626,N_1144,N_1220);
and U2627 (N_2627,N_1421,N_640);
xor U2628 (N_2628,N_859,N_106);
nor U2629 (N_2629,N_631,N_1075);
and U2630 (N_2630,N_631,N_657);
and U2631 (N_2631,N_1265,N_673);
or U2632 (N_2632,N_482,N_255);
and U2633 (N_2633,N_94,N_412);
or U2634 (N_2634,N_30,N_373);
nand U2635 (N_2635,N_846,N_642);
nor U2636 (N_2636,N_1299,N_750);
nor U2637 (N_2637,N_1470,N_453);
nand U2638 (N_2638,N_482,N_716);
nand U2639 (N_2639,N_73,N_264);
and U2640 (N_2640,N_326,N_331);
and U2641 (N_2641,N_1126,N_1104);
and U2642 (N_2642,N_1085,N_1261);
nor U2643 (N_2643,N_244,N_1327);
or U2644 (N_2644,N_582,N_578);
nor U2645 (N_2645,N_658,N_1006);
and U2646 (N_2646,N_238,N_961);
or U2647 (N_2647,N_1139,N_892);
nand U2648 (N_2648,N_1229,N_1109);
or U2649 (N_2649,N_43,N_578);
or U2650 (N_2650,N_199,N_473);
nand U2651 (N_2651,N_1126,N_443);
or U2652 (N_2652,N_328,N_1054);
and U2653 (N_2653,N_1211,N_276);
and U2654 (N_2654,N_1347,N_1376);
nand U2655 (N_2655,N_30,N_957);
and U2656 (N_2656,N_271,N_1261);
and U2657 (N_2657,N_970,N_521);
and U2658 (N_2658,N_1088,N_1073);
or U2659 (N_2659,N_938,N_117);
nand U2660 (N_2660,N_607,N_1395);
nor U2661 (N_2661,N_1281,N_534);
and U2662 (N_2662,N_1021,N_1250);
nor U2663 (N_2663,N_120,N_802);
and U2664 (N_2664,N_1247,N_303);
nor U2665 (N_2665,N_512,N_894);
and U2666 (N_2666,N_1299,N_590);
or U2667 (N_2667,N_626,N_1286);
nor U2668 (N_2668,N_383,N_455);
and U2669 (N_2669,N_61,N_1364);
or U2670 (N_2670,N_1273,N_1174);
nand U2671 (N_2671,N_318,N_967);
and U2672 (N_2672,N_862,N_937);
and U2673 (N_2673,N_981,N_447);
nor U2674 (N_2674,N_751,N_1332);
or U2675 (N_2675,N_396,N_1150);
nor U2676 (N_2676,N_797,N_554);
nor U2677 (N_2677,N_927,N_1479);
nand U2678 (N_2678,N_408,N_67);
or U2679 (N_2679,N_594,N_800);
or U2680 (N_2680,N_1085,N_35);
nand U2681 (N_2681,N_1402,N_72);
nand U2682 (N_2682,N_447,N_630);
or U2683 (N_2683,N_354,N_724);
nand U2684 (N_2684,N_456,N_207);
nor U2685 (N_2685,N_143,N_524);
or U2686 (N_2686,N_1455,N_328);
and U2687 (N_2687,N_443,N_1353);
or U2688 (N_2688,N_1369,N_905);
and U2689 (N_2689,N_919,N_1084);
nor U2690 (N_2690,N_65,N_421);
or U2691 (N_2691,N_1498,N_755);
and U2692 (N_2692,N_468,N_1178);
nor U2693 (N_2693,N_814,N_1423);
nor U2694 (N_2694,N_1473,N_1255);
nand U2695 (N_2695,N_1134,N_674);
or U2696 (N_2696,N_1287,N_1419);
and U2697 (N_2697,N_355,N_0);
nand U2698 (N_2698,N_819,N_338);
and U2699 (N_2699,N_274,N_1469);
nand U2700 (N_2700,N_1004,N_1235);
nor U2701 (N_2701,N_1332,N_215);
nand U2702 (N_2702,N_1323,N_73);
or U2703 (N_2703,N_291,N_516);
nand U2704 (N_2704,N_547,N_1455);
nand U2705 (N_2705,N_788,N_1263);
nor U2706 (N_2706,N_928,N_470);
and U2707 (N_2707,N_528,N_428);
or U2708 (N_2708,N_263,N_187);
xor U2709 (N_2709,N_423,N_841);
and U2710 (N_2710,N_954,N_1495);
nor U2711 (N_2711,N_718,N_955);
nand U2712 (N_2712,N_283,N_462);
or U2713 (N_2713,N_101,N_1419);
nor U2714 (N_2714,N_609,N_1450);
nor U2715 (N_2715,N_216,N_1486);
and U2716 (N_2716,N_1434,N_8);
nand U2717 (N_2717,N_550,N_906);
and U2718 (N_2718,N_435,N_382);
xor U2719 (N_2719,N_866,N_220);
nand U2720 (N_2720,N_1259,N_884);
nand U2721 (N_2721,N_1386,N_1314);
nor U2722 (N_2722,N_480,N_375);
nor U2723 (N_2723,N_122,N_132);
or U2724 (N_2724,N_1424,N_1029);
nand U2725 (N_2725,N_67,N_1482);
or U2726 (N_2726,N_699,N_109);
and U2727 (N_2727,N_218,N_1242);
or U2728 (N_2728,N_1248,N_43);
nand U2729 (N_2729,N_522,N_743);
nand U2730 (N_2730,N_609,N_1267);
or U2731 (N_2731,N_901,N_382);
or U2732 (N_2732,N_635,N_663);
nor U2733 (N_2733,N_179,N_1324);
or U2734 (N_2734,N_1047,N_771);
or U2735 (N_2735,N_1289,N_421);
nand U2736 (N_2736,N_1006,N_556);
nor U2737 (N_2737,N_183,N_1300);
nor U2738 (N_2738,N_139,N_1289);
or U2739 (N_2739,N_1433,N_875);
nor U2740 (N_2740,N_445,N_758);
or U2741 (N_2741,N_4,N_1077);
and U2742 (N_2742,N_476,N_89);
and U2743 (N_2743,N_681,N_572);
or U2744 (N_2744,N_675,N_807);
nor U2745 (N_2745,N_708,N_444);
xnor U2746 (N_2746,N_633,N_127);
nor U2747 (N_2747,N_224,N_708);
nor U2748 (N_2748,N_387,N_637);
and U2749 (N_2749,N_1189,N_248);
or U2750 (N_2750,N_1221,N_466);
xor U2751 (N_2751,N_798,N_344);
and U2752 (N_2752,N_978,N_1311);
nor U2753 (N_2753,N_196,N_1150);
nand U2754 (N_2754,N_1337,N_236);
nand U2755 (N_2755,N_96,N_791);
nor U2756 (N_2756,N_746,N_1100);
and U2757 (N_2757,N_1391,N_1159);
and U2758 (N_2758,N_849,N_105);
or U2759 (N_2759,N_599,N_607);
nand U2760 (N_2760,N_205,N_343);
or U2761 (N_2761,N_304,N_478);
or U2762 (N_2762,N_1145,N_727);
nand U2763 (N_2763,N_689,N_440);
and U2764 (N_2764,N_532,N_1413);
nand U2765 (N_2765,N_541,N_1163);
nand U2766 (N_2766,N_49,N_457);
nor U2767 (N_2767,N_384,N_963);
nor U2768 (N_2768,N_548,N_196);
and U2769 (N_2769,N_695,N_875);
or U2770 (N_2770,N_453,N_644);
nand U2771 (N_2771,N_44,N_48);
nor U2772 (N_2772,N_8,N_1491);
or U2773 (N_2773,N_1232,N_799);
nand U2774 (N_2774,N_869,N_1063);
or U2775 (N_2775,N_239,N_864);
or U2776 (N_2776,N_25,N_213);
or U2777 (N_2777,N_411,N_1135);
and U2778 (N_2778,N_1164,N_1261);
nand U2779 (N_2779,N_1360,N_3);
and U2780 (N_2780,N_1275,N_1456);
nand U2781 (N_2781,N_52,N_1175);
and U2782 (N_2782,N_629,N_1122);
or U2783 (N_2783,N_1399,N_1305);
or U2784 (N_2784,N_1171,N_216);
or U2785 (N_2785,N_643,N_1442);
nand U2786 (N_2786,N_198,N_74);
or U2787 (N_2787,N_156,N_915);
or U2788 (N_2788,N_626,N_126);
or U2789 (N_2789,N_242,N_1494);
nand U2790 (N_2790,N_149,N_976);
and U2791 (N_2791,N_338,N_162);
or U2792 (N_2792,N_320,N_454);
or U2793 (N_2793,N_140,N_1490);
nor U2794 (N_2794,N_427,N_5);
nor U2795 (N_2795,N_517,N_916);
or U2796 (N_2796,N_324,N_782);
and U2797 (N_2797,N_1376,N_615);
and U2798 (N_2798,N_599,N_878);
nor U2799 (N_2799,N_628,N_433);
or U2800 (N_2800,N_885,N_1481);
and U2801 (N_2801,N_153,N_835);
nor U2802 (N_2802,N_277,N_311);
and U2803 (N_2803,N_946,N_170);
nand U2804 (N_2804,N_477,N_22);
or U2805 (N_2805,N_1311,N_901);
and U2806 (N_2806,N_397,N_494);
and U2807 (N_2807,N_920,N_827);
nor U2808 (N_2808,N_229,N_670);
or U2809 (N_2809,N_519,N_735);
and U2810 (N_2810,N_423,N_864);
nor U2811 (N_2811,N_771,N_661);
and U2812 (N_2812,N_1218,N_444);
nor U2813 (N_2813,N_374,N_161);
nor U2814 (N_2814,N_1349,N_120);
and U2815 (N_2815,N_395,N_840);
or U2816 (N_2816,N_782,N_419);
or U2817 (N_2817,N_551,N_120);
nor U2818 (N_2818,N_844,N_1206);
nand U2819 (N_2819,N_340,N_1016);
nand U2820 (N_2820,N_611,N_35);
and U2821 (N_2821,N_310,N_1005);
nand U2822 (N_2822,N_644,N_665);
or U2823 (N_2823,N_783,N_1269);
and U2824 (N_2824,N_297,N_355);
nand U2825 (N_2825,N_553,N_124);
nand U2826 (N_2826,N_637,N_718);
or U2827 (N_2827,N_1332,N_142);
nor U2828 (N_2828,N_1440,N_272);
or U2829 (N_2829,N_1067,N_126);
nor U2830 (N_2830,N_14,N_807);
nand U2831 (N_2831,N_743,N_1127);
and U2832 (N_2832,N_421,N_802);
nor U2833 (N_2833,N_475,N_281);
nor U2834 (N_2834,N_533,N_563);
nand U2835 (N_2835,N_407,N_942);
or U2836 (N_2836,N_432,N_1235);
nor U2837 (N_2837,N_575,N_1290);
nor U2838 (N_2838,N_377,N_969);
nand U2839 (N_2839,N_178,N_172);
nor U2840 (N_2840,N_1404,N_1245);
or U2841 (N_2841,N_1331,N_1418);
nor U2842 (N_2842,N_501,N_172);
and U2843 (N_2843,N_1105,N_171);
nor U2844 (N_2844,N_1309,N_254);
or U2845 (N_2845,N_115,N_231);
or U2846 (N_2846,N_92,N_152);
or U2847 (N_2847,N_556,N_166);
nand U2848 (N_2848,N_1229,N_682);
nand U2849 (N_2849,N_345,N_537);
and U2850 (N_2850,N_775,N_253);
nor U2851 (N_2851,N_734,N_490);
nor U2852 (N_2852,N_573,N_61);
nand U2853 (N_2853,N_1265,N_1159);
or U2854 (N_2854,N_1443,N_41);
nor U2855 (N_2855,N_350,N_426);
and U2856 (N_2856,N_201,N_11);
or U2857 (N_2857,N_265,N_1457);
nor U2858 (N_2858,N_788,N_819);
xnor U2859 (N_2859,N_912,N_296);
nand U2860 (N_2860,N_1133,N_1159);
nand U2861 (N_2861,N_287,N_325);
and U2862 (N_2862,N_613,N_32);
and U2863 (N_2863,N_299,N_127);
nand U2864 (N_2864,N_1201,N_1279);
nor U2865 (N_2865,N_368,N_447);
and U2866 (N_2866,N_685,N_1384);
or U2867 (N_2867,N_455,N_1020);
nand U2868 (N_2868,N_656,N_851);
nand U2869 (N_2869,N_1276,N_1394);
or U2870 (N_2870,N_747,N_902);
nor U2871 (N_2871,N_1458,N_752);
or U2872 (N_2872,N_496,N_1408);
and U2873 (N_2873,N_889,N_1460);
nand U2874 (N_2874,N_156,N_436);
and U2875 (N_2875,N_183,N_716);
or U2876 (N_2876,N_1163,N_9);
or U2877 (N_2877,N_1380,N_429);
and U2878 (N_2878,N_495,N_1376);
nand U2879 (N_2879,N_818,N_510);
nand U2880 (N_2880,N_601,N_600);
nand U2881 (N_2881,N_1238,N_18);
xor U2882 (N_2882,N_1018,N_1057);
and U2883 (N_2883,N_993,N_1016);
and U2884 (N_2884,N_845,N_37);
xnor U2885 (N_2885,N_1025,N_854);
nand U2886 (N_2886,N_785,N_657);
and U2887 (N_2887,N_641,N_1325);
nor U2888 (N_2888,N_127,N_1115);
and U2889 (N_2889,N_787,N_1128);
nand U2890 (N_2890,N_859,N_162);
nor U2891 (N_2891,N_372,N_786);
or U2892 (N_2892,N_761,N_1115);
xnor U2893 (N_2893,N_917,N_981);
and U2894 (N_2894,N_571,N_616);
and U2895 (N_2895,N_808,N_856);
nor U2896 (N_2896,N_1403,N_1424);
nor U2897 (N_2897,N_694,N_1041);
nand U2898 (N_2898,N_152,N_946);
nand U2899 (N_2899,N_388,N_1);
and U2900 (N_2900,N_22,N_803);
or U2901 (N_2901,N_755,N_362);
and U2902 (N_2902,N_1376,N_1345);
and U2903 (N_2903,N_594,N_79);
and U2904 (N_2904,N_785,N_580);
nor U2905 (N_2905,N_220,N_674);
and U2906 (N_2906,N_1177,N_707);
or U2907 (N_2907,N_1023,N_1414);
nand U2908 (N_2908,N_753,N_824);
nor U2909 (N_2909,N_697,N_835);
and U2910 (N_2910,N_840,N_709);
and U2911 (N_2911,N_1349,N_767);
nand U2912 (N_2912,N_827,N_1154);
and U2913 (N_2913,N_1278,N_1431);
nand U2914 (N_2914,N_708,N_1102);
and U2915 (N_2915,N_441,N_1058);
or U2916 (N_2916,N_984,N_767);
or U2917 (N_2917,N_76,N_1480);
nor U2918 (N_2918,N_1150,N_1099);
or U2919 (N_2919,N_308,N_898);
nor U2920 (N_2920,N_558,N_421);
or U2921 (N_2921,N_776,N_1297);
and U2922 (N_2922,N_1073,N_274);
nor U2923 (N_2923,N_1415,N_1493);
or U2924 (N_2924,N_1309,N_1113);
nand U2925 (N_2925,N_470,N_213);
nand U2926 (N_2926,N_814,N_627);
or U2927 (N_2927,N_1458,N_635);
and U2928 (N_2928,N_174,N_254);
or U2929 (N_2929,N_520,N_1423);
nand U2930 (N_2930,N_488,N_735);
or U2931 (N_2931,N_629,N_178);
or U2932 (N_2932,N_302,N_1315);
and U2933 (N_2933,N_1125,N_706);
nor U2934 (N_2934,N_1478,N_621);
and U2935 (N_2935,N_630,N_198);
or U2936 (N_2936,N_858,N_1150);
and U2937 (N_2937,N_430,N_1348);
nor U2938 (N_2938,N_48,N_176);
and U2939 (N_2939,N_1462,N_323);
xor U2940 (N_2940,N_1067,N_1270);
and U2941 (N_2941,N_711,N_6);
and U2942 (N_2942,N_1145,N_434);
nor U2943 (N_2943,N_115,N_730);
and U2944 (N_2944,N_965,N_342);
and U2945 (N_2945,N_54,N_826);
and U2946 (N_2946,N_285,N_989);
nor U2947 (N_2947,N_1091,N_294);
nor U2948 (N_2948,N_695,N_352);
nand U2949 (N_2949,N_797,N_899);
nor U2950 (N_2950,N_1259,N_304);
and U2951 (N_2951,N_228,N_1323);
nor U2952 (N_2952,N_1061,N_612);
and U2953 (N_2953,N_1403,N_521);
or U2954 (N_2954,N_1433,N_657);
and U2955 (N_2955,N_473,N_351);
or U2956 (N_2956,N_1423,N_257);
or U2957 (N_2957,N_900,N_940);
nor U2958 (N_2958,N_1276,N_1470);
and U2959 (N_2959,N_1103,N_52);
nand U2960 (N_2960,N_173,N_513);
nor U2961 (N_2961,N_1183,N_1398);
and U2962 (N_2962,N_435,N_432);
nor U2963 (N_2963,N_520,N_1327);
nand U2964 (N_2964,N_1309,N_1152);
nor U2965 (N_2965,N_4,N_289);
or U2966 (N_2966,N_1321,N_64);
nor U2967 (N_2967,N_706,N_714);
nor U2968 (N_2968,N_1451,N_840);
and U2969 (N_2969,N_1145,N_167);
or U2970 (N_2970,N_255,N_568);
nand U2971 (N_2971,N_968,N_682);
nand U2972 (N_2972,N_579,N_731);
and U2973 (N_2973,N_308,N_1461);
or U2974 (N_2974,N_1201,N_1492);
and U2975 (N_2975,N_879,N_1242);
or U2976 (N_2976,N_334,N_1173);
or U2977 (N_2977,N_487,N_1026);
nand U2978 (N_2978,N_539,N_281);
and U2979 (N_2979,N_730,N_1105);
or U2980 (N_2980,N_417,N_454);
nor U2981 (N_2981,N_366,N_513);
or U2982 (N_2982,N_170,N_1479);
and U2983 (N_2983,N_1394,N_1091);
xor U2984 (N_2984,N_717,N_24);
or U2985 (N_2985,N_299,N_125);
nand U2986 (N_2986,N_699,N_763);
nor U2987 (N_2987,N_492,N_724);
nand U2988 (N_2988,N_1137,N_1208);
or U2989 (N_2989,N_531,N_39);
nand U2990 (N_2990,N_1275,N_1215);
or U2991 (N_2991,N_1021,N_1232);
xor U2992 (N_2992,N_854,N_939);
and U2993 (N_2993,N_556,N_1420);
nand U2994 (N_2994,N_497,N_1127);
xor U2995 (N_2995,N_146,N_903);
or U2996 (N_2996,N_1225,N_273);
or U2997 (N_2997,N_693,N_235);
nor U2998 (N_2998,N_337,N_443);
nor U2999 (N_2999,N_349,N_1011);
and U3000 (N_3000,N_1981,N_1706);
or U3001 (N_3001,N_2476,N_2608);
or U3002 (N_3002,N_2940,N_1880);
nand U3003 (N_3003,N_2686,N_2403);
and U3004 (N_3004,N_2302,N_2550);
nor U3005 (N_3005,N_2086,N_1814);
nand U3006 (N_3006,N_2062,N_2372);
and U3007 (N_3007,N_1543,N_2484);
or U3008 (N_3008,N_1996,N_2161);
or U3009 (N_3009,N_2059,N_2091);
or U3010 (N_3010,N_1863,N_2728);
nand U3011 (N_3011,N_1529,N_2173);
nand U3012 (N_3012,N_2245,N_2343);
nor U3013 (N_3013,N_1786,N_1868);
nor U3014 (N_3014,N_2603,N_2075);
or U3015 (N_3015,N_2650,N_1993);
and U3016 (N_3016,N_2396,N_2363);
nor U3017 (N_3017,N_2146,N_2624);
or U3018 (N_3018,N_2300,N_2283);
and U3019 (N_3019,N_1979,N_2406);
nand U3020 (N_3020,N_2911,N_2811);
and U3021 (N_3021,N_1772,N_2371);
nor U3022 (N_3022,N_2839,N_2357);
nor U3023 (N_3023,N_2899,N_2276);
nor U3024 (N_3024,N_2362,N_1956);
or U3025 (N_3025,N_2392,N_2916);
and U3026 (N_3026,N_1554,N_2596);
or U3027 (N_3027,N_2769,N_2452);
and U3028 (N_3028,N_2174,N_1600);
and U3029 (N_3029,N_1566,N_2050);
nand U3030 (N_3030,N_1716,N_2642);
nand U3031 (N_3031,N_2522,N_2006);
nor U3032 (N_3032,N_2255,N_1746);
nor U3033 (N_3033,N_2206,N_2387);
or U3034 (N_3034,N_1944,N_1684);
and U3035 (N_3035,N_2260,N_2195);
nor U3036 (N_3036,N_1589,N_2320);
or U3037 (N_3037,N_2984,N_2758);
nand U3038 (N_3038,N_1699,N_1753);
and U3039 (N_3039,N_1774,N_1740);
or U3040 (N_3040,N_2253,N_2151);
nand U3041 (N_3041,N_1526,N_2943);
and U3042 (N_3042,N_2474,N_1731);
nand U3043 (N_3043,N_1888,N_1663);
nand U3044 (N_3044,N_2582,N_2717);
or U3045 (N_3045,N_1704,N_1884);
nor U3046 (N_3046,N_2103,N_1816);
nand U3047 (N_3047,N_2511,N_2945);
and U3048 (N_3048,N_2077,N_2118);
nand U3049 (N_3049,N_1895,N_2877);
nor U3050 (N_3050,N_1667,N_1946);
xnor U3051 (N_3051,N_2785,N_1949);
and U3052 (N_3052,N_1604,N_2823);
and U3053 (N_3053,N_2532,N_1922);
and U3054 (N_3054,N_2274,N_2663);
or U3055 (N_3055,N_2386,N_2616);
nand U3056 (N_3056,N_1782,N_2031);
nor U3057 (N_3057,N_1661,N_2678);
nor U3058 (N_3058,N_2776,N_2808);
and U3059 (N_3059,N_2819,N_2487);
and U3060 (N_3060,N_2322,N_2506);
nand U3061 (N_3061,N_1668,N_2165);
nand U3062 (N_3062,N_2617,N_1641);
xor U3063 (N_3063,N_1867,N_2157);
nand U3064 (N_3064,N_2925,N_2346);
and U3065 (N_3065,N_1727,N_2671);
and U3066 (N_3066,N_2598,N_1797);
nor U3067 (N_3067,N_2572,N_1999);
and U3068 (N_3068,N_2459,N_2036);
nand U3069 (N_3069,N_2304,N_2604);
xnor U3070 (N_3070,N_2820,N_2424);
nor U3071 (N_3071,N_2583,N_1788);
nand U3072 (N_3072,N_2350,N_2869);
or U3073 (N_3073,N_1758,N_2429);
nor U3074 (N_3074,N_2637,N_2883);
or U3075 (N_3075,N_1528,N_2106);
nand U3076 (N_3076,N_1843,N_2766);
nand U3077 (N_3077,N_2149,N_2134);
and U3078 (N_3078,N_2521,N_2166);
nand U3079 (N_3079,N_1771,N_2740);
or U3080 (N_3080,N_2779,N_2690);
nor U3081 (N_3081,N_1921,N_2222);
nand U3082 (N_3082,N_2992,N_2147);
nor U3083 (N_3083,N_2181,N_2189);
or U3084 (N_3084,N_2012,N_1990);
and U3085 (N_3085,N_1714,N_1871);
or U3086 (N_3086,N_2793,N_2310);
or U3087 (N_3087,N_2438,N_2090);
or U3088 (N_3088,N_1682,N_2798);
nand U3089 (N_3089,N_1739,N_2337);
nor U3090 (N_3090,N_2767,N_2319);
or U3091 (N_3091,N_2141,N_2379);
nor U3092 (N_3092,N_2131,N_1718);
and U3093 (N_3093,N_1586,N_2998);
or U3094 (N_3094,N_2230,N_1961);
nor U3095 (N_3095,N_1966,N_2441);
or U3096 (N_3096,N_1992,N_2982);
and U3097 (N_3097,N_2145,N_2205);
or U3098 (N_3098,N_1562,N_1627);
nor U3099 (N_3099,N_1953,N_2607);
nand U3100 (N_3100,N_1693,N_2332);
nor U3101 (N_3101,N_1834,N_2965);
nor U3102 (N_3102,N_2067,N_1577);
nand U3103 (N_3103,N_2207,N_2672);
nor U3104 (N_3104,N_2780,N_2339);
nand U3105 (N_3105,N_1665,N_1896);
nor U3106 (N_3106,N_1831,N_2082);
and U3107 (N_3107,N_2196,N_2803);
xnor U3108 (N_3108,N_2004,N_2570);
or U3109 (N_3109,N_2411,N_2962);
nand U3110 (N_3110,N_1901,N_2390);
and U3111 (N_3111,N_1929,N_2997);
nand U3112 (N_3112,N_2810,N_1752);
xor U3113 (N_3113,N_1964,N_1859);
or U3114 (N_3114,N_2226,N_1733);
nor U3115 (N_3115,N_2680,N_1556);
nor U3116 (N_3116,N_1524,N_2950);
nand U3117 (N_3117,N_2266,N_1507);
nand U3118 (N_3118,N_1555,N_2132);
and U3119 (N_3119,N_1862,N_1748);
nand U3120 (N_3120,N_1702,N_2317);
nand U3121 (N_3121,N_1813,N_1829);
and U3122 (N_3122,N_2546,N_2289);
nor U3123 (N_3123,N_2257,N_2581);
nor U3124 (N_3124,N_2073,N_2405);
and U3125 (N_3125,N_2023,N_1887);
or U3126 (N_3126,N_2898,N_2177);
nand U3127 (N_3127,N_1621,N_1502);
nand U3128 (N_3128,N_1781,N_2731);
nor U3129 (N_3129,N_1613,N_2739);
and U3130 (N_3130,N_1710,N_2845);
nor U3131 (N_3131,N_2960,N_1672);
nand U3132 (N_3132,N_1991,N_2952);
and U3133 (N_3133,N_1801,N_2730);
nor U3134 (N_3134,N_1989,N_2273);
nand U3135 (N_3135,N_2171,N_2977);
nand U3136 (N_3136,N_2436,N_2626);
nor U3137 (N_3137,N_2391,N_2264);
and U3138 (N_3138,N_2555,N_2024);
and U3139 (N_3139,N_1516,N_1840);
nand U3140 (N_3140,N_1910,N_2400);
or U3141 (N_3141,N_2590,N_2974);
and U3142 (N_3142,N_1764,N_2233);
or U3143 (N_3143,N_2609,N_2243);
and U3144 (N_3144,N_2432,N_2102);
or U3145 (N_3145,N_2854,N_2790);
nand U3146 (N_3146,N_2834,N_2968);
nor U3147 (N_3147,N_1546,N_1988);
nor U3148 (N_3148,N_1552,N_2172);
nand U3149 (N_3149,N_2928,N_1755);
nand U3150 (N_3150,N_1547,N_2540);
xnor U3151 (N_3151,N_2762,N_2634);
nor U3152 (N_3152,N_1845,N_2721);
and U3153 (N_3153,N_2847,N_2996);
nor U3154 (N_3154,N_2880,N_2744);
nand U3155 (N_3155,N_1965,N_1730);
or U3156 (N_3156,N_2882,N_2185);
or U3157 (N_3157,N_2236,N_2385);
nor U3158 (N_3158,N_1579,N_2860);
or U3159 (N_3159,N_1626,N_2765);
nand U3160 (N_3160,N_1928,N_2755);
or U3161 (N_3161,N_2413,N_2682);
xor U3162 (N_3162,N_2323,N_2813);
or U3163 (N_3163,N_2365,N_2802);
nor U3164 (N_3164,N_1905,N_2098);
xnor U3165 (N_3165,N_2846,N_2211);
nor U3166 (N_3166,N_1823,N_1970);
nand U3167 (N_3167,N_2515,N_2115);
nor U3168 (N_3168,N_1924,N_2833);
and U3169 (N_3169,N_1977,N_2223);
nand U3170 (N_3170,N_2081,N_2001);
nor U3171 (N_3171,N_2787,N_2559);
or U3172 (N_3172,N_2922,N_1864);
and U3173 (N_3173,N_2116,N_2043);
nand U3174 (N_3174,N_1550,N_2100);
and U3175 (N_3175,N_1588,N_2704);
and U3176 (N_3176,N_2577,N_2473);
and U3177 (N_3177,N_2294,N_1968);
nand U3178 (N_3178,N_2058,N_2221);
nand U3179 (N_3179,N_1837,N_2921);
and U3180 (N_3180,N_2451,N_2130);
and U3181 (N_3181,N_2752,N_1670);
nor U3182 (N_3182,N_1776,N_1942);
and U3183 (N_3183,N_1914,N_2942);
and U3184 (N_3184,N_2258,N_1899);
nor U3185 (N_3185,N_2886,N_2771);
nand U3186 (N_3186,N_2093,N_2543);
or U3187 (N_3187,N_2589,N_2303);
and U3188 (N_3188,N_2821,N_2011);
nand U3189 (N_3189,N_1872,N_2993);
xnor U3190 (N_3190,N_2623,N_1923);
nand U3191 (N_3191,N_2139,N_2137);
nor U3192 (N_3192,N_2014,N_2485);
nand U3193 (N_3193,N_2085,N_2250);
or U3194 (N_3194,N_1701,N_2468);
xor U3195 (N_3195,N_2120,N_1724);
or U3196 (N_3196,N_2913,N_1817);
nand U3197 (N_3197,N_2972,N_2510);
nand U3198 (N_3198,N_2295,N_1590);
nand U3199 (N_3199,N_2770,N_2374);
and U3200 (N_3200,N_2469,N_1892);
nand U3201 (N_3201,N_1582,N_2931);
nor U3202 (N_3202,N_2696,N_1518);
or U3203 (N_3203,N_2007,N_1595);
or U3204 (N_3204,N_1612,N_1792);
and U3205 (N_3205,N_2265,N_2076);
and U3206 (N_3206,N_1631,N_2318);
nor U3207 (N_3207,N_1911,N_2584);
or U3208 (N_3208,N_2450,N_2158);
nor U3209 (N_3209,N_2618,N_2687);
and U3210 (N_3210,N_2707,N_1646);
nor U3211 (N_3211,N_2733,N_2649);
or U3212 (N_3212,N_2791,N_2627);
and U3213 (N_3213,N_1508,N_2108);
and U3214 (N_3214,N_2015,N_2517);
nand U3215 (N_3215,N_1794,N_2939);
nand U3216 (N_3216,N_2868,N_2805);
nand U3217 (N_3217,N_2738,N_2800);
and U3218 (N_3218,N_2852,N_1960);
and U3219 (N_3219,N_2194,N_2751);
and U3220 (N_3220,N_1602,N_1737);
nand U3221 (N_3221,N_2150,N_1997);
xnor U3222 (N_3222,N_2615,N_2366);
and U3223 (N_3223,N_2660,N_2336);
and U3224 (N_3224,N_1688,N_1622);
nand U3225 (N_3225,N_2900,N_1918);
nand U3226 (N_3226,N_2261,N_1711);
and U3227 (N_3227,N_2849,N_1900);
nand U3228 (N_3228,N_2259,N_2838);
or U3229 (N_3229,N_2159,N_1994);
nor U3230 (N_3230,N_2252,N_2280);
nor U3231 (N_3231,N_2092,N_2639);
nand U3232 (N_3232,N_1917,N_2685);
nor U3233 (N_3233,N_2453,N_1935);
or U3234 (N_3234,N_2673,N_2488);
nor U3235 (N_3235,N_2279,N_2674);
nor U3236 (N_3236,N_2599,N_2269);
nor U3237 (N_3237,N_2560,N_2224);
nor U3238 (N_3238,N_2836,N_2442);
nor U3239 (N_3239,N_2064,N_2143);
nand U3240 (N_3240,N_2580,N_1599);
and U3241 (N_3241,N_1683,N_2830);
and U3242 (N_3242,N_2632,N_2551);
nand U3243 (N_3243,N_1765,N_1898);
xor U3244 (N_3244,N_2241,N_2544);
and U3245 (N_3245,N_1882,N_2478);
nand U3246 (N_3246,N_2710,N_1705);
nor U3247 (N_3247,N_1879,N_2489);
nand U3248 (N_3248,N_2270,N_2029);
nor U3249 (N_3249,N_1975,N_1958);
nor U3250 (N_3250,N_2645,N_2713);
and U3251 (N_3251,N_2352,N_1926);
nand U3252 (N_3252,N_2953,N_2017);
or U3253 (N_3253,N_1652,N_1793);
nand U3254 (N_3254,N_2742,N_2594);
and U3255 (N_3255,N_2349,N_2375);
and U3256 (N_3256,N_2286,N_2504);
nor U3257 (N_3257,N_2575,N_2421);
nand U3258 (N_3258,N_2622,N_2954);
nor U3259 (N_3259,N_1608,N_1870);
nor U3260 (N_3260,N_1544,N_1983);
nand U3261 (N_3261,N_2030,N_2325);
or U3262 (N_3262,N_2725,N_2219);
or U3263 (N_3263,N_1973,N_2518);
nand U3264 (N_3264,N_1656,N_2531);
and U3265 (N_3265,N_1632,N_1743);
or U3266 (N_3266,N_2809,N_1597);
nand U3267 (N_3267,N_2536,N_2423);
nor U3268 (N_3268,N_1617,N_2465);
nand U3269 (N_3269,N_2112,N_2154);
or U3270 (N_3270,N_1619,N_2587);
nor U3271 (N_3271,N_2446,N_2268);
nand U3272 (N_3272,N_2360,N_2493);
or U3273 (N_3273,N_1854,N_2825);
nor U3274 (N_3274,N_2949,N_2121);
nand U3275 (N_3275,N_1594,N_2525);
or U3276 (N_3276,N_1649,N_2653);
nand U3277 (N_3277,N_1607,N_2367);
and U3278 (N_3278,N_1745,N_2419);
nor U3279 (N_3279,N_2991,N_2907);
and U3280 (N_3280,N_2657,N_2702);
or U3281 (N_3281,N_1936,N_2549);
nor U3282 (N_3282,N_2711,N_1603);
or U3283 (N_3283,N_2985,N_2351);
and U3284 (N_3284,N_2398,N_1985);
and U3285 (N_3285,N_2435,N_2373);
or U3286 (N_3286,N_1674,N_2724);
and U3287 (N_3287,N_2281,N_2018);
or U3288 (N_3288,N_2315,N_1698);
nand U3289 (N_3289,N_1809,N_1509);
or U3290 (N_3290,N_2843,N_1967);
or U3291 (N_3291,N_2547,N_2123);
and U3292 (N_3292,N_2698,N_1653);
nand U3293 (N_3293,N_2792,N_2815);
or U3294 (N_3294,N_2213,N_2407);
nor U3295 (N_3295,N_1534,N_1648);
nor U3296 (N_3296,N_2864,N_2142);
and U3297 (N_3297,N_1841,N_1742);
and U3298 (N_3298,N_2688,N_1651);
nor U3299 (N_3299,N_2995,N_1568);
nand U3300 (N_3300,N_2329,N_1978);
nor U3301 (N_3301,N_1757,N_2313);
nand U3302 (N_3302,N_2901,N_2973);
nand U3303 (N_3303,N_2291,N_2937);
nand U3304 (N_3304,N_1932,N_2908);
xnor U3305 (N_3305,N_2037,N_2060);
nand U3306 (N_3306,N_2079,N_2923);
and U3307 (N_3307,N_1886,N_2884);
or U3308 (N_3308,N_2025,N_2503);
or U3309 (N_3309,N_2670,N_1720);
nor U3310 (N_3310,N_2558,N_2826);
nand U3311 (N_3311,N_1869,N_2119);
nor U3312 (N_3312,N_1606,N_2795);
xnor U3313 (N_3313,N_1520,N_1707);
nand U3314 (N_3314,N_2113,N_1703);
or U3315 (N_3315,N_1940,N_2369);
and U3316 (N_3316,N_2669,N_2620);
nand U3317 (N_3317,N_2046,N_2244);
and U3318 (N_3318,N_2797,N_2969);
and U3319 (N_3319,N_1678,N_2975);
nor U3320 (N_3320,N_2679,N_2914);
and U3321 (N_3321,N_1647,N_1931);
or U3322 (N_3322,N_2736,N_2160);
or U3323 (N_3323,N_1618,N_2238);
nand U3324 (N_3324,N_2723,N_2818);
nand U3325 (N_3325,N_2388,N_2104);
and U3326 (N_3326,N_2210,N_1954);
nor U3327 (N_3327,N_2978,N_1934);
and U3328 (N_3328,N_2548,N_1734);
nor U3329 (N_3329,N_1624,N_2463);
and U3330 (N_3330,N_2801,N_2187);
nand U3331 (N_3331,N_2472,N_2324);
and U3332 (N_3332,N_1824,N_1645);
nand U3333 (N_3333,N_2824,N_2905);
nand U3334 (N_3334,N_2695,N_1835);
or U3335 (N_3335,N_2344,N_1655);
nor U3336 (N_3336,N_2122,N_1679);
nand U3337 (N_3337,N_2799,N_2648);
and U3338 (N_3338,N_2296,N_2111);
and U3339 (N_3339,N_2353,N_2389);
nand U3340 (N_3340,N_1511,N_2885);
nand U3341 (N_3341,N_2527,N_1874);
xnor U3342 (N_3342,N_2875,N_1728);
nor U3343 (N_3343,N_2410,N_2920);
and U3344 (N_3344,N_2612,N_2855);
and U3345 (N_3345,N_1717,N_2545);
xor U3346 (N_3346,N_1536,N_1723);
nor U3347 (N_3347,N_1769,N_1609);
nor U3348 (N_3348,N_1943,N_2164);
or U3349 (N_3349,N_2292,N_1738);
nand U3350 (N_3350,N_1969,N_2867);
nand U3351 (N_3351,N_1735,N_1766);
nor U3352 (N_3352,N_1548,N_1807);
nor U3353 (N_3353,N_2537,N_1659);
nor U3354 (N_3354,N_2010,N_1584);
nor U3355 (N_3355,N_2988,N_2193);
and U3356 (N_3356,N_2894,N_2715);
nor U3357 (N_3357,N_2862,N_2109);
and U3358 (N_3358,N_1838,N_2097);
or U3359 (N_3359,N_1732,N_2202);
or U3360 (N_3360,N_1768,N_2301);
xnor U3361 (N_3361,N_2976,N_2041);
and U3362 (N_3362,N_1686,N_2628);
nand U3363 (N_3363,N_2022,N_2591);
and U3364 (N_3364,N_2354,N_2910);
or U3365 (N_3365,N_2807,N_2418);
nor U3366 (N_3366,N_2753,N_2056);
or U3367 (N_3367,N_1971,N_2856);
or U3368 (N_3368,N_1572,N_2298);
nand U3369 (N_3369,N_2870,N_2057);
nor U3370 (N_3370,N_1815,N_1551);
xnor U3371 (N_3371,N_2876,N_2393);
nor U3372 (N_3372,N_2055,N_2307);
or U3373 (N_3373,N_2078,N_1877);
and U3374 (N_3374,N_2231,N_1637);
and U3375 (N_3375,N_1787,N_2404);
and U3376 (N_3376,N_2709,N_2831);
or U3377 (N_3377,N_1540,N_2044);
and U3378 (N_3378,N_2080,N_1522);
nand U3379 (N_3379,N_2415,N_1856);
or U3380 (N_3380,N_2027,N_1643);
nand U3381 (N_3381,N_2578,N_2267);
or U3382 (N_3382,N_2667,N_2052);
or U3383 (N_3383,N_2455,N_2593);
nand U3384 (N_3384,N_2471,N_2416);
and U3385 (N_3385,N_1636,N_1847);
nand U3386 (N_3386,N_2033,N_2606);
nand U3387 (N_3387,N_2936,N_2290);
and U3388 (N_3388,N_2448,N_2186);
and U3389 (N_3389,N_2288,N_2859);
or U3390 (N_3390,N_2198,N_2722);
and U3391 (N_3391,N_2735,N_1947);
and U3392 (N_3392,N_1848,N_2072);
nand U3393 (N_3393,N_1553,N_2458);
nand U3394 (N_3394,N_2734,N_2359);
or U3395 (N_3395,N_2538,N_2275);
and U3396 (N_3396,N_1860,N_2948);
or U3397 (N_3397,N_2720,N_2378);
nor U3398 (N_3398,N_2249,N_1798);
nor U3399 (N_3399,N_1567,N_2523);
nand U3400 (N_3400,N_1885,N_1938);
nor U3401 (N_3401,N_1865,N_2401);
or U3402 (N_3402,N_1819,N_2184);
nor U3403 (N_3403,N_1980,N_1598);
or U3404 (N_3404,N_2214,N_2228);
nor U3405 (N_3405,N_1601,N_2964);
nor U3406 (N_3406,N_2381,N_2941);
and U3407 (N_3407,N_2032,N_2534);
nor U3408 (N_3408,N_2412,N_1976);
and U3409 (N_3409,N_2906,N_2666);
nor U3410 (N_3410,N_1821,N_1912);
nand U3411 (N_3411,N_1515,N_2494);
nand U3412 (N_3412,N_2498,N_1532);
or U3413 (N_3413,N_2595,N_2764);
and U3414 (N_3414,N_1749,N_2271);
and U3415 (N_3415,N_2110,N_1583);
or U3416 (N_3416,N_1736,N_2066);
nand U3417 (N_3417,N_2557,N_2837);
or U3418 (N_3418,N_2089,N_1666);
and U3419 (N_3419,N_2505,N_2528);
nor U3420 (N_3420,N_1941,N_1842);
or U3421 (N_3421,N_2701,N_2358);
nand U3422 (N_3422,N_1952,N_1571);
or U3423 (N_3423,N_2621,N_2567);
nor U3424 (N_3424,N_2760,N_2661);
nand U3425 (N_3425,N_2083,N_2850);
nor U3426 (N_3426,N_2892,N_2576);
or U3427 (N_3427,N_1564,N_2225);
nand U3428 (N_3428,N_2611,N_2482);
and U3429 (N_3429,N_1713,N_2840);
and U3430 (N_3430,N_1542,N_2491);
nor U3431 (N_3431,N_2464,N_2246);
xnor U3432 (N_3432,N_1610,N_1616);
and U3433 (N_3433,N_2425,N_2169);
nand U3434 (N_3434,N_1527,N_1592);
nor U3435 (N_3435,N_1689,N_1687);
nor U3436 (N_3436,N_2574,N_1987);
or U3437 (N_3437,N_2430,N_2692);
nor U3438 (N_3438,N_2857,N_1825);
and U3439 (N_3439,N_2308,N_2930);
and U3440 (N_3440,N_1875,N_2422);
or U3441 (N_3441,N_2705,N_1839);
nor U3442 (N_3442,N_2665,N_2140);
nor U3443 (N_3443,N_2507,N_1907);
or U3444 (N_3444,N_2239,N_1846);
or U3445 (N_3445,N_2873,N_2812);
and U3446 (N_3446,N_1537,N_1640);
or U3447 (N_3447,N_1541,N_2817);
and U3448 (N_3448,N_2640,N_1681);
and U3449 (N_3449,N_2851,N_2314);
or U3450 (N_3450,N_2509,N_2651);
nand U3451 (N_3451,N_1623,N_2775);
and U3452 (N_3452,N_2168,N_2437);
and U3453 (N_3453,N_2566,N_2554);
nand U3454 (N_3454,N_1692,N_1796);
nand U3455 (N_3455,N_2084,N_1916);
nand U3456 (N_3456,N_2061,N_2912);
or U3457 (N_3457,N_2781,N_2105);
and U3458 (N_3458,N_2242,N_2989);
nand U3459 (N_3459,N_1530,N_2979);
or U3460 (N_3460,N_2216,N_1799);
or U3461 (N_3461,N_2944,N_2417);
nor U3462 (N_3462,N_2646,N_2716);
nor U3463 (N_3463,N_2853,N_2778);
nand U3464 (N_3464,N_2946,N_2201);
nor U3465 (N_3465,N_1857,N_1504);
and U3466 (N_3466,N_2321,N_2335);
nor U3467 (N_3467,N_2099,N_2597);
and U3468 (N_3468,N_2287,N_2457);
nor U3469 (N_3469,N_1658,N_2539);
or U3470 (N_3470,N_1828,N_2756);
nand U3471 (N_3471,N_1789,N_2535);
nor U3472 (N_3472,N_2655,N_1712);
and U3473 (N_3473,N_2934,N_2774);
nand U3474 (N_3474,N_2208,N_1959);
and U3475 (N_3475,N_2204,N_2714);
nor U3476 (N_3476,N_2356,N_1767);
nor U3477 (N_3477,N_2094,N_2285);
nor U3478 (N_3478,N_2330,N_1673);
or U3479 (N_3479,N_1500,N_1822);
nand U3480 (N_3480,N_2444,N_1750);
nor U3481 (N_3481,N_1811,N_2786);
or U3482 (N_3482,N_2163,N_2040);
nand U3483 (N_3483,N_2247,N_2042);
nand U3484 (N_3484,N_1691,N_1625);
xnor U3485 (N_3485,N_2917,N_2519);
nor U3486 (N_3486,N_1662,N_2124);
nand U3487 (N_3487,N_2563,N_1826);
nand U3488 (N_3488,N_2772,N_2420);
nor U3489 (N_3489,N_2585,N_2395);
and U3490 (N_3490,N_2384,N_1933);
and U3491 (N_3491,N_2605,N_2835);
xnor U3492 (N_3492,N_2684,N_2200);
or U3493 (N_3493,N_1760,N_1756);
or U3494 (N_3494,N_2256,N_2377);
or U3495 (N_3495,N_2971,N_1574);
nand U3496 (N_3496,N_2034,N_2697);
and U3497 (N_3497,N_2376,N_2828);
nand U3498 (N_3498,N_2888,N_1777);
nand U3499 (N_3499,N_2980,N_2483);
or U3500 (N_3500,N_2592,N_2647);
or U3501 (N_3501,N_2879,N_2903);
nor U3502 (N_3502,N_2477,N_1995);
nor U3503 (N_3503,N_2848,N_2345);
and U3504 (N_3504,N_2520,N_2529);
nand U3505 (N_3505,N_1919,N_2470);
nor U3506 (N_3506,N_2619,N_1844);
nand U3507 (N_3507,N_2175,N_1611);
nor U3508 (N_3508,N_2887,N_2138);
or U3509 (N_3509,N_1517,N_1881);
and U3510 (N_3510,N_1820,N_2095);
nor U3511 (N_3511,N_1675,N_2761);
or U3512 (N_3512,N_1523,N_2983);
or U3513 (N_3513,N_2794,N_2129);
or U3514 (N_3514,N_2866,N_2447);
or U3515 (N_3515,N_1974,N_2179);
nand U3516 (N_3516,N_2631,N_1873);
or U3517 (N_3517,N_2297,N_2492);
and U3518 (N_3518,N_1909,N_2915);
and U3519 (N_3519,N_1581,N_1897);
nand U3520 (N_3520,N_2955,N_2746);
nor U3521 (N_3521,N_2712,N_1915);
nor U3522 (N_3522,N_1696,N_2564);
xor U3523 (N_3523,N_1657,N_1615);
nand U3524 (N_3524,N_1513,N_2569);
nand U3525 (N_3525,N_2003,N_2101);
or U3526 (N_3526,N_2565,N_2747);
nand U3527 (N_3527,N_2155,N_2254);
nor U3528 (N_3528,N_1593,N_2918);
and U3529 (N_3529,N_1903,N_2659);
or U3530 (N_3530,N_1721,N_1563);
and U3531 (N_3531,N_1501,N_2878);
nor U3532 (N_3532,N_2541,N_1808);
and U3533 (N_3533,N_1573,N_2654);
nor U3534 (N_3534,N_1889,N_2427);
and U3535 (N_3535,N_2891,N_1803);
nor U3536 (N_3536,N_2051,N_2729);
or U3537 (N_3537,N_2338,N_2328);
and U3538 (N_3538,N_1982,N_2426);
nand U3539 (N_3539,N_1894,N_2562);
and U3540 (N_3540,N_2635,N_2533);
or U3541 (N_3541,N_1937,N_2508);
nand U3542 (N_3542,N_2601,N_2128);
or U3543 (N_3543,N_2125,N_2176);
and U3544 (N_3544,N_2341,N_1866);
nand U3545 (N_3545,N_1510,N_2827);
and U3546 (N_3546,N_2361,N_2788);
nand U3547 (N_3547,N_2490,N_1853);
nor U3548 (N_3548,N_1855,N_2759);
and U3549 (N_3549,N_2745,N_1986);
nor U3550 (N_3550,N_2049,N_2087);
nand U3551 (N_3551,N_2402,N_2394);
and U3552 (N_3552,N_2987,N_2144);
and U3553 (N_3553,N_2136,N_2737);
or U3554 (N_3554,N_2234,N_1800);
or U3555 (N_3555,N_2524,N_2636);
and U3556 (N_3556,N_2552,N_1587);
and U3557 (N_3557,N_2197,N_2063);
or U3558 (N_3558,N_1715,N_1694);
and U3559 (N_3559,N_2240,N_2935);
or U3560 (N_3560,N_2496,N_1726);
nor U3561 (N_3561,N_2832,N_2668);
nand U3562 (N_3562,N_1580,N_1677);
or U3563 (N_3563,N_2841,N_2568);
and U3564 (N_3564,N_2383,N_1654);
and U3565 (N_3565,N_1784,N_2263);
nor U3566 (N_3566,N_2191,N_2904);
nor U3567 (N_3567,N_2135,N_2718);
and U3568 (N_3568,N_1700,N_2188);
or U3569 (N_3569,N_2629,N_2305);
nor U3570 (N_3570,N_1560,N_2248);
nand U3571 (N_3571,N_1906,N_2573);
or U3572 (N_3572,N_2986,N_2467);
nand U3573 (N_3573,N_2414,N_1506);
nor U3574 (N_3574,N_1676,N_2126);
nand U3575 (N_3575,N_2306,N_2959);
xor U3576 (N_3576,N_2212,N_2192);
nand U3577 (N_3577,N_2932,N_2881);
nand U3578 (N_3578,N_2215,N_1972);
nor U3579 (N_3579,N_2272,N_1950);
xnor U3580 (N_3580,N_2178,N_2431);
or U3581 (N_3581,N_2571,N_2777);
nor U3582 (N_3582,N_2961,N_1852);
nor U3583 (N_3583,N_2293,N_2162);
and U3584 (N_3584,N_2021,N_1512);
nor U3585 (N_3585,N_2630,N_1836);
or U3586 (N_3586,N_1697,N_1629);
nor U3587 (N_3587,N_1963,N_1531);
nand U3588 (N_3588,N_1570,N_2958);
nand U3589 (N_3589,N_2152,N_2114);
or U3590 (N_3590,N_2658,N_2153);
xor U3591 (N_3591,N_2784,N_2005);
and U3592 (N_3592,N_2726,N_1519);
nand U3593 (N_3593,N_1741,N_2251);
or U3594 (N_3594,N_2071,N_2553);
nor U3595 (N_3595,N_2499,N_1639);
nand U3596 (N_3596,N_1925,N_1770);
nor U3597 (N_3597,N_1920,N_1827);
and U3598 (N_3598,N_1945,N_2380);
nor U3599 (N_3599,N_1810,N_2028);
nand U3600 (N_3600,N_1533,N_2683);
nand U3601 (N_3601,N_2677,N_2727);
nand U3602 (N_3602,N_2662,N_2397);
or U3603 (N_3603,N_2641,N_1754);
or U3604 (N_3604,N_2203,N_2804);
or U3605 (N_3605,N_1635,N_2782);
or U3606 (N_3606,N_2443,N_2902);
nand U3607 (N_3607,N_2235,N_2190);
nor U3608 (N_3608,N_2966,N_2951);
or U3609 (N_3609,N_1628,N_2237);
nor U3610 (N_3610,N_2719,N_1818);
nor U3611 (N_3611,N_2497,N_2990);
nor U3612 (N_3612,N_2816,N_2045);
nand U3613 (N_3613,N_1805,N_1893);
nand U3614 (N_3614,N_2284,N_1591);
and U3615 (N_3615,N_1549,N_2020);
or U3616 (N_3616,N_1791,N_2822);
nor U3617 (N_3617,N_1883,N_1775);
nand U3618 (N_3618,N_2643,N_2074);
or U3619 (N_3619,N_1539,N_2602);
nand U3620 (N_3620,N_2096,N_2806);
nand U3621 (N_3621,N_2008,N_2994);
and U3622 (N_3622,N_1725,N_2743);
nor U3623 (N_3623,N_2947,N_2262);
nor U3624 (N_3624,N_1759,N_2048);
nor U3625 (N_3625,N_2889,N_1790);
or U3626 (N_3626,N_1927,N_2530);
nor U3627 (N_3627,N_2861,N_2183);
nand U3628 (N_3628,N_2334,N_2579);
nand U3629 (N_3629,N_1669,N_2462);
nor U3630 (N_3630,N_2664,N_1795);
or U3631 (N_3631,N_1578,N_1762);
and U3632 (N_3632,N_1747,N_1890);
nor U3633 (N_3633,N_2127,N_1505);
and U3634 (N_3634,N_2676,N_2501);
nor U3635 (N_3635,N_2039,N_2000);
xor U3636 (N_3636,N_2117,N_1596);
or U3637 (N_3637,N_1783,N_2613);
nor U3638 (N_3638,N_2331,N_2068);
nor U3639 (N_3639,N_2232,N_2500);
nand U3640 (N_3640,N_1830,N_2454);
and U3641 (N_3641,N_2316,N_1948);
or U3642 (N_3642,N_2512,N_2633);
nand U3643 (N_3643,N_1763,N_2741);
nor U3644 (N_3644,N_2481,N_1802);
nor U3645 (N_3645,N_2088,N_2299);
and U3646 (N_3646,N_2513,N_1614);
or U3647 (N_3647,N_2070,N_2382);
or U3648 (N_3648,N_1575,N_2750);
nand U3649 (N_3649,N_2656,N_2644);
or U3650 (N_3650,N_1876,N_2844);
and U3651 (N_3651,N_2456,N_2897);
nor U3652 (N_3652,N_1833,N_1962);
nand U3653 (N_3653,N_2019,N_2054);
or U3654 (N_3654,N_2600,N_2326);
and U3655 (N_3655,N_1850,N_2542);
nand U3656 (N_3656,N_2327,N_1545);
nand U3657 (N_3657,N_1955,N_1729);
or U3658 (N_3658,N_2924,N_2342);
or U3659 (N_3659,N_2445,N_1535);
nand U3660 (N_3660,N_2348,N_2783);
nor U3661 (N_3661,N_2170,N_1806);
or U3662 (N_3662,N_2890,N_2561);
or U3663 (N_3663,N_2754,N_2625);
nor U3664 (N_3664,N_1538,N_2133);
and U3665 (N_3665,N_2970,N_2689);
nor U3666 (N_3666,N_2814,N_2956);
or U3667 (N_3667,N_2675,N_2227);
and U3668 (N_3668,N_2399,N_1861);
and U3669 (N_3669,N_1804,N_2874);
or U3670 (N_3670,N_2277,N_2789);
and U3671 (N_3671,N_1722,N_1773);
nand U3672 (N_3672,N_1858,N_1779);
or U3673 (N_3673,N_1576,N_1744);
and U3674 (N_3674,N_2167,N_1908);
or U3675 (N_3675,N_2526,N_1695);
or U3676 (N_3676,N_2872,N_2309);
and U3677 (N_3677,N_2218,N_2768);
nor U3678 (N_3678,N_2433,N_1812);
and U3679 (N_3679,N_2016,N_2434);
nor U3680 (N_3680,N_2516,N_1951);
or U3681 (N_3681,N_2895,N_2475);
and U3682 (N_3682,N_1851,N_1557);
nand U3683 (N_3683,N_1902,N_2749);
nand U3684 (N_3684,N_2614,N_1514);
nor U3685 (N_3685,N_2927,N_2333);
nand U3686 (N_3686,N_2556,N_2460);
and U3687 (N_3687,N_1633,N_2829);
nand U3688 (N_3688,N_1709,N_2871);
nor U3689 (N_3689,N_2514,N_2909);
nand U3690 (N_3690,N_1939,N_2355);
and U3691 (N_3691,N_1521,N_2486);
and U3692 (N_3692,N_1559,N_2863);
or U3693 (N_3693,N_2026,N_2865);
nor U3694 (N_3694,N_1569,N_2893);
and U3695 (N_3695,N_2708,N_2035);
nor U3696 (N_3696,N_2703,N_2002);
nor U3697 (N_3697,N_2009,N_1671);
nor U3698 (N_3698,N_2347,N_2311);
nor U3699 (N_3699,N_1585,N_2929);
nand U3700 (N_3700,N_1650,N_2842);
or U3701 (N_3701,N_2999,N_2773);
or U3702 (N_3702,N_2278,N_1998);
nor U3703 (N_3703,N_2694,N_2706);
or U3704 (N_3704,N_1690,N_2981);
nand U3705 (N_3705,N_2610,N_1620);
or U3706 (N_3706,N_2652,N_1930);
nor U3707 (N_3707,N_2681,N_2340);
or U3708 (N_3708,N_2408,N_2282);
nor U3709 (N_3709,N_1761,N_1957);
nand U3710 (N_3710,N_2700,N_2638);
nand U3711 (N_3711,N_2370,N_2479);
and U3712 (N_3712,N_1634,N_1558);
and U3713 (N_3713,N_2926,N_2763);
or U3714 (N_3714,N_1638,N_2038);
nor U3715 (N_3715,N_2858,N_1849);
xor U3716 (N_3716,N_2495,N_1891);
nor U3717 (N_3717,N_1751,N_2461);
nor U3718 (N_3718,N_1785,N_2069);
nor U3719 (N_3719,N_2963,N_2693);
nor U3720 (N_3720,N_2229,N_2957);
and U3721 (N_3721,N_1503,N_2967);
nor U3722 (N_3722,N_2938,N_2586);
nand U3723 (N_3723,N_2449,N_2699);
nor U3724 (N_3724,N_1719,N_1780);
nand U3725 (N_3725,N_1525,N_2047);
and U3726 (N_3726,N_2440,N_2796);
or U3727 (N_3727,N_1664,N_2896);
and U3728 (N_3728,N_1984,N_2180);
nand U3729 (N_3729,N_1561,N_1778);
nand U3730 (N_3730,N_1913,N_1708);
nor U3731 (N_3731,N_2439,N_2312);
nand U3732 (N_3732,N_2428,N_2466);
nor U3733 (N_3733,N_2148,N_2217);
nor U3734 (N_3734,N_2209,N_2065);
and U3735 (N_3735,N_1630,N_1644);
nor U3736 (N_3736,N_1565,N_2156);
or U3737 (N_3737,N_2409,N_1904);
nor U3738 (N_3738,N_2502,N_2757);
and U3739 (N_3739,N_2691,N_1685);
and U3740 (N_3740,N_2480,N_2368);
nand U3741 (N_3741,N_1605,N_1832);
nand U3742 (N_3742,N_2933,N_2364);
or U3743 (N_3743,N_2107,N_1680);
nand U3744 (N_3744,N_2199,N_2588);
nor U3745 (N_3745,N_1878,N_1660);
and U3746 (N_3746,N_2182,N_2732);
or U3747 (N_3747,N_2053,N_2013);
nand U3748 (N_3748,N_1642,N_2220);
nor U3749 (N_3749,N_2919,N_2748);
nand U3750 (N_3750,N_1577,N_2193);
and U3751 (N_3751,N_2603,N_1635);
nor U3752 (N_3752,N_1949,N_2360);
nor U3753 (N_3753,N_2800,N_1747);
nor U3754 (N_3754,N_1520,N_2852);
nand U3755 (N_3755,N_1904,N_2873);
nand U3756 (N_3756,N_1922,N_2472);
and U3757 (N_3757,N_2856,N_2748);
or U3758 (N_3758,N_1717,N_1999);
or U3759 (N_3759,N_2321,N_2368);
and U3760 (N_3760,N_2173,N_2634);
nor U3761 (N_3761,N_2940,N_2101);
and U3762 (N_3762,N_2561,N_1847);
nand U3763 (N_3763,N_1809,N_2335);
and U3764 (N_3764,N_1693,N_1572);
nor U3765 (N_3765,N_2640,N_2176);
or U3766 (N_3766,N_2278,N_2323);
or U3767 (N_3767,N_2416,N_2813);
or U3768 (N_3768,N_1601,N_1514);
and U3769 (N_3769,N_2666,N_2417);
and U3770 (N_3770,N_2434,N_1563);
nand U3771 (N_3771,N_2566,N_1535);
or U3772 (N_3772,N_1904,N_2164);
xnor U3773 (N_3773,N_2699,N_1542);
nor U3774 (N_3774,N_1884,N_2569);
or U3775 (N_3775,N_2115,N_2599);
nand U3776 (N_3776,N_2421,N_2387);
and U3777 (N_3777,N_1755,N_1843);
nand U3778 (N_3778,N_1598,N_2327);
nand U3779 (N_3779,N_2611,N_2260);
and U3780 (N_3780,N_2243,N_2661);
nand U3781 (N_3781,N_1948,N_1584);
or U3782 (N_3782,N_1783,N_1955);
nor U3783 (N_3783,N_1847,N_2048);
or U3784 (N_3784,N_2093,N_1917);
nor U3785 (N_3785,N_2726,N_2593);
nand U3786 (N_3786,N_2502,N_2619);
nor U3787 (N_3787,N_2332,N_1653);
nor U3788 (N_3788,N_1526,N_2907);
nor U3789 (N_3789,N_1882,N_1505);
nor U3790 (N_3790,N_2743,N_1682);
and U3791 (N_3791,N_1973,N_2789);
nor U3792 (N_3792,N_2568,N_1509);
nor U3793 (N_3793,N_2565,N_1699);
nand U3794 (N_3794,N_1789,N_2864);
and U3795 (N_3795,N_1734,N_1737);
nor U3796 (N_3796,N_2562,N_1988);
nor U3797 (N_3797,N_1550,N_2507);
nor U3798 (N_3798,N_1615,N_2276);
or U3799 (N_3799,N_1734,N_2027);
xnor U3800 (N_3800,N_2593,N_2666);
nor U3801 (N_3801,N_1954,N_2417);
nand U3802 (N_3802,N_2052,N_2765);
nor U3803 (N_3803,N_2680,N_2471);
or U3804 (N_3804,N_1961,N_1609);
xor U3805 (N_3805,N_2677,N_1855);
nor U3806 (N_3806,N_1985,N_1818);
and U3807 (N_3807,N_1610,N_2103);
and U3808 (N_3808,N_1874,N_2834);
or U3809 (N_3809,N_2837,N_2359);
and U3810 (N_3810,N_2190,N_2304);
or U3811 (N_3811,N_1953,N_2148);
nor U3812 (N_3812,N_2037,N_2081);
nand U3813 (N_3813,N_2615,N_2980);
and U3814 (N_3814,N_1561,N_2767);
or U3815 (N_3815,N_1916,N_2495);
nor U3816 (N_3816,N_2623,N_1864);
nand U3817 (N_3817,N_2133,N_2665);
nor U3818 (N_3818,N_2587,N_2458);
nand U3819 (N_3819,N_1543,N_2990);
and U3820 (N_3820,N_2862,N_2575);
or U3821 (N_3821,N_2273,N_1816);
and U3822 (N_3822,N_2479,N_1537);
or U3823 (N_3823,N_1588,N_2825);
nand U3824 (N_3824,N_1595,N_2925);
nand U3825 (N_3825,N_2977,N_1594);
nand U3826 (N_3826,N_2424,N_2219);
or U3827 (N_3827,N_2350,N_1947);
xor U3828 (N_3828,N_2844,N_1644);
nand U3829 (N_3829,N_1730,N_2724);
or U3830 (N_3830,N_2188,N_1968);
nor U3831 (N_3831,N_2765,N_2857);
nor U3832 (N_3832,N_2349,N_2906);
and U3833 (N_3833,N_1954,N_1581);
or U3834 (N_3834,N_2852,N_2342);
or U3835 (N_3835,N_2673,N_2124);
or U3836 (N_3836,N_1710,N_1919);
or U3837 (N_3837,N_1861,N_2514);
nand U3838 (N_3838,N_2860,N_2712);
or U3839 (N_3839,N_2640,N_2408);
nand U3840 (N_3840,N_2193,N_1592);
or U3841 (N_3841,N_1731,N_2161);
or U3842 (N_3842,N_2085,N_1630);
or U3843 (N_3843,N_1546,N_1606);
nand U3844 (N_3844,N_1508,N_2078);
or U3845 (N_3845,N_2706,N_2815);
and U3846 (N_3846,N_2627,N_2242);
nand U3847 (N_3847,N_2882,N_1786);
and U3848 (N_3848,N_2251,N_1904);
or U3849 (N_3849,N_2398,N_2052);
nand U3850 (N_3850,N_1825,N_2587);
xnor U3851 (N_3851,N_1610,N_2303);
nand U3852 (N_3852,N_2754,N_1554);
nor U3853 (N_3853,N_2716,N_1665);
and U3854 (N_3854,N_2698,N_2136);
or U3855 (N_3855,N_2082,N_2889);
and U3856 (N_3856,N_2125,N_1997);
or U3857 (N_3857,N_2363,N_1500);
or U3858 (N_3858,N_1576,N_2624);
nand U3859 (N_3859,N_1919,N_2363);
nor U3860 (N_3860,N_2405,N_2291);
and U3861 (N_3861,N_2320,N_2887);
or U3862 (N_3862,N_1755,N_2399);
and U3863 (N_3863,N_2523,N_1823);
and U3864 (N_3864,N_1664,N_1636);
nor U3865 (N_3865,N_2090,N_1736);
and U3866 (N_3866,N_2637,N_2202);
or U3867 (N_3867,N_2943,N_2557);
nand U3868 (N_3868,N_2837,N_1538);
nor U3869 (N_3869,N_1736,N_2798);
nand U3870 (N_3870,N_1685,N_1872);
or U3871 (N_3871,N_2688,N_2889);
or U3872 (N_3872,N_2659,N_2564);
or U3873 (N_3873,N_2562,N_1629);
nor U3874 (N_3874,N_2393,N_2811);
and U3875 (N_3875,N_1963,N_1639);
or U3876 (N_3876,N_2445,N_2810);
nand U3877 (N_3877,N_2517,N_1508);
or U3878 (N_3878,N_2510,N_2303);
and U3879 (N_3879,N_2550,N_2476);
or U3880 (N_3880,N_2063,N_1764);
nor U3881 (N_3881,N_2209,N_2583);
nand U3882 (N_3882,N_2859,N_2231);
nand U3883 (N_3883,N_1756,N_2177);
nor U3884 (N_3884,N_1522,N_1630);
nor U3885 (N_3885,N_1874,N_1559);
xnor U3886 (N_3886,N_1964,N_1664);
nand U3887 (N_3887,N_1814,N_1576);
nand U3888 (N_3888,N_2690,N_1882);
nand U3889 (N_3889,N_2338,N_2436);
nor U3890 (N_3890,N_1659,N_2523);
nor U3891 (N_3891,N_1575,N_2565);
nand U3892 (N_3892,N_2752,N_2199);
nor U3893 (N_3893,N_1510,N_1695);
nand U3894 (N_3894,N_2175,N_1787);
nor U3895 (N_3895,N_1765,N_2687);
nand U3896 (N_3896,N_2420,N_2471);
xnor U3897 (N_3897,N_1838,N_1648);
xor U3898 (N_3898,N_2273,N_2750);
or U3899 (N_3899,N_2476,N_2776);
nand U3900 (N_3900,N_2112,N_2815);
and U3901 (N_3901,N_1674,N_1879);
nor U3902 (N_3902,N_2569,N_2631);
or U3903 (N_3903,N_1505,N_2136);
nor U3904 (N_3904,N_2999,N_2769);
nand U3905 (N_3905,N_2720,N_1580);
nor U3906 (N_3906,N_2988,N_2543);
nand U3907 (N_3907,N_1502,N_1529);
nor U3908 (N_3908,N_1952,N_1757);
nand U3909 (N_3909,N_2016,N_1853);
nor U3910 (N_3910,N_2636,N_1526);
and U3911 (N_3911,N_1728,N_2867);
nor U3912 (N_3912,N_1777,N_2788);
or U3913 (N_3913,N_1649,N_2348);
and U3914 (N_3914,N_2735,N_2164);
nand U3915 (N_3915,N_2677,N_2828);
or U3916 (N_3916,N_2472,N_1812);
or U3917 (N_3917,N_1740,N_2716);
or U3918 (N_3918,N_2783,N_2394);
or U3919 (N_3919,N_2547,N_1778);
nand U3920 (N_3920,N_1708,N_1998);
nand U3921 (N_3921,N_1622,N_2363);
nand U3922 (N_3922,N_1604,N_2071);
or U3923 (N_3923,N_1816,N_1928);
and U3924 (N_3924,N_1655,N_1997);
or U3925 (N_3925,N_2033,N_2097);
nand U3926 (N_3926,N_2829,N_2272);
nand U3927 (N_3927,N_2681,N_2295);
or U3928 (N_3928,N_1874,N_2336);
or U3929 (N_3929,N_1759,N_2974);
or U3930 (N_3930,N_1953,N_2366);
nor U3931 (N_3931,N_2950,N_2344);
nand U3932 (N_3932,N_2608,N_1586);
nor U3933 (N_3933,N_2606,N_2730);
or U3934 (N_3934,N_1647,N_2030);
or U3935 (N_3935,N_1653,N_2123);
nor U3936 (N_3936,N_2840,N_2554);
nor U3937 (N_3937,N_1841,N_2463);
or U3938 (N_3938,N_2729,N_2653);
or U3939 (N_3939,N_2932,N_2506);
nor U3940 (N_3940,N_2199,N_2099);
nor U3941 (N_3941,N_1842,N_2007);
and U3942 (N_3942,N_2056,N_2823);
nand U3943 (N_3943,N_2868,N_2020);
or U3944 (N_3944,N_2055,N_2935);
nand U3945 (N_3945,N_2580,N_2197);
and U3946 (N_3946,N_2932,N_2943);
or U3947 (N_3947,N_2520,N_2918);
and U3948 (N_3948,N_1592,N_2595);
nor U3949 (N_3949,N_1545,N_2883);
nor U3950 (N_3950,N_1508,N_1932);
nand U3951 (N_3951,N_2721,N_1612);
or U3952 (N_3952,N_2190,N_2807);
or U3953 (N_3953,N_1507,N_1564);
nor U3954 (N_3954,N_2759,N_2278);
nand U3955 (N_3955,N_1821,N_2079);
nand U3956 (N_3956,N_2655,N_2924);
xnor U3957 (N_3957,N_1549,N_1614);
nand U3958 (N_3958,N_2318,N_2455);
nor U3959 (N_3959,N_1582,N_2497);
and U3960 (N_3960,N_2805,N_2109);
or U3961 (N_3961,N_2854,N_2330);
or U3962 (N_3962,N_2409,N_2094);
nand U3963 (N_3963,N_2574,N_2354);
nor U3964 (N_3964,N_1524,N_1542);
nand U3965 (N_3965,N_2531,N_2920);
xor U3966 (N_3966,N_2708,N_2829);
and U3967 (N_3967,N_1570,N_2043);
nor U3968 (N_3968,N_2000,N_2571);
nor U3969 (N_3969,N_2153,N_2365);
nand U3970 (N_3970,N_2204,N_2377);
or U3971 (N_3971,N_1995,N_2325);
nand U3972 (N_3972,N_2258,N_2882);
nor U3973 (N_3973,N_1672,N_2980);
nand U3974 (N_3974,N_2478,N_1642);
or U3975 (N_3975,N_2179,N_2877);
or U3976 (N_3976,N_2074,N_2815);
or U3977 (N_3977,N_1605,N_1970);
nand U3978 (N_3978,N_2988,N_1608);
or U3979 (N_3979,N_2933,N_2133);
nand U3980 (N_3980,N_2476,N_2044);
nand U3981 (N_3981,N_2664,N_1985);
or U3982 (N_3982,N_1781,N_2243);
or U3983 (N_3983,N_2405,N_2461);
or U3984 (N_3984,N_2991,N_1549);
or U3985 (N_3985,N_2341,N_2780);
nor U3986 (N_3986,N_2521,N_2150);
or U3987 (N_3987,N_2484,N_2493);
or U3988 (N_3988,N_2303,N_1533);
nand U3989 (N_3989,N_2667,N_2026);
nand U3990 (N_3990,N_2176,N_2591);
and U3991 (N_3991,N_2795,N_1562);
and U3992 (N_3992,N_2215,N_2134);
nand U3993 (N_3993,N_2166,N_1657);
xor U3994 (N_3994,N_2554,N_2729);
nor U3995 (N_3995,N_2662,N_2856);
nand U3996 (N_3996,N_2184,N_2396);
nor U3997 (N_3997,N_2393,N_2854);
nand U3998 (N_3998,N_2825,N_2968);
and U3999 (N_3999,N_2582,N_2380);
and U4000 (N_4000,N_1840,N_2027);
and U4001 (N_4001,N_2308,N_2379);
nand U4002 (N_4002,N_2339,N_2404);
and U4003 (N_4003,N_1520,N_1926);
nor U4004 (N_4004,N_2396,N_2466);
nor U4005 (N_4005,N_2835,N_2077);
xnor U4006 (N_4006,N_1926,N_2810);
or U4007 (N_4007,N_2058,N_2690);
and U4008 (N_4008,N_2452,N_2192);
and U4009 (N_4009,N_2701,N_1771);
or U4010 (N_4010,N_1590,N_1682);
nand U4011 (N_4011,N_1633,N_1872);
xnor U4012 (N_4012,N_2218,N_1805);
and U4013 (N_4013,N_2129,N_2132);
or U4014 (N_4014,N_2586,N_1808);
nor U4015 (N_4015,N_2439,N_1513);
and U4016 (N_4016,N_2212,N_1972);
and U4017 (N_4017,N_2669,N_1768);
and U4018 (N_4018,N_2644,N_1877);
nor U4019 (N_4019,N_1575,N_2546);
nand U4020 (N_4020,N_1930,N_2230);
nor U4021 (N_4021,N_1937,N_2566);
or U4022 (N_4022,N_2781,N_1650);
nand U4023 (N_4023,N_2893,N_2011);
nand U4024 (N_4024,N_1937,N_2132);
nand U4025 (N_4025,N_1900,N_2431);
and U4026 (N_4026,N_1794,N_2646);
nor U4027 (N_4027,N_2694,N_2743);
nand U4028 (N_4028,N_2507,N_1937);
or U4029 (N_4029,N_1859,N_2614);
and U4030 (N_4030,N_1501,N_1964);
or U4031 (N_4031,N_1524,N_2003);
nor U4032 (N_4032,N_2789,N_1530);
nor U4033 (N_4033,N_2234,N_2260);
and U4034 (N_4034,N_2611,N_2591);
nand U4035 (N_4035,N_2531,N_2806);
nand U4036 (N_4036,N_2136,N_2975);
nand U4037 (N_4037,N_2944,N_2412);
nor U4038 (N_4038,N_2628,N_2316);
nand U4039 (N_4039,N_2363,N_2007);
or U4040 (N_4040,N_1514,N_2806);
nand U4041 (N_4041,N_2698,N_2908);
or U4042 (N_4042,N_2025,N_2017);
and U4043 (N_4043,N_1602,N_2284);
and U4044 (N_4044,N_1553,N_2587);
nand U4045 (N_4045,N_2805,N_2316);
or U4046 (N_4046,N_2088,N_1616);
nand U4047 (N_4047,N_2466,N_2790);
nand U4048 (N_4048,N_1643,N_2380);
xor U4049 (N_4049,N_1940,N_2656);
nor U4050 (N_4050,N_2316,N_2017);
and U4051 (N_4051,N_2457,N_1748);
and U4052 (N_4052,N_2593,N_2716);
nor U4053 (N_4053,N_2545,N_2937);
or U4054 (N_4054,N_2087,N_2929);
nand U4055 (N_4055,N_2412,N_1926);
or U4056 (N_4056,N_1952,N_2134);
xnor U4057 (N_4057,N_2427,N_2458);
nor U4058 (N_4058,N_2420,N_1974);
and U4059 (N_4059,N_1713,N_2303);
and U4060 (N_4060,N_1668,N_2458);
nand U4061 (N_4061,N_1553,N_2076);
nor U4062 (N_4062,N_1763,N_2012);
nand U4063 (N_4063,N_1816,N_2040);
and U4064 (N_4064,N_2340,N_2707);
nand U4065 (N_4065,N_2372,N_2832);
nor U4066 (N_4066,N_2674,N_2513);
nand U4067 (N_4067,N_1726,N_1938);
and U4068 (N_4068,N_2160,N_1846);
or U4069 (N_4069,N_1520,N_1875);
and U4070 (N_4070,N_2789,N_1826);
nand U4071 (N_4071,N_2310,N_2685);
and U4072 (N_4072,N_1961,N_1909);
and U4073 (N_4073,N_1656,N_1699);
nand U4074 (N_4074,N_2358,N_2789);
nand U4075 (N_4075,N_2182,N_1543);
or U4076 (N_4076,N_2024,N_2200);
or U4077 (N_4077,N_1927,N_2082);
or U4078 (N_4078,N_2406,N_2511);
and U4079 (N_4079,N_2632,N_2532);
or U4080 (N_4080,N_2976,N_1616);
nor U4081 (N_4081,N_1887,N_2586);
or U4082 (N_4082,N_2936,N_2763);
nand U4083 (N_4083,N_1928,N_1926);
nor U4084 (N_4084,N_1707,N_2618);
nor U4085 (N_4085,N_1735,N_2150);
xor U4086 (N_4086,N_2168,N_1745);
and U4087 (N_4087,N_2495,N_2636);
nor U4088 (N_4088,N_1946,N_2664);
and U4089 (N_4089,N_2224,N_1798);
and U4090 (N_4090,N_2140,N_2351);
and U4091 (N_4091,N_2347,N_2180);
nor U4092 (N_4092,N_1561,N_2315);
nand U4093 (N_4093,N_1766,N_1616);
nand U4094 (N_4094,N_2508,N_2048);
nand U4095 (N_4095,N_1649,N_2209);
or U4096 (N_4096,N_2385,N_2513);
nand U4097 (N_4097,N_2927,N_2975);
and U4098 (N_4098,N_2160,N_2882);
or U4099 (N_4099,N_2525,N_2681);
or U4100 (N_4100,N_2030,N_2372);
or U4101 (N_4101,N_1784,N_2226);
nor U4102 (N_4102,N_2238,N_1587);
nor U4103 (N_4103,N_2427,N_2242);
nand U4104 (N_4104,N_2753,N_2072);
and U4105 (N_4105,N_1567,N_2058);
and U4106 (N_4106,N_2190,N_2623);
nand U4107 (N_4107,N_2642,N_2088);
or U4108 (N_4108,N_1710,N_2035);
or U4109 (N_4109,N_1592,N_2766);
nand U4110 (N_4110,N_2406,N_2870);
xnor U4111 (N_4111,N_2144,N_2301);
nand U4112 (N_4112,N_2285,N_2066);
nand U4113 (N_4113,N_1915,N_2393);
nor U4114 (N_4114,N_2668,N_1811);
and U4115 (N_4115,N_2791,N_1757);
and U4116 (N_4116,N_1747,N_1881);
or U4117 (N_4117,N_1743,N_2008);
xor U4118 (N_4118,N_2927,N_1622);
and U4119 (N_4119,N_2482,N_2607);
nor U4120 (N_4120,N_2106,N_2014);
nand U4121 (N_4121,N_2980,N_2072);
nor U4122 (N_4122,N_2483,N_2078);
nand U4123 (N_4123,N_2011,N_1897);
or U4124 (N_4124,N_2178,N_2082);
nand U4125 (N_4125,N_1548,N_1817);
and U4126 (N_4126,N_1599,N_2521);
or U4127 (N_4127,N_2253,N_1744);
and U4128 (N_4128,N_2907,N_1580);
or U4129 (N_4129,N_1731,N_1898);
xor U4130 (N_4130,N_2661,N_2726);
and U4131 (N_4131,N_2350,N_1554);
nor U4132 (N_4132,N_2066,N_2377);
nand U4133 (N_4133,N_2506,N_1999);
and U4134 (N_4134,N_1650,N_2100);
and U4135 (N_4135,N_2610,N_2429);
or U4136 (N_4136,N_1852,N_1762);
nand U4137 (N_4137,N_1940,N_2868);
and U4138 (N_4138,N_2369,N_2479);
nor U4139 (N_4139,N_1940,N_1889);
and U4140 (N_4140,N_2503,N_1727);
nor U4141 (N_4141,N_2499,N_2531);
or U4142 (N_4142,N_2549,N_2061);
and U4143 (N_4143,N_1575,N_2250);
and U4144 (N_4144,N_2587,N_2744);
and U4145 (N_4145,N_2738,N_1886);
or U4146 (N_4146,N_1554,N_1993);
or U4147 (N_4147,N_2459,N_1620);
nor U4148 (N_4148,N_2558,N_2466);
and U4149 (N_4149,N_2961,N_1914);
nor U4150 (N_4150,N_2073,N_2130);
nor U4151 (N_4151,N_2443,N_1540);
and U4152 (N_4152,N_2929,N_1713);
nor U4153 (N_4153,N_2424,N_2252);
and U4154 (N_4154,N_1567,N_2037);
nor U4155 (N_4155,N_1532,N_1784);
or U4156 (N_4156,N_2799,N_1821);
xnor U4157 (N_4157,N_1649,N_2732);
or U4158 (N_4158,N_2718,N_1965);
nor U4159 (N_4159,N_1614,N_2177);
or U4160 (N_4160,N_2007,N_2463);
or U4161 (N_4161,N_2163,N_2417);
or U4162 (N_4162,N_2696,N_2572);
and U4163 (N_4163,N_2446,N_1962);
or U4164 (N_4164,N_2204,N_2319);
nor U4165 (N_4165,N_2310,N_1679);
or U4166 (N_4166,N_2784,N_1712);
nor U4167 (N_4167,N_2742,N_2054);
nand U4168 (N_4168,N_2042,N_2412);
nand U4169 (N_4169,N_2934,N_1985);
and U4170 (N_4170,N_2904,N_2872);
and U4171 (N_4171,N_1847,N_2219);
and U4172 (N_4172,N_1592,N_2738);
nor U4173 (N_4173,N_1563,N_2464);
and U4174 (N_4174,N_2107,N_2066);
and U4175 (N_4175,N_2574,N_1906);
or U4176 (N_4176,N_2149,N_1621);
nor U4177 (N_4177,N_1882,N_2032);
and U4178 (N_4178,N_2096,N_2340);
nor U4179 (N_4179,N_2127,N_2453);
nor U4180 (N_4180,N_2689,N_1983);
or U4181 (N_4181,N_1521,N_2634);
or U4182 (N_4182,N_2842,N_2993);
nor U4183 (N_4183,N_2032,N_2596);
and U4184 (N_4184,N_2783,N_2089);
and U4185 (N_4185,N_2403,N_1510);
or U4186 (N_4186,N_1584,N_2432);
or U4187 (N_4187,N_1612,N_2327);
and U4188 (N_4188,N_1729,N_1719);
nor U4189 (N_4189,N_1884,N_2446);
and U4190 (N_4190,N_1548,N_2905);
nor U4191 (N_4191,N_1770,N_2243);
and U4192 (N_4192,N_2924,N_1896);
nor U4193 (N_4193,N_2370,N_2519);
or U4194 (N_4194,N_1858,N_2096);
or U4195 (N_4195,N_2391,N_2460);
and U4196 (N_4196,N_2854,N_2848);
or U4197 (N_4197,N_2177,N_2172);
nand U4198 (N_4198,N_2004,N_2190);
and U4199 (N_4199,N_2552,N_1633);
or U4200 (N_4200,N_1710,N_1691);
or U4201 (N_4201,N_2365,N_1501);
or U4202 (N_4202,N_1866,N_2446);
and U4203 (N_4203,N_1699,N_2749);
xnor U4204 (N_4204,N_2192,N_1740);
or U4205 (N_4205,N_2669,N_2089);
xnor U4206 (N_4206,N_2076,N_2424);
nor U4207 (N_4207,N_1874,N_2061);
or U4208 (N_4208,N_2686,N_1652);
or U4209 (N_4209,N_2393,N_1687);
xor U4210 (N_4210,N_2763,N_2286);
or U4211 (N_4211,N_2350,N_2515);
and U4212 (N_4212,N_1514,N_2405);
nand U4213 (N_4213,N_2518,N_2942);
and U4214 (N_4214,N_2094,N_2063);
nand U4215 (N_4215,N_2547,N_2971);
nand U4216 (N_4216,N_1925,N_2413);
nand U4217 (N_4217,N_2500,N_2627);
and U4218 (N_4218,N_2751,N_1900);
nand U4219 (N_4219,N_1844,N_2339);
nor U4220 (N_4220,N_2668,N_2800);
nand U4221 (N_4221,N_2629,N_1698);
and U4222 (N_4222,N_2942,N_2163);
xnor U4223 (N_4223,N_2470,N_1938);
or U4224 (N_4224,N_2021,N_1593);
nor U4225 (N_4225,N_2236,N_1526);
and U4226 (N_4226,N_2410,N_2846);
or U4227 (N_4227,N_1890,N_2945);
or U4228 (N_4228,N_2753,N_2956);
or U4229 (N_4229,N_1904,N_1696);
xor U4230 (N_4230,N_2765,N_2647);
or U4231 (N_4231,N_2808,N_2054);
nor U4232 (N_4232,N_1652,N_1917);
or U4233 (N_4233,N_2362,N_2222);
or U4234 (N_4234,N_2373,N_2697);
and U4235 (N_4235,N_1807,N_1797);
or U4236 (N_4236,N_2211,N_1667);
nor U4237 (N_4237,N_2817,N_2500);
nor U4238 (N_4238,N_2339,N_1662);
nor U4239 (N_4239,N_1949,N_2868);
or U4240 (N_4240,N_2223,N_2381);
or U4241 (N_4241,N_1902,N_2193);
or U4242 (N_4242,N_2987,N_1823);
xnor U4243 (N_4243,N_1541,N_1544);
nand U4244 (N_4244,N_1757,N_2305);
and U4245 (N_4245,N_2709,N_2420);
or U4246 (N_4246,N_2686,N_2117);
and U4247 (N_4247,N_2183,N_2860);
nor U4248 (N_4248,N_2596,N_2842);
nand U4249 (N_4249,N_2892,N_2027);
nand U4250 (N_4250,N_2440,N_2342);
and U4251 (N_4251,N_1568,N_1517);
nand U4252 (N_4252,N_1516,N_1933);
or U4253 (N_4253,N_2347,N_1872);
nor U4254 (N_4254,N_2925,N_2680);
nand U4255 (N_4255,N_2264,N_1668);
nor U4256 (N_4256,N_1631,N_2156);
or U4257 (N_4257,N_2128,N_1899);
nand U4258 (N_4258,N_2810,N_1912);
or U4259 (N_4259,N_2517,N_1939);
nor U4260 (N_4260,N_2806,N_2408);
or U4261 (N_4261,N_1786,N_1980);
nor U4262 (N_4262,N_2641,N_2171);
xnor U4263 (N_4263,N_1578,N_2246);
and U4264 (N_4264,N_1697,N_2656);
nor U4265 (N_4265,N_2783,N_2362);
nor U4266 (N_4266,N_2253,N_2500);
and U4267 (N_4267,N_2954,N_2818);
or U4268 (N_4268,N_2619,N_2990);
nand U4269 (N_4269,N_2767,N_2191);
and U4270 (N_4270,N_2855,N_1620);
and U4271 (N_4271,N_2236,N_1538);
nor U4272 (N_4272,N_2864,N_1592);
and U4273 (N_4273,N_1694,N_1958);
nor U4274 (N_4274,N_2581,N_1889);
or U4275 (N_4275,N_2391,N_2832);
nand U4276 (N_4276,N_2938,N_1675);
or U4277 (N_4277,N_2705,N_2101);
and U4278 (N_4278,N_2796,N_2865);
and U4279 (N_4279,N_2667,N_2017);
or U4280 (N_4280,N_2922,N_2811);
nor U4281 (N_4281,N_2353,N_1706);
nand U4282 (N_4282,N_2374,N_2799);
or U4283 (N_4283,N_2988,N_1594);
nand U4284 (N_4284,N_2364,N_1705);
nor U4285 (N_4285,N_1625,N_1554);
xor U4286 (N_4286,N_2869,N_2367);
nand U4287 (N_4287,N_1553,N_2745);
nor U4288 (N_4288,N_2839,N_2952);
nand U4289 (N_4289,N_2214,N_2071);
nand U4290 (N_4290,N_2858,N_2391);
nand U4291 (N_4291,N_1650,N_2435);
nor U4292 (N_4292,N_1771,N_2915);
or U4293 (N_4293,N_1918,N_1823);
nor U4294 (N_4294,N_2679,N_2425);
or U4295 (N_4295,N_2985,N_1653);
nand U4296 (N_4296,N_1910,N_1500);
nor U4297 (N_4297,N_2528,N_2243);
or U4298 (N_4298,N_2439,N_1812);
or U4299 (N_4299,N_2988,N_2268);
or U4300 (N_4300,N_1503,N_2304);
xnor U4301 (N_4301,N_1976,N_1843);
and U4302 (N_4302,N_2099,N_2884);
or U4303 (N_4303,N_1669,N_2665);
and U4304 (N_4304,N_2293,N_1974);
or U4305 (N_4305,N_1875,N_2948);
and U4306 (N_4306,N_1989,N_2237);
and U4307 (N_4307,N_2479,N_2455);
or U4308 (N_4308,N_1571,N_2150);
nor U4309 (N_4309,N_1711,N_2461);
nor U4310 (N_4310,N_2306,N_2122);
or U4311 (N_4311,N_2734,N_1579);
nor U4312 (N_4312,N_2652,N_2237);
and U4313 (N_4313,N_2617,N_2374);
and U4314 (N_4314,N_1660,N_2512);
nor U4315 (N_4315,N_2864,N_2205);
or U4316 (N_4316,N_1895,N_2580);
or U4317 (N_4317,N_1864,N_1967);
or U4318 (N_4318,N_1891,N_2436);
or U4319 (N_4319,N_2482,N_1757);
nand U4320 (N_4320,N_2311,N_2968);
nor U4321 (N_4321,N_2061,N_2207);
and U4322 (N_4322,N_2265,N_2763);
and U4323 (N_4323,N_1956,N_2375);
and U4324 (N_4324,N_2694,N_2393);
or U4325 (N_4325,N_2185,N_2674);
and U4326 (N_4326,N_1996,N_1734);
and U4327 (N_4327,N_1984,N_2233);
or U4328 (N_4328,N_2812,N_2524);
or U4329 (N_4329,N_1766,N_2777);
nand U4330 (N_4330,N_2791,N_1732);
or U4331 (N_4331,N_1537,N_2287);
or U4332 (N_4332,N_1824,N_2691);
nand U4333 (N_4333,N_2170,N_2750);
nand U4334 (N_4334,N_2307,N_1689);
and U4335 (N_4335,N_2600,N_1912);
nor U4336 (N_4336,N_1919,N_2465);
nor U4337 (N_4337,N_2375,N_1796);
nand U4338 (N_4338,N_2500,N_2350);
nand U4339 (N_4339,N_1955,N_2018);
or U4340 (N_4340,N_2329,N_1770);
nor U4341 (N_4341,N_2379,N_2122);
xor U4342 (N_4342,N_2313,N_2945);
nor U4343 (N_4343,N_2284,N_2015);
and U4344 (N_4344,N_2684,N_1718);
nand U4345 (N_4345,N_1606,N_1570);
nor U4346 (N_4346,N_1547,N_2906);
nand U4347 (N_4347,N_2512,N_2037);
nand U4348 (N_4348,N_1827,N_2407);
and U4349 (N_4349,N_2732,N_2313);
and U4350 (N_4350,N_2564,N_1973);
or U4351 (N_4351,N_1627,N_1855);
and U4352 (N_4352,N_2902,N_2940);
nand U4353 (N_4353,N_1670,N_1939);
and U4354 (N_4354,N_1965,N_2213);
and U4355 (N_4355,N_2483,N_1798);
nor U4356 (N_4356,N_2088,N_2849);
or U4357 (N_4357,N_1582,N_2109);
nor U4358 (N_4358,N_2052,N_1567);
and U4359 (N_4359,N_2731,N_2467);
and U4360 (N_4360,N_1679,N_2791);
or U4361 (N_4361,N_1837,N_2842);
nor U4362 (N_4362,N_1604,N_2266);
xnor U4363 (N_4363,N_1696,N_2683);
and U4364 (N_4364,N_1994,N_1654);
and U4365 (N_4365,N_2841,N_2202);
or U4366 (N_4366,N_2221,N_1893);
or U4367 (N_4367,N_2910,N_2248);
or U4368 (N_4368,N_1795,N_2354);
and U4369 (N_4369,N_2438,N_2801);
or U4370 (N_4370,N_2935,N_1756);
nand U4371 (N_4371,N_2399,N_2951);
and U4372 (N_4372,N_1879,N_2128);
or U4373 (N_4373,N_1764,N_2191);
nor U4374 (N_4374,N_1660,N_2148);
nand U4375 (N_4375,N_1985,N_1715);
nor U4376 (N_4376,N_2434,N_2033);
nor U4377 (N_4377,N_1503,N_2475);
nand U4378 (N_4378,N_2004,N_2924);
or U4379 (N_4379,N_2384,N_2580);
xnor U4380 (N_4380,N_2620,N_1706);
and U4381 (N_4381,N_2340,N_2935);
nand U4382 (N_4382,N_2710,N_2984);
or U4383 (N_4383,N_2583,N_2354);
or U4384 (N_4384,N_1617,N_2880);
or U4385 (N_4385,N_2179,N_2826);
nor U4386 (N_4386,N_1947,N_2666);
nor U4387 (N_4387,N_1755,N_2284);
or U4388 (N_4388,N_2839,N_2877);
nor U4389 (N_4389,N_1918,N_2722);
or U4390 (N_4390,N_2594,N_1687);
nor U4391 (N_4391,N_2976,N_2670);
or U4392 (N_4392,N_2702,N_1648);
nand U4393 (N_4393,N_2698,N_2646);
nor U4394 (N_4394,N_2355,N_2845);
nand U4395 (N_4395,N_1690,N_1508);
nor U4396 (N_4396,N_2464,N_2728);
and U4397 (N_4397,N_2505,N_2606);
or U4398 (N_4398,N_2254,N_2522);
nor U4399 (N_4399,N_1500,N_2629);
nor U4400 (N_4400,N_2283,N_2406);
or U4401 (N_4401,N_2935,N_2778);
or U4402 (N_4402,N_2199,N_1924);
xor U4403 (N_4403,N_2973,N_2838);
nor U4404 (N_4404,N_1962,N_2874);
and U4405 (N_4405,N_2820,N_1844);
or U4406 (N_4406,N_2583,N_2930);
or U4407 (N_4407,N_1516,N_1605);
nand U4408 (N_4408,N_1899,N_2724);
nor U4409 (N_4409,N_2076,N_2626);
nor U4410 (N_4410,N_2383,N_2941);
or U4411 (N_4411,N_2887,N_2323);
nor U4412 (N_4412,N_1762,N_2206);
and U4413 (N_4413,N_1637,N_2980);
nor U4414 (N_4414,N_2285,N_1776);
or U4415 (N_4415,N_2761,N_2063);
and U4416 (N_4416,N_1618,N_2352);
nand U4417 (N_4417,N_1525,N_2885);
xnor U4418 (N_4418,N_1868,N_1768);
or U4419 (N_4419,N_2812,N_2834);
nand U4420 (N_4420,N_2431,N_2330);
nand U4421 (N_4421,N_2296,N_1723);
and U4422 (N_4422,N_1940,N_1926);
or U4423 (N_4423,N_1868,N_1860);
and U4424 (N_4424,N_2219,N_1854);
nor U4425 (N_4425,N_1982,N_1804);
nand U4426 (N_4426,N_1612,N_2034);
xnor U4427 (N_4427,N_1673,N_1743);
or U4428 (N_4428,N_2670,N_1993);
nand U4429 (N_4429,N_2458,N_2486);
and U4430 (N_4430,N_1970,N_1984);
nor U4431 (N_4431,N_1909,N_2188);
nand U4432 (N_4432,N_1876,N_2813);
xnor U4433 (N_4433,N_1649,N_2713);
or U4434 (N_4434,N_2990,N_1952);
nor U4435 (N_4435,N_1505,N_2638);
or U4436 (N_4436,N_2477,N_1574);
or U4437 (N_4437,N_1848,N_1948);
or U4438 (N_4438,N_1897,N_1750);
nor U4439 (N_4439,N_2541,N_2222);
and U4440 (N_4440,N_2008,N_2144);
or U4441 (N_4441,N_2372,N_2484);
nand U4442 (N_4442,N_2302,N_2380);
nand U4443 (N_4443,N_2518,N_2188);
or U4444 (N_4444,N_2015,N_1768);
nor U4445 (N_4445,N_2239,N_1734);
nand U4446 (N_4446,N_2067,N_1936);
nor U4447 (N_4447,N_1941,N_1829);
and U4448 (N_4448,N_1531,N_1700);
nor U4449 (N_4449,N_2100,N_2726);
and U4450 (N_4450,N_2155,N_2166);
or U4451 (N_4451,N_2345,N_1958);
nand U4452 (N_4452,N_2119,N_1953);
nand U4453 (N_4453,N_1914,N_2987);
nand U4454 (N_4454,N_2880,N_2112);
nor U4455 (N_4455,N_2799,N_2476);
nor U4456 (N_4456,N_2855,N_2794);
nor U4457 (N_4457,N_2374,N_1637);
or U4458 (N_4458,N_2828,N_1971);
nor U4459 (N_4459,N_2932,N_1578);
or U4460 (N_4460,N_2837,N_1556);
nand U4461 (N_4461,N_2250,N_1777);
and U4462 (N_4462,N_1792,N_1922);
nand U4463 (N_4463,N_1538,N_1738);
and U4464 (N_4464,N_1517,N_2225);
nor U4465 (N_4465,N_2891,N_1548);
nand U4466 (N_4466,N_1889,N_2922);
and U4467 (N_4467,N_1941,N_1504);
or U4468 (N_4468,N_1890,N_2231);
and U4469 (N_4469,N_1988,N_2652);
nor U4470 (N_4470,N_2391,N_2121);
and U4471 (N_4471,N_2404,N_1923);
xnor U4472 (N_4472,N_1961,N_1578);
nand U4473 (N_4473,N_2568,N_1745);
or U4474 (N_4474,N_2190,N_2482);
or U4475 (N_4475,N_2365,N_2294);
or U4476 (N_4476,N_2523,N_2307);
nor U4477 (N_4477,N_2498,N_1614);
and U4478 (N_4478,N_2482,N_1927);
and U4479 (N_4479,N_1960,N_2053);
nor U4480 (N_4480,N_2752,N_2532);
and U4481 (N_4481,N_2426,N_2125);
nand U4482 (N_4482,N_2597,N_2915);
and U4483 (N_4483,N_1642,N_1579);
or U4484 (N_4484,N_1798,N_2490);
or U4485 (N_4485,N_2462,N_2135);
or U4486 (N_4486,N_2691,N_2233);
nand U4487 (N_4487,N_2291,N_2756);
and U4488 (N_4488,N_1817,N_1794);
nor U4489 (N_4489,N_1736,N_2264);
nor U4490 (N_4490,N_2721,N_2126);
and U4491 (N_4491,N_1518,N_2908);
nor U4492 (N_4492,N_2336,N_1991);
and U4493 (N_4493,N_2692,N_2347);
and U4494 (N_4494,N_2207,N_1720);
or U4495 (N_4495,N_2492,N_2393);
nand U4496 (N_4496,N_2499,N_2038);
or U4497 (N_4497,N_2871,N_2789);
nor U4498 (N_4498,N_1649,N_2053);
nand U4499 (N_4499,N_1962,N_2688);
and U4500 (N_4500,N_3590,N_3873);
and U4501 (N_4501,N_4494,N_4393);
nor U4502 (N_4502,N_3445,N_4458);
and U4503 (N_4503,N_4209,N_3777);
or U4504 (N_4504,N_3058,N_4235);
nor U4505 (N_4505,N_3377,N_3392);
nand U4506 (N_4506,N_3533,N_3512);
nand U4507 (N_4507,N_4288,N_3783);
nor U4508 (N_4508,N_4077,N_3913);
and U4509 (N_4509,N_4130,N_3492);
nand U4510 (N_4510,N_3004,N_3971);
nor U4511 (N_4511,N_3963,N_3162);
and U4512 (N_4512,N_4182,N_3115);
or U4513 (N_4513,N_3321,N_3060);
and U4514 (N_4514,N_3081,N_3651);
nor U4515 (N_4515,N_4283,N_3928);
nor U4516 (N_4516,N_3523,N_3107);
xor U4517 (N_4517,N_4020,N_4426);
or U4518 (N_4518,N_3704,N_3008);
nand U4519 (N_4519,N_3369,N_4065);
nor U4520 (N_4520,N_3310,N_4059);
and U4521 (N_4521,N_3046,N_3847);
nor U4522 (N_4522,N_3420,N_4286);
nor U4523 (N_4523,N_3840,N_4015);
or U4524 (N_4524,N_3832,N_4388);
and U4525 (N_4525,N_3553,N_4369);
nand U4526 (N_4526,N_4372,N_3750);
nand U4527 (N_4527,N_4166,N_4448);
nand U4528 (N_4528,N_4136,N_3375);
nand U4529 (N_4529,N_3209,N_4128);
nor U4530 (N_4530,N_3159,N_4127);
nand U4531 (N_4531,N_3453,N_3430);
or U4532 (N_4532,N_3902,N_3466);
or U4533 (N_4533,N_3341,N_3603);
nand U4534 (N_4534,N_3338,N_3127);
xor U4535 (N_4535,N_4217,N_3964);
or U4536 (N_4536,N_3614,N_3161);
nand U4537 (N_4537,N_3906,N_3484);
nor U4538 (N_4538,N_3637,N_3677);
nand U4539 (N_4539,N_3988,N_3226);
and U4540 (N_4540,N_3950,N_4213);
or U4541 (N_4541,N_4281,N_3549);
nor U4542 (N_4542,N_3361,N_3569);
and U4543 (N_4543,N_3708,N_3731);
nand U4544 (N_4544,N_3752,N_3176);
nor U4545 (N_4545,N_3979,N_3554);
nor U4546 (N_4546,N_3811,N_4304);
or U4547 (N_4547,N_4186,N_3397);
or U4548 (N_4548,N_3556,N_4463);
or U4549 (N_4549,N_3471,N_3674);
or U4550 (N_4550,N_3507,N_3922);
and U4551 (N_4551,N_3409,N_4107);
and U4552 (N_4552,N_3411,N_3374);
and U4553 (N_4553,N_4353,N_3244);
xnor U4554 (N_4554,N_4267,N_4345);
and U4555 (N_4555,N_3695,N_4334);
and U4556 (N_4556,N_3951,N_4421);
or U4557 (N_4557,N_4265,N_3596);
or U4558 (N_4558,N_3080,N_3742);
or U4559 (N_4559,N_3618,N_3510);
and U4560 (N_4560,N_3932,N_3679);
or U4561 (N_4561,N_3927,N_3770);
or U4562 (N_4562,N_3406,N_3221);
or U4563 (N_4563,N_4483,N_4306);
nand U4564 (N_4564,N_3433,N_3224);
and U4565 (N_4565,N_3359,N_4462);
nor U4566 (N_4566,N_4461,N_3710);
and U4567 (N_4567,N_4432,N_3790);
nand U4568 (N_4568,N_3091,N_3636);
nand U4569 (N_4569,N_3442,N_3855);
nand U4570 (N_4570,N_3942,N_3625);
nand U4571 (N_4571,N_4338,N_4366);
nand U4572 (N_4572,N_3707,N_4208);
or U4573 (N_4573,N_3875,N_3588);
nor U4574 (N_4574,N_3681,N_4444);
and U4575 (N_4575,N_4046,N_4332);
and U4576 (N_4576,N_3228,N_3427);
nor U4577 (N_4577,N_3506,N_3144);
or U4578 (N_4578,N_4425,N_4001);
nand U4579 (N_4579,N_3938,N_3878);
nor U4580 (N_4580,N_3771,N_3986);
nand U4581 (N_4581,N_3535,N_3388);
nor U4582 (N_4582,N_3308,N_4187);
or U4583 (N_4583,N_3952,N_3468);
nor U4584 (N_4584,N_3945,N_3493);
nor U4585 (N_4585,N_3895,N_4126);
nor U4586 (N_4586,N_4245,N_3068);
and U4587 (N_4587,N_4274,N_3123);
or U4588 (N_4588,N_4105,N_4409);
nor U4589 (N_4589,N_4019,N_3714);
or U4590 (N_4590,N_3311,N_4446);
and U4591 (N_4591,N_3076,N_4460);
nand U4592 (N_4592,N_4358,N_3273);
or U4593 (N_4593,N_3548,N_4493);
nor U4594 (N_4594,N_3086,N_4325);
and U4595 (N_4595,N_3524,N_3142);
and U4596 (N_4596,N_3276,N_3877);
or U4597 (N_4597,N_3562,N_3488);
or U4598 (N_4598,N_3326,N_3269);
nand U4599 (N_4599,N_3872,N_4045);
xnor U4600 (N_4600,N_3935,N_3670);
nor U4601 (N_4601,N_3264,N_3717);
nand U4602 (N_4602,N_3027,N_3051);
nor U4603 (N_4603,N_3190,N_3732);
nand U4604 (N_4604,N_3067,N_3376);
or U4605 (N_4605,N_3546,N_4103);
nand U4606 (N_4606,N_3734,N_3110);
or U4607 (N_4607,N_4148,N_4254);
nand U4608 (N_4608,N_4113,N_3678);
nor U4609 (N_4609,N_4043,N_3331);
xor U4610 (N_4610,N_3421,N_3156);
and U4611 (N_4611,N_4296,N_4453);
nor U4612 (N_4612,N_3786,N_3703);
and U4613 (N_4613,N_3826,N_3059);
and U4614 (N_4614,N_3090,N_3933);
nand U4615 (N_4615,N_3197,N_3911);
or U4616 (N_4616,N_3976,N_3461);
nand U4617 (N_4617,N_3767,N_4007);
nand U4618 (N_4618,N_4106,N_3617);
and U4619 (N_4619,N_3463,N_4496);
xor U4620 (N_4620,N_3093,N_3633);
and U4621 (N_4621,N_4034,N_3040);
nor U4622 (N_4622,N_3381,N_3622);
or U4623 (N_4623,N_4331,N_4029);
and U4624 (N_4624,N_3812,N_4210);
and U4625 (N_4625,N_4144,N_4039);
and U4626 (N_4626,N_3599,N_3712);
nand U4627 (N_4627,N_3275,N_3793);
and U4628 (N_4628,N_3494,N_3036);
nor U4629 (N_4629,N_3281,N_3543);
or U4630 (N_4630,N_3644,N_3440);
and U4631 (N_4631,N_4230,N_3481);
or U4632 (N_4632,N_3020,N_4356);
nor U4633 (N_4633,N_3789,N_3830);
or U4634 (N_4634,N_3843,N_3274);
nor U4635 (N_4635,N_4359,N_3667);
nor U4636 (N_4636,N_3333,N_3045);
nor U4637 (N_4637,N_3073,N_3721);
nor U4638 (N_4638,N_3191,N_3758);
nand U4639 (N_4639,N_3129,N_4112);
and U4640 (N_4640,N_3555,N_4261);
and U4641 (N_4641,N_4134,N_3307);
or U4642 (N_4642,N_3330,N_3682);
nand U4643 (N_4643,N_3470,N_4394);
or U4644 (N_4644,N_3283,N_3684);
nor U4645 (N_4645,N_3836,N_3192);
nor U4646 (N_4646,N_3739,N_3854);
nand U4647 (N_4647,N_4390,N_3859);
nor U4648 (N_4648,N_3043,N_4035);
and U4649 (N_4649,N_4398,N_4347);
nand U4650 (N_4650,N_3738,N_4317);
nor U4651 (N_4651,N_4195,N_4350);
or U4652 (N_4652,N_3993,N_4289);
or U4653 (N_4653,N_4290,N_3200);
or U4654 (N_4654,N_3848,N_3842);
nand U4655 (N_4655,N_3315,N_3921);
or U4656 (N_4656,N_3720,N_3566);
or U4657 (N_4657,N_3038,N_4312);
nor U4658 (N_4658,N_3317,N_4156);
xnor U4659 (N_4659,N_3831,N_3598);
or U4660 (N_4660,N_4455,N_3052);
nor U4661 (N_4661,N_3821,N_4205);
and U4662 (N_4662,N_3671,N_3133);
nor U4663 (N_4663,N_3278,N_4294);
and U4664 (N_4664,N_3939,N_4054);
nand U4665 (N_4665,N_3962,N_3177);
nand U4666 (N_4666,N_4361,N_4420);
nand U4667 (N_4667,N_3019,N_3743);
nor U4668 (N_4668,N_4298,N_4440);
or U4669 (N_4669,N_3905,N_3313);
or U4670 (N_4670,N_4246,N_3595);
nand U4671 (N_4671,N_4164,N_4439);
nor U4672 (N_4672,N_3336,N_4469);
and U4673 (N_4673,N_3711,N_3585);
nor U4674 (N_4674,N_4407,N_3474);
nand U4675 (N_4675,N_3629,N_3893);
nand U4676 (N_4676,N_4087,N_4070);
or U4677 (N_4677,N_3072,N_3353);
and U4678 (N_4678,N_3343,N_4419);
or U4679 (N_4679,N_3582,N_3578);
and U4680 (N_4680,N_3716,N_4081);
or U4681 (N_4681,N_3640,N_3661);
nand U4682 (N_4682,N_3763,N_3458);
or U4683 (N_4683,N_3202,N_3610);
nand U4684 (N_4684,N_3092,N_3815);
nand U4685 (N_4685,N_3672,N_4078);
nor U4686 (N_4686,N_3121,N_4477);
and U4687 (N_4687,N_3356,N_3982);
and U4688 (N_4688,N_4495,N_3607);
xor U4689 (N_4689,N_4049,N_4129);
nand U4690 (N_4690,N_3733,N_4048);
nor U4691 (N_4691,N_3592,N_3655);
nand U4692 (N_4692,N_3113,N_4473);
nor U4693 (N_4693,N_4285,N_3689);
or U4694 (N_4694,N_3220,N_3728);
nand U4695 (N_4695,N_3953,N_3680);
and U4696 (N_4696,N_3163,N_3784);
nor U4697 (N_4697,N_3094,N_3218);
xnor U4698 (N_4698,N_4231,N_3522);
and U4699 (N_4699,N_3865,N_3242);
or U4700 (N_4700,N_3642,N_3627);
nand U4701 (N_4701,N_3340,N_4228);
and U4702 (N_4702,N_4063,N_4275);
nor U4703 (N_4703,N_3062,N_3508);
or U4704 (N_4704,N_3444,N_4189);
nor U4705 (N_4705,N_4486,N_4397);
and U4706 (N_4706,N_3150,N_3550);
and U4707 (N_4707,N_3850,N_4427);
nand U4708 (N_4708,N_4499,N_4023);
xor U4709 (N_4709,N_3407,N_4219);
xnor U4710 (N_4710,N_3424,N_3478);
and U4711 (N_4711,N_4382,N_4423);
and U4712 (N_4712,N_4307,N_4239);
nor U4713 (N_4713,N_3065,N_3926);
or U4714 (N_4714,N_4266,N_4165);
or U4715 (N_4715,N_3233,N_3037);
nand U4716 (N_4716,N_3663,N_4215);
or U4717 (N_4717,N_3247,N_3243);
and U4718 (N_4718,N_4222,N_3455);
and U4719 (N_4719,N_3903,N_3268);
and U4720 (N_4720,N_4279,N_3454);
and U4721 (N_4721,N_4237,N_4472);
nor U4722 (N_4722,N_3542,N_3064);
or U4723 (N_4723,N_3217,N_3529);
or U4724 (N_4724,N_3312,N_3897);
nor U4725 (N_4725,N_3839,N_3885);
or U4726 (N_4726,N_3262,N_3013);
and U4727 (N_4727,N_3074,N_3152);
or U4728 (N_4728,N_4346,N_4027);
nor U4729 (N_4729,N_4056,N_3305);
and U4730 (N_4730,N_4389,N_3309);
nor U4731 (N_4731,N_3143,N_4096);
and U4732 (N_4732,N_3766,N_3955);
nor U4733 (N_4733,N_4280,N_4441);
nand U4734 (N_4734,N_3441,N_3929);
xor U4735 (N_4735,N_3509,N_3146);
and U4736 (N_4736,N_3082,N_3571);
or U4737 (N_4737,N_3560,N_3531);
nand U4738 (N_4738,N_3735,N_4058);
and U4739 (N_4739,N_4102,N_3999);
or U4740 (N_4740,N_3360,N_3213);
nand U4741 (N_4741,N_4211,N_3085);
nor U4742 (N_4742,N_3638,N_4248);
nand U4743 (N_4743,N_4138,N_4158);
nor U4744 (N_4744,N_4308,N_4411);
nand U4745 (N_4745,N_3547,N_3722);
and U4746 (N_4746,N_3889,N_3423);
nand U4747 (N_4747,N_3975,N_4395);
and U4748 (N_4748,N_4492,N_3327);
nor U4749 (N_4749,N_3241,N_3501);
xor U4750 (N_4750,N_4040,N_3000);
nor U4751 (N_4751,N_3861,N_3657);
nor U4752 (N_4752,N_3851,N_3099);
nor U4753 (N_4753,N_3324,N_4482);
or U4754 (N_4754,N_3391,N_3545);
and U4755 (N_4755,N_4172,N_3316);
or U4756 (N_4756,N_3114,N_3892);
nor U4757 (N_4757,N_3486,N_4471);
nor U4758 (N_4758,N_3904,N_4270);
or U4759 (N_4759,N_3367,N_3477);
and U4760 (N_4760,N_4028,N_3061);
nand U4761 (N_4761,N_3573,N_3210);
xnor U4762 (N_4762,N_3565,N_3239);
nand U4763 (N_4763,N_3139,N_3961);
or U4764 (N_4764,N_3803,N_3172);
nand U4765 (N_4765,N_3325,N_3683);
nor U4766 (N_4766,N_3487,N_4170);
nor U4767 (N_4767,N_3613,N_4375);
nand U4768 (N_4768,N_3888,N_4227);
and U4769 (N_4769,N_3809,N_4169);
nand U4770 (N_4770,N_3828,N_4116);
nor U4771 (N_4771,N_3901,N_3880);
nand U4772 (N_4772,N_3186,N_3624);
or U4773 (N_4773,N_3697,N_3694);
nand U4774 (N_4774,N_4089,N_4475);
nor U4775 (N_4775,N_3398,N_3660);
nor U4776 (N_4776,N_4354,N_3833);
nand U4777 (N_4777,N_4363,N_3688);
nand U4778 (N_4778,N_4319,N_4161);
and U4779 (N_4779,N_3016,N_3586);
or U4780 (N_4780,N_4497,N_3112);
or U4781 (N_4781,N_3457,N_3352);
or U4782 (N_4782,N_3118,N_3447);
nand U4783 (N_4783,N_3414,N_3724);
or U4784 (N_4784,N_3718,N_3799);
and U4785 (N_4785,N_3997,N_3621);
nor U4786 (N_4786,N_4467,N_4362);
or U4787 (N_4787,N_3606,N_3084);
or U4788 (N_4788,N_3778,N_3800);
and U4789 (N_4789,N_3609,N_4073);
and U4790 (N_4790,N_4329,N_3154);
and U4791 (N_4791,N_3966,N_3580);
nand U4792 (N_4792,N_3286,N_4097);
nor U4793 (N_4793,N_4111,N_3483);
or U4794 (N_4794,N_3298,N_3775);
or U4795 (N_4795,N_4154,N_3857);
nand U4796 (N_4796,N_4125,N_3160);
and U4797 (N_4797,N_4255,N_3591);
nand U4798 (N_4798,N_4250,N_4424);
nor U4799 (N_4799,N_3881,N_3318);
nand U4800 (N_4800,N_3299,N_3169);
nand U4801 (N_4801,N_3124,N_3260);
nand U4802 (N_4802,N_3277,N_3504);
and U4803 (N_4803,N_3796,N_4021);
nor U4804 (N_4804,N_4218,N_4271);
and U4805 (N_4805,N_3314,N_3496);
nand U4806 (N_4806,N_3475,N_4149);
nor U4807 (N_4807,N_3413,N_4032);
or U4808 (N_4808,N_4099,N_4282);
nand U4809 (N_4809,N_3515,N_3643);
nor U4810 (N_4810,N_3737,N_3106);
or U4811 (N_4811,N_3010,N_3329);
nor U4812 (N_4812,N_3132,N_3028);
xor U4813 (N_4813,N_3368,N_4234);
or U4814 (N_4814,N_4314,N_4117);
or U4815 (N_4815,N_4036,N_4190);
nand U4816 (N_4816,N_4413,N_4091);
and U4817 (N_4817,N_3692,N_3048);
nor U4818 (N_4818,N_3476,N_3157);
and U4819 (N_4819,N_3017,N_3141);
and U4820 (N_4820,N_3593,N_3602);
nor U4821 (N_4821,N_3165,N_3647);
nor U4822 (N_4822,N_3557,N_3229);
nor U4823 (N_4823,N_4431,N_3188);
and U4824 (N_4824,N_3673,N_4339);
nor U4825 (N_4825,N_3205,N_3151);
and U4826 (N_4826,N_3705,N_3910);
and U4827 (N_4827,N_4405,N_3379);
nand U4828 (N_4828,N_3254,N_3234);
or U4829 (N_4829,N_3490,N_4171);
nand U4830 (N_4830,N_3285,N_3395);
nor U4831 (N_4831,N_4026,N_3594);
nor U4832 (N_4832,N_3887,N_4468);
xnor U4833 (N_4833,N_4079,N_4067);
nand U4834 (N_4834,N_3105,N_3404);
nor U4835 (N_4835,N_4202,N_4253);
nor U4836 (N_4836,N_4229,N_3943);
and U4837 (N_4837,N_3267,N_4061);
or U4838 (N_4838,N_3448,N_3443);
and U4839 (N_4839,N_4256,N_4155);
nor U4840 (N_4840,N_3874,N_3972);
and U4841 (N_4841,N_3119,N_4086);
nor U4842 (N_4842,N_3741,N_4092);
and U4843 (N_4843,N_4051,N_3498);
and U4844 (N_4844,N_3479,N_4016);
and U4845 (N_4845,N_3236,N_3339);
nor U4846 (N_4846,N_3033,N_4068);
nand U4847 (N_4847,N_3351,N_3656);
or U4848 (N_4848,N_4022,N_3023);
nand U4849 (N_4849,N_3173,N_4074);
nor U4850 (N_4850,N_3527,N_3265);
and U4851 (N_4851,N_3863,N_3335);
nor U4852 (N_4852,N_4249,N_3100);
nand U4853 (N_4853,N_3551,N_3302);
nand U4854 (N_4854,N_3794,N_3054);
nand U4855 (N_4855,N_4216,N_3171);
nand U4856 (N_4856,N_3194,N_4474);
nand U4857 (N_4857,N_3473,N_3422);
nand U4858 (N_4858,N_4260,N_3412);
nand U4859 (N_4859,N_3604,N_3467);
nor U4860 (N_4860,N_4320,N_3511);
nor U4861 (N_4861,N_3373,N_3378);
nand U4862 (N_4862,N_3130,N_3528);
and U4863 (N_4863,N_3956,N_4287);
nand U4864 (N_4864,N_4371,N_3958);
and U4865 (N_4865,N_3012,N_3460);
nand U4866 (N_4866,N_4122,N_4142);
and U4867 (N_4867,N_3787,N_4044);
or U4868 (N_4868,N_3978,N_4031);
nand U4869 (N_4869,N_3025,N_3754);
nor U4870 (N_4870,N_3250,N_4006);
or U4871 (N_4871,N_3615,N_4429);
or U4872 (N_4872,N_3416,N_4447);
or U4873 (N_4873,N_3292,N_4069);
or U4874 (N_4874,N_3280,N_3184);
and U4875 (N_4875,N_3805,N_4030);
and U4876 (N_4876,N_3860,N_3801);
nand U4877 (N_4877,N_3259,N_3561);
nand U4878 (N_4878,N_3007,N_4373);
nor U4879 (N_4879,N_3185,N_4037);
nor U4880 (N_4880,N_3204,N_4151);
or U4881 (N_4881,N_4072,N_3539);
xnor U4882 (N_4882,N_3410,N_3856);
and U4883 (N_4883,N_3886,N_4140);
xnor U4884 (N_4884,N_4163,N_3841);
and U4885 (N_4885,N_3289,N_4118);
nor U4886 (N_4886,N_4197,N_3713);
and U4887 (N_4887,N_3415,N_3931);
nor U4888 (N_4888,N_4365,N_3853);
nand U4889 (N_4889,N_3253,N_3567);
or U4890 (N_4890,N_4115,N_3348);
and U4891 (N_4891,N_3075,N_3845);
nand U4892 (N_4892,N_3869,N_3349);
or U4893 (N_4893,N_4490,N_4152);
or U4894 (N_4894,N_4109,N_3516);
and U4895 (N_4895,N_3053,N_3700);
nand U4896 (N_4896,N_3896,N_4196);
nand U4897 (N_4897,N_3252,N_3179);
nor U4898 (N_4898,N_4342,N_3153);
nand U4899 (N_4899,N_4203,N_3917);
nand U4900 (N_4900,N_3266,N_3029);
and U4901 (N_4901,N_3662,N_3757);
nor U4902 (N_4902,N_4381,N_4009);
and U4903 (N_4903,N_4327,N_3773);
and U4904 (N_4904,N_3563,N_3998);
or U4905 (N_4905,N_3987,N_4387);
and U4906 (N_4906,N_3354,N_3125);
nand U4907 (N_4907,N_3520,N_3852);
nor U4908 (N_4908,N_3089,N_4082);
nand U4909 (N_4909,N_3047,N_4487);
and U4910 (N_4910,N_3919,N_3482);
and U4911 (N_4911,N_3898,N_3762);
nand U4912 (N_4912,N_3727,N_4370);
or U4913 (N_4913,N_3034,N_4360);
nor U4914 (N_4914,N_3729,N_3320);
nand U4915 (N_4915,N_4053,N_4348);
nand U4916 (N_4916,N_3227,N_3894);
nand U4917 (N_4917,N_3148,N_4247);
and U4918 (N_4918,N_3147,N_4185);
and U4919 (N_4919,N_3925,N_3049);
nand U4920 (N_4920,N_3039,N_4276);
and U4921 (N_4921,N_3837,N_3564);
and U4922 (N_4922,N_3175,N_4445);
or U4923 (N_4923,N_3282,N_3429);
nor U4924 (N_4924,N_4143,N_4180);
nor U4925 (N_4925,N_3018,N_3446);
and U4926 (N_4926,N_3134,N_3583);
nor U4927 (N_4927,N_3077,N_3916);
nor U4928 (N_4928,N_3182,N_3989);
or U4929 (N_4929,N_3288,N_3669);
and U4930 (N_4930,N_3214,N_3180);
and U4931 (N_4931,N_4402,N_3109);
and U4932 (N_4932,N_4349,N_4038);
and U4933 (N_4933,N_3044,N_4326);
and U4934 (N_4934,N_4406,N_3011);
nand U4935 (N_4935,N_3884,N_3968);
or U4936 (N_4936,N_3649,N_3385);
or U4937 (N_4937,N_3178,N_3005);
and U4938 (N_4938,N_3306,N_4062);
or U4939 (N_4939,N_3568,N_3364);
and U4940 (N_4940,N_3350,N_3690);
and U4941 (N_4941,N_3070,N_3170);
or U4942 (N_4942,N_4221,N_3417);
and U4943 (N_4943,N_4491,N_4017);
nor U4944 (N_4944,N_3208,N_3383);
and U4945 (N_4945,N_3452,N_3332);
nand U4946 (N_4946,N_3371,N_3817);
nand U4947 (N_4947,N_3756,N_4452);
nand U4948 (N_4948,N_3459,N_4415);
and U4949 (N_4949,N_3736,N_4378);
or U4950 (N_4950,N_3795,N_4258);
or U4951 (N_4951,N_4408,N_3135);
nor U4952 (N_4952,N_3189,N_4013);
nand U4953 (N_4953,N_3296,N_4098);
or U4954 (N_4954,N_3405,N_3702);
or U4955 (N_4955,N_3347,N_4272);
nand U4956 (N_4956,N_3866,N_3232);
or U4957 (N_4957,N_3879,N_4414);
nor U4958 (N_4958,N_4412,N_3992);
nor U4959 (N_4959,N_3589,N_4418);
and U4960 (N_4960,N_4416,N_4318);
or U4961 (N_4961,N_3605,N_3503);
or U4962 (N_4962,N_4392,N_4002);
nor U4963 (N_4963,N_3726,N_3394);
or U4964 (N_4964,N_3449,N_3995);
or U4965 (N_4965,N_3934,N_3537);
and U4966 (N_4966,N_3425,N_4174);
or U4967 (N_4967,N_4324,N_3900);
and U4968 (N_4968,N_3518,N_3864);
and U4969 (N_4969,N_3552,N_3820);
and U4970 (N_4970,N_4456,N_3665);
and U4971 (N_4971,N_3814,N_3965);
nand U4972 (N_4972,N_4454,N_3095);
nor U4973 (N_4973,N_3977,N_3193);
nand U4974 (N_4974,N_3434,N_3030);
nor U4975 (N_4975,N_4252,N_4223);
nor U4976 (N_4976,N_3382,N_3301);
nand U4977 (N_4977,N_3323,N_4135);
and U4978 (N_4978,N_3293,N_3149);
nand U4979 (N_4979,N_3969,N_3626);
nor U4980 (N_4980,N_3823,N_4090);
nand U4981 (N_4981,N_4438,N_3973);
and U4982 (N_4982,N_4242,N_3936);
and U4983 (N_4983,N_3914,N_4052);
or U4984 (N_4984,N_3066,N_3485);
nand U4985 (N_4985,N_3436,N_4297);
nor U4986 (N_4986,N_3211,N_3723);
nand U4987 (N_4987,N_3380,N_3818);
nor U4988 (N_4988,N_3650,N_3181);
nand U4989 (N_4989,N_4241,N_3263);
nor U4990 (N_4990,N_3055,N_4139);
or U4991 (N_4991,N_3513,N_3970);
nand U4992 (N_4992,N_4018,N_4012);
and U4993 (N_4993,N_4101,N_3120);
or U4994 (N_4994,N_4259,N_4316);
and U4995 (N_4995,N_3098,N_4264);
nand U4996 (N_4996,N_4145,N_4367);
nand U4997 (N_4997,N_3006,N_3456);
nor U4998 (N_4998,N_4273,N_3122);
nand U4999 (N_4999,N_3785,N_3437);
nor U5000 (N_5000,N_3536,N_3428);
or U5001 (N_5001,N_4100,N_3664);
and U5002 (N_5002,N_4141,N_3319);
or U5003 (N_5003,N_4075,N_3947);
or U5004 (N_5004,N_4480,N_3835);
xor U5005 (N_5005,N_4047,N_4243);
nand U5006 (N_5006,N_4268,N_3168);
and U5007 (N_5007,N_3868,N_4465);
or U5008 (N_5008,N_3384,N_4064);
and U5009 (N_5009,N_3808,N_3816);
and U5010 (N_5010,N_4340,N_3623);
or U5011 (N_5011,N_4124,N_3579);
or U5012 (N_5012,N_3740,N_3063);
nand U5013 (N_5013,N_3908,N_3641);
and U5014 (N_5014,N_4336,N_3450);
nor U5015 (N_5015,N_3807,N_3372);
nor U5016 (N_5016,N_4333,N_4178);
and U5017 (N_5017,N_4313,N_4042);
or U5018 (N_5018,N_4167,N_3284);
nor U5019 (N_5019,N_3363,N_4291);
or U5020 (N_5020,N_3990,N_4435);
nor U5021 (N_5021,N_3631,N_3035);
nand U5022 (N_5022,N_3419,N_3648);
nand U5023 (N_5023,N_3581,N_4168);
nand U5024 (N_5024,N_4132,N_4341);
or U5025 (N_5025,N_4476,N_3985);
nor U5026 (N_5026,N_3608,N_3538);
and U5027 (N_5027,N_3056,N_3923);
nand U5028 (N_5028,N_3116,N_3101);
and U5029 (N_5029,N_4437,N_3559);
and U5030 (N_5030,N_3014,N_4457);
nor U5031 (N_5031,N_3451,N_3540);
and U5032 (N_5032,N_3701,N_3439);
nor U5033 (N_5033,N_4449,N_3230);
nand U5034 (N_5034,N_3261,N_3838);
or U5035 (N_5035,N_3827,N_4263);
and U5036 (N_5036,N_3270,N_3195);
or U5037 (N_5037,N_3003,N_3867);
nor U5038 (N_5038,N_3300,N_3810);
nand U5039 (N_5039,N_4104,N_3201);
and U5040 (N_5040,N_3251,N_4114);
nor U5041 (N_5041,N_3587,N_3876);
or U5042 (N_5042,N_3279,N_3924);
and U5043 (N_5043,N_3654,N_3645);
nor U5044 (N_5044,N_3145,N_3071);
or U5045 (N_5045,N_3031,N_3915);
nand U5046 (N_5046,N_4150,N_3525);
and U5047 (N_5047,N_4430,N_3772);
nor U5048 (N_5048,N_3078,N_3844);
or U5049 (N_5049,N_3572,N_4311);
and U5050 (N_5050,N_3517,N_3346);
or U5051 (N_5051,N_3994,N_3240);
nand U5052 (N_5052,N_4198,N_4071);
and U5053 (N_5053,N_4428,N_4120);
nand U5054 (N_5054,N_4379,N_3207);
nor U5055 (N_5055,N_3108,N_3822);
or U5056 (N_5056,N_4183,N_3597);
nand U5057 (N_5057,N_3131,N_4284);
or U5058 (N_5058,N_4330,N_4083);
nand U5059 (N_5059,N_3140,N_3203);
or U5060 (N_5060,N_4303,N_3303);
nand U5061 (N_5061,N_3957,N_4485);
or U5062 (N_5062,N_4309,N_3357);
and U5063 (N_5063,N_3646,N_4299);
or U5064 (N_5064,N_3497,N_3521);
or U5065 (N_5065,N_4193,N_3781);
nand U5066 (N_5066,N_3666,N_3749);
nand U5067 (N_5067,N_3575,N_4033);
and U5068 (N_5068,N_4206,N_3981);
nor U5069 (N_5069,N_3138,N_4300);
nand U5070 (N_5070,N_4204,N_4137);
nor U5071 (N_5071,N_3980,N_4383);
xor U5072 (N_5072,N_3001,N_3402);
nor U5073 (N_5073,N_3918,N_3883);
or U5074 (N_5074,N_3730,N_4443);
or U5075 (N_5075,N_4391,N_4175);
nor U5076 (N_5076,N_3015,N_4123);
nand U5077 (N_5077,N_3231,N_3791);
nand U5078 (N_5078,N_3746,N_4293);
or U5079 (N_5079,N_3804,N_4364);
or U5080 (N_5080,N_3087,N_4050);
nor U5081 (N_5081,N_4224,N_3235);
and U5082 (N_5082,N_3959,N_4403);
and U5083 (N_5083,N_3760,N_4131);
nor U5084 (N_5084,N_4489,N_4160);
nor U5085 (N_5085,N_3526,N_4240);
nand U5086 (N_5086,N_4377,N_3693);
and U5087 (N_5087,N_4214,N_3909);
nand U5088 (N_5088,N_3619,N_3755);
nand U5089 (N_5089,N_3370,N_4434);
nand U5090 (N_5090,N_3944,N_3639);
or U5091 (N_5091,N_3954,N_3745);
nand U5092 (N_5092,N_4302,N_3237);
nor U5093 (N_5093,N_3937,N_3334);
nand U5094 (N_5094,N_4442,N_3136);
nand U5095 (N_5095,N_3686,N_4212);
nor U5096 (N_5096,N_4344,N_3653);
nor U5097 (N_5097,N_3083,N_3769);
nor U5098 (N_5098,N_3246,N_4385);
and U5099 (N_5099,N_3570,N_3255);
nand U5100 (N_5100,N_3344,N_4386);
nor U5101 (N_5101,N_3577,N_3813);
and U5102 (N_5102,N_3502,N_3500);
nor U5103 (N_5103,N_3870,N_4080);
and U5104 (N_5104,N_3126,N_3418);
nand U5105 (N_5105,N_4003,N_4004);
and U5106 (N_5106,N_4233,N_3780);
or U5107 (N_5107,N_4368,N_3825);
nor U5108 (N_5108,N_3399,N_3659);
and U5109 (N_5109,N_3687,N_3215);
or U5110 (N_5110,N_4417,N_3393);
or U5111 (N_5111,N_4119,N_4177);
and U5112 (N_5112,N_3222,N_3069);
and U5113 (N_5113,N_3882,N_3304);
nor U5114 (N_5114,N_3258,N_3362);
nand U5115 (N_5115,N_3691,N_3212);
nand U5116 (N_5116,N_3706,N_3164);
and U5117 (N_5117,N_3635,N_4436);
nand U5118 (N_5118,N_3634,N_3891);
or U5119 (N_5119,N_4066,N_4184);
or U5120 (N_5120,N_3797,N_3675);
nor U5121 (N_5121,N_3198,N_3824);
or U5122 (N_5122,N_4176,N_4010);
nand U5123 (N_5123,N_3753,N_4055);
nand U5124 (N_5124,N_4085,N_4301);
or U5125 (N_5125,N_4257,N_3534);
or U5126 (N_5126,N_3532,N_3628);
nand U5127 (N_5127,N_3779,N_3183);
or U5128 (N_5128,N_4133,N_3996);
nand U5129 (N_5129,N_4410,N_4376);
nor U5130 (N_5130,N_3249,N_3322);
nor U5131 (N_5131,N_3342,N_4146);
nand U5132 (N_5132,N_4484,N_3009);
nor U5133 (N_5133,N_3519,N_3616);
nor U5134 (N_5134,N_3103,N_4110);
and U5135 (N_5135,N_3668,N_3057);
or U5136 (N_5136,N_4262,N_3696);
nor U5137 (N_5137,N_3652,N_3438);
or U5138 (N_5138,N_3505,N_3600);
or U5139 (N_5139,N_3751,N_3685);
nand U5140 (N_5140,N_3846,N_4466);
or U5141 (N_5141,N_4157,N_3365);
nor U5142 (N_5142,N_3223,N_3199);
or U5143 (N_5143,N_4352,N_3256);
nand U5144 (N_5144,N_4433,N_3248);
or U5145 (N_5145,N_3469,N_3948);
nor U5146 (N_5146,N_4251,N_3432);
nor U5147 (N_5147,N_4201,N_4464);
and U5148 (N_5148,N_4008,N_3907);
and U5149 (N_5149,N_3291,N_3584);
nor U5150 (N_5150,N_3403,N_3974);
and U5151 (N_5151,N_4236,N_3819);
and U5152 (N_5152,N_3967,N_4481);
or U5153 (N_5153,N_3941,N_3174);
nor U5154 (N_5154,N_3464,N_3155);
nand U5155 (N_5155,N_4292,N_3401);
or U5156 (N_5156,N_3097,N_4200);
and U5157 (N_5157,N_3699,N_3788);
nand U5158 (N_5158,N_3802,N_4011);
or U5159 (N_5159,N_3530,N_3219);
or U5160 (N_5160,N_4191,N_3495);
nand U5161 (N_5161,N_4401,N_3849);
and U5162 (N_5162,N_3960,N_3491);
nand U5163 (N_5163,N_4194,N_3946);
or U5164 (N_5164,N_3890,N_3297);
or U5165 (N_5165,N_3386,N_3544);
and U5166 (N_5166,N_4188,N_3940);
nand U5167 (N_5167,N_3630,N_4323);
nor U5168 (N_5168,N_3930,N_3002);
nand U5169 (N_5169,N_3782,N_4343);
nor U5170 (N_5170,N_3022,N_3764);
and U5171 (N_5171,N_3287,N_4295);
and U5172 (N_5172,N_3026,N_4076);
or U5173 (N_5173,N_3858,N_3480);
nand U5174 (N_5174,N_3366,N_3725);
nor U5175 (N_5175,N_4450,N_4269);
nand U5176 (N_5176,N_4310,N_3991);
or U5177 (N_5177,N_3166,N_4244);
nand U5178 (N_5178,N_4121,N_3983);
or U5179 (N_5179,N_3834,N_4088);
nand U5180 (N_5180,N_3216,N_4153);
nand U5181 (N_5181,N_4315,N_4488);
nor U5182 (N_5182,N_3196,N_4277);
nor U5183 (N_5183,N_4057,N_4173);
nor U5184 (N_5184,N_3472,N_3272);
or U5185 (N_5185,N_4384,N_4238);
nor U5186 (N_5186,N_3206,N_3576);
or U5187 (N_5187,N_3396,N_4060);
or U5188 (N_5188,N_4024,N_3111);
or U5189 (N_5189,N_3158,N_3709);
nor U5190 (N_5190,N_4328,N_4400);
or U5191 (N_5191,N_3611,N_3290);
nor U5192 (N_5192,N_3387,N_4095);
and U5193 (N_5193,N_3096,N_3104);
nand U5194 (N_5194,N_3759,N_3294);
nand U5195 (N_5195,N_3024,N_4226);
nand U5196 (N_5196,N_4207,N_3358);
nor U5197 (N_5197,N_3088,N_4199);
and U5198 (N_5198,N_3032,N_4278);
nand U5199 (N_5199,N_4005,N_3719);
and U5200 (N_5200,N_3798,N_3612);
nand U5201 (N_5201,N_3862,N_4374);
nor U5202 (N_5202,N_3829,N_4159);
and U5203 (N_5203,N_3462,N_3041);
or U5204 (N_5204,N_4162,N_3328);
nand U5205 (N_5205,N_4225,N_4321);
nor U5206 (N_5206,N_3345,N_3601);
and U5207 (N_5207,N_3632,N_3400);
and U5208 (N_5208,N_3984,N_3871);
nand U5209 (N_5209,N_3271,N_4220);
nor U5210 (N_5210,N_4396,N_3776);
nor U5211 (N_5211,N_3658,N_4014);
nand U5212 (N_5212,N_3408,N_4084);
or U5213 (N_5213,N_3390,N_4380);
nand U5214 (N_5214,N_4355,N_4305);
nand U5215 (N_5215,N_3489,N_3187);
and U5216 (N_5216,N_3137,N_4357);
and U5217 (N_5217,N_3117,N_3238);
or U5218 (N_5218,N_4470,N_3920);
nor U5219 (N_5219,N_3744,N_3245);
and U5220 (N_5220,N_3765,N_4094);
nand U5221 (N_5221,N_3257,N_4399);
or U5222 (N_5222,N_3806,N_4041);
and U5223 (N_5223,N_4322,N_4478);
or U5224 (N_5224,N_3574,N_4337);
or U5225 (N_5225,N_4179,N_3514);
and U5226 (N_5226,N_4498,N_4108);
or U5227 (N_5227,N_3761,N_3079);
nand U5228 (N_5228,N_3389,N_3747);
nand U5229 (N_5229,N_3768,N_3792);
nor U5230 (N_5230,N_3912,N_3295);
nand U5231 (N_5231,N_4192,N_3167);
or U5232 (N_5232,N_4351,N_4147);
nor U5233 (N_5233,N_4232,N_3748);
nor U5234 (N_5234,N_4451,N_3541);
nor U5235 (N_5235,N_4422,N_3102);
and U5236 (N_5236,N_3715,N_3431);
or U5237 (N_5237,N_3426,N_4459);
or U5238 (N_5238,N_4093,N_3050);
nand U5239 (N_5239,N_3899,N_3465);
nand U5240 (N_5240,N_3558,N_4025);
nor U5241 (N_5241,N_4335,N_3774);
or U5242 (N_5242,N_3042,N_4000);
nor U5243 (N_5243,N_3225,N_3698);
or U5244 (N_5244,N_3620,N_3435);
nand U5245 (N_5245,N_3337,N_4404);
or U5246 (N_5246,N_4181,N_3499);
nand U5247 (N_5247,N_3021,N_3949);
nand U5248 (N_5248,N_3355,N_4479);
nand U5249 (N_5249,N_3128,N_3676);
nand U5250 (N_5250,N_4160,N_4046);
or U5251 (N_5251,N_4037,N_3795);
nand U5252 (N_5252,N_3401,N_3086);
or U5253 (N_5253,N_3566,N_4263);
nand U5254 (N_5254,N_3430,N_3708);
nor U5255 (N_5255,N_3678,N_3058);
nor U5256 (N_5256,N_3658,N_3256);
or U5257 (N_5257,N_3716,N_4026);
nand U5258 (N_5258,N_4061,N_3154);
nor U5259 (N_5259,N_4011,N_3801);
nand U5260 (N_5260,N_4405,N_3579);
or U5261 (N_5261,N_3664,N_4177);
nor U5262 (N_5262,N_3178,N_4248);
nor U5263 (N_5263,N_4034,N_3433);
and U5264 (N_5264,N_4064,N_3244);
nor U5265 (N_5265,N_4415,N_3851);
or U5266 (N_5266,N_3741,N_3500);
or U5267 (N_5267,N_4492,N_3381);
nand U5268 (N_5268,N_4381,N_3309);
and U5269 (N_5269,N_3267,N_4253);
or U5270 (N_5270,N_3641,N_3782);
or U5271 (N_5271,N_4180,N_3122);
or U5272 (N_5272,N_4098,N_3664);
nand U5273 (N_5273,N_3930,N_4140);
or U5274 (N_5274,N_4101,N_3508);
or U5275 (N_5275,N_3999,N_3961);
and U5276 (N_5276,N_3413,N_3986);
and U5277 (N_5277,N_4354,N_3525);
nand U5278 (N_5278,N_3874,N_3169);
nor U5279 (N_5279,N_4001,N_3150);
or U5280 (N_5280,N_3159,N_3911);
nand U5281 (N_5281,N_4156,N_3988);
nor U5282 (N_5282,N_3486,N_3345);
nor U5283 (N_5283,N_3771,N_3183);
nand U5284 (N_5284,N_3694,N_4452);
xnor U5285 (N_5285,N_3227,N_4380);
and U5286 (N_5286,N_3282,N_3487);
or U5287 (N_5287,N_3967,N_4298);
or U5288 (N_5288,N_3579,N_3673);
nor U5289 (N_5289,N_4060,N_3308);
nor U5290 (N_5290,N_3227,N_3187);
or U5291 (N_5291,N_3228,N_3686);
nand U5292 (N_5292,N_3414,N_3250);
or U5293 (N_5293,N_4427,N_4291);
or U5294 (N_5294,N_3990,N_3130);
and U5295 (N_5295,N_3055,N_3376);
nor U5296 (N_5296,N_3461,N_4366);
or U5297 (N_5297,N_4347,N_4499);
and U5298 (N_5298,N_3464,N_3633);
nand U5299 (N_5299,N_3971,N_3442);
nor U5300 (N_5300,N_3481,N_4130);
nor U5301 (N_5301,N_3958,N_4322);
or U5302 (N_5302,N_3405,N_4145);
or U5303 (N_5303,N_3184,N_3984);
nand U5304 (N_5304,N_4261,N_3530);
nor U5305 (N_5305,N_3101,N_3643);
xor U5306 (N_5306,N_4244,N_3583);
nor U5307 (N_5307,N_4140,N_3940);
or U5308 (N_5308,N_3660,N_3589);
and U5309 (N_5309,N_4206,N_3517);
or U5310 (N_5310,N_3222,N_4182);
and U5311 (N_5311,N_3445,N_3980);
or U5312 (N_5312,N_4083,N_4248);
or U5313 (N_5313,N_4120,N_3309);
or U5314 (N_5314,N_4156,N_4255);
nor U5315 (N_5315,N_3091,N_4127);
or U5316 (N_5316,N_4105,N_3206);
nor U5317 (N_5317,N_3252,N_4320);
or U5318 (N_5318,N_3643,N_3884);
nor U5319 (N_5319,N_3187,N_4127);
nor U5320 (N_5320,N_3239,N_3095);
and U5321 (N_5321,N_3910,N_3566);
and U5322 (N_5322,N_3911,N_3745);
and U5323 (N_5323,N_4451,N_3845);
nor U5324 (N_5324,N_3509,N_4412);
or U5325 (N_5325,N_4124,N_3850);
nor U5326 (N_5326,N_3779,N_3932);
nor U5327 (N_5327,N_3731,N_3867);
nand U5328 (N_5328,N_3957,N_3624);
nor U5329 (N_5329,N_3105,N_4468);
and U5330 (N_5330,N_4065,N_4471);
nand U5331 (N_5331,N_3110,N_4253);
and U5332 (N_5332,N_4343,N_3468);
nand U5333 (N_5333,N_3601,N_3179);
or U5334 (N_5334,N_3511,N_3752);
and U5335 (N_5335,N_3004,N_3767);
and U5336 (N_5336,N_4295,N_3722);
and U5337 (N_5337,N_4005,N_3159);
nor U5338 (N_5338,N_3286,N_3517);
or U5339 (N_5339,N_4286,N_3897);
or U5340 (N_5340,N_4224,N_4335);
nor U5341 (N_5341,N_4283,N_4297);
nor U5342 (N_5342,N_3354,N_3237);
nor U5343 (N_5343,N_3588,N_4094);
nor U5344 (N_5344,N_3395,N_3476);
nor U5345 (N_5345,N_3041,N_3378);
nand U5346 (N_5346,N_4032,N_3053);
or U5347 (N_5347,N_4497,N_3926);
and U5348 (N_5348,N_4156,N_3604);
and U5349 (N_5349,N_4383,N_3426);
and U5350 (N_5350,N_3566,N_3903);
nand U5351 (N_5351,N_3473,N_3414);
nand U5352 (N_5352,N_3776,N_3219);
nand U5353 (N_5353,N_3640,N_3928);
xor U5354 (N_5354,N_3614,N_3485);
and U5355 (N_5355,N_4349,N_4347);
or U5356 (N_5356,N_3253,N_3595);
nor U5357 (N_5357,N_3274,N_4041);
nand U5358 (N_5358,N_4286,N_3381);
or U5359 (N_5359,N_4282,N_3606);
nor U5360 (N_5360,N_3344,N_4315);
or U5361 (N_5361,N_3337,N_3539);
nand U5362 (N_5362,N_4498,N_3058);
xor U5363 (N_5363,N_3009,N_3187);
and U5364 (N_5364,N_4394,N_3070);
nand U5365 (N_5365,N_4420,N_3572);
and U5366 (N_5366,N_3065,N_3867);
or U5367 (N_5367,N_3389,N_4009);
xor U5368 (N_5368,N_3667,N_3425);
nand U5369 (N_5369,N_4420,N_3745);
and U5370 (N_5370,N_3981,N_3099);
and U5371 (N_5371,N_4177,N_4439);
and U5372 (N_5372,N_3933,N_3300);
nand U5373 (N_5373,N_4002,N_4151);
nand U5374 (N_5374,N_3485,N_3544);
and U5375 (N_5375,N_3521,N_3184);
xnor U5376 (N_5376,N_3223,N_4127);
or U5377 (N_5377,N_4471,N_3571);
nand U5378 (N_5378,N_3366,N_3287);
nor U5379 (N_5379,N_4478,N_3695);
and U5380 (N_5380,N_3845,N_3286);
nor U5381 (N_5381,N_3901,N_3573);
and U5382 (N_5382,N_3769,N_4110);
nor U5383 (N_5383,N_3637,N_3085);
or U5384 (N_5384,N_3458,N_4193);
and U5385 (N_5385,N_3124,N_3428);
and U5386 (N_5386,N_3888,N_3428);
nand U5387 (N_5387,N_3627,N_3803);
or U5388 (N_5388,N_4396,N_3159);
nor U5389 (N_5389,N_3429,N_3279);
nand U5390 (N_5390,N_4148,N_3466);
nand U5391 (N_5391,N_3278,N_4110);
or U5392 (N_5392,N_4006,N_4302);
or U5393 (N_5393,N_3239,N_3895);
nand U5394 (N_5394,N_3886,N_3751);
nor U5395 (N_5395,N_3810,N_3241);
and U5396 (N_5396,N_3552,N_4433);
and U5397 (N_5397,N_3775,N_3214);
and U5398 (N_5398,N_3178,N_3828);
and U5399 (N_5399,N_4125,N_4304);
nand U5400 (N_5400,N_3540,N_3614);
nand U5401 (N_5401,N_4263,N_3524);
and U5402 (N_5402,N_3812,N_3787);
and U5403 (N_5403,N_3123,N_4003);
nand U5404 (N_5404,N_4073,N_3159);
or U5405 (N_5405,N_4336,N_3538);
nand U5406 (N_5406,N_4175,N_3180);
and U5407 (N_5407,N_4152,N_3031);
and U5408 (N_5408,N_3319,N_3926);
nor U5409 (N_5409,N_4048,N_4441);
and U5410 (N_5410,N_4230,N_3258);
or U5411 (N_5411,N_4338,N_4304);
nor U5412 (N_5412,N_3535,N_3847);
or U5413 (N_5413,N_3577,N_3529);
nand U5414 (N_5414,N_3673,N_3281);
nand U5415 (N_5415,N_3918,N_3613);
or U5416 (N_5416,N_3573,N_4029);
and U5417 (N_5417,N_3969,N_3445);
nand U5418 (N_5418,N_3899,N_3782);
or U5419 (N_5419,N_4347,N_3689);
nand U5420 (N_5420,N_3243,N_3149);
nor U5421 (N_5421,N_3710,N_3065);
nor U5422 (N_5422,N_3192,N_3419);
nor U5423 (N_5423,N_3480,N_4123);
and U5424 (N_5424,N_4285,N_3535);
nor U5425 (N_5425,N_3662,N_3777);
and U5426 (N_5426,N_4301,N_3096);
and U5427 (N_5427,N_3423,N_4411);
nand U5428 (N_5428,N_3453,N_3174);
and U5429 (N_5429,N_4389,N_4111);
or U5430 (N_5430,N_3183,N_3552);
nand U5431 (N_5431,N_4310,N_3257);
and U5432 (N_5432,N_3487,N_3490);
nor U5433 (N_5433,N_4044,N_3683);
nand U5434 (N_5434,N_4136,N_4444);
and U5435 (N_5435,N_4189,N_3716);
or U5436 (N_5436,N_3920,N_4172);
nand U5437 (N_5437,N_3882,N_4162);
and U5438 (N_5438,N_4357,N_4068);
and U5439 (N_5439,N_3025,N_4158);
or U5440 (N_5440,N_3155,N_3419);
and U5441 (N_5441,N_3547,N_3236);
or U5442 (N_5442,N_3283,N_3703);
and U5443 (N_5443,N_3075,N_3342);
and U5444 (N_5444,N_3968,N_3861);
and U5445 (N_5445,N_3061,N_4220);
nor U5446 (N_5446,N_4126,N_3586);
or U5447 (N_5447,N_3919,N_3114);
nand U5448 (N_5448,N_3391,N_3017);
nand U5449 (N_5449,N_4430,N_4370);
nor U5450 (N_5450,N_4179,N_3450);
nor U5451 (N_5451,N_3931,N_3734);
nand U5452 (N_5452,N_4357,N_4418);
or U5453 (N_5453,N_4286,N_3120);
and U5454 (N_5454,N_4220,N_3173);
and U5455 (N_5455,N_3984,N_3495);
nand U5456 (N_5456,N_3038,N_3899);
nor U5457 (N_5457,N_3916,N_3534);
and U5458 (N_5458,N_4242,N_4326);
nor U5459 (N_5459,N_3127,N_3909);
nand U5460 (N_5460,N_3263,N_3514);
nor U5461 (N_5461,N_3156,N_3084);
nand U5462 (N_5462,N_3023,N_3801);
or U5463 (N_5463,N_3632,N_4353);
nor U5464 (N_5464,N_3622,N_3758);
or U5465 (N_5465,N_4322,N_4114);
nand U5466 (N_5466,N_3317,N_3290);
or U5467 (N_5467,N_3878,N_3473);
or U5468 (N_5468,N_3831,N_4392);
and U5469 (N_5469,N_3358,N_3150);
and U5470 (N_5470,N_3877,N_3631);
and U5471 (N_5471,N_4354,N_3402);
and U5472 (N_5472,N_3988,N_3726);
or U5473 (N_5473,N_3215,N_3010);
nand U5474 (N_5474,N_3958,N_4370);
nand U5475 (N_5475,N_3714,N_4131);
nand U5476 (N_5476,N_4083,N_4288);
and U5477 (N_5477,N_3989,N_4309);
nor U5478 (N_5478,N_4061,N_3896);
nand U5479 (N_5479,N_3128,N_4456);
nor U5480 (N_5480,N_3709,N_4369);
nor U5481 (N_5481,N_4001,N_4225);
nand U5482 (N_5482,N_3686,N_4436);
or U5483 (N_5483,N_3889,N_3154);
and U5484 (N_5484,N_3008,N_3854);
nand U5485 (N_5485,N_3648,N_4175);
nor U5486 (N_5486,N_3946,N_3755);
or U5487 (N_5487,N_4401,N_3123);
nor U5488 (N_5488,N_3276,N_4311);
nand U5489 (N_5489,N_4441,N_4149);
and U5490 (N_5490,N_3953,N_3683);
and U5491 (N_5491,N_3118,N_3146);
and U5492 (N_5492,N_4164,N_3246);
xor U5493 (N_5493,N_3538,N_3751);
nand U5494 (N_5494,N_3623,N_3860);
and U5495 (N_5495,N_4127,N_3873);
nor U5496 (N_5496,N_3011,N_3131);
and U5497 (N_5497,N_3405,N_4485);
nor U5498 (N_5498,N_3421,N_3268);
and U5499 (N_5499,N_3284,N_4312);
and U5500 (N_5500,N_3543,N_3068);
and U5501 (N_5501,N_3233,N_3163);
nor U5502 (N_5502,N_3138,N_4037);
nor U5503 (N_5503,N_3621,N_4124);
nand U5504 (N_5504,N_4005,N_4432);
and U5505 (N_5505,N_3708,N_3628);
nor U5506 (N_5506,N_3342,N_4133);
nor U5507 (N_5507,N_3791,N_3957);
and U5508 (N_5508,N_3866,N_3582);
and U5509 (N_5509,N_4355,N_3008);
or U5510 (N_5510,N_3104,N_4195);
nand U5511 (N_5511,N_3709,N_3771);
and U5512 (N_5512,N_4154,N_3489);
and U5513 (N_5513,N_3883,N_4293);
and U5514 (N_5514,N_4391,N_3181);
and U5515 (N_5515,N_4126,N_3904);
nand U5516 (N_5516,N_4097,N_3936);
nor U5517 (N_5517,N_3642,N_3333);
nand U5518 (N_5518,N_4140,N_3224);
nor U5519 (N_5519,N_4178,N_3841);
nand U5520 (N_5520,N_3209,N_3301);
or U5521 (N_5521,N_4120,N_4272);
nand U5522 (N_5522,N_3589,N_3432);
and U5523 (N_5523,N_3006,N_3514);
nand U5524 (N_5524,N_4065,N_4323);
and U5525 (N_5525,N_3865,N_3914);
nor U5526 (N_5526,N_4139,N_3568);
nor U5527 (N_5527,N_4191,N_3007);
or U5528 (N_5528,N_3342,N_4216);
or U5529 (N_5529,N_4069,N_4041);
nand U5530 (N_5530,N_3885,N_4215);
or U5531 (N_5531,N_3113,N_3887);
and U5532 (N_5532,N_3961,N_3565);
or U5533 (N_5533,N_3461,N_3223);
nor U5534 (N_5534,N_4365,N_3460);
and U5535 (N_5535,N_4229,N_3745);
nor U5536 (N_5536,N_3412,N_4137);
or U5537 (N_5537,N_3086,N_3489);
nand U5538 (N_5538,N_3964,N_3065);
nand U5539 (N_5539,N_3964,N_3166);
nor U5540 (N_5540,N_3503,N_3212);
and U5541 (N_5541,N_3835,N_3371);
nand U5542 (N_5542,N_4208,N_3732);
and U5543 (N_5543,N_3877,N_4282);
nand U5544 (N_5544,N_3925,N_4414);
nor U5545 (N_5545,N_3284,N_3313);
nor U5546 (N_5546,N_4320,N_3956);
and U5547 (N_5547,N_3826,N_3528);
and U5548 (N_5548,N_3385,N_4025);
nand U5549 (N_5549,N_3514,N_3949);
or U5550 (N_5550,N_3371,N_3441);
nor U5551 (N_5551,N_3697,N_3628);
nor U5552 (N_5552,N_4497,N_3995);
nor U5553 (N_5553,N_3303,N_3968);
nor U5554 (N_5554,N_4359,N_3465);
nand U5555 (N_5555,N_3003,N_3363);
or U5556 (N_5556,N_3040,N_3102);
or U5557 (N_5557,N_3194,N_4169);
or U5558 (N_5558,N_4253,N_3636);
nor U5559 (N_5559,N_4177,N_3872);
and U5560 (N_5560,N_4321,N_4095);
and U5561 (N_5561,N_4204,N_3498);
nor U5562 (N_5562,N_4349,N_3583);
xor U5563 (N_5563,N_3243,N_3861);
nand U5564 (N_5564,N_3476,N_3618);
or U5565 (N_5565,N_4152,N_3205);
or U5566 (N_5566,N_4294,N_4310);
nor U5567 (N_5567,N_4363,N_3220);
nand U5568 (N_5568,N_3722,N_3873);
nor U5569 (N_5569,N_3094,N_3226);
nor U5570 (N_5570,N_3642,N_3370);
and U5571 (N_5571,N_3184,N_4253);
nor U5572 (N_5572,N_4464,N_4080);
and U5573 (N_5573,N_3018,N_3136);
nand U5574 (N_5574,N_3533,N_4480);
and U5575 (N_5575,N_3380,N_3830);
nand U5576 (N_5576,N_4191,N_3705);
nor U5577 (N_5577,N_3235,N_4267);
and U5578 (N_5578,N_4334,N_3100);
and U5579 (N_5579,N_3640,N_3678);
nor U5580 (N_5580,N_3939,N_3620);
nor U5581 (N_5581,N_3948,N_4142);
or U5582 (N_5582,N_3367,N_3889);
nor U5583 (N_5583,N_4292,N_4185);
or U5584 (N_5584,N_3851,N_4463);
or U5585 (N_5585,N_4446,N_3289);
or U5586 (N_5586,N_4398,N_3429);
nor U5587 (N_5587,N_3544,N_4100);
and U5588 (N_5588,N_3201,N_3373);
nor U5589 (N_5589,N_3003,N_4362);
nand U5590 (N_5590,N_3587,N_4000);
nor U5591 (N_5591,N_3097,N_4043);
or U5592 (N_5592,N_3852,N_4224);
or U5593 (N_5593,N_3636,N_3817);
or U5594 (N_5594,N_4198,N_4258);
and U5595 (N_5595,N_3670,N_3253);
or U5596 (N_5596,N_3141,N_4172);
nand U5597 (N_5597,N_3783,N_3629);
or U5598 (N_5598,N_3162,N_3664);
or U5599 (N_5599,N_3259,N_3055);
nor U5600 (N_5600,N_3182,N_4450);
and U5601 (N_5601,N_3084,N_3146);
and U5602 (N_5602,N_3856,N_4399);
nand U5603 (N_5603,N_3987,N_3058);
or U5604 (N_5604,N_4498,N_3130);
and U5605 (N_5605,N_4218,N_4095);
nand U5606 (N_5606,N_3697,N_3970);
nor U5607 (N_5607,N_4471,N_4474);
nor U5608 (N_5608,N_3992,N_3864);
nor U5609 (N_5609,N_4052,N_3029);
and U5610 (N_5610,N_3709,N_4414);
nor U5611 (N_5611,N_3402,N_3860);
or U5612 (N_5612,N_3328,N_4462);
nor U5613 (N_5613,N_4477,N_3554);
nand U5614 (N_5614,N_3105,N_3483);
and U5615 (N_5615,N_3829,N_4389);
nand U5616 (N_5616,N_3122,N_3794);
nand U5617 (N_5617,N_3023,N_3049);
xnor U5618 (N_5618,N_4032,N_4209);
xor U5619 (N_5619,N_3341,N_3371);
nand U5620 (N_5620,N_3668,N_3210);
nor U5621 (N_5621,N_4445,N_3475);
nor U5622 (N_5622,N_4085,N_3279);
nor U5623 (N_5623,N_3312,N_3328);
or U5624 (N_5624,N_4098,N_3578);
nand U5625 (N_5625,N_3329,N_3289);
or U5626 (N_5626,N_3205,N_4387);
or U5627 (N_5627,N_3281,N_4348);
or U5628 (N_5628,N_3407,N_4332);
and U5629 (N_5629,N_3909,N_3341);
nand U5630 (N_5630,N_4014,N_4103);
and U5631 (N_5631,N_4242,N_4419);
or U5632 (N_5632,N_4045,N_4120);
nand U5633 (N_5633,N_4057,N_3160);
nand U5634 (N_5634,N_3838,N_3299);
nor U5635 (N_5635,N_3793,N_3677);
and U5636 (N_5636,N_3224,N_3822);
or U5637 (N_5637,N_3248,N_4153);
nor U5638 (N_5638,N_3177,N_3859);
and U5639 (N_5639,N_4341,N_4328);
or U5640 (N_5640,N_3955,N_3991);
and U5641 (N_5641,N_4252,N_3258);
nand U5642 (N_5642,N_3748,N_3048);
nor U5643 (N_5643,N_3736,N_3518);
nand U5644 (N_5644,N_3905,N_3688);
nor U5645 (N_5645,N_4399,N_4393);
nand U5646 (N_5646,N_4463,N_3256);
nor U5647 (N_5647,N_3852,N_3382);
nand U5648 (N_5648,N_4106,N_3979);
nand U5649 (N_5649,N_3535,N_3113);
nand U5650 (N_5650,N_3290,N_4055);
nor U5651 (N_5651,N_3058,N_4200);
nor U5652 (N_5652,N_4081,N_3931);
or U5653 (N_5653,N_4328,N_4457);
nand U5654 (N_5654,N_4486,N_3088);
nand U5655 (N_5655,N_3857,N_4330);
nor U5656 (N_5656,N_4386,N_4047);
and U5657 (N_5657,N_3738,N_4267);
or U5658 (N_5658,N_4372,N_3639);
nand U5659 (N_5659,N_4442,N_3157);
or U5660 (N_5660,N_3361,N_3263);
or U5661 (N_5661,N_4317,N_3780);
and U5662 (N_5662,N_4327,N_3270);
and U5663 (N_5663,N_3711,N_3643);
nor U5664 (N_5664,N_3593,N_4031);
nand U5665 (N_5665,N_4447,N_3370);
and U5666 (N_5666,N_4351,N_3142);
nor U5667 (N_5667,N_3380,N_3343);
nand U5668 (N_5668,N_3085,N_4233);
or U5669 (N_5669,N_4430,N_4255);
or U5670 (N_5670,N_3688,N_3560);
nand U5671 (N_5671,N_4154,N_3950);
or U5672 (N_5672,N_4244,N_3870);
and U5673 (N_5673,N_3664,N_3446);
nor U5674 (N_5674,N_4054,N_4497);
or U5675 (N_5675,N_3728,N_4484);
nor U5676 (N_5676,N_3908,N_4246);
nor U5677 (N_5677,N_3807,N_4412);
and U5678 (N_5678,N_3500,N_3247);
and U5679 (N_5679,N_4476,N_4175);
nand U5680 (N_5680,N_4494,N_4296);
nor U5681 (N_5681,N_4043,N_3709);
nand U5682 (N_5682,N_4293,N_3323);
nand U5683 (N_5683,N_3377,N_4212);
nand U5684 (N_5684,N_3410,N_3853);
or U5685 (N_5685,N_3915,N_3402);
nand U5686 (N_5686,N_3679,N_4365);
and U5687 (N_5687,N_4004,N_3859);
or U5688 (N_5688,N_4381,N_4157);
and U5689 (N_5689,N_3635,N_3712);
xor U5690 (N_5690,N_4185,N_4029);
nor U5691 (N_5691,N_4039,N_4050);
xor U5692 (N_5692,N_3281,N_4154);
nor U5693 (N_5693,N_3592,N_3675);
and U5694 (N_5694,N_4232,N_3541);
or U5695 (N_5695,N_4380,N_4368);
and U5696 (N_5696,N_4474,N_3516);
nor U5697 (N_5697,N_3656,N_3616);
nor U5698 (N_5698,N_3893,N_3339);
or U5699 (N_5699,N_3550,N_3460);
xnor U5700 (N_5700,N_4491,N_3715);
and U5701 (N_5701,N_4065,N_4330);
and U5702 (N_5702,N_3397,N_4302);
or U5703 (N_5703,N_4315,N_3649);
xnor U5704 (N_5704,N_4196,N_4005);
nor U5705 (N_5705,N_3286,N_3062);
nor U5706 (N_5706,N_3784,N_3960);
and U5707 (N_5707,N_3576,N_4373);
and U5708 (N_5708,N_3002,N_3430);
nand U5709 (N_5709,N_4174,N_3815);
or U5710 (N_5710,N_3767,N_3164);
nor U5711 (N_5711,N_4333,N_3467);
and U5712 (N_5712,N_4123,N_3935);
or U5713 (N_5713,N_3715,N_3528);
or U5714 (N_5714,N_3945,N_3923);
nor U5715 (N_5715,N_3829,N_3481);
nand U5716 (N_5716,N_3896,N_3812);
nand U5717 (N_5717,N_3536,N_3457);
or U5718 (N_5718,N_4349,N_4240);
and U5719 (N_5719,N_3743,N_4206);
nor U5720 (N_5720,N_3837,N_3860);
or U5721 (N_5721,N_4469,N_3234);
nor U5722 (N_5722,N_3286,N_3713);
nor U5723 (N_5723,N_3348,N_3451);
and U5724 (N_5724,N_3872,N_3578);
nor U5725 (N_5725,N_4017,N_3954);
nand U5726 (N_5726,N_3477,N_3173);
nand U5727 (N_5727,N_3904,N_4410);
and U5728 (N_5728,N_3623,N_4178);
nor U5729 (N_5729,N_3334,N_4125);
nor U5730 (N_5730,N_3702,N_3517);
nand U5731 (N_5731,N_3291,N_3939);
and U5732 (N_5732,N_3398,N_4124);
nor U5733 (N_5733,N_3425,N_4362);
nor U5734 (N_5734,N_3765,N_3883);
and U5735 (N_5735,N_3526,N_4301);
or U5736 (N_5736,N_3370,N_3969);
and U5737 (N_5737,N_3369,N_3328);
nor U5738 (N_5738,N_4387,N_3235);
nor U5739 (N_5739,N_3486,N_4298);
or U5740 (N_5740,N_3888,N_3279);
nand U5741 (N_5741,N_3377,N_4385);
nor U5742 (N_5742,N_3495,N_3486);
nand U5743 (N_5743,N_3275,N_3200);
or U5744 (N_5744,N_3387,N_4164);
nor U5745 (N_5745,N_4103,N_3075);
nand U5746 (N_5746,N_3311,N_4235);
and U5747 (N_5747,N_3530,N_3496);
or U5748 (N_5748,N_4088,N_4294);
nor U5749 (N_5749,N_4333,N_3313);
or U5750 (N_5750,N_3345,N_3403);
nand U5751 (N_5751,N_3917,N_3419);
and U5752 (N_5752,N_3461,N_4046);
and U5753 (N_5753,N_4497,N_3546);
xor U5754 (N_5754,N_3394,N_3829);
nand U5755 (N_5755,N_4198,N_3631);
or U5756 (N_5756,N_4278,N_3051);
nor U5757 (N_5757,N_3919,N_3231);
nand U5758 (N_5758,N_3507,N_4029);
nor U5759 (N_5759,N_4444,N_3522);
or U5760 (N_5760,N_3776,N_4337);
and U5761 (N_5761,N_3417,N_4443);
nor U5762 (N_5762,N_3458,N_4389);
and U5763 (N_5763,N_4027,N_3800);
nand U5764 (N_5764,N_3109,N_3103);
and U5765 (N_5765,N_3420,N_3506);
and U5766 (N_5766,N_3615,N_3935);
and U5767 (N_5767,N_3624,N_4467);
and U5768 (N_5768,N_4147,N_3047);
and U5769 (N_5769,N_3443,N_4132);
nor U5770 (N_5770,N_3434,N_4064);
or U5771 (N_5771,N_4270,N_4375);
and U5772 (N_5772,N_4259,N_4211);
and U5773 (N_5773,N_4395,N_3954);
or U5774 (N_5774,N_4134,N_3700);
nor U5775 (N_5775,N_3188,N_3720);
nand U5776 (N_5776,N_3892,N_3665);
nor U5777 (N_5777,N_4405,N_4348);
nor U5778 (N_5778,N_3408,N_3231);
and U5779 (N_5779,N_3061,N_3752);
nor U5780 (N_5780,N_4097,N_3853);
and U5781 (N_5781,N_3306,N_4382);
nand U5782 (N_5782,N_3058,N_4490);
and U5783 (N_5783,N_3492,N_3955);
and U5784 (N_5784,N_3695,N_3397);
nor U5785 (N_5785,N_3910,N_4409);
nand U5786 (N_5786,N_4425,N_4390);
and U5787 (N_5787,N_3665,N_3119);
nand U5788 (N_5788,N_3520,N_3427);
or U5789 (N_5789,N_3258,N_4094);
nor U5790 (N_5790,N_4142,N_3952);
xnor U5791 (N_5791,N_3783,N_3612);
nand U5792 (N_5792,N_3739,N_3022);
nand U5793 (N_5793,N_3772,N_4293);
or U5794 (N_5794,N_3286,N_3019);
nor U5795 (N_5795,N_4112,N_3211);
and U5796 (N_5796,N_3257,N_4058);
and U5797 (N_5797,N_4493,N_3881);
or U5798 (N_5798,N_3646,N_4482);
xnor U5799 (N_5799,N_3392,N_4014);
nor U5800 (N_5800,N_3286,N_3189);
nor U5801 (N_5801,N_3626,N_4082);
and U5802 (N_5802,N_3741,N_3311);
nand U5803 (N_5803,N_3756,N_3201);
nor U5804 (N_5804,N_3318,N_3578);
nor U5805 (N_5805,N_4035,N_3042);
nand U5806 (N_5806,N_3096,N_3456);
or U5807 (N_5807,N_3176,N_3698);
nand U5808 (N_5808,N_3338,N_3496);
nor U5809 (N_5809,N_4464,N_4409);
and U5810 (N_5810,N_4144,N_3750);
nor U5811 (N_5811,N_4343,N_3296);
or U5812 (N_5812,N_3642,N_3413);
and U5813 (N_5813,N_3435,N_3105);
nand U5814 (N_5814,N_4318,N_3270);
and U5815 (N_5815,N_3694,N_4151);
and U5816 (N_5816,N_3489,N_3102);
nor U5817 (N_5817,N_4287,N_4080);
nor U5818 (N_5818,N_3155,N_3752);
and U5819 (N_5819,N_3177,N_4279);
nand U5820 (N_5820,N_3639,N_4323);
nor U5821 (N_5821,N_3673,N_4207);
nand U5822 (N_5822,N_4361,N_3776);
or U5823 (N_5823,N_3375,N_3950);
and U5824 (N_5824,N_4495,N_3663);
nor U5825 (N_5825,N_3401,N_3766);
nand U5826 (N_5826,N_4190,N_3883);
xor U5827 (N_5827,N_3454,N_3033);
xor U5828 (N_5828,N_3034,N_4123);
nor U5829 (N_5829,N_3918,N_3074);
nor U5830 (N_5830,N_4148,N_4390);
or U5831 (N_5831,N_3437,N_4272);
nand U5832 (N_5832,N_4207,N_4376);
or U5833 (N_5833,N_3943,N_4189);
and U5834 (N_5834,N_3816,N_3488);
and U5835 (N_5835,N_3639,N_3638);
and U5836 (N_5836,N_3858,N_3008);
nand U5837 (N_5837,N_4017,N_4246);
nand U5838 (N_5838,N_3854,N_4253);
nor U5839 (N_5839,N_4431,N_4484);
nor U5840 (N_5840,N_4399,N_3098);
nand U5841 (N_5841,N_3204,N_4298);
xor U5842 (N_5842,N_3173,N_3628);
or U5843 (N_5843,N_3307,N_3546);
nand U5844 (N_5844,N_3792,N_3760);
or U5845 (N_5845,N_3512,N_4233);
or U5846 (N_5846,N_3784,N_4435);
nand U5847 (N_5847,N_4495,N_3438);
nand U5848 (N_5848,N_3516,N_4401);
and U5849 (N_5849,N_3021,N_3922);
and U5850 (N_5850,N_4280,N_4087);
nand U5851 (N_5851,N_3823,N_3255);
nand U5852 (N_5852,N_4418,N_4131);
nand U5853 (N_5853,N_3312,N_3561);
xor U5854 (N_5854,N_3969,N_3950);
nand U5855 (N_5855,N_3341,N_3781);
nand U5856 (N_5856,N_3154,N_3689);
nor U5857 (N_5857,N_3832,N_3132);
nand U5858 (N_5858,N_4163,N_3360);
nand U5859 (N_5859,N_4369,N_3703);
nand U5860 (N_5860,N_4271,N_4285);
or U5861 (N_5861,N_3340,N_4047);
and U5862 (N_5862,N_4469,N_3008);
nand U5863 (N_5863,N_3563,N_3018);
nand U5864 (N_5864,N_3283,N_4310);
nand U5865 (N_5865,N_3927,N_4472);
or U5866 (N_5866,N_3781,N_3090);
nor U5867 (N_5867,N_4279,N_4453);
nand U5868 (N_5868,N_3527,N_3955);
nor U5869 (N_5869,N_3212,N_3781);
nor U5870 (N_5870,N_3573,N_4225);
nor U5871 (N_5871,N_3763,N_4281);
or U5872 (N_5872,N_3204,N_3369);
nand U5873 (N_5873,N_4344,N_3248);
nor U5874 (N_5874,N_4352,N_4091);
nand U5875 (N_5875,N_4363,N_4388);
and U5876 (N_5876,N_3543,N_3348);
nor U5877 (N_5877,N_4293,N_3274);
nand U5878 (N_5878,N_4219,N_3902);
and U5879 (N_5879,N_4048,N_4401);
and U5880 (N_5880,N_3913,N_3656);
or U5881 (N_5881,N_4101,N_4464);
nor U5882 (N_5882,N_4274,N_3197);
nor U5883 (N_5883,N_3288,N_3033);
nor U5884 (N_5884,N_3526,N_3299);
or U5885 (N_5885,N_3848,N_4364);
and U5886 (N_5886,N_3350,N_4434);
nor U5887 (N_5887,N_4354,N_4160);
or U5888 (N_5888,N_3674,N_3093);
nand U5889 (N_5889,N_3316,N_3115);
nand U5890 (N_5890,N_4041,N_4282);
and U5891 (N_5891,N_4365,N_4162);
and U5892 (N_5892,N_4355,N_4164);
nand U5893 (N_5893,N_3943,N_3101);
nand U5894 (N_5894,N_3923,N_4165);
nand U5895 (N_5895,N_3058,N_3119);
nand U5896 (N_5896,N_4325,N_3844);
or U5897 (N_5897,N_4049,N_3458);
nor U5898 (N_5898,N_3567,N_4272);
or U5899 (N_5899,N_4478,N_3321);
or U5900 (N_5900,N_4290,N_4371);
nor U5901 (N_5901,N_3062,N_3713);
nor U5902 (N_5902,N_3456,N_3075);
nand U5903 (N_5903,N_4350,N_3738);
and U5904 (N_5904,N_3329,N_4445);
or U5905 (N_5905,N_3259,N_3968);
xor U5906 (N_5906,N_3511,N_3408);
nor U5907 (N_5907,N_3852,N_3980);
nor U5908 (N_5908,N_3119,N_3772);
and U5909 (N_5909,N_4401,N_3676);
and U5910 (N_5910,N_3772,N_3258);
and U5911 (N_5911,N_3262,N_3465);
nand U5912 (N_5912,N_3641,N_4015);
nor U5913 (N_5913,N_3625,N_3514);
nor U5914 (N_5914,N_3673,N_3667);
or U5915 (N_5915,N_3464,N_4322);
nand U5916 (N_5916,N_4405,N_3024);
nor U5917 (N_5917,N_3399,N_3232);
xor U5918 (N_5918,N_3814,N_4175);
and U5919 (N_5919,N_3729,N_3525);
or U5920 (N_5920,N_3832,N_3618);
and U5921 (N_5921,N_3940,N_3080);
and U5922 (N_5922,N_3334,N_3164);
and U5923 (N_5923,N_3105,N_4439);
nor U5924 (N_5924,N_3722,N_4094);
nand U5925 (N_5925,N_4305,N_3784);
nor U5926 (N_5926,N_3453,N_3271);
xnor U5927 (N_5927,N_4290,N_3190);
nand U5928 (N_5928,N_3806,N_4282);
and U5929 (N_5929,N_3322,N_4386);
nor U5930 (N_5930,N_4451,N_3003);
and U5931 (N_5931,N_4217,N_4362);
nand U5932 (N_5932,N_3396,N_3104);
or U5933 (N_5933,N_4164,N_3014);
nand U5934 (N_5934,N_3053,N_3519);
nor U5935 (N_5935,N_3971,N_4492);
and U5936 (N_5936,N_3753,N_3721);
or U5937 (N_5937,N_3702,N_3271);
nor U5938 (N_5938,N_3188,N_3288);
or U5939 (N_5939,N_4144,N_3433);
xor U5940 (N_5940,N_3377,N_4194);
nand U5941 (N_5941,N_3631,N_3846);
or U5942 (N_5942,N_4434,N_3515);
and U5943 (N_5943,N_3450,N_3931);
or U5944 (N_5944,N_4173,N_3977);
nand U5945 (N_5945,N_3376,N_3632);
nand U5946 (N_5946,N_4322,N_3105);
nand U5947 (N_5947,N_3853,N_3763);
nand U5948 (N_5948,N_3332,N_4165);
or U5949 (N_5949,N_3576,N_4004);
and U5950 (N_5950,N_3746,N_4450);
nor U5951 (N_5951,N_3535,N_4154);
or U5952 (N_5952,N_3074,N_3916);
and U5953 (N_5953,N_4369,N_3817);
nand U5954 (N_5954,N_4264,N_3818);
or U5955 (N_5955,N_3476,N_3299);
xor U5956 (N_5956,N_3175,N_3769);
nor U5957 (N_5957,N_3747,N_4495);
nand U5958 (N_5958,N_4319,N_3502);
or U5959 (N_5959,N_3616,N_3082);
nand U5960 (N_5960,N_3793,N_4039);
nand U5961 (N_5961,N_3955,N_3839);
nor U5962 (N_5962,N_4382,N_3429);
and U5963 (N_5963,N_3370,N_3470);
nand U5964 (N_5964,N_3480,N_3694);
nand U5965 (N_5965,N_3925,N_4209);
and U5966 (N_5966,N_3257,N_4267);
nor U5967 (N_5967,N_3776,N_4090);
and U5968 (N_5968,N_3654,N_3025);
nand U5969 (N_5969,N_3586,N_4314);
or U5970 (N_5970,N_3775,N_3895);
or U5971 (N_5971,N_3635,N_3997);
and U5972 (N_5972,N_4328,N_3113);
and U5973 (N_5973,N_3801,N_3068);
nand U5974 (N_5974,N_3360,N_3090);
nor U5975 (N_5975,N_3122,N_4211);
nand U5976 (N_5976,N_4031,N_3638);
nor U5977 (N_5977,N_4477,N_3041);
nor U5978 (N_5978,N_3439,N_4191);
or U5979 (N_5979,N_3701,N_3730);
nand U5980 (N_5980,N_4119,N_3026);
nor U5981 (N_5981,N_4078,N_3915);
or U5982 (N_5982,N_3911,N_3133);
nand U5983 (N_5983,N_4309,N_3729);
and U5984 (N_5984,N_3395,N_4046);
nor U5985 (N_5985,N_4206,N_4147);
or U5986 (N_5986,N_4195,N_3982);
nor U5987 (N_5987,N_4172,N_3223);
nand U5988 (N_5988,N_3347,N_4124);
nand U5989 (N_5989,N_4199,N_3872);
and U5990 (N_5990,N_4039,N_3479);
or U5991 (N_5991,N_3643,N_3288);
nand U5992 (N_5992,N_3691,N_3437);
and U5993 (N_5993,N_3257,N_3236);
and U5994 (N_5994,N_3557,N_3107);
and U5995 (N_5995,N_3020,N_4182);
or U5996 (N_5996,N_3239,N_3820);
or U5997 (N_5997,N_3136,N_4005);
nand U5998 (N_5998,N_3626,N_3797);
nor U5999 (N_5999,N_3598,N_3795);
or U6000 (N_6000,N_5158,N_5085);
and U6001 (N_6001,N_5156,N_4552);
nor U6002 (N_6002,N_4597,N_5954);
nor U6003 (N_6003,N_5846,N_5637);
or U6004 (N_6004,N_4503,N_5262);
nand U6005 (N_6005,N_4847,N_5609);
and U6006 (N_6006,N_5576,N_5256);
or U6007 (N_6007,N_5558,N_5688);
nand U6008 (N_6008,N_4828,N_5932);
or U6009 (N_6009,N_5300,N_5916);
and U6010 (N_6010,N_4730,N_5957);
nand U6011 (N_6011,N_5818,N_5137);
and U6012 (N_6012,N_5090,N_4733);
nor U6013 (N_6013,N_5853,N_5810);
nand U6014 (N_6014,N_4893,N_4599);
nor U6015 (N_6015,N_5131,N_5623);
nand U6016 (N_6016,N_5759,N_4740);
or U6017 (N_6017,N_5923,N_4727);
nor U6018 (N_6018,N_5612,N_5074);
or U6019 (N_6019,N_5313,N_5679);
or U6020 (N_6020,N_5439,N_4765);
nor U6021 (N_6021,N_5726,N_5010);
and U6022 (N_6022,N_5038,N_4735);
nand U6023 (N_6023,N_5646,N_5870);
and U6024 (N_6024,N_5253,N_5906);
nor U6025 (N_6025,N_5662,N_5023);
nand U6026 (N_6026,N_5036,N_5845);
nand U6027 (N_6027,N_5015,N_5761);
nand U6028 (N_6028,N_5033,N_5611);
nor U6029 (N_6029,N_5482,N_5016);
or U6030 (N_6030,N_5035,N_4671);
nand U6031 (N_6031,N_5488,N_5054);
nand U6032 (N_6032,N_4659,N_5392);
and U6033 (N_6033,N_4941,N_5711);
nand U6034 (N_6034,N_4983,N_4592);
and U6035 (N_6035,N_5095,N_4668);
nor U6036 (N_6036,N_4926,N_5433);
or U6037 (N_6037,N_5370,N_4664);
nor U6038 (N_6038,N_5922,N_5438);
and U6039 (N_6039,N_5776,N_4981);
nand U6040 (N_6040,N_5804,N_4624);
or U6041 (N_6041,N_5465,N_4761);
nor U6042 (N_6042,N_4631,N_5700);
and U6043 (N_6043,N_5094,N_4561);
and U6044 (N_6044,N_4897,N_5007);
nand U6045 (N_6045,N_4793,N_5964);
or U6046 (N_6046,N_5871,N_5334);
and U6047 (N_6047,N_4999,N_5258);
nor U6048 (N_6048,N_4822,N_5725);
nor U6049 (N_6049,N_4850,N_5824);
nor U6050 (N_6050,N_5049,N_5037);
or U6051 (N_6051,N_5944,N_5750);
and U6052 (N_6052,N_5467,N_4694);
nand U6053 (N_6053,N_4997,N_5398);
nor U6054 (N_6054,N_5254,N_5765);
or U6055 (N_6055,N_5430,N_5595);
nand U6056 (N_6056,N_5435,N_5244);
nand U6057 (N_6057,N_5155,N_5476);
nand U6058 (N_6058,N_5118,N_5089);
nand U6059 (N_6059,N_5802,N_5250);
or U6060 (N_6060,N_5971,N_5738);
and U6061 (N_6061,N_5167,N_4688);
nand U6062 (N_6062,N_4809,N_5494);
nand U6063 (N_6063,N_4900,N_4549);
nand U6064 (N_6064,N_5998,N_5841);
and U6065 (N_6065,N_5934,N_5891);
nand U6066 (N_6066,N_5615,N_5247);
and U6067 (N_6067,N_4589,N_5717);
nand U6068 (N_6068,N_4584,N_4689);
and U6069 (N_6069,N_5358,N_4810);
or U6070 (N_6070,N_5575,N_5983);
or U6071 (N_6071,N_4917,N_4598);
nor U6072 (N_6072,N_5965,N_4633);
or U6073 (N_6073,N_5703,N_5315);
nand U6074 (N_6074,N_5625,N_5568);
or U6075 (N_6075,N_5865,N_4530);
and U6076 (N_6076,N_4968,N_5390);
and U6077 (N_6077,N_5894,N_5861);
nor U6078 (N_6078,N_5563,N_4988);
or U6079 (N_6079,N_5276,N_5626);
nor U6080 (N_6080,N_4800,N_5753);
or U6081 (N_6081,N_5839,N_4881);
or U6082 (N_6082,N_5102,N_5082);
nand U6083 (N_6083,N_5422,N_4557);
nor U6084 (N_6084,N_4879,N_4690);
nand U6085 (N_6085,N_5748,N_5365);
nor U6086 (N_6086,N_4936,N_4617);
and U6087 (N_6087,N_4675,N_4885);
nand U6088 (N_6088,N_4665,N_5855);
nor U6089 (N_6089,N_5526,N_5681);
and U6090 (N_6090,N_5063,N_4839);
and U6091 (N_6091,N_5421,N_5785);
nor U6092 (N_6092,N_5064,N_4798);
or U6093 (N_6093,N_5402,N_5831);
nand U6094 (N_6094,N_4512,N_4529);
or U6095 (N_6095,N_5573,N_5309);
nand U6096 (N_6096,N_5863,N_5455);
or U6097 (N_6097,N_5992,N_5875);
nor U6098 (N_6098,N_4860,N_4628);
or U6099 (N_6099,N_5683,N_5006);
or U6100 (N_6100,N_5990,N_5589);
or U6101 (N_6101,N_5565,N_4851);
nor U6102 (N_6102,N_5661,N_5552);
nand U6103 (N_6103,N_5508,N_5580);
or U6104 (N_6104,N_4612,N_5379);
nand U6105 (N_6105,N_4776,N_4823);
or U6106 (N_6106,N_5788,N_5705);
or U6107 (N_6107,N_5440,N_4952);
nand U6108 (N_6108,N_5252,N_4801);
and U6109 (N_6109,N_5867,N_4666);
or U6110 (N_6110,N_5574,N_5296);
nor U6111 (N_6111,N_5341,N_5933);
xnor U6112 (N_6112,N_5235,N_5004);
nor U6113 (N_6113,N_5175,N_5086);
nor U6114 (N_6114,N_4869,N_5275);
nand U6115 (N_6115,N_5851,N_5177);
nand U6116 (N_6116,N_5666,N_5278);
or U6117 (N_6117,N_5525,N_4836);
and U6118 (N_6118,N_4741,N_5745);
nand U6119 (N_6119,N_4635,N_5671);
nor U6120 (N_6120,N_5701,N_5409);
nand U6121 (N_6121,N_4901,N_5687);
nor U6122 (N_6122,N_5635,N_4891);
or U6123 (N_6123,N_4804,N_5585);
nand U6124 (N_6124,N_4830,N_5081);
or U6125 (N_6125,N_5113,N_4928);
nand U6126 (N_6126,N_5133,N_5521);
or U6127 (N_6127,N_5047,N_5862);
and U6128 (N_6128,N_5075,N_5881);
or U6129 (N_6129,N_5491,N_5187);
or U6130 (N_6130,N_5767,N_5647);
nand U6131 (N_6131,N_5996,N_5678);
nand U6132 (N_6132,N_4616,N_5034);
nor U6133 (N_6133,N_5069,N_4710);
nor U6134 (N_6134,N_5271,N_5413);
or U6135 (N_6135,N_5099,N_5215);
or U6136 (N_6136,N_4626,N_4532);
nor U6137 (N_6137,N_5393,N_5273);
and U6138 (N_6138,N_5970,N_5660);
nand U6139 (N_6139,N_5925,N_5196);
or U6140 (N_6140,N_4718,N_5578);
or U6141 (N_6141,N_4760,N_5436);
and U6142 (N_6142,N_5559,N_5835);
nand U6143 (N_6143,N_5060,N_5210);
nor U6144 (N_6144,N_5537,N_4551);
or U6145 (N_6145,N_5968,N_4536);
nand U6146 (N_6146,N_4591,N_4590);
nand U6147 (N_6147,N_4511,N_4656);
or U6148 (N_6148,N_4709,N_5652);
and U6149 (N_6149,N_5415,N_5386);
nor U6150 (N_6150,N_5193,N_5050);
nor U6151 (N_6151,N_5424,N_5805);
nand U6152 (N_6152,N_4622,N_5773);
nor U6153 (N_6153,N_4946,N_4767);
and U6154 (N_6154,N_5694,N_4751);
nand U6155 (N_6155,N_5551,N_5527);
nand U6156 (N_6156,N_5170,N_5189);
nor U6157 (N_6157,N_4764,N_5361);
or U6158 (N_6158,N_5103,N_5909);
nor U6159 (N_6159,N_4802,N_5985);
and U6160 (N_6160,N_5307,N_5493);
or U6161 (N_6161,N_4782,N_5115);
nor U6162 (N_6162,N_4962,N_5326);
or U6163 (N_6163,N_4636,N_5344);
or U6164 (N_6164,N_4747,N_4570);
and U6165 (N_6165,N_5993,N_5257);
nor U6166 (N_6166,N_5728,N_5472);
or U6167 (N_6167,N_4501,N_4819);
and U6168 (N_6168,N_4898,N_5766);
nor U6169 (N_6169,N_4995,N_4517);
nor U6170 (N_6170,N_5991,N_5668);
or U6171 (N_6171,N_4867,N_4522);
or U6172 (N_6172,N_4657,N_5684);
or U6173 (N_6173,N_4533,N_5443);
nor U6174 (N_6174,N_4976,N_5594);
and U6175 (N_6175,N_5907,N_5640);
xor U6176 (N_6176,N_5619,N_5718);
and U6177 (N_6177,N_5483,N_5447);
nor U6178 (N_6178,N_5106,N_4837);
and U6179 (N_6179,N_5799,N_5363);
nor U6180 (N_6180,N_5534,N_4854);
or U6181 (N_6181,N_5351,N_4534);
nor U6182 (N_6182,N_4775,N_5446);
and U6183 (N_6183,N_5966,N_4874);
nand U6184 (N_6184,N_4527,N_5471);
or U6185 (N_6185,N_4623,N_4965);
or U6186 (N_6186,N_5530,N_5065);
nor U6187 (N_6187,N_5984,N_4609);
nand U6188 (N_6188,N_5887,N_5227);
and U6189 (N_6189,N_5211,N_5066);
or U6190 (N_6190,N_5259,N_4621);
nor U6191 (N_6191,N_5653,N_5739);
and U6192 (N_6192,N_5204,N_4739);
or U6193 (N_6193,N_4920,N_5588);
nor U6194 (N_6194,N_4580,N_5457);
nand U6195 (N_6195,N_5444,N_4725);
or U6196 (N_6196,N_5762,N_4648);
and U6197 (N_6197,N_4519,N_5132);
nor U6198 (N_6198,N_5473,N_5495);
nand U6199 (N_6199,N_4896,N_4955);
nor U6200 (N_6200,N_5502,N_5280);
and U6201 (N_6201,N_5866,N_4732);
or U6202 (N_6202,N_4913,N_5655);
or U6203 (N_6203,N_5892,N_4959);
nand U6204 (N_6204,N_5453,N_5190);
or U6205 (N_6205,N_5771,N_4514);
nand U6206 (N_6206,N_4607,N_5667);
and U6207 (N_6207,N_5590,N_4707);
or U6208 (N_6208,N_5607,N_5041);
or U6209 (N_6209,N_5868,N_4510);
nand U6210 (N_6210,N_5289,N_5009);
nand U6211 (N_6211,N_5736,N_5889);
nor U6212 (N_6212,N_4771,N_5591);
nor U6213 (N_6213,N_5543,N_4556);
nand U6214 (N_6214,N_4957,N_5032);
nor U6215 (N_6215,N_5121,N_5740);
and U6216 (N_6216,N_4611,N_5019);
nor U6217 (N_6217,N_5481,N_5270);
nor U6218 (N_6218,N_5790,N_4980);
and U6219 (N_6219,N_4708,N_5396);
nand U6220 (N_6220,N_5397,N_4978);
nor U6221 (N_6221,N_5228,N_5223);
and U6222 (N_6222,N_4562,N_4729);
or U6223 (N_6223,N_4832,N_4588);
nor U6224 (N_6224,N_5618,N_5821);
or U6225 (N_6225,N_5973,N_5333);
nor U6226 (N_6226,N_5939,N_5729);
or U6227 (N_6227,N_5389,N_4660);
and U6228 (N_6228,N_4878,N_5381);
or U6229 (N_6229,N_5355,N_4606);
nor U6230 (N_6230,N_4960,N_5305);
xor U6231 (N_6231,N_4964,N_5179);
nand U6232 (N_6232,N_5786,N_5431);
nor U6233 (N_6233,N_5913,N_5140);
nor U6234 (N_6234,N_5336,N_5027);
or U6235 (N_6235,N_5169,N_5956);
nand U6236 (N_6236,N_4742,N_4676);
nor U6237 (N_6237,N_5428,N_5100);
or U6238 (N_6238,N_5876,N_5423);
nand U6239 (N_6239,N_5345,N_5621);
and U6240 (N_6240,N_5741,N_5632);
xor U6241 (N_6241,N_4903,N_5849);
or U6242 (N_6242,N_5459,N_5936);
and U6243 (N_6243,N_4994,N_5878);
nor U6244 (N_6244,N_5260,N_4788);
or U6245 (N_6245,N_4655,N_4686);
and U6246 (N_6246,N_5942,N_5859);
nand U6247 (N_6247,N_5564,N_5012);
nor U6248 (N_6248,N_5157,N_4772);
nand U6249 (N_6249,N_5627,N_4778);
or U6250 (N_6250,N_5480,N_5756);
or U6251 (N_6251,N_5828,N_4949);
or U6252 (N_6252,N_5644,N_5292);
and U6253 (N_6253,N_4565,N_5524);
nand U6254 (N_6254,N_5138,N_4963);
and U6255 (N_6255,N_4989,N_4774);
nand U6256 (N_6256,N_5221,N_4546);
nand U6257 (N_6257,N_5731,N_4834);
nor U6258 (N_6258,N_5324,N_5418);
or U6259 (N_6259,N_5201,N_4572);
or U6260 (N_6260,N_4757,N_4639);
or U6261 (N_6261,N_4567,N_5689);
and U6262 (N_6262,N_5205,N_5555);
nor U6263 (N_6263,N_4814,N_5323);
and U6264 (N_6264,N_5910,N_5322);
nand U6265 (N_6265,N_5056,N_4991);
or U6266 (N_6266,N_4560,N_4605);
and U6267 (N_6267,N_5164,N_4642);
nand U6268 (N_6268,N_5067,N_5371);
or U6269 (N_6269,N_5125,N_5994);
and U6270 (N_6270,N_4791,N_5874);
nor U6271 (N_6271,N_5407,N_4558);
and U6272 (N_6272,N_5793,N_5403);
and U6273 (N_6273,N_5148,N_5634);
nand U6274 (N_6274,N_5293,N_4614);
or U6275 (N_6275,N_5057,N_5380);
nand U6276 (N_6276,N_5335,N_5707);
xor U6277 (N_6277,N_4559,N_5497);
nor U6278 (N_6278,N_5274,N_4603);
or U6279 (N_6279,N_4803,N_5918);
nand U6280 (N_6280,N_5721,N_5116);
xor U6281 (N_6281,N_5781,N_5893);
nand U6282 (N_6282,N_5837,N_4696);
and U6283 (N_6283,N_5515,N_4883);
nor U6284 (N_6284,N_4578,N_5958);
and U6285 (N_6285,N_4669,N_5988);
nand U6286 (N_6286,N_5022,N_5226);
nor U6287 (N_6287,N_4973,N_5429);
nor U6288 (N_6288,N_5829,N_4706);
or U6289 (N_6289,N_5977,N_4835);
or U6290 (N_6290,N_5325,N_4922);
or U6291 (N_6291,N_4911,N_4613);
and U6292 (N_6292,N_4647,N_5774);
and U6293 (N_6293,N_5822,N_5489);
nor U6294 (N_6294,N_5107,N_5570);
nor U6295 (N_6295,N_4744,N_5416);
nand U6296 (N_6296,N_5927,N_5195);
and U6297 (N_6297,N_5921,N_5528);
or U6298 (N_6298,N_5329,N_5359);
nand U6299 (N_6299,N_4939,N_4638);
nand U6300 (N_6300,N_4826,N_5174);
nand U6301 (N_6301,N_5680,N_4700);
nand U6302 (N_6302,N_4855,N_4750);
nand U6303 (N_6303,N_4521,N_5940);
or U6304 (N_6304,N_4784,N_4990);
and U6305 (N_6305,N_5648,N_4912);
and U6306 (N_6306,N_4754,N_5224);
or U6307 (N_6307,N_4977,N_5354);
and U6308 (N_6308,N_4852,N_5499);
and U6309 (N_6309,N_5061,N_5505);
and U6310 (N_6310,N_4672,N_5789);
and U6311 (N_6311,N_5111,N_4792);
or U6312 (N_6312,N_5070,N_5279);
nor U6313 (N_6313,N_4697,N_4610);
and U6314 (N_6314,N_5943,N_5979);
nor U6315 (N_6315,N_5542,N_5364);
nor U6316 (N_6316,N_5531,N_5306);
nor U6317 (N_6317,N_5030,N_5506);
or U6318 (N_6318,N_4927,N_5147);
nand U6319 (N_6319,N_5059,N_5243);
nand U6320 (N_6320,N_4644,N_4880);
nor U6321 (N_6321,N_4890,N_4745);
nand U6322 (N_6322,N_4843,N_5842);
and U6323 (N_6323,N_5484,N_5732);
nor U6324 (N_6324,N_5911,N_4889);
and U6325 (N_6325,N_4538,N_5477);
and U6326 (N_6326,N_5475,N_5240);
or U6327 (N_6327,N_5523,N_5490);
and U6328 (N_6328,N_5544,N_4691);
nor U6329 (N_6329,N_5955,N_5860);
and U6330 (N_6330,N_4789,N_4717);
and U6331 (N_6331,N_4719,N_5161);
nand U6332 (N_6332,N_5599,N_5895);
nand U6333 (N_6333,N_5929,N_4820);
nand U6334 (N_6334,N_4619,N_4579);
nor U6335 (N_6335,N_4865,N_5451);
and U6336 (N_6336,N_5154,N_5952);
or U6337 (N_6337,N_5743,N_5562);
xor U6338 (N_6338,N_4513,N_4544);
or U6339 (N_6339,N_5328,N_5775);
nand U6340 (N_6340,N_5046,N_4554);
nor U6341 (N_6341,N_5975,N_5385);
nor U6342 (N_6342,N_5468,N_5083);
or U6343 (N_6343,N_4526,N_5522);
or U6344 (N_6344,N_4970,N_5222);
nor U6345 (N_6345,N_5659,N_4569);
or U6346 (N_6346,N_5784,N_5657);
and U6347 (N_6347,N_4692,N_5803);
and U6348 (N_6348,N_5225,N_5062);
nor U6349 (N_6349,N_5299,N_5649);
nor U6350 (N_6350,N_5624,N_5545);
nand U6351 (N_6351,N_5520,N_5031);
nor U6352 (N_6352,N_5613,N_5281);
or U6353 (N_6353,N_4918,N_5087);
xnor U6354 (N_6354,N_4705,N_4866);
nor U6355 (N_6355,N_5935,N_5606);
nor U6356 (N_6356,N_5685,N_5610);
and U6357 (N_6357,N_5742,N_4915);
nand U6358 (N_6358,N_4755,N_5304);
or U6359 (N_6359,N_4724,N_4781);
or U6360 (N_6360,N_5536,N_5213);
and U6361 (N_6361,N_4674,N_5598);
nor U6362 (N_6362,N_5924,N_4722);
or U6363 (N_6363,N_4811,N_5643);
and U6364 (N_6364,N_5233,N_5639);
nor U6365 (N_6365,N_4884,N_4673);
nand U6366 (N_6366,N_5556,N_5084);
and U6367 (N_6367,N_5414,N_5191);
and U6368 (N_6368,N_4892,N_5282);
or U6369 (N_6369,N_4736,N_5885);
nor U6370 (N_6370,N_5614,N_5744);
or U6371 (N_6371,N_5764,N_5360);
or U6372 (N_6372,N_5946,N_5630);
nand U6373 (N_6373,N_5230,N_4799);
and U6374 (N_6374,N_5708,N_4919);
nor U6375 (N_6375,N_5567,N_4662);
and U6376 (N_6376,N_5093,N_4974);
xnor U6377 (N_6377,N_4594,N_4726);
nand U6378 (N_6378,N_5128,N_5173);
nor U6379 (N_6379,N_4541,N_5974);
nor U6380 (N_6380,N_5417,N_5832);
nor U6381 (N_6381,N_5631,N_5723);
nand U6382 (N_6382,N_5026,N_5561);
or U6383 (N_6383,N_4773,N_5989);
nor U6384 (N_6384,N_4816,N_4678);
or U6385 (N_6385,N_4882,N_5622);
and U6386 (N_6386,N_5816,N_4844);
nand U6387 (N_6387,N_5665,N_5209);
nand U6388 (N_6388,N_5504,N_5456);
nor U6389 (N_6389,N_5586,N_4721);
and U6390 (N_6390,N_4779,N_5176);
and U6391 (N_6391,N_4524,N_4753);
nand U6392 (N_6392,N_5572,N_4738);
nor U6393 (N_6393,N_5884,N_4502);
or U6394 (N_6394,N_5104,N_4966);
nor U6395 (N_6395,N_5999,N_4743);
or U6396 (N_6396,N_5814,N_5404);
nand U6397 (N_6397,N_4758,N_4979);
nand U6398 (N_6398,N_4806,N_5145);
nor U6399 (N_6399,N_5168,N_5899);
or U6400 (N_6400,N_5068,N_5986);
nor U6401 (N_6401,N_4637,N_4861);
and U6402 (N_6402,N_5352,N_5419);
or U6403 (N_6403,N_5602,N_5003);
nand U6404 (N_6404,N_4573,N_5709);
and U6405 (N_6405,N_5265,N_5603);
and U6406 (N_6406,N_5327,N_5937);
and U6407 (N_6407,N_5620,N_5461);
or U6408 (N_6408,N_4703,N_5654);
nand U6409 (N_6409,N_5693,N_4734);
nor U6410 (N_6410,N_5020,N_4871);
nand U6411 (N_6411,N_5079,N_5458);
and U6412 (N_6412,N_5880,N_5827);
and U6413 (N_6413,N_5587,N_4749);
nand U6414 (N_6414,N_5124,N_5510);
nand U6415 (N_6415,N_5577,N_4998);
or U6416 (N_6416,N_5264,N_4608);
or U6417 (N_6417,N_4701,N_4907);
nor U6418 (N_6418,N_5864,N_5288);
or U6419 (N_6419,N_5088,N_5900);
nand U6420 (N_6420,N_4818,N_5848);
nand U6421 (N_6421,N_5162,N_5638);
or U6422 (N_6422,N_5199,N_4658);
or U6423 (N_6423,N_5912,N_5658);
or U6424 (N_6424,N_5291,N_4575);
and U6425 (N_6425,N_5149,N_5972);
and U6426 (N_6426,N_4595,N_5317);
nor U6427 (N_6427,N_4582,N_4704);
or U6428 (N_6428,N_5830,N_4996);
nor U6429 (N_6429,N_5408,N_4716);
nand U6430 (N_6430,N_4842,N_5812);
or U6431 (N_6431,N_5406,N_4650);
nor U6432 (N_6432,N_5501,N_5284);
nand U6433 (N_6433,N_4645,N_5486);
or U6434 (N_6434,N_5532,N_5077);
or U6435 (N_6435,N_5601,N_5263);
or U6436 (N_6436,N_4542,N_4571);
nand U6437 (N_6437,N_5350,N_5673);
and U6438 (N_6438,N_4956,N_5337);
or U6439 (N_6439,N_4543,N_4825);
or U6440 (N_6440,N_5847,N_5600);
and U6441 (N_6441,N_5377,N_5220);
or U6442 (N_6442,N_4653,N_4540);
nand U6443 (N_6443,N_4600,N_4947);
nand U6444 (N_6444,N_4785,N_5792);
nor U6445 (N_6445,N_5783,N_5246);
nand U6446 (N_6446,N_4935,N_4766);
and U6447 (N_6447,N_5682,N_5134);
and U6448 (N_6448,N_5114,N_4577);
nor U6449 (N_6449,N_4961,N_5734);
nor U6450 (N_6450,N_5616,N_5206);
nor U6451 (N_6451,N_4943,N_5126);
or U6452 (N_6452,N_5159,N_4585);
xnor U6453 (N_6453,N_5582,N_4862);
nand U6454 (N_6454,N_5208,N_5312);
and U6455 (N_6455,N_5139,N_5375);
nor U6456 (N_6456,N_4942,N_5931);
and U6457 (N_6457,N_5277,N_5400);
or U6458 (N_6458,N_5098,N_5549);
and U6459 (N_6459,N_5838,N_5078);
and U6460 (N_6460,N_5342,N_4993);
or U6461 (N_6461,N_5980,N_5513);
and U6462 (N_6462,N_4790,N_5242);
nor U6463 (N_6463,N_5928,N_4634);
nor U6464 (N_6464,N_5698,N_5941);
nor U6465 (N_6465,N_4905,N_4923);
or U6466 (N_6466,N_5782,N_4987);
nand U6467 (N_6467,N_4940,N_5963);
and U6468 (N_6468,N_5091,N_4858);
or U6469 (N_6469,N_4849,N_5695);
nor U6470 (N_6470,N_4831,N_4731);
or U6471 (N_6471,N_4953,N_5185);
nor U6472 (N_6472,N_5981,N_5755);
nand U6473 (N_6473,N_5150,N_5704);
or U6474 (N_6474,N_4870,N_5463);
and U6475 (N_6475,N_5770,N_5778);
nand U6476 (N_6476,N_4563,N_5691);
and U6477 (N_6477,N_4649,N_5163);
or U6478 (N_6478,N_5730,N_5540);
or U6479 (N_6479,N_5011,N_5000);
or U6480 (N_6480,N_5583,N_5496);
nor U6481 (N_6481,N_4508,N_4916);
nand U6482 (N_6482,N_5710,N_4746);
nand U6483 (N_6483,N_5153,N_4887);
and U6484 (N_6484,N_4972,N_4895);
or U6485 (N_6485,N_5642,N_5432);
and U6486 (N_6486,N_4520,N_4714);
and U6487 (N_6487,N_5391,N_4728);
and U6488 (N_6488,N_5427,N_5197);
nor U6489 (N_6489,N_4507,N_4627);
or U6490 (N_6490,N_5207,N_5897);
and U6491 (N_6491,N_5285,N_4812);
and U6492 (N_6492,N_5772,N_5593);
nand U6493 (N_6493,N_4643,N_5298);
and U6494 (N_6494,N_5401,N_4762);
nand U6495 (N_6495,N_4992,N_5130);
nor U6496 (N_6496,N_5362,N_4576);
and U6497 (N_6497,N_5706,N_4948);
or U6498 (N_6498,N_5470,N_5951);
nand U6499 (N_6499,N_5960,N_5042);
or U6500 (N_6500,N_5109,N_5119);
or U6501 (N_6501,N_4632,N_5071);
nor U6502 (N_6502,N_5498,N_4518);
nor U6503 (N_6503,N_5656,N_4528);
xnor U6504 (N_6504,N_5272,N_5791);
and U6505 (N_6505,N_4566,N_4906);
nand U6506 (N_6506,N_4568,N_4699);
nor U6507 (N_6507,N_5819,N_5395);
or U6508 (N_6508,N_4652,N_5017);
or U6509 (N_6509,N_5872,N_5366);
or U6510 (N_6510,N_5092,N_5249);
nor U6511 (N_6511,N_5357,N_4715);
and U6512 (N_6512,N_5604,N_5569);
nand U6513 (N_6513,N_4537,N_5953);
and U6514 (N_6514,N_5901,N_4768);
nand U6515 (N_6515,N_5464,N_5546);
nand U6516 (N_6516,N_5374,N_5557);
nand U6517 (N_6517,N_5025,N_5519);
and U6518 (N_6518,N_5348,N_5123);
or U6519 (N_6519,N_5382,N_4661);
or U6520 (N_6520,N_5080,N_5171);
nor U6521 (N_6521,N_4525,N_4564);
and U6522 (N_6522,N_4693,N_5807);
nor U6523 (N_6523,N_5840,N_4505);
nor U6524 (N_6524,N_5978,N_5663);
nor U6525 (N_6525,N_5127,N_4640);
nor U6526 (N_6526,N_5696,N_5232);
nor U6527 (N_6527,N_4856,N_5117);
nand U6528 (N_6528,N_5541,N_5768);
and U6529 (N_6529,N_5800,N_5437);
or U6530 (N_6530,N_5203,N_5919);
and U6531 (N_6531,N_5650,N_5314);
or U6532 (N_6532,N_5823,N_4824);
and U6533 (N_6533,N_5160,N_5969);
nor U6534 (N_6534,N_4813,N_5487);
xnor U6535 (N_6535,N_4574,N_4888);
or U6536 (N_6536,N_5538,N_5412);
or U6537 (N_6537,N_5686,N_4548);
and U6538 (N_6538,N_5474,N_5372);
nor U6539 (N_6539,N_5045,N_5479);
nor U6540 (N_6540,N_5218,N_4506);
nor U6541 (N_6541,N_5055,N_5617);
nor U6542 (N_6542,N_4930,N_5308);
nor U6543 (N_6543,N_5141,N_5320);
nor U6544 (N_6544,N_5028,N_5890);
nor U6545 (N_6545,N_4797,N_5198);
nand U6546 (N_6546,N_5714,N_4945);
nor U6547 (N_6547,N_5566,N_5388);
and U6548 (N_6548,N_5194,N_5758);
nand U6549 (N_6549,N_4763,N_5539);
or U6550 (N_6550,N_5511,N_4698);
or U6551 (N_6551,N_5261,N_5787);
nor U6552 (N_6552,N_4969,N_5883);
and U6553 (N_6553,N_5722,N_5949);
nand U6554 (N_6554,N_4827,N_5399);
nor U6555 (N_6555,N_4954,N_4681);
or U6556 (N_6556,N_5995,N_5096);
or U6557 (N_6557,N_4786,N_4759);
and U6558 (N_6558,N_4685,N_4944);
nor U6559 (N_6559,N_5675,N_4902);
and U6560 (N_6560,N_4670,N_4925);
and U6561 (N_6561,N_5267,N_5434);
nor U6562 (N_6562,N_5449,N_5869);
nand U6563 (N_6563,N_4817,N_4641);
nor U6564 (N_6564,N_5735,N_4654);
nor U6565 (N_6565,N_5982,N_5760);
and U6566 (N_6566,N_4875,N_4683);
nand U6567 (N_6567,N_5503,N_5553);
or U6568 (N_6568,N_5769,N_5383);
nand U6569 (N_6569,N_5441,N_4958);
and U6570 (N_6570,N_4535,N_5676);
and U6571 (N_6571,N_5733,N_5316);
or U6572 (N_6572,N_4752,N_5347);
nor U6573 (N_6573,N_5005,N_5592);
nand U6574 (N_6574,N_5727,N_5948);
or U6575 (N_6575,N_5798,N_5460);
or U6576 (N_6576,N_5002,N_5795);
or U6577 (N_6577,N_5237,N_5353);
nor U6578 (N_6578,N_5879,N_4795);
and U6579 (N_6579,N_5697,N_4848);
xnor U6580 (N_6580,N_5394,N_5346);
nor U6581 (N_6581,N_5844,N_5959);
nand U6582 (N_6582,N_4931,N_5420);
and U6583 (N_6583,N_4770,N_5651);
and U6584 (N_6584,N_4986,N_4821);
nand U6585 (N_6585,N_5692,N_5013);
or U6586 (N_6586,N_5142,N_4646);
or U6587 (N_6587,N_5410,N_5873);
nor U6588 (N_6588,N_5636,N_4924);
or U6589 (N_6589,N_5008,N_5677);
nor U6590 (N_6590,N_4846,N_5182);
and U6591 (N_6591,N_5165,N_5597);
or U6592 (N_6592,N_5251,N_5255);
nand U6593 (N_6593,N_5967,N_5229);
nor U6594 (N_6594,N_5516,N_5311);
nand U6595 (N_6595,N_5283,N_4794);
and U6596 (N_6596,N_5645,N_4845);
nor U6597 (N_6597,N_5571,N_5101);
or U6598 (N_6598,N_4531,N_5245);
nor U6599 (N_6599,N_5850,N_5076);
nand U6600 (N_6600,N_4840,N_5843);
and U6601 (N_6601,N_5896,N_4829);
nand U6602 (N_6602,N_5373,N_5796);
and U6603 (N_6603,N_4748,N_4971);
and U6604 (N_6604,N_5806,N_4910);
and U6605 (N_6605,N_4586,N_4787);
or U6606 (N_6606,N_4876,N_5720);
and U6607 (N_6607,N_5269,N_5122);
nor U6608 (N_6608,N_5178,N_4886);
nand U6609 (N_6609,N_5330,N_5001);
nand U6610 (N_6610,N_5166,N_4872);
xnor U6611 (N_6611,N_5836,N_4808);
or U6612 (N_6612,N_5926,N_5018);
nand U6613 (N_6613,N_4539,N_4682);
nand U6614 (N_6614,N_5340,N_5405);
or U6615 (N_6615,N_5719,N_4516);
nand U6616 (N_6616,N_4841,N_4593);
nor U6617 (N_6617,N_5297,N_5039);
or U6618 (N_6618,N_5833,N_5920);
nor U6619 (N_6619,N_5053,N_5462);
or U6620 (N_6620,N_5310,N_4509);
nor U6621 (N_6621,N_5605,N_5231);
nand U6622 (N_6622,N_5533,N_5529);
nand U6623 (N_6623,N_4515,N_4680);
nor U6624 (N_6624,N_4838,N_5445);
nor U6625 (N_6625,N_4663,N_4602);
xor U6626 (N_6626,N_5813,N_4904);
nor U6627 (N_6627,N_4863,N_5794);
and U6628 (N_6628,N_4937,N_5181);
nor U6629 (N_6629,N_4909,N_5641);
nand U6630 (N_6630,N_5904,N_5331);
nand U6631 (N_6631,N_5903,N_5136);
nor U6632 (N_6632,N_4967,N_4687);
nor U6633 (N_6633,N_4857,N_5302);
nor U6634 (N_6634,N_5239,N_5188);
or U6635 (N_6635,N_5815,N_5987);
nor U6636 (N_6636,N_5633,N_5338);
nor U6637 (N_6637,N_5024,N_5669);
nor U6638 (N_6638,N_4618,N_5048);
nand U6639 (N_6639,N_5518,N_5367);
or U6640 (N_6640,N_5608,N_5947);
or U6641 (N_6641,N_5411,N_5550);
and U6642 (N_6642,N_5110,N_5852);
and U6643 (N_6643,N_4807,N_4713);
nand U6644 (N_6644,N_5192,N_5777);
nand U6645 (N_6645,N_4982,N_5146);
and U6646 (N_6646,N_4581,N_5749);
nor U6647 (N_6647,N_5801,N_5143);
nor U6648 (N_6648,N_5961,N_4873);
nand U6649 (N_6649,N_5286,N_5200);
and U6650 (N_6650,N_4985,N_4864);
or U6651 (N_6651,N_4975,N_5715);
nand U6652 (N_6652,N_5180,N_5584);
and U6653 (N_6653,N_4695,N_4583);
or U6654 (N_6654,N_4780,N_5339);
nand U6655 (N_6655,N_4677,N_5450);
nand U6656 (N_6656,N_5780,N_5266);
nand U6657 (N_6657,N_5426,N_5674);
nor U6658 (N_6658,N_5135,N_5757);
nand U6659 (N_6659,N_4684,N_5811);
nand U6660 (N_6660,N_5287,N_5184);
nand U6661 (N_6661,N_5144,N_5858);
nand U6662 (N_6662,N_4667,N_5712);
and U6663 (N_6663,N_5294,N_5500);
and U6664 (N_6664,N_5214,N_5478);
nand U6665 (N_6665,N_4951,N_5172);
nor U6666 (N_6666,N_4929,N_5690);
nand U6667 (N_6667,N_5303,N_5517);
or U6668 (N_6668,N_5236,N_4523);
nor U6669 (N_6669,N_5120,N_5507);
nor U6670 (N_6670,N_4894,N_5664);
or U6671 (N_6671,N_5917,N_4550);
or U6672 (N_6672,N_5581,N_4651);
nand U6673 (N_6673,N_5763,N_5052);
nand U6674 (N_6674,N_4615,N_5183);
or U6675 (N_6675,N_5856,N_5629);
nand U6676 (N_6676,N_4853,N_5857);
and U6677 (N_6677,N_5186,N_5809);
nor U6678 (N_6678,N_5318,N_5825);
and U6679 (N_6679,N_5976,N_5535);
and U6680 (N_6680,N_5043,N_5915);
nor U6681 (N_6681,N_4796,N_4899);
or U6682 (N_6682,N_5129,N_5234);
nor U6683 (N_6683,N_5509,N_5746);
nand U6684 (N_6684,N_4500,N_5751);
or U6685 (N_6685,N_4504,N_4723);
and U6686 (N_6686,N_4877,N_4921);
nand U6687 (N_6687,N_5152,N_5997);
nor U6688 (N_6688,N_5492,N_5882);
nor U6689 (N_6689,N_5295,N_5826);
or U6690 (N_6690,N_5097,N_5212);
or U6691 (N_6691,N_5241,N_5699);
nand U6692 (N_6692,N_5877,N_5108);
nor U6693 (N_6693,N_4547,N_4783);
and U6694 (N_6694,N_5014,N_5886);
and U6695 (N_6695,N_5902,N_5151);
nand U6696 (N_6696,N_4833,N_5051);
nand U6697 (N_6697,N_4934,N_5548);
nand U6698 (N_6698,N_5378,N_4604);
or U6699 (N_6699,N_5112,N_5817);
or U6700 (N_6700,N_5332,N_5469);
or U6701 (N_6701,N_5724,N_5702);
nor U6702 (N_6702,N_4805,N_5387);
nor U6703 (N_6703,N_5021,N_5290);
and U6704 (N_6704,N_5930,N_5716);
or U6705 (N_6705,N_4950,N_5238);
and U6706 (N_6706,N_5219,N_4545);
and U6707 (N_6707,N_5452,N_5105);
or U6708 (N_6708,N_5672,N_5898);
or U6709 (N_6709,N_5514,N_5448);
nor U6710 (N_6710,N_4914,N_4868);
or U6711 (N_6711,N_5073,N_5376);
nand U6712 (N_6712,N_5834,N_5747);
nand U6713 (N_6713,N_5321,N_5072);
nand U6714 (N_6714,N_5779,N_5216);
and U6715 (N_6715,N_5058,N_4908);
nor U6716 (N_6716,N_5217,N_4702);
nand U6717 (N_6717,N_5356,N_5554);
nor U6718 (N_6718,N_4737,N_5888);
and U6719 (N_6719,N_4630,N_5914);
nand U6720 (N_6720,N_5945,N_4679);
nor U6721 (N_6721,N_5905,N_5752);
or U6722 (N_6722,N_5369,N_4625);
or U6723 (N_6723,N_5670,N_4777);
nand U6724 (N_6724,N_5029,N_5349);
nand U6725 (N_6725,N_4601,N_5044);
or U6726 (N_6726,N_5384,N_5754);
nor U6727 (N_6727,N_5579,N_5797);
nor U6728 (N_6728,N_5547,N_5854);
and U6729 (N_6729,N_4933,N_5713);
nand U6730 (N_6730,N_5908,N_5938);
nand U6731 (N_6731,N_5628,N_4932);
and U6732 (N_6732,N_5425,N_4555);
nand U6733 (N_6733,N_4553,N_5442);
nor U6734 (N_6734,N_4587,N_4984);
nand U6735 (N_6735,N_5596,N_5319);
and U6736 (N_6736,N_4769,N_5950);
nand U6737 (N_6737,N_4596,N_5737);
nor U6738 (N_6738,N_5040,N_4620);
xor U6739 (N_6739,N_4938,N_4756);
and U6740 (N_6740,N_4711,N_5343);
nand U6741 (N_6741,N_5368,N_4629);
and U6742 (N_6742,N_5202,N_5301);
and U6743 (N_6743,N_4815,N_5808);
nand U6744 (N_6744,N_4712,N_5454);
xor U6745 (N_6745,N_5512,N_4859);
xor U6746 (N_6746,N_5560,N_5268);
or U6747 (N_6747,N_5962,N_5485);
xnor U6748 (N_6748,N_5466,N_5248);
nor U6749 (N_6749,N_5820,N_4720);
xor U6750 (N_6750,N_4507,N_4626);
and U6751 (N_6751,N_4958,N_5537);
nor U6752 (N_6752,N_5456,N_4723);
nand U6753 (N_6753,N_5883,N_4988);
and U6754 (N_6754,N_5557,N_5086);
and U6755 (N_6755,N_5702,N_5749);
nor U6756 (N_6756,N_4890,N_5762);
or U6757 (N_6757,N_5368,N_5217);
and U6758 (N_6758,N_5958,N_5646);
nand U6759 (N_6759,N_5218,N_5357);
nor U6760 (N_6760,N_5062,N_5456);
nor U6761 (N_6761,N_4993,N_5318);
or U6762 (N_6762,N_5336,N_5400);
and U6763 (N_6763,N_5630,N_5663);
and U6764 (N_6764,N_4954,N_4968);
and U6765 (N_6765,N_5230,N_4891);
and U6766 (N_6766,N_5089,N_4700);
and U6767 (N_6767,N_5738,N_5393);
nor U6768 (N_6768,N_4777,N_4600);
and U6769 (N_6769,N_5093,N_4869);
or U6770 (N_6770,N_5725,N_4634);
nand U6771 (N_6771,N_5546,N_5473);
nand U6772 (N_6772,N_5218,N_5702);
and U6773 (N_6773,N_4996,N_5561);
nand U6774 (N_6774,N_5485,N_5233);
nor U6775 (N_6775,N_4852,N_5589);
xor U6776 (N_6776,N_5243,N_5536);
or U6777 (N_6777,N_5209,N_5141);
nor U6778 (N_6778,N_5275,N_4613);
and U6779 (N_6779,N_4996,N_5350);
or U6780 (N_6780,N_5967,N_5937);
and U6781 (N_6781,N_5288,N_5472);
and U6782 (N_6782,N_5672,N_5656);
nor U6783 (N_6783,N_5647,N_5132);
nand U6784 (N_6784,N_5231,N_5088);
nor U6785 (N_6785,N_4891,N_4731);
nand U6786 (N_6786,N_4714,N_4935);
nor U6787 (N_6787,N_5009,N_4999);
or U6788 (N_6788,N_4645,N_5585);
and U6789 (N_6789,N_4779,N_5326);
nor U6790 (N_6790,N_4508,N_5816);
nor U6791 (N_6791,N_5321,N_4673);
nor U6792 (N_6792,N_5048,N_5354);
or U6793 (N_6793,N_5756,N_5074);
nand U6794 (N_6794,N_5734,N_5269);
nor U6795 (N_6795,N_5627,N_5966);
or U6796 (N_6796,N_5524,N_5485);
and U6797 (N_6797,N_5672,N_4585);
nand U6798 (N_6798,N_5546,N_4831);
or U6799 (N_6799,N_5468,N_5340);
nor U6800 (N_6800,N_4940,N_5873);
or U6801 (N_6801,N_5986,N_4647);
or U6802 (N_6802,N_5674,N_5841);
or U6803 (N_6803,N_4848,N_4595);
nand U6804 (N_6804,N_5732,N_4915);
nor U6805 (N_6805,N_4727,N_5208);
nor U6806 (N_6806,N_4842,N_5608);
or U6807 (N_6807,N_5391,N_4897);
or U6808 (N_6808,N_4761,N_5903);
nor U6809 (N_6809,N_5088,N_5549);
and U6810 (N_6810,N_4522,N_5185);
nand U6811 (N_6811,N_4910,N_5042);
or U6812 (N_6812,N_5213,N_5451);
nor U6813 (N_6813,N_4622,N_5711);
nand U6814 (N_6814,N_5400,N_4664);
nor U6815 (N_6815,N_5010,N_5195);
and U6816 (N_6816,N_4576,N_4646);
and U6817 (N_6817,N_5323,N_4732);
nor U6818 (N_6818,N_4567,N_5336);
and U6819 (N_6819,N_5047,N_5071);
nor U6820 (N_6820,N_5511,N_5830);
nor U6821 (N_6821,N_5107,N_4701);
nor U6822 (N_6822,N_4657,N_5174);
and U6823 (N_6823,N_4769,N_4576);
nand U6824 (N_6824,N_5304,N_4815);
or U6825 (N_6825,N_5852,N_5659);
nor U6826 (N_6826,N_5023,N_5955);
and U6827 (N_6827,N_4945,N_5881);
nor U6828 (N_6828,N_5051,N_4901);
nand U6829 (N_6829,N_5368,N_4533);
or U6830 (N_6830,N_4964,N_4710);
or U6831 (N_6831,N_5594,N_5269);
and U6832 (N_6832,N_4963,N_4882);
and U6833 (N_6833,N_5084,N_5627);
nor U6834 (N_6834,N_5633,N_5245);
nand U6835 (N_6835,N_5677,N_5383);
and U6836 (N_6836,N_5783,N_5726);
xor U6837 (N_6837,N_5512,N_5060);
and U6838 (N_6838,N_5787,N_5908);
nand U6839 (N_6839,N_4716,N_5879);
xnor U6840 (N_6840,N_4943,N_4768);
and U6841 (N_6841,N_4628,N_4539);
nand U6842 (N_6842,N_5190,N_5321);
or U6843 (N_6843,N_4851,N_5378);
nand U6844 (N_6844,N_5966,N_4834);
and U6845 (N_6845,N_4626,N_5578);
nor U6846 (N_6846,N_5427,N_5082);
and U6847 (N_6847,N_5935,N_4586);
and U6848 (N_6848,N_5518,N_5067);
or U6849 (N_6849,N_5457,N_5769);
and U6850 (N_6850,N_5728,N_5910);
nor U6851 (N_6851,N_5431,N_5541);
nand U6852 (N_6852,N_5785,N_5064);
or U6853 (N_6853,N_5316,N_5087);
nand U6854 (N_6854,N_5189,N_5866);
and U6855 (N_6855,N_5893,N_4986);
nor U6856 (N_6856,N_5997,N_4693);
nand U6857 (N_6857,N_4569,N_4850);
xor U6858 (N_6858,N_5929,N_5214);
nand U6859 (N_6859,N_5958,N_4913);
nor U6860 (N_6860,N_5573,N_5256);
or U6861 (N_6861,N_4936,N_4695);
nor U6862 (N_6862,N_5237,N_4868);
nand U6863 (N_6863,N_5630,N_4828);
nor U6864 (N_6864,N_5555,N_4873);
nand U6865 (N_6865,N_5512,N_5858);
and U6866 (N_6866,N_5053,N_5187);
nand U6867 (N_6867,N_4610,N_4857);
nor U6868 (N_6868,N_5990,N_4600);
nor U6869 (N_6869,N_5886,N_5737);
nand U6870 (N_6870,N_5683,N_5871);
and U6871 (N_6871,N_5543,N_5408);
or U6872 (N_6872,N_5358,N_4713);
nor U6873 (N_6873,N_5752,N_4887);
or U6874 (N_6874,N_4669,N_4939);
or U6875 (N_6875,N_5624,N_5800);
xor U6876 (N_6876,N_5438,N_5322);
nor U6877 (N_6877,N_4710,N_5272);
and U6878 (N_6878,N_5098,N_5919);
nand U6879 (N_6879,N_5281,N_5497);
xnor U6880 (N_6880,N_5969,N_4711);
and U6881 (N_6881,N_5437,N_5502);
nand U6882 (N_6882,N_5818,N_5186);
nor U6883 (N_6883,N_5944,N_4993);
nor U6884 (N_6884,N_5785,N_5859);
nor U6885 (N_6885,N_5343,N_4629);
and U6886 (N_6886,N_5258,N_5289);
nand U6887 (N_6887,N_5780,N_5014);
nand U6888 (N_6888,N_5739,N_5456);
or U6889 (N_6889,N_5327,N_5557);
and U6890 (N_6890,N_4580,N_5174);
and U6891 (N_6891,N_5348,N_4852);
nand U6892 (N_6892,N_5309,N_5693);
or U6893 (N_6893,N_5316,N_5839);
and U6894 (N_6894,N_5219,N_5659);
or U6895 (N_6895,N_5397,N_5659);
nor U6896 (N_6896,N_5972,N_5682);
or U6897 (N_6897,N_5663,N_5139);
or U6898 (N_6898,N_5192,N_5841);
and U6899 (N_6899,N_5861,N_5096);
or U6900 (N_6900,N_5095,N_4776);
or U6901 (N_6901,N_5220,N_5841);
and U6902 (N_6902,N_5841,N_4562);
nor U6903 (N_6903,N_5760,N_5331);
and U6904 (N_6904,N_4643,N_4974);
nor U6905 (N_6905,N_4680,N_5234);
or U6906 (N_6906,N_4637,N_5623);
nor U6907 (N_6907,N_4856,N_4542);
nand U6908 (N_6908,N_5362,N_5491);
xor U6909 (N_6909,N_5300,N_4669);
nor U6910 (N_6910,N_5351,N_5635);
nor U6911 (N_6911,N_4699,N_5175);
or U6912 (N_6912,N_4651,N_5977);
nand U6913 (N_6913,N_5903,N_4974);
nor U6914 (N_6914,N_5921,N_5231);
nor U6915 (N_6915,N_4906,N_5755);
and U6916 (N_6916,N_5584,N_5099);
nand U6917 (N_6917,N_5433,N_4716);
and U6918 (N_6918,N_5189,N_5724);
nand U6919 (N_6919,N_5271,N_5140);
or U6920 (N_6920,N_4801,N_5852);
and U6921 (N_6921,N_5197,N_4751);
nor U6922 (N_6922,N_5394,N_5584);
and U6923 (N_6923,N_5452,N_5810);
nand U6924 (N_6924,N_5840,N_5502);
or U6925 (N_6925,N_5336,N_5216);
nand U6926 (N_6926,N_5253,N_5572);
and U6927 (N_6927,N_4830,N_5234);
or U6928 (N_6928,N_5093,N_5384);
or U6929 (N_6929,N_4971,N_5699);
and U6930 (N_6930,N_4880,N_5375);
nand U6931 (N_6931,N_4657,N_4720);
or U6932 (N_6932,N_5755,N_5822);
nand U6933 (N_6933,N_4544,N_5291);
and U6934 (N_6934,N_5488,N_4510);
nand U6935 (N_6935,N_5971,N_5899);
or U6936 (N_6936,N_4648,N_4622);
nand U6937 (N_6937,N_5549,N_4525);
and U6938 (N_6938,N_5674,N_4749);
nand U6939 (N_6939,N_5645,N_5732);
nand U6940 (N_6940,N_5849,N_5240);
or U6941 (N_6941,N_5182,N_5502);
or U6942 (N_6942,N_4514,N_4548);
nor U6943 (N_6943,N_5531,N_5559);
nor U6944 (N_6944,N_5628,N_5875);
and U6945 (N_6945,N_5422,N_4735);
nor U6946 (N_6946,N_5008,N_5449);
or U6947 (N_6947,N_4834,N_5375);
and U6948 (N_6948,N_5734,N_5470);
and U6949 (N_6949,N_5284,N_5898);
or U6950 (N_6950,N_5199,N_5594);
or U6951 (N_6951,N_5727,N_5489);
and U6952 (N_6952,N_4776,N_4807);
nor U6953 (N_6953,N_4599,N_5393);
or U6954 (N_6954,N_5212,N_4910);
xor U6955 (N_6955,N_5708,N_5515);
or U6956 (N_6956,N_5393,N_5166);
or U6957 (N_6957,N_4721,N_5254);
nor U6958 (N_6958,N_4516,N_5427);
nor U6959 (N_6959,N_4611,N_4871);
and U6960 (N_6960,N_5499,N_5442);
and U6961 (N_6961,N_4660,N_4944);
and U6962 (N_6962,N_5969,N_4633);
nand U6963 (N_6963,N_5198,N_4869);
nor U6964 (N_6964,N_4539,N_5804);
or U6965 (N_6965,N_4713,N_4598);
or U6966 (N_6966,N_5688,N_5734);
or U6967 (N_6967,N_4558,N_5865);
or U6968 (N_6968,N_5144,N_5280);
and U6969 (N_6969,N_4922,N_5488);
nor U6970 (N_6970,N_5500,N_5019);
xnor U6971 (N_6971,N_5339,N_5851);
nor U6972 (N_6972,N_4666,N_5541);
nor U6973 (N_6973,N_5914,N_5145);
nand U6974 (N_6974,N_5218,N_5937);
and U6975 (N_6975,N_5693,N_5743);
or U6976 (N_6976,N_5270,N_5243);
nand U6977 (N_6977,N_5959,N_5182);
nand U6978 (N_6978,N_5856,N_4796);
nand U6979 (N_6979,N_5127,N_4730);
or U6980 (N_6980,N_4738,N_5802);
or U6981 (N_6981,N_4759,N_4580);
nand U6982 (N_6982,N_4995,N_5742);
nor U6983 (N_6983,N_5746,N_4520);
nor U6984 (N_6984,N_5324,N_5420);
nand U6985 (N_6985,N_4726,N_5589);
and U6986 (N_6986,N_4593,N_5308);
nor U6987 (N_6987,N_5265,N_4825);
and U6988 (N_6988,N_5149,N_4713);
nand U6989 (N_6989,N_5510,N_5316);
and U6990 (N_6990,N_5605,N_5254);
nor U6991 (N_6991,N_4803,N_4942);
nor U6992 (N_6992,N_5941,N_5019);
and U6993 (N_6993,N_4723,N_5538);
or U6994 (N_6994,N_5457,N_4687);
nor U6995 (N_6995,N_4789,N_5040);
nor U6996 (N_6996,N_4723,N_4951);
and U6997 (N_6997,N_5192,N_5649);
nor U6998 (N_6998,N_4542,N_4782);
or U6999 (N_6999,N_5317,N_4553);
nand U7000 (N_7000,N_5235,N_4786);
nor U7001 (N_7001,N_4857,N_5693);
and U7002 (N_7002,N_5998,N_5187);
or U7003 (N_7003,N_5282,N_5004);
and U7004 (N_7004,N_5623,N_5636);
nor U7005 (N_7005,N_5552,N_5358);
or U7006 (N_7006,N_4710,N_4619);
or U7007 (N_7007,N_4997,N_4960);
and U7008 (N_7008,N_4645,N_5492);
nand U7009 (N_7009,N_5907,N_5633);
or U7010 (N_7010,N_4689,N_4822);
or U7011 (N_7011,N_5792,N_5678);
nand U7012 (N_7012,N_5040,N_5809);
nor U7013 (N_7013,N_5320,N_4630);
or U7014 (N_7014,N_5865,N_5092);
or U7015 (N_7015,N_5690,N_5483);
and U7016 (N_7016,N_5707,N_5952);
nand U7017 (N_7017,N_5392,N_5280);
and U7018 (N_7018,N_5990,N_4832);
or U7019 (N_7019,N_5764,N_5155);
xor U7020 (N_7020,N_5930,N_5420);
and U7021 (N_7021,N_5682,N_5037);
and U7022 (N_7022,N_5233,N_4599);
nand U7023 (N_7023,N_5714,N_5949);
and U7024 (N_7024,N_5200,N_4980);
or U7025 (N_7025,N_4932,N_5097);
or U7026 (N_7026,N_5736,N_5536);
and U7027 (N_7027,N_5731,N_4622);
nand U7028 (N_7028,N_5723,N_4752);
nor U7029 (N_7029,N_5713,N_4989);
and U7030 (N_7030,N_5115,N_5346);
nand U7031 (N_7031,N_5792,N_5980);
nor U7032 (N_7032,N_4606,N_5499);
nor U7033 (N_7033,N_5480,N_5122);
nor U7034 (N_7034,N_5581,N_5292);
nand U7035 (N_7035,N_4871,N_4705);
nand U7036 (N_7036,N_5014,N_5971);
nand U7037 (N_7037,N_5622,N_5398);
nor U7038 (N_7038,N_5108,N_4933);
or U7039 (N_7039,N_5374,N_5901);
or U7040 (N_7040,N_4881,N_5125);
nand U7041 (N_7041,N_4753,N_5929);
and U7042 (N_7042,N_5284,N_4714);
nor U7043 (N_7043,N_5140,N_5105);
or U7044 (N_7044,N_5429,N_4949);
nand U7045 (N_7045,N_5584,N_4652);
nor U7046 (N_7046,N_5152,N_5817);
nor U7047 (N_7047,N_5543,N_4516);
nor U7048 (N_7048,N_5679,N_4952);
nor U7049 (N_7049,N_4821,N_5013);
nand U7050 (N_7050,N_4746,N_5662);
or U7051 (N_7051,N_5528,N_5881);
nor U7052 (N_7052,N_4727,N_4637);
and U7053 (N_7053,N_5405,N_5505);
nor U7054 (N_7054,N_5444,N_4967);
and U7055 (N_7055,N_4647,N_4696);
or U7056 (N_7056,N_5326,N_4512);
or U7057 (N_7057,N_5798,N_4806);
or U7058 (N_7058,N_5473,N_5933);
nor U7059 (N_7059,N_4980,N_5961);
or U7060 (N_7060,N_4898,N_4741);
or U7061 (N_7061,N_5179,N_4516);
or U7062 (N_7062,N_5646,N_5566);
nor U7063 (N_7063,N_4599,N_5406);
or U7064 (N_7064,N_5849,N_5287);
and U7065 (N_7065,N_4848,N_4880);
nand U7066 (N_7066,N_5257,N_4961);
nor U7067 (N_7067,N_5093,N_5449);
nand U7068 (N_7068,N_5008,N_5127);
or U7069 (N_7069,N_5036,N_5157);
and U7070 (N_7070,N_5290,N_4764);
xor U7071 (N_7071,N_4891,N_4810);
nor U7072 (N_7072,N_4743,N_4868);
or U7073 (N_7073,N_5312,N_4854);
nor U7074 (N_7074,N_5443,N_4950);
or U7075 (N_7075,N_4660,N_5559);
nor U7076 (N_7076,N_4541,N_4671);
nor U7077 (N_7077,N_4970,N_5089);
or U7078 (N_7078,N_4695,N_4806);
nor U7079 (N_7079,N_4677,N_5859);
nand U7080 (N_7080,N_5355,N_5637);
xnor U7081 (N_7081,N_5177,N_4949);
xnor U7082 (N_7082,N_4998,N_5405);
and U7083 (N_7083,N_5755,N_5086);
nor U7084 (N_7084,N_5497,N_4747);
nand U7085 (N_7085,N_5478,N_4707);
nand U7086 (N_7086,N_4561,N_5512);
nand U7087 (N_7087,N_5080,N_5609);
or U7088 (N_7088,N_5383,N_4542);
or U7089 (N_7089,N_5796,N_5320);
and U7090 (N_7090,N_4873,N_4587);
nand U7091 (N_7091,N_4612,N_5183);
nand U7092 (N_7092,N_4741,N_4868);
nor U7093 (N_7093,N_5091,N_5337);
and U7094 (N_7094,N_5847,N_5288);
nand U7095 (N_7095,N_5772,N_4889);
nor U7096 (N_7096,N_5284,N_5671);
xnor U7097 (N_7097,N_4609,N_5380);
nand U7098 (N_7098,N_5498,N_5365);
and U7099 (N_7099,N_5592,N_5435);
nor U7100 (N_7100,N_4940,N_5294);
or U7101 (N_7101,N_5187,N_5476);
xnor U7102 (N_7102,N_4588,N_5408);
or U7103 (N_7103,N_4977,N_5413);
or U7104 (N_7104,N_4916,N_4785);
or U7105 (N_7105,N_4800,N_5825);
nand U7106 (N_7106,N_5286,N_5051);
nand U7107 (N_7107,N_4698,N_4878);
and U7108 (N_7108,N_4944,N_5866);
nand U7109 (N_7109,N_5603,N_4884);
and U7110 (N_7110,N_5191,N_5830);
nand U7111 (N_7111,N_4730,N_4781);
nor U7112 (N_7112,N_5024,N_5757);
nand U7113 (N_7113,N_4713,N_4660);
or U7114 (N_7114,N_4712,N_5147);
and U7115 (N_7115,N_5558,N_4647);
xnor U7116 (N_7116,N_5351,N_4980);
nor U7117 (N_7117,N_5481,N_5201);
or U7118 (N_7118,N_5456,N_5224);
and U7119 (N_7119,N_5555,N_5655);
or U7120 (N_7120,N_4586,N_5165);
and U7121 (N_7121,N_5785,N_4520);
nor U7122 (N_7122,N_5336,N_4813);
nor U7123 (N_7123,N_5839,N_4700);
and U7124 (N_7124,N_5799,N_4877);
nor U7125 (N_7125,N_5719,N_4544);
or U7126 (N_7126,N_5933,N_4736);
xnor U7127 (N_7127,N_5903,N_5285);
nand U7128 (N_7128,N_5700,N_4504);
nand U7129 (N_7129,N_4888,N_5205);
nand U7130 (N_7130,N_5803,N_5365);
nor U7131 (N_7131,N_4718,N_5210);
or U7132 (N_7132,N_5485,N_5963);
or U7133 (N_7133,N_5781,N_4787);
nand U7134 (N_7134,N_4943,N_4911);
and U7135 (N_7135,N_4808,N_5311);
or U7136 (N_7136,N_5271,N_5469);
or U7137 (N_7137,N_5202,N_4736);
and U7138 (N_7138,N_5125,N_5022);
nand U7139 (N_7139,N_5972,N_5572);
and U7140 (N_7140,N_4801,N_4918);
nor U7141 (N_7141,N_4598,N_5881);
and U7142 (N_7142,N_5202,N_5226);
or U7143 (N_7143,N_5064,N_5408);
nor U7144 (N_7144,N_5660,N_5931);
and U7145 (N_7145,N_5862,N_5266);
or U7146 (N_7146,N_5457,N_5191);
or U7147 (N_7147,N_4978,N_5800);
and U7148 (N_7148,N_5594,N_4648);
or U7149 (N_7149,N_5839,N_5905);
nor U7150 (N_7150,N_5658,N_4786);
nand U7151 (N_7151,N_4793,N_5431);
or U7152 (N_7152,N_5561,N_4918);
xnor U7153 (N_7153,N_5195,N_5484);
nor U7154 (N_7154,N_5728,N_5523);
nor U7155 (N_7155,N_5543,N_5332);
or U7156 (N_7156,N_5658,N_5439);
or U7157 (N_7157,N_5455,N_5133);
nor U7158 (N_7158,N_4968,N_4800);
nor U7159 (N_7159,N_4544,N_5093);
or U7160 (N_7160,N_5594,N_5170);
nand U7161 (N_7161,N_5983,N_4518);
nand U7162 (N_7162,N_4823,N_5675);
or U7163 (N_7163,N_5219,N_4970);
or U7164 (N_7164,N_5390,N_4617);
and U7165 (N_7165,N_4573,N_4966);
xor U7166 (N_7166,N_5702,N_5318);
or U7167 (N_7167,N_5242,N_4923);
nand U7168 (N_7168,N_5774,N_5137);
nand U7169 (N_7169,N_5851,N_5972);
nand U7170 (N_7170,N_4807,N_4679);
or U7171 (N_7171,N_4707,N_4765);
or U7172 (N_7172,N_4585,N_5194);
and U7173 (N_7173,N_4879,N_4547);
or U7174 (N_7174,N_5674,N_5548);
and U7175 (N_7175,N_4733,N_5666);
nand U7176 (N_7176,N_4804,N_4886);
nor U7177 (N_7177,N_4928,N_5321);
and U7178 (N_7178,N_5453,N_5620);
nor U7179 (N_7179,N_4821,N_5074);
and U7180 (N_7180,N_5721,N_5948);
nand U7181 (N_7181,N_5897,N_4817);
or U7182 (N_7182,N_5267,N_5594);
and U7183 (N_7183,N_5612,N_5909);
nand U7184 (N_7184,N_5815,N_5326);
or U7185 (N_7185,N_5061,N_5128);
nand U7186 (N_7186,N_5672,N_5561);
or U7187 (N_7187,N_5985,N_5162);
nand U7188 (N_7188,N_5410,N_5845);
nor U7189 (N_7189,N_5163,N_4607);
xnor U7190 (N_7190,N_5480,N_5485);
or U7191 (N_7191,N_4808,N_4818);
or U7192 (N_7192,N_5413,N_4561);
nand U7193 (N_7193,N_5342,N_5202);
nand U7194 (N_7194,N_5261,N_5861);
nand U7195 (N_7195,N_5568,N_5355);
nand U7196 (N_7196,N_4582,N_5147);
xnor U7197 (N_7197,N_4669,N_4680);
nor U7198 (N_7198,N_5715,N_4928);
or U7199 (N_7199,N_5536,N_5860);
or U7200 (N_7200,N_4757,N_4743);
nand U7201 (N_7201,N_5625,N_5378);
or U7202 (N_7202,N_4557,N_5463);
nor U7203 (N_7203,N_5347,N_5149);
nor U7204 (N_7204,N_5017,N_4851);
or U7205 (N_7205,N_5071,N_5039);
nand U7206 (N_7206,N_4549,N_5098);
nand U7207 (N_7207,N_5367,N_5379);
and U7208 (N_7208,N_5364,N_5821);
or U7209 (N_7209,N_5876,N_4783);
or U7210 (N_7210,N_5516,N_5616);
or U7211 (N_7211,N_4974,N_4713);
nor U7212 (N_7212,N_5736,N_5532);
and U7213 (N_7213,N_4877,N_4675);
nand U7214 (N_7214,N_5713,N_5965);
or U7215 (N_7215,N_5945,N_4792);
and U7216 (N_7216,N_5781,N_4785);
nand U7217 (N_7217,N_4850,N_4965);
and U7218 (N_7218,N_4531,N_5168);
and U7219 (N_7219,N_5506,N_5741);
or U7220 (N_7220,N_5722,N_5959);
and U7221 (N_7221,N_5654,N_5236);
or U7222 (N_7222,N_5700,N_5894);
nand U7223 (N_7223,N_5518,N_5955);
nand U7224 (N_7224,N_5861,N_5280);
or U7225 (N_7225,N_5452,N_4683);
or U7226 (N_7226,N_5124,N_5493);
nand U7227 (N_7227,N_5483,N_4893);
nand U7228 (N_7228,N_4955,N_4629);
and U7229 (N_7229,N_4647,N_5849);
nor U7230 (N_7230,N_5995,N_5391);
or U7231 (N_7231,N_5940,N_5728);
and U7232 (N_7232,N_5478,N_4965);
nor U7233 (N_7233,N_5539,N_5334);
nor U7234 (N_7234,N_5118,N_5932);
or U7235 (N_7235,N_5832,N_4976);
nand U7236 (N_7236,N_4908,N_4949);
xnor U7237 (N_7237,N_5795,N_5299);
nand U7238 (N_7238,N_4707,N_5117);
nor U7239 (N_7239,N_5612,N_5672);
nor U7240 (N_7240,N_5575,N_4645);
nand U7241 (N_7241,N_5015,N_5582);
nor U7242 (N_7242,N_4528,N_5677);
nor U7243 (N_7243,N_5779,N_5874);
nand U7244 (N_7244,N_5995,N_4947);
and U7245 (N_7245,N_5639,N_5309);
or U7246 (N_7246,N_5306,N_5319);
nand U7247 (N_7247,N_5181,N_5300);
nor U7248 (N_7248,N_5639,N_5728);
nor U7249 (N_7249,N_5607,N_5886);
or U7250 (N_7250,N_5465,N_5569);
nand U7251 (N_7251,N_5984,N_4689);
and U7252 (N_7252,N_5472,N_5732);
nand U7253 (N_7253,N_4751,N_4815);
nor U7254 (N_7254,N_4542,N_5354);
or U7255 (N_7255,N_4960,N_5505);
nand U7256 (N_7256,N_5064,N_5885);
and U7257 (N_7257,N_4552,N_4846);
nand U7258 (N_7258,N_5877,N_5460);
or U7259 (N_7259,N_5368,N_5670);
and U7260 (N_7260,N_5020,N_5110);
nor U7261 (N_7261,N_5242,N_5607);
or U7262 (N_7262,N_4584,N_4503);
nand U7263 (N_7263,N_4784,N_5163);
and U7264 (N_7264,N_4850,N_5286);
and U7265 (N_7265,N_5017,N_5942);
nor U7266 (N_7266,N_4721,N_5402);
nor U7267 (N_7267,N_5207,N_5749);
nand U7268 (N_7268,N_5116,N_5917);
nor U7269 (N_7269,N_4712,N_4750);
nand U7270 (N_7270,N_4992,N_5323);
xor U7271 (N_7271,N_5277,N_5796);
nand U7272 (N_7272,N_4524,N_4639);
or U7273 (N_7273,N_4769,N_5599);
or U7274 (N_7274,N_4999,N_5626);
nand U7275 (N_7275,N_5635,N_4857);
nor U7276 (N_7276,N_4941,N_5367);
and U7277 (N_7277,N_5690,N_4520);
nand U7278 (N_7278,N_5820,N_5961);
nand U7279 (N_7279,N_4723,N_4985);
nor U7280 (N_7280,N_5953,N_4775);
and U7281 (N_7281,N_4797,N_5147);
or U7282 (N_7282,N_5577,N_5355);
and U7283 (N_7283,N_4998,N_4679);
nor U7284 (N_7284,N_5180,N_5567);
or U7285 (N_7285,N_5943,N_5521);
and U7286 (N_7286,N_5836,N_4536);
nor U7287 (N_7287,N_4821,N_5854);
nor U7288 (N_7288,N_5414,N_5418);
or U7289 (N_7289,N_5552,N_4932);
and U7290 (N_7290,N_5073,N_5128);
and U7291 (N_7291,N_5120,N_4675);
and U7292 (N_7292,N_4833,N_5044);
nor U7293 (N_7293,N_4629,N_5348);
and U7294 (N_7294,N_5970,N_4872);
nand U7295 (N_7295,N_5001,N_5924);
nor U7296 (N_7296,N_5723,N_4613);
and U7297 (N_7297,N_5130,N_5185);
or U7298 (N_7298,N_5057,N_5083);
nor U7299 (N_7299,N_5446,N_5094);
nor U7300 (N_7300,N_5804,N_5679);
nand U7301 (N_7301,N_5132,N_5290);
or U7302 (N_7302,N_5255,N_4841);
or U7303 (N_7303,N_4950,N_5503);
nand U7304 (N_7304,N_5149,N_5760);
or U7305 (N_7305,N_4935,N_4841);
nand U7306 (N_7306,N_4731,N_5601);
or U7307 (N_7307,N_5130,N_4983);
and U7308 (N_7308,N_5399,N_4648);
and U7309 (N_7309,N_4801,N_5413);
nand U7310 (N_7310,N_4969,N_5045);
and U7311 (N_7311,N_5970,N_4504);
or U7312 (N_7312,N_5679,N_5867);
and U7313 (N_7313,N_5997,N_5470);
nor U7314 (N_7314,N_5652,N_5233);
or U7315 (N_7315,N_4717,N_5753);
nand U7316 (N_7316,N_4609,N_5901);
nand U7317 (N_7317,N_5677,N_4642);
and U7318 (N_7318,N_5862,N_4612);
nor U7319 (N_7319,N_4690,N_5559);
or U7320 (N_7320,N_4508,N_4940);
nand U7321 (N_7321,N_5298,N_5761);
nor U7322 (N_7322,N_5855,N_5081);
nand U7323 (N_7323,N_5953,N_5191);
and U7324 (N_7324,N_5251,N_5936);
or U7325 (N_7325,N_4729,N_5788);
or U7326 (N_7326,N_5574,N_5615);
nand U7327 (N_7327,N_5785,N_5456);
nand U7328 (N_7328,N_4877,N_5864);
and U7329 (N_7329,N_5088,N_4687);
nand U7330 (N_7330,N_5405,N_5127);
or U7331 (N_7331,N_5983,N_4731);
nand U7332 (N_7332,N_4677,N_4585);
nand U7333 (N_7333,N_5670,N_5964);
and U7334 (N_7334,N_5796,N_5704);
xnor U7335 (N_7335,N_5320,N_5400);
nor U7336 (N_7336,N_5910,N_5727);
or U7337 (N_7337,N_5232,N_5763);
nand U7338 (N_7338,N_5068,N_5526);
or U7339 (N_7339,N_5900,N_4879);
nor U7340 (N_7340,N_5559,N_5809);
or U7341 (N_7341,N_4917,N_5382);
nand U7342 (N_7342,N_5270,N_5928);
and U7343 (N_7343,N_4619,N_5414);
nor U7344 (N_7344,N_5069,N_5742);
or U7345 (N_7345,N_4686,N_5116);
nand U7346 (N_7346,N_5671,N_5283);
and U7347 (N_7347,N_4634,N_5489);
nor U7348 (N_7348,N_5093,N_5839);
nor U7349 (N_7349,N_4690,N_4651);
nor U7350 (N_7350,N_4774,N_5572);
or U7351 (N_7351,N_5958,N_4542);
nand U7352 (N_7352,N_5005,N_5429);
or U7353 (N_7353,N_4606,N_5248);
and U7354 (N_7354,N_5319,N_4768);
nor U7355 (N_7355,N_5804,N_5212);
or U7356 (N_7356,N_5763,N_4731);
nand U7357 (N_7357,N_4708,N_5470);
xor U7358 (N_7358,N_4799,N_4719);
and U7359 (N_7359,N_5701,N_4683);
and U7360 (N_7360,N_5436,N_4845);
or U7361 (N_7361,N_5447,N_5682);
or U7362 (N_7362,N_4525,N_5451);
and U7363 (N_7363,N_5220,N_5916);
and U7364 (N_7364,N_5695,N_5680);
xnor U7365 (N_7365,N_5530,N_5170);
or U7366 (N_7366,N_5522,N_5817);
or U7367 (N_7367,N_5877,N_4511);
nand U7368 (N_7368,N_4867,N_4734);
and U7369 (N_7369,N_5355,N_5772);
nor U7370 (N_7370,N_5258,N_4721);
nand U7371 (N_7371,N_4987,N_4784);
nor U7372 (N_7372,N_4868,N_5502);
nor U7373 (N_7373,N_5682,N_5657);
and U7374 (N_7374,N_5165,N_5578);
nor U7375 (N_7375,N_4525,N_5664);
xor U7376 (N_7376,N_4587,N_4819);
nand U7377 (N_7377,N_5456,N_4512);
and U7378 (N_7378,N_4613,N_4764);
or U7379 (N_7379,N_5072,N_5636);
xnor U7380 (N_7380,N_5038,N_5205);
xnor U7381 (N_7381,N_5375,N_5658);
or U7382 (N_7382,N_5553,N_4957);
nor U7383 (N_7383,N_4556,N_5359);
nand U7384 (N_7384,N_5700,N_5514);
nand U7385 (N_7385,N_5769,N_5873);
nor U7386 (N_7386,N_5045,N_4798);
nor U7387 (N_7387,N_4863,N_5943);
nand U7388 (N_7388,N_5730,N_5990);
and U7389 (N_7389,N_4759,N_4668);
xor U7390 (N_7390,N_4823,N_4576);
nand U7391 (N_7391,N_5426,N_5074);
or U7392 (N_7392,N_4797,N_5702);
nand U7393 (N_7393,N_4538,N_5807);
nand U7394 (N_7394,N_5902,N_5968);
or U7395 (N_7395,N_5972,N_4821);
nor U7396 (N_7396,N_5714,N_4918);
nand U7397 (N_7397,N_4623,N_5469);
nand U7398 (N_7398,N_5864,N_4803);
nor U7399 (N_7399,N_5457,N_5583);
nor U7400 (N_7400,N_5145,N_5660);
or U7401 (N_7401,N_5002,N_5230);
nand U7402 (N_7402,N_4753,N_5370);
nor U7403 (N_7403,N_5652,N_5441);
nor U7404 (N_7404,N_5857,N_5603);
nand U7405 (N_7405,N_5055,N_4749);
or U7406 (N_7406,N_4510,N_5087);
nand U7407 (N_7407,N_5023,N_4508);
xnor U7408 (N_7408,N_5187,N_4658);
or U7409 (N_7409,N_5283,N_4980);
or U7410 (N_7410,N_4652,N_5256);
nor U7411 (N_7411,N_5666,N_4668);
nand U7412 (N_7412,N_4761,N_5170);
or U7413 (N_7413,N_5743,N_4730);
and U7414 (N_7414,N_5694,N_5425);
and U7415 (N_7415,N_5050,N_5505);
xnor U7416 (N_7416,N_4817,N_5520);
nor U7417 (N_7417,N_4757,N_5955);
and U7418 (N_7418,N_5682,N_5692);
nor U7419 (N_7419,N_5388,N_5473);
or U7420 (N_7420,N_5166,N_4774);
and U7421 (N_7421,N_5890,N_5093);
nor U7422 (N_7422,N_4982,N_5282);
nand U7423 (N_7423,N_5488,N_5928);
or U7424 (N_7424,N_5296,N_4693);
and U7425 (N_7425,N_5524,N_5498);
nand U7426 (N_7426,N_5561,N_4844);
and U7427 (N_7427,N_5683,N_4937);
or U7428 (N_7428,N_4565,N_4574);
and U7429 (N_7429,N_5214,N_4596);
nand U7430 (N_7430,N_5257,N_5511);
and U7431 (N_7431,N_5590,N_5463);
nand U7432 (N_7432,N_5612,N_5619);
and U7433 (N_7433,N_5494,N_5059);
and U7434 (N_7434,N_5006,N_5426);
nand U7435 (N_7435,N_5053,N_5082);
or U7436 (N_7436,N_5411,N_5376);
nand U7437 (N_7437,N_5545,N_5131);
nand U7438 (N_7438,N_5765,N_5324);
or U7439 (N_7439,N_4524,N_4746);
and U7440 (N_7440,N_4737,N_4935);
nand U7441 (N_7441,N_5565,N_5964);
xor U7442 (N_7442,N_5710,N_5462);
nor U7443 (N_7443,N_5884,N_5498);
nand U7444 (N_7444,N_4975,N_5338);
nor U7445 (N_7445,N_4695,N_4532);
or U7446 (N_7446,N_5568,N_5941);
xor U7447 (N_7447,N_5049,N_5567);
and U7448 (N_7448,N_4805,N_5441);
nor U7449 (N_7449,N_5526,N_4835);
or U7450 (N_7450,N_4880,N_5053);
or U7451 (N_7451,N_5102,N_4670);
nor U7452 (N_7452,N_4590,N_5498);
nand U7453 (N_7453,N_4888,N_5267);
nand U7454 (N_7454,N_4990,N_5186);
and U7455 (N_7455,N_4890,N_4988);
or U7456 (N_7456,N_5678,N_5970);
nand U7457 (N_7457,N_5902,N_5457);
xnor U7458 (N_7458,N_5561,N_5864);
or U7459 (N_7459,N_5474,N_5742);
nand U7460 (N_7460,N_5463,N_5656);
or U7461 (N_7461,N_4650,N_5471);
or U7462 (N_7462,N_5555,N_5007);
nand U7463 (N_7463,N_5683,N_5012);
nand U7464 (N_7464,N_5718,N_5952);
nor U7465 (N_7465,N_5593,N_5470);
nand U7466 (N_7466,N_5030,N_4856);
or U7467 (N_7467,N_5506,N_4589);
nor U7468 (N_7468,N_5902,N_4922);
and U7469 (N_7469,N_5197,N_5631);
nand U7470 (N_7470,N_5498,N_5303);
nand U7471 (N_7471,N_5714,N_5645);
nand U7472 (N_7472,N_5614,N_5538);
nor U7473 (N_7473,N_5910,N_4714);
nand U7474 (N_7474,N_5514,N_4671);
nand U7475 (N_7475,N_4633,N_4823);
nand U7476 (N_7476,N_5544,N_4763);
nand U7477 (N_7477,N_4608,N_5048);
nor U7478 (N_7478,N_4943,N_4710);
or U7479 (N_7479,N_4760,N_5942);
nand U7480 (N_7480,N_5895,N_5055);
or U7481 (N_7481,N_4641,N_5300);
nor U7482 (N_7482,N_5848,N_5183);
or U7483 (N_7483,N_5863,N_5049);
and U7484 (N_7484,N_5662,N_4969);
or U7485 (N_7485,N_5899,N_5184);
or U7486 (N_7486,N_5144,N_5497);
nand U7487 (N_7487,N_5526,N_5713);
nand U7488 (N_7488,N_5556,N_5608);
or U7489 (N_7489,N_5704,N_5572);
nand U7490 (N_7490,N_5364,N_5610);
and U7491 (N_7491,N_5314,N_4649);
nor U7492 (N_7492,N_4833,N_5279);
nor U7493 (N_7493,N_5393,N_5588);
nand U7494 (N_7494,N_4630,N_5626);
and U7495 (N_7495,N_4732,N_5642);
nor U7496 (N_7496,N_5495,N_5941);
or U7497 (N_7497,N_4973,N_5164);
and U7498 (N_7498,N_5665,N_5646);
and U7499 (N_7499,N_5351,N_5470);
nand U7500 (N_7500,N_6476,N_6717);
and U7501 (N_7501,N_6895,N_6602);
or U7502 (N_7502,N_6204,N_7366);
or U7503 (N_7503,N_6990,N_6233);
nand U7504 (N_7504,N_6004,N_6086);
nor U7505 (N_7505,N_6122,N_7058);
nand U7506 (N_7506,N_7340,N_6860);
or U7507 (N_7507,N_7190,N_6845);
nor U7508 (N_7508,N_6520,N_6667);
nand U7509 (N_7509,N_6182,N_6152);
nand U7510 (N_7510,N_6832,N_6688);
nor U7511 (N_7511,N_6188,N_6931);
or U7512 (N_7512,N_6171,N_6342);
nor U7513 (N_7513,N_7361,N_6043);
xor U7514 (N_7514,N_7370,N_7164);
nor U7515 (N_7515,N_7010,N_6428);
nand U7516 (N_7516,N_6438,N_6799);
nand U7517 (N_7517,N_6450,N_6183);
nor U7518 (N_7518,N_6258,N_6032);
nand U7519 (N_7519,N_6570,N_6942);
and U7520 (N_7520,N_6973,N_6261);
nor U7521 (N_7521,N_6844,N_6246);
nand U7522 (N_7522,N_6376,N_6142);
nor U7523 (N_7523,N_6927,N_6083);
nor U7524 (N_7524,N_6680,N_6935);
and U7525 (N_7525,N_6684,N_7193);
nand U7526 (N_7526,N_6611,N_7292);
or U7527 (N_7527,N_6074,N_7279);
and U7528 (N_7528,N_6414,N_6196);
nor U7529 (N_7529,N_6389,N_6528);
nand U7530 (N_7530,N_6820,N_6898);
or U7531 (N_7531,N_7336,N_6180);
and U7532 (N_7532,N_6908,N_6195);
nand U7533 (N_7533,N_7048,N_6561);
and U7534 (N_7534,N_6480,N_7159);
nor U7535 (N_7535,N_6417,N_6581);
or U7536 (N_7536,N_7427,N_7020);
nand U7537 (N_7537,N_6771,N_6535);
nor U7538 (N_7538,N_6344,N_6569);
nand U7539 (N_7539,N_6185,N_7355);
and U7540 (N_7540,N_6802,N_7071);
or U7541 (N_7541,N_6787,N_6076);
nor U7542 (N_7542,N_7166,N_7109);
nand U7543 (N_7543,N_6698,N_6465);
nor U7544 (N_7544,N_6782,N_6282);
nand U7545 (N_7545,N_7022,N_7456);
nand U7546 (N_7546,N_6231,N_6404);
or U7547 (N_7547,N_6328,N_6783);
or U7548 (N_7548,N_6606,N_7354);
and U7549 (N_7549,N_6523,N_7154);
or U7550 (N_7550,N_7283,N_6037);
or U7551 (N_7551,N_6518,N_6347);
and U7552 (N_7552,N_6403,N_7247);
or U7553 (N_7553,N_6592,N_7063);
and U7554 (N_7554,N_7088,N_6909);
and U7555 (N_7555,N_6538,N_7296);
nor U7556 (N_7556,N_6358,N_6884);
nor U7557 (N_7557,N_6988,N_6761);
nand U7558 (N_7558,N_6863,N_6541);
or U7559 (N_7559,N_7358,N_6811);
xor U7560 (N_7560,N_6686,N_6390);
and U7561 (N_7561,N_7294,N_6841);
nor U7562 (N_7562,N_6387,N_6406);
nand U7563 (N_7563,N_6490,N_6558);
nor U7564 (N_7564,N_6409,N_7242);
or U7565 (N_7565,N_6093,N_6367);
nor U7566 (N_7566,N_6290,N_6621);
or U7567 (N_7567,N_7441,N_6678);
nor U7568 (N_7568,N_6851,N_6760);
nor U7569 (N_7569,N_7330,N_6842);
and U7570 (N_7570,N_7188,N_6830);
nor U7571 (N_7571,N_6508,N_6716);
or U7572 (N_7572,N_6587,N_7332);
nor U7573 (N_7573,N_7449,N_6469);
nor U7574 (N_7574,N_6970,N_7203);
xnor U7575 (N_7575,N_7012,N_6694);
nand U7576 (N_7576,N_6110,N_7468);
and U7577 (N_7577,N_6997,N_6619);
nor U7578 (N_7578,N_6781,N_7389);
or U7579 (N_7579,N_7240,N_7001);
and U7580 (N_7580,N_7393,N_7318);
or U7581 (N_7581,N_6399,N_7017);
nand U7582 (N_7582,N_6666,N_6738);
and U7583 (N_7583,N_7249,N_6145);
nor U7584 (N_7584,N_7440,N_6922);
or U7585 (N_7585,N_6325,N_7356);
nand U7586 (N_7586,N_6013,N_7281);
nor U7587 (N_7587,N_7268,N_7400);
and U7588 (N_7588,N_6912,N_6579);
nand U7589 (N_7589,N_7375,N_7421);
nor U7590 (N_7590,N_7253,N_6094);
xnor U7591 (N_7591,N_7107,N_7021);
or U7592 (N_7592,N_6641,N_7298);
and U7593 (N_7593,N_7181,N_7313);
and U7594 (N_7594,N_6045,N_7350);
nand U7595 (N_7595,N_7404,N_6607);
or U7596 (N_7596,N_6192,N_7192);
nand U7597 (N_7597,N_7187,N_6048);
or U7598 (N_7598,N_6910,N_6430);
nor U7599 (N_7599,N_7202,N_6179);
and U7600 (N_7600,N_6939,N_6797);
and U7601 (N_7601,N_6646,N_6457);
and U7602 (N_7602,N_6664,N_6493);
or U7603 (N_7603,N_7429,N_6130);
or U7604 (N_7604,N_7300,N_6373);
and U7605 (N_7605,N_6872,N_6352);
nor U7606 (N_7606,N_6253,N_7446);
or U7607 (N_7607,N_6107,N_6022);
or U7608 (N_7608,N_6451,N_6634);
and U7609 (N_7609,N_6527,N_7078);
xor U7610 (N_7610,N_6434,N_6727);
and U7611 (N_7611,N_6156,N_6251);
nand U7612 (N_7612,N_6768,N_7291);
and U7613 (N_7613,N_6335,N_7027);
nor U7614 (N_7614,N_6598,N_7487);
nand U7615 (N_7615,N_6303,N_7386);
nand U7616 (N_7616,N_6464,N_7056);
and U7617 (N_7617,N_7096,N_6275);
or U7618 (N_7618,N_6386,N_6645);
nand U7619 (N_7619,N_6916,N_6766);
and U7620 (N_7620,N_6172,N_7475);
nand U7621 (N_7621,N_7444,N_6098);
nor U7622 (N_7622,N_6502,N_6315);
and U7623 (N_7623,N_6370,N_6856);
nor U7624 (N_7624,N_7224,N_6175);
nand U7625 (N_7625,N_7038,N_6263);
nand U7626 (N_7626,N_6147,N_7273);
nand U7627 (N_7627,N_7485,N_7138);
nand U7628 (N_7628,N_6273,N_7211);
and U7629 (N_7629,N_7099,N_6416);
nor U7630 (N_7630,N_6374,N_7070);
or U7631 (N_7631,N_6255,N_6546);
and U7632 (N_7632,N_6683,N_6774);
nand U7633 (N_7633,N_7033,N_6550);
nor U7634 (N_7634,N_6560,N_7156);
nor U7635 (N_7635,N_6993,N_6720);
nor U7636 (N_7636,N_6571,N_6998);
or U7637 (N_7637,N_6333,N_6862);
xnor U7638 (N_7638,N_6801,N_6216);
nand U7639 (N_7639,N_7112,N_6050);
nand U7640 (N_7640,N_7225,N_7266);
nand U7641 (N_7641,N_7359,N_6087);
nand U7642 (N_7642,N_7477,N_6620);
nor U7643 (N_7643,N_6792,N_7293);
or U7644 (N_7644,N_6260,N_6522);
nand U7645 (N_7645,N_6248,N_6690);
nand U7646 (N_7646,N_7116,N_6169);
or U7647 (N_7647,N_7371,N_6769);
nand U7648 (N_7648,N_6135,N_6882);
nand U7649 (N_7649,N_6963,N_7275);
nand U7650 (N_7650,N_6512,N_7260);
and U7651 (N_7651,N_6208,N_6285);
xnor U7652 (N_7652,N_6366,N_6869);
or U7653 (N_7653,N_6498,N_7245);
or U7654 (N_7654,N_7310,N_7448);
nor U7655 (N_7655,N_7008,N_6915);
nor U7656 (N_7656,N_6548,N_6578);
nor U7657 (N_7657,N_6547,N_6937);
nand U7658 (N_7658,N_6456,N_7437);
and U7659 (N_7659,N_6016,N_7305);
or U7660 (N_7660,N_6066,N_6831);
and U7661 (N_7661,N_6757,N_6239);
and U7662 (N_7662,N_7277,N_7082);
or U7663 (N_7663,N_6405,N_7458);
nor U7664 (N_7664,N_6818,N_6987);
nor U7665 (N_7665,N_6529,N_6848);
nand U7666 (N_7666,N_6711,N_6858);
and U7667 (N_7667,N_6170,N_6116);
and U7668 (N_7668,N_7496,N_7480);
nor U7669 (N_7669,N_7050,N_6868);
or U7670 (N_7670,N_7396,N_7373);
nor U7671 (N_7671,N_7029,N_6123);
nand U7672 (N_7672,N_7307,N_6299);
nand U7673 (N_7673,N_7433,N_6778);
and U7674 (N_7674,N_6254,N_7288);
or U7675 (N_7675,N_7367,N_6633);
and U7676 (N_7676,N_6266,N_6015);
xnor U7677 (N_7677,N_6815,N_6234);
and U7678 (N_7678,N_6616,N_7465);
nand U7679 (N_7679,N_6064,N_6637);
or U7680 (N_7680,N_7199,N_6724);
and U7681 (N_7681,N_7047,N_6789);
and U7682 (N_7682,N_6980,N_6207);
nor U7683 (N_7683,N_7093,N_6256);
and U7684 (N_7684,N_6610,N_7484);
nand U7685 (N_7685,N_7152,N_7334);
or U7686 (N_7686,N_6454,N_6336);
nor U7687 (N_7687,N_7113,N_6886);
or U7688 (N_7688,N_7117,N_6929);
nor U7689 (N_7689,N_7322,N_7114);
and U7690 (N_7690,N_7476,N_6654);
nor U7691 (N_7691,N_6038,N_6348);
nor U7692 (N_7692,N_6455,N_7325);
nand U7693 (N_7693,N_6120,N_6201);
nand U7694 (N_7694,N_6971,N_6906);
and U7695 (N_7695,N_7143,N_7349);
nor U7696 (N_7696,N_6785,N_6095);
nand U7697 (N_7697,N_6096,N_7431);
and U7698 (N_7698,N_6959,N_6599);
nand U7699 (N_7699,N_7258,N_6642);
nand U7700 (N_7700,N_6375,N_7009);
or U7701 (N_7701,N_6613,N_6264);
or U7702 (N_7702,N_7119,N_6458);
or U7703 (N_7703,N_6805,N_7309);
nand U7704 (N_7704,N_7103,N_7158);
nand U7705 (N_7705,N_6850,N_6791);
or U7706 (N_7706,N_6262,N_7360);
xnor U7707 (N_7707,N_6867,N_7388);
nand U7708 (N_7708,N_6776,N_6446);
nand U7709 (N_7709,N_6426,N_6310);
and U7710 (N_7710,N_6632,N_7072);
nand U7711 (N_7711,N_7092,N_6187);
or U7712 (N_7712,N_7347,N_6154);
nand U7713 (N_7713,N_6878,N_6121);
or U7714 (N_7714,N_7066,N_7422);
nor U7715 (N_7715,N_7214,N_6810);
or U7716 (N_7716,N_6693,N_7241);
and U7717 (N_7717,N_6473,N_7206);
nor U7718 (N_7718,N_6343,N_6111);
nand U7719 (N_7719,N_6272,N_6584);
nor U7720 (N_7720,N_7416,N_6492);
and U7721 (N_7721,N_7074,N_6274);
and U7722 (N_7722,N_7323,N_6025);
and U7723 (N_7723,N_6617,N_6806);
nand U7724 (N_7724,N_7368,N_7230);
nand U7725 (N_7725,N_7172,N_7381);
or U7726 (N_7726,N_7348,N_7052);
xor U7727 (N_7727,N_7491,N_6871);
nor U7728 (N_7728,N_7398,N_6758);
nand U7729 (N_7729,N_6813,N_6018);
or U7730 (N_7730,N_7329,N_6651);
nand U7731 (N_7731,N_6166,N_7216);
and U7732 (N_7732,N_7053,N_7221);
nand U7733 (N_7733,N_7423,N_7196);
nand U7734 (N_7734,N_6674,N_6008);
and U7735 (N_7735,N_6790,N_6072);
and U7736 (N_7736,N_6091,N_7357);
nor U7737 (N_7737,N_7418,N_6224);
or U7738 (N_7738,N_7057,N_7326);
nand U7739 (N_7739,N_6807,N_6999);
nand U7740 (N_7740,N_7068,N_6977);
and U7741 (N_7741,N_7083,N_7262);
nor U7742 (N_7742,N_7462,N_6662);
and U7743 (N_7743,N_6301,N_7351);
nand U7744 (N_7744,N_6919,N_6835);
nand U7745 (N_7745,N_6148,N_6322);
nor U7746 (N_7746,N_7271,N_7383);
nor U7747 (N_7747,N_6955,N_6829);
and U7748 (N_7748,N_7498,N_7343);
or U7749 (N_7749,N_6411,N_7013);
or U7750 (N_7750,N_7365,N_7101);
nand U7751 (N_7751,N_6483,N_7165);
or U7752 (N_7752,N_7231,N_6005);
or U7753 (N_7753,N_6568,N_6106);
or U7754 (N_7754,N_6612,N_6267);
nor U7755 (N_7755,N_6975,N_6276);
nand U7756 (N_7756,N_7451,N_7474);
or U7757 (N_7757,N_7136,N_6109);
nand U7758 (N_7758,N_6055,N_7233);
nand U7759 (N_7759,N_6989,N_6311);
nor U7760 (N_7760,N_6509,N_7081);
nand U7761 (N_7761,N_6767,N_7454);
or U7762 (N_7762,N_6640,N_6903);
and U7763 (N_7763,N_7380,N_7178);
nand U7764 (N_7764,N_6961,N_7424);
or U7765 (N_7765,N_6719,N_7183);
and U7766 (N_7766,N_6992,N_6294);
or U7767 (N_7767,N_7302,N_6515);
nand U7768 (N_7768,N_6199,N_7274);
xor U7769 (N_7769,N_6097,N_7376);
or U7770 (N_7770,N_7150,N_6883);
or U7771 (N_7771,N_6444,N_7362);
nor U7772 (N_7772,N_6108,N_6158);
nand U7773 (N_7773,N_6764,N_6614);
and U7774 (N_7774,N_6452,N_6046);
or U7775 (N_7775,N_6215,N_6735);
nor U7776 (N_7776,N_6163,N_7130);
or U7777 (N_7777,N_7142,N_6533);
or U7778 (N_7778,N_6174,N_7110);
nor U7779 (N_7779,N_6388,N_7133);
nand U7780 (N_7780,N_6567,N_7000);
nor U7781 (N_7781,N_7229,N_7426);
or U7782 (N_7782,N_6269,N_6542);
nand U7783 (N_7783,N_6855,N_6349);
nor U7784 (N_7784,N_6329,N_7301);
or U7785 (N_7785,N_6630,N_6427);
or U7786 (N_7786,N_6917,N_7067);
nand U7787 (N_7787,N_7025,N_7397);
and U7788 (N_7788,N_6326,N_7189);
or U7789 (N_7789,N_7186,N_6756);
and U7790 (N_7790,N_6398,N_6749);
and U7791 (N_7791,N_6759,N_7147);
and U7792 (N_7792,N_6713,N_7146);
and U7793 (N_7793,N_6880,N_6876);
nor U7794 (N_7794,N_6583,N_6226);
nor U7795 (N_7795,N_6437,N_6419);
nand U7796 (N_7796,N_6624,N_6345);
nor U7797 (N_7797,N_6877,N_7314);
nor U7798 (N_7798,N_6151,N_6468);
nand U7799 (N_7799,N_7238,N_6237);
nand U7800 (N_7800,N_6115,N_6031);
nand U7801 (N_7801,N_6138,N_7153);
or U7802 (N_7802,N_6676,N_6176);
nand U7803 (N_7803,N_7410,N_7471);
or U7804 (N_7804,N_6751,N_7256);
nor U7805 (N_7805,N_6968,N_6944);
or U7806 (N_7806,N_7155,N_6816);
or U7807 (N_7807,N_6647,N_6178);
nor U7808 (N_7808,N_6306,N_7200);
or U7809 (N_7809,N_6576,N_6320);
nand U7810 (N_7810,N_6291,N_6259);
or U7811 (N_7811,N_7261,N_7129);
nor U7812 (N_7812,N_6780,N_6773);
and U7813 (N_7813,N_6270,N_7195);
nand U7814 (N_7814,N_6295,N_7406);
or U7815 (N_7815,N_7399,N_6209);
or U7816 (N_7816,N_6679,N_6580);
and U7817 (N_7817,N_7269,N_6162);
nand U7818 (N_7818,N_6383,N_6639);
nor U7819 (N_7819,N_6257,N_7126);
nand U7820 (N_7820,N_7272,N_6822);
xor U7821 (N_7821,N_7168,N_6695);
and U7822 (N_7822,N_6460,N_6415);
nor U7823 (N_7823,N_6012,N_7045);
and U7824 (N_7824,N_6706,N_7377);
nor U7825 (N_7825,N_7144,N_6672);
and U7826 (N_7826,N_6649,N_7091);
nor U7827 (N_7827,N_7387,N_7478);
and U7828 (N_7828,N_6365,N_7205);
or U7829 (N_7829,N_6021,N_7341);
or U7830 (N_7830,N_6881,N_7044);
and U7831 (N_7831,N_6181,N_7308);
nor U7832 (N_7832,N_6134,N_7075);
nor U7833 (N_7833,N_6566,N_6228);
or U7834 (N_7834,N_7284,N_7213);
and U7835 (N_7835,N_7479,N_7122);
and U7836 (N_7836,N_6265,N_6689);
and U7837 (N_7837,N_6305,N_7411);
nor U7838 (N_7838,N_7095,N_7304);
nor U7839 (N_7839,N_6938,N_6413);
xor U7840 (N_7840,N_7134,N_6324);
and U7841 (N_7841,N_6041,N_6957);
nand U7842 (N_7842,N_6605,N_6934);
nor U7843 (N_7843,N_7461,N_6748);
or U7844 (N_7844,N_6284,N_6962);
nor U7845 (N_7845,N_6371,N_6047);
and U7846 (N_7846,N_7264,N_6788);
or U7847 (N_7847,N_7467,N_7353);
nor U7848 (N_7848,N_6594,N_7450);
or U7849 (N_7849,N_7391,N_6839);
or U7850 (N_7850,N_6960,N_6067);
or U7851 (N_7851,N_6236,N_7392);
nor U7852 (N_7852,N_7255,N_7335);
nand U7853 (N_7853,N_6506,N_7097);
nor U7854 (N_7854,N_6117,N_7016);
or U7855 (N_7855,N_6754,N_6368);
nor U7856 (N_7856,N_6623,N_6472);
nand U7857 (N_7857,N_6369,N_6551);
nand U7858 (N_7858,N_6191,N_6139);
or U7859 (N_7859,N_6817,N_6755);
nand U7860 (N_7860,N_7132,N_6673);
nor U7861 (N_7861,N_7111,N_6625);
and U7862 (N_7862,N_6396,N_6668);
or U7863 (N_7863,N_6608,N_7311);
nand U7864 (N_7864,N_7106,N_7197);
and U7865 (N_7865,N_6481,N_6384);
or U7866 (N_7866,N_7338,N_7179);
xor U7867 (N_7867,N_6786,N_6534);
nor U7868 (N_7868,N_6340,N_6924);
or U7869 (N_7869,N_6077,N_6459);
nand U7870 (N_7870,N_7403,N_6491);
and U7871 (N_7871,N_6597,N_7289);
and U7872 (N_7872,N_6995,N_6210);
or U7873 (N_7873,N_7402,N_6586);
nand U7874 (N_7874,N_6526,N_6190);
nor U7875 (N_7875,N_6770,N_6219);
nand U7876 (N_7876,N_7163,N_6699);
and U7877 (N_7877,N_7087,N_7115);
nand U7878 (N_7878,N_7015,N_6467);
and U7879 (N_7879,N_6033,N_7472);
nand U7880 (N_7880,N_6669,N_7379);
nor U7881 (N_7881,N_7018,N_7243);
or U7882 (N_7882,N_7488,N_6794);
or U7883 (N_7883,N_6966,N_7145);
and U7884 (N_7884,N_6080,N_7135);
and U7885 (N_7885,N_7085,N_7297);
nand U7886 (N_7886,N_6814,N_7079);
or U7887 (N_7887,N_7259,N_6238);
nand U7888 (N_7888,N_6800,N_6068);
and U7889 (N_7889,N_7464,N_6144);
and U7890 (N_7890,N_6317,N_6900);
nand U7891 (N_7891,N_6061,N_6391);
nor U7892 (N_7892,N_7108,N_7290);
nand U7893 (N_7893,N_6394,N_6557);
nor U7894 (N_7894,N_6671,N_6300);
and U7895 (N_7895,N_6380,N_6562);
nor U7896 (N_7896,N_6921,N_7263);
and U7897 (N_7897,N_6826,N_6332);
and U7898 (N_7898,N_6381,N_6421);
nand U7899 (N_7899,N_7276,N_6081);
nand U7900 (N_7900,N_6575,N_7445);
and U7901 (N_7901,N_7042,N_6979);
nand U7902 (N_7902,N_6408,N_7002);
and U7903 (N_7903,N_6359,N_6743);
and U7904 (N_7904,N_6946,N_7251);
nor U7905 (N_7905,N_6379,N_6752);
nand U7906 (N_7906,N_6153,N_7140);
or U7907 (N_7907,N_7385,N_6304);
or U7908 (N_7908,N_7473,N_6126);
and U7909 (N_7909,N_6189,N_6334);
nand U7910 (N_7910,N_6420,N_6000);
nor U7911 (N_7911,N_6429,N_7191);
and U7912 (N_7912,N_6319,N_7287);
nand U7913 (N_7913,N_6745,N_6875);
xnor U7914 (N_7914,N_6737,N_6951);
nand U7915 (N_7915,N_6099,N_7234);
and U7916 (N_7916,N_6517,N_7223);
nor U7917 (N_7917,N_6911,N_6039);
nor U7918 (N_7918,N_6722,N_6137);
or U7919 (N_7919,N_7345,N_7415);
or U7920 (N_7920,N_6351,N_7267);
nand U7921 (N_7921,N_6035,N_6354);
xor U7922 (N_7922,N_6707,N_6531);
nor U7923 (N_7923,N_6014,N_6511);
nor U7924 (N_7924,N_6034,N_7428);
and U7925 (N_7925,N_6206,N_7011);
and U7926 (N_7926,N_6119,N_6161);
nand U7927 (N_7927,N_6339,N_6574);
nor U7928 (N_7928,N_6297,N_7442);
and U7929 (N_7929,N_6622,N_6364);
nand U7930 (N_7930,N_6073,N_6484);
and U7931 (N_7931,N_6941,N_6833);
and U7932 (N_7932,N_6244,N_6721);
nor U7933 (N_7933,N_6360,N_7139);
nand U7934 (N_7934,N_7104,N_6225);
or U7935 (N_7935,N_6958,N_6313);
nand U7936 (N_7936,N_7059,N_6796);
nor U7937 (N_7937,N_6412,N_6603);
or U7938 (N_7938,N_7306,N_6658);
nand U7939 (N_7939,N_7346,N_6540);
nor U7940 (N_7940,N_7469,N_6292);
nor U7941 (N_7941,N_6353,N_7080);
nor U7942 (N_7942,N_6078,N_7014);
or U7943 (N_7943,N_6505,N_7043);
and U7944 (N_7944,N_6357,N_7098);
nand U7945 (N_7945,N_7089,N_6981);
nand U7946 (N_7946,N_6435,N_6131);
nor U7947 (N_7947,N_7204,N_6956);
or U7948 (N_7948,N_7303,N_6213);
or U7949 (N_7949,N_6400,N_6840);
nor U7950 (N_7950,N_6590,N_7118);
or U7951 (N_7951,N_6657,N_6710);
xnor U7952 (N_7952,N_6991,N_6023);
nor U7953 (N_7953,N_6986,N_6585);
nand U7954 (N_7954,N_6482,N_7065);
and U7955 (N_7955,N_7169,N_7160);
or U7956 (N_7956,N_7086,N_6949);
nor U7957 (N_7957,N_6217,N_6950);
or U7958 (N_7958,N_7174,N_6936);
nor U7959 (N_7959,N_7395,N_6277);
nand U7960 (N_7960,N_7436,N_6132);
and U7961 (N_7961,N_7034,N_6221);
and U7962 (N_7962,N_6020,N_6879);
xor U7963 (N_7963,N_6894,N_7209);
nor U7964 (N_7964,N_6947,N_6202);
nand U7965 (N_7965,N_7201,N_7212);
or U7966 (N_7966,N_7320,N_6984);
or U7967 (N_7967,N_6513,N_6499);
and U7968 (N_7968,N_7319,N_7447);
xnor U7969 (N_7969,N_6113,N_7407);
and U7970 (N_7970,N_7124,N_7270);
or U7971 (N_7971,N_6925,N_6160);
or U7972 (N_7972,N_6448,N_7019);
and U7973 (N_7973,N_6441,N_7299);
nor U7974 (N_7974,N_6982,N_6905);
nor U7975 (N_7975,N_7278,N_6762);
or U7976 (N_7976,N_6027,N_7344);
or U7977 (N_7977,N_7049,N_6024);
nand U7978 (N_7978,N_6082,N_6065);
nand U7979 (N_7979,N_6338,N_6363);
or U7980 (N_7980,N_6280,N_6744);
nor U7981 (N_7981,N_6197,N_7054);
or U7982 (N_7982,N_6205,N_6084);
xor U7983 (N_7983,N_7497,N_7384);
or U7984 (N_7984,N_7250,N_6864);
nor U7985 (N_7985,N_6596,N_7459);
nor U7986 (N_7986,N_6974,N_6337);
or U7987 (N_7987,N_6165,N_6193);
and U7988 (N_7988,N_6825,N_6545);
xnor U7989 (N_7989,N_6914,N_6051);
or U7990 (N_7990,N_6173,N_6410);
nor U7991 (N_7991,N_6677,N_6635);
xnor U7992 (N_7992,N_6857,N_7162);
and U7993 (N_7993,N_6659,N_6595);
or U7994 (N_7994,N_6742,N_7420);
nor U7995 (N_7995,N_7128,N_7363);
and U7996 (N_7996,N_6069,N_7470);
nor U7997 (N_7997,N_6443,N_6049);
nand U7998 (N_7998,N_6740,N_6874);
or U7999 (N_7999,N_7149,N_6985);
or U8000 (N_8000,N_6652,N_6889);
nor U8001 (N_8001,N_6837,N_6885);
or U8002 (N_8002,N_7032,N_7131);
xnor U8003 (N_8003,N_6725,N_7265);
nand U8004 (N_8004,N_6397,N_6356);
nor U8005 (N_8005,N_7492,N_6488);
or U8006 (N_8006,N_6953,N_7024);
nand U8007 (N_8007,N_7102,N_6440);
nor U8008 (N_8008,N_6103,N_7226);
or U8009 (N_8009,N_6819,N_7452);
nand U8010 (N_8010,N_6824,N_6891);
nand U8011 (N_8011,N_6661,N_6062);
and U8012 (N_8012,N_7499,N_6186);
nor U8013 (N_8013,N_6660,N_6923);
and U8014 (N_8014,N_6009,N_6793);
nor U8015 (N_8015,N_6203,N_6888);
nand U8016 (N_8016,N_7208,N_6006);
or U8017 (N_8017,N_6362,N_6804);
nor U8018 (N_8018,N_6167,N_6507);
or U8019 (N_8019,N_6474,N_6395);
xor U8020 (N_8020,N_6920,N_6736);
and U8021 (N_8021,N_7175,N_7490);
and U8022 (N_8022,N_7409,N_6983);
xnor U8023 (N_8023,N_7023,N_7295);
nor U8024 (N_8024,N_6530,N_7486);
nand U8025 (N_8025,N_6779,N_7222);
and U8026 (N_8026,N_6112,N_6795);
or U8027 (N_8027,N_6141,N_7041);
and U8028 (N_8028,N_6715,N_6164);
or U8029 (N_8029,N_7430,N_6432);
and U8030 (N_8030,N_7046,N_7286);
and U8031 (N_8031,N_6127,N_6836);
or U8032 (N_8032,N_6964,N_6220);
nor U8033 (N_8033,N_7061,N_6198);
nor U8034 (N_8034,N_6893,N_6449);
or U8035 (N_8035,N_6784,N_6537);
nand U8036 (N_8036,N_6510,N_6593);
or U8037 (N_8037,N_6685,N_7494);
nand U8038 (N_8038,N_6495,N_6128);
or U8039 (N_8039,N_6289,N_7039);
nor U8040 (N_8040,N_6439,N_6808);
or U8041 (N_8041,N_7090,N_6442);
nand U8042 (N_8042,N_6615,N_6242);
and U8043 (N_8043,N_6556,N_7460);
and U8044 (N_8044,N_6314,N_6071);
or U8045 (N_8045,N_6462,N_6114);
nand U8046 (N_8046,N_6591,N_6393);
or U8047 (N_8047,N_7177,N_6431);
nand U8048 (N_8048,N_6572,N_6003);
nor U8049 (N_8049,N_6503,N_6070);
or U8050 (N_8050,N_6007,N_6129);
nand U8051 (N_8051,N_6775,N_7414);
or U8052 (N_8052,N_6681,N_7328);
nand U8053 (N_8053,N_6227,N_6682);
nor U8054 (N_8054,N_6296,N_6054);
or U8055 (N_8055,N_7121,N_6089);
and U8056 (N_8056,N_7084,N_7248);
or U8057 (N_8057,N_6124,N_6854);
nand U8058 (N_8058,N_6828,N_6627);
and U8059 (N_8059,N_6247,N_6053);
and U8060 (N_8060,N_6327,N_6870);
or U8061 (N_8061,N_6288,N_6954);
nor U8062 (N_8062,N_7419,N_7035);
nor U8063 (N_8063,N_6536,N_6629);
nor U8064 (N_8064,N_6240,N_6026);
or U8065 (N_8065,N_6655,N_7185);
nor U8066 (N_8066,N_6445,N_6286);
nand U8067 (N_8067,N_6730,N_6063);
or U8068 (N_8068,N_6543,N_6524);
and U8069 (N_8069,N_7382,N_6928);
nor U8070 (N_8070,N_6407,N_6090);
and U8071 (N_8071,N_6803,N_7137);
and U8072 (N_8072,N_7228,N_7062);
and U8073 (N_8073,N_6618,N_7466);
nor U8074 (N_8074,N_6709,N_6899);
nand U8075 (N_8075,N_7434,N_6478);
and U8076 (N_8076,N_6118,N_7167);
nand U8077 (N_8077,N_6029,N_6425);
nor U8078 (N_8078,N_6890,N_6700);
and U8079 (N_8079,N_7438,N_6241);
and U8080 (N_8080,N_6401,N_7030);
nor U8081 (N_8081,N_6577,N_7184);
or U8082 (N_8082,N_6056,N_6346);
or U8083 (N_8083,N_6168,N_7483);
nor U8084 (N_8084,N_6687,N_6157);
and U8085 (N_8085,N_7040,N_6133);
and U8086 (N_8086,N_7182,N_6330);
nand U8087 (N_8087,N_6691,N_7312);
nand U8088 (N_8088,N_7401,N_6044);
nand U8089 (N_8089,N_6553,N_7324);
and U8090 (N_8090,N_6750,N_6692);
nor U8091 (N_8091,N_6812,N_7246);
or U8092 (N_8092,N_6943,N_6422);
nor U8093 (N_8093,N_6555,N_6485);
nor U8094 (N_8094,N_6865,N_6626);
and U8095 (N_8095,N_7236,N_6212);
nand U8096 (N_8096,N_6670,N_6732);
or U8097 (N_8097,N_6731,N_6487);
nor U8098 (N_8098,N_6609,N_6554);
nand U8099 (N_8099,N_6901,N_6463);
and U8100 (N_8100,N_6470,N_6827);
nor U8101 (N_8101,N_6972,N_6656);
nand U8102 (N_8102,N_7482,N_6777);
and U8103 (N_8103,N_6696,N_6847);
and U8104 (N_8104,N_6424,N_6036);
and U8105 (N_8105,N_6475,N_6861);
and U8106 (N_8106,N_6323,N_6809);
or U8107 (N_8107,N_7005,N_6521);
or U8108 (N_8108,N_7364,N_7235);
nand U8109 (N_8109,N_6466,N_6940);
or U8110 (N_8110,N_6897,N_6321);
and U8111 (N_8111,N_7028,N_7413);
nor U8112 (N_8112,N_6092,N_6516);
or U8113 (N_8113,N_6628,N_6926);
nor U8114 (N_8114,N_6281,N_6497);
nor U8115 (N_8115,N_7315,N_6309);
and U8116 (N_8116,N_7170,N_6638);
or U8117 (N_8117,N_7232,N_7031);
nand U8118 (N_8118,N_6159,N_7125);
nor U8119 (N_8119,N_7003,N_6896);
and U8120 (N_8120,N_6232,N_6125);
nand U8121 (N_8121,N_6268,N_6222);
or U8122 (N_8122,N_6525,N_6849);
nand U8123 (N_8123,N_6714,N_6494);
and U8124 (N_8124,N_7105,N_6866);
nand U8125 (N_8125,N_6734,N_7151);
or U8126 (N_8126,N_7237,N_6675);
and U8127 (N_8127,N_6479,N_6563);
and U8128 (N_8128,N_6361,N_6763);
or U8129 (N_8129,N_7219,N_6589);
nor U8130 (N_8130,N_6418,N_7317);
and U8131 (N_8131,N_7453,N_6377);
nor U8132 (N_8132,N_7408,N_6823);
and U8133 (N_8133,N_7443,N_7161);
nor U8134 (N_8134,N_6042,N_7390);
and U8135 (N_8135,N_6100,N_6705);
or U8136 (N_8136,N_6136,N_6316);
nor U8137 (N_8137,N_6648,N_6283);
and U8138 (N_8138,N_6994,N_6500);
and U8139 (N_8139,N_7210,N_6703);
nor U8140 (N_8140,N_6287,N_6948);
nand U8141 (N_8141,N_6532,N_7352);
nor U8142 (N_8142,N_6298,N_6741);
or U8143 (N_8143,N_6278,N_6057);
and U8144 (N_8144,N_7180,N_7285);
nor U8145 (N_8145,N_6105,N_6052);
and U8146 (N_8146,N_6718,N_6088);
or U8147 (N_8147,N_6002,N_6355);
and U8148 (N_8148,N_6271,N_6588);
nand U8149 (N_8149,N_6501,N_6230);
or U8150 (N_8150,N_7171,N_7457);
and U8151 (N_8151,N_6728,N_6017);
nand U8152 (N_8152,N_6821,N_7055);
and U8153 (N_8153,N_6650,N_7489);
and U8154 (N_8154,N_6486,N_7417);
nand U8155 (N_8155,N_6601,N_7069);
or U8156 (N_8156,N_7077,N_6907);
and U8157 (N_8157,N_6746,N_6218);
or U8158 (N_8158,N_7076,N_7006);
nor U8159 (N_8159,N_6200,N_6447);
and U8160 (N_8160,N_7120,N_7339);
and U8161 (N_8161,N_6544,N_6040);
or U8162 (N_8162,N_6211,N_6382);
nand U8163 (N_8163,N_7157,N_6902);
or U8164 (N_8164,N_6489,N_6636);
nor U8165 (N_8165,N_6372,N_7331);
or U8166 (N_8166,N_7141,N_6729);
or U8167 (N_8167,N_6058,N_6101);
nor U8168 (N_8168,N_7051,N_7337);
nor U8169 (N_8169,N_6631,N_7060);
or U8170 (N_8170,N_6798,N_6933);
and U8171 (N_8171,N_6559,N_6697);
and U8172 (N_8172,N_6194,N_6385);
or U8173 (N_8173,N_6564,N_6723);
and U8174 (N_8174,N_6834,N_6229);
nand U8175 (N_8175,N_7333,N_6461);
nand U8176 (N_8176,N_7254,N_6708);
nand U8177 (N_8177,N_7094,N_7342);
and U8178 (N_8178,N_6028,N_6030);
nor U8179 (N_8179,N_6085,N_6712);
and U8180 (N_8180,N_6843,N_7455);
nor U8181 (N_8181,N_6307,N_7217);
nor U8182 (N_8182,N_6918,N_7207);
nor U8183 (N_8183,N_7004,N_6838);
nand U8184 (N_8184,N_7037,N_6665);
or U8185 (N_8185,N_7495,N_6539);
and U8186 (N_8186,N_6245,N_6726);
nand U8187 (N_8187,N_7227,N_6945);
and U8188 (N_8188,N_6150,N_6249);
nor U8189 (N_8189,N_6976,N_6552);
nor U8190 (N_8190,N_6653,N_6140);
or U8191 (N_8191,N_6996,N_6739);
or U8192 (N_8192,N_6293,N_7215);
nand U8193 (N_8193,N_7252,N_7394);
nor U8194 (N_8194,N_6582,N_7244);
nor U8195 (N_8195,N_6514,N_6573);
and U8196 (N_8196,N_6302,N_7220);
nor U8197 (N_8197,N_7481,N_6969);
or U8198 (N_8198,N_6279,N_7073);
nor U8199 (N_8199,N_6423,N_7036);
nor U8200 (N_8200,N_6146,N_6978);
nand U8201 (N_8201,N_6177,N_6102);
xnor U8202 (N_8202,N_6565,N_6308);
nor U8203 (N_8203,N_6549,N_7493);
nor U8204 (N_8204,N_6350,N_7173);
and U8205 (N_8205,N_6859,N_6019);
nor U8206 (N_8206,N_6104,N_7148);
or U8207 (N_8207,N_7198,N_6747);
or U8208 (N_8208,N_6331,N_7282);
and U8209 (N_8209,N_6887,N_7435);
nor U8210 (N_8210,N_6001,N_6235);
or U8211 (N_8211,N_6155,N_6341);
or U8212 (N_8212,N_6312,N_6853);
nor U8213 (N_8213,N_6223,N_7463);
nand U8214 (N_8214,N_6433,N_6060);
or U8215 (N_8215,N_7127,N_6243);
or U8216 (N_8216,N_7412,N_7405);
nor U8217 (N_8217,N_7374,N_6600);
and U8218 (N_8218,N_7316,N_7425);
and U8219 (N_8219,N_6250,N_7378);
xor U8220 (N_8220,N_6184,N_7432);
or U8221 (N_8221,N_6904,N_6643);
or U8222 (N_8222,N_7026,N_6932);
or U8223 (N_8223,N_6967,N_6873);
nor U8224 (N_8224,N_6477,N_6010);
nand U8225 (N_8225,N_6471,N_6846);
or U8226 (N_8226,N_7064,N_6392);
or U8227 (N_8227,N_6496,N_7327);
and U8228 (N_8228,N_7439,N_6252);
or U8229 (N_8229,N_6059,N_6011);
or U8230 (N_8230,N_6965,N_6453);
nor U8231 (N_8231,N_6772,N_7239);
nor U8232 (N_8232,N_7123,N_6402);
nand U8233 (N_8233,N_7100,N_6852);
nand U8234 (N_8234,N_6702,N_6149);
and U8235 (N_8235,N_7257,N_6753);
or U8236 (N_8236,N_6519,N_6892);
xnor U8237 (N_8237,N_7280,N_6504);
and U8238 (N_8238,N_6436,N_6079);
nand U8239 (N_8239,N_6930,N_6143);
and U8240 (N_8240,N_6765,N_6644);
nor U8241 (N_8241,N_7369,N_7321);
and U8242 (N_8242,N_6704,N_6075);
nand U8243 (N_8243,N_6378,N_7007);
and U8244 (N_8244,N_6318,N_7372);
or U8245 (N_8245,N_7176,N_6952);
xnor U8246 (N_8246,N_6214,N_6913);
or U8247 (N_8247,N_6733,N_7194);
or U8248 (N_8248,N_6604,N_6701);
and U8249 (N_8249,N_6663,N_7218);
xor U8250 (N_8250,N_7050,N_6337);
xor U8251 (N_8251,N_6739,N_6463);
nand U8252 (N_8252,N_6135,N_7005);
nor U8253 (N_8253,N_6931,N_7111);
or U8254 (N_8254,N_7305,N_6130);
and U8255 (N_8255,N_6039,N_6999);
nor U8256 (N_8256,N_6485,N_7209);
nand U8257 (N_8257,N_7205,N_6833);
nor U8258 (N_8258,N_6552,N_7023);
and U8259 (N_8259,N_6509,N_7020);
and U8260 (N_8260,N_7020,N_6635);
or U8261 (N_8261,N_7152,N_7214);
nand U8262 (N_8262,N_6752,N_6173);
nor U8263 (N_8263,N_6541,N_7344);
nand U8264 (N_8264,N_6785,N_6585);
nor U8265 (N_8265,N_7131,N_6072);
and U8266 (N_8266,N_6046,N_6129);
and U8267 (N_8267,N_6974,N_6491);
and U8268 (N_8268,N_6874,N_7045);
nand U8269 (N_8269,N_7152,N_7016);
and U8270 (N_8270,N_6985,N_7476);
or U8271 (N_8271,N_7038,N_6633);
nand U8272 (N_8272,N_7065,N_6583);
or U8273 (N_8273,N_6802,N_6325);
nor U8274 (N_8274,N_6578,N_6227);
nor U8275 (N_8275,N_6646,N_6606);
and U8276 (N_8276,N_6191,N_7446);
and U8277 (N_8277,N_6952,N_6704);
nand U8278 (N_8278,N_6067,N_6788);
and U8279 (N_8279,N_7457,N_6848);
nor U8280 (N_8280,N_6841,N_7158);
nand U8281 (N_8281,N_7192,N_6134);
xnor U8282 (N_8282,N_7254,N_7187);
nor U8283 (N_8283,N_7409,N_6740);
or U8284 (N_8284,N_6299,N_6874);
nand U8285 (N_8285,N_6249,N_6600);
or U8286 (N_8286,N_6244,N_6373);
or U8287 (N_8287,N_6472,N_7428);
nand U8288 (N_8288,N_6446,N_6892);
nor U8289 (N_8289,N_7265,N_7392);
and U8290 (N_8290,N_6392,N_6453);
or U8291 (N_8291,N_7260,N_6189);
nand U8292 (N_8292,N_7007,N_6065);
nor U8293 (N_8293,N_6711,N_6237);
nor U8294 (N_8294,N_7115,N_6695);
nor U8295 (N_8295,N_7061,N_6005);
or U8296 (N_8296,N_7125,N_6750);
nor U8297 (N_8297,N_6074,N_7027);
nor U8298 (N_8298,N_7335,N_6527);
or U8299 (N_8299,N_7393,N_6354);
and U8300 (N_8300,N_6457,N_6193);
nor U8301 (N_8301,N_7128,N_6792);
or U8302 (N_8302,N_6653,N_7165);
or U8303 (N_8303,N_6070,N_7087);
nor U8304 (N_8304,N_6040,N_6456);
and U8305 (N_8305,N_6530,N_6437);
nor U8306 (N_8306,N_6726,N_7169);
xnor U8307 (N_8307,N_6883,N_7048);
or U8308 (N_8308,N_6617,N_6469);
or U8309 (N_8309,N_6735,N_6666);
nor U8310 (N_8310,N_7457,N_7272);
and U8311 (N_8311,N_6718,N_7029);
nor U8312 (N_8312,N_7011,N_7266);
and U8313 (N_8313,N_6549,N_7191);
nor U8314 (N_8314,N_6593,N_6125);
nand U8315 (N_8315,N_7334,N_6541);
and U8316 (N_8316,N_7327,N_7277);
nor U8317 (N_8317,N_6043,N_7108);
nor U8318 (N_8318,N_6702,N_6516);
and U8319 (N_8319,N_6440,N_7082);
nand U8320 (N_8320,N_6689,N_7442);
nand U8321 (N_8321,N_6326,N_7377);
or U8322 (N_8322,N_7240,N_7267);
or U8323 (N_8323,N_7409,N_6947);
or U8324 (N_8324,N_6976,N_6090);
nand U8325 (N_8325,N_6134,N_6708);
nor U8326 (N_8326,N_6892,N_6669);
and U8327 (N_8327,N_6318,N_6306);
or U8328 (N_8328,N_7348,N_6522);
or U8329 (N_8329,N_7066,N_7053);
and U8330 (N_8330,N_6360,N_7050);
nor U8331 (N_8331,N_7395,N_7147);
and U8332 (N_8332,N_6456,N_7240);
nand U8333 (N_8333,N_6168,N_7280);
and U8334 (N_8334,N_6064,N_6626);
and U8335 (N_8335,N_7466,N_6826);
nor U8336 (N_8336,N_6954,N_7302);
and U8337 (N_8337,N_6432,N_6323);
nor U8338 (N_8338,N_6091,N_6627);
nor U8339 (N_8339,N_6576,N_7024);
or U8340 (N_8340,N_6632,N_6682);
nor U8341 (N_8341,N_6766,N_6910);
nand U8342 (N_8342,N_7220,N_6116);
xor U8343 (N_8343,N_6058,N_7238);
or U8344 (N_8344,N_6691,N_7487);
and U8345 (N_8345,N_6902,N_7265);
and U8346 (N_8346,N_6109,N_6807);
nand U8347 (N_8347,N_7062,N_6151);
nor U8348 (N_8348,N_6734,N_6604);
nand U8349 (N_8349,N_6744,N_6354);
nand U8350 (N_8350,N_6301,N_7348);
and U8351 (N_8351,N_6510,N_6149);
nor U8352 (N_8352,N_6669,N_7043);
nor U8353 (N_8353,N_6709,N_6739);
or U8354 (N_8354,N_7292,N_6002);
nand U8355 (N_8355,N_7448,N_6274);
nand U8356 (N_8356,N_7348,N_6896);
and U8357 (N_8357,N_6467,N_6797);
nand U8358 (N_8358,N_6588,N_6403);
nor U8359 (N_8359,N_6563,N_6608);
nor U8360 (N_8360,N_7420,N_7110);
or U8361 (N_8361,N_6207,N_6436);
nand U8362 (N_8362,N_7346,N_7031);
or U8363 (N_8363,N_6121,N_7023);
or U8364 (N_8364,N_7438,N_6296);
nand U8365 (N_8365,N_6713,N_6934);
or U8366 (N_8366,N_6367,N_6730);
xnor U8367 (N_8367,N_6115,N_6843);
and U8368 (N_8368,N_6999,N_6537);
and U8369 (N_8369,N_6215,N_6053);
nor U8370 (N_8370,N_6932,N_7080);
nor U8371 (N_8371,N_6320,N_6055);
nand U8372 (N_8372,N_6218,N_7458);
or U8373 (N_8373,N_6828,N_6320);
and U8374 (N_8374,N_7204,N_6865);
nand U8375 (N_8375,N_6888,N_7460);
or U8376 (N_8376,N_7318,N_6945);
and U8377 (N_8377,N_7331,N_6797);
or U8378 (N_8378,N_6532,N_6831);
or U8379 (N_8379,N_6300,N_7087);
nor U8380 (N_8380,N_7067,N_7282);
nand U8381 (N_8381,N_6161,N_6112);
and U8382 (N_8382,N_6579,N_6487);
or U8383 (N_8383,N_6321,N_6960);
nor U8384 (N_8384,N_6211,N_6695);
nor U8385 (N_8385,N_6946,N_6849);
and U8386 (N_8386,N_6566,N_7360);
nand U8387 (N_8387,N_6427,N_6013);
nand U8388 (N_8388,N_6705,N_6585);
nand U8389 (N_8389,N_7187,N_6047);
or U8390 (N_8390,N_6077,N_7481);
or U8391 (N_8391,N_6584,N_6006);
nand U8392 (N_8392,N_7136,N_7233);
nand U8393 (N_8393,N_7317,N_6668);
nor U8394 (N_8394,N_7280,N_7495);
or U8395 (N_8395,N_6516,N_6808);
and U8396 (N_8396,N_7465,N_7477);
and U8397 (N_8397,N_7189,N_7043);
and U8398 (N_8398,N_6285,N_7114);
and U8399 (N_8399,N_6995,N_6573);
or U8400 (N_8400,N_7066,N_7468);
nor U8401 (N_8401,N_7043,N_6677);
or U8402 (N_8402,N_7096,N_6250);
nand U8403 (N_8403,N_6542,N_6674);
nand U8404 (N_8404,N_6717,N_7080);
nand U8405 (N_8405,N_7046,N_6687);
xor U8406 (N_8406,N_6399,N_6716);
and U8407 (N_8407,N_6329,N_6324);
or U8408 (N_8408,N_6411,N_6783);
and U8409 (N_8409,N_7217,N_6251);
nand U8410 (N_8410,N_6307,N_6578);
nor U8411 (N_8411,N_6658,N_6439);
or U8412 (N_8412,N_6199,N_6146);
nand U8413 (N_8413,N_6025,N_7477);
nand U8414 (N_8414,N_6744,N_6562);
nand U8415 (N_8415,N_6314,N_6671);
and U8416 (N_8416,N_7317,N_7018);
or U8417 (N_8417,N_7224,N_7120);
nor U8418 (N_8418,N_7062,N_6299);
nor U8419 (N_8419,N_6190,N_7389);
nor U8420 (N_8420,N_6964,N_6374);
nor U8421 (N_8421,N_7162,N_6398);
nand U8422 (N_8422,N_7090,N_7128);
nand U8423 (N_8423,N_7348,N_6198);
nor U8424 (N_8424,N_7307,N_6683);
nor U8425 (N_8425,N_6683,N_6974);
nor U8426 (N_8426,N_7085,N_6962);
and U8427 (N_8427,N_6696,N_6163);
nand U8428 (N_8428,N_6251,N_6523);
or U8429 (N_8429,N_7298,N_6504);
nand U8430 (N_8430,N_6674,N_6970);
nand U8431 (N_8431,N_6804,N_6233);
nand U8432 (N_8432,N_6366,N_7313);
or U8433 (N_8433,N_6595,N_6628);
xnor U8434 (N_8434,N_6327,N_6479);
nor U8435 (N_8435,N_6870,N_6115);
and U8436 (N_8436,N_6888,N_7188);
nor U8437 (N_8437,N_6340,N_6048);
or U8438 (N_8438,N_6442,N_6378);
and U8439 (N_8439,N_6950,N_6192);
xnor U8440 (N_8440,N_7474,N_6499);
and U8441 (N_8441,N_7078,N_7216);
nand U8442 (N_8442,N_6077,N_6245);
nand U8443 (N_8443,N_6399,N_6352);
nor U8444 (N_8444,N_6375,N_6308);
nand U8445 (N_8445,N_6872,N_6772);
and U8446 (N_8446,N_7370,N_6238);
or U8447 (N_8447,N_6312,N_7316);
and U8448 (N_8448,N_7036,N_7435);
nor U8449 (N_8449,N_7049,N_7205);
and U8450 (N_8450,N_6388,N_6066);
and U8451 (N_8451,N_6688,N_6645);
nand U8452 (N_8452,N_6268,N_6374);
and U8453 (N_8453,N_6211,N_7188);
nor U8454 (N_8454,N_6606,N_6092);
nor U8455 (N_8455,N_6591,N_6419);
and U8456 (N_8456,N_6970,N_6256);
and U8457 (N_8457,N_6650,N_6038);
or U8458 (N_8458,N_7289,N_6240);
or U8459 (N_8459,N_6234,N_6362);
xor U8460 (N_8460,N_7202,N_6097);
nand U8461 (N_8461,N_6736,N_7330);
nand U8462 (N_8462,N_7089,N_7014);
nand U8463 (N_8463,N_6067,N_7463);
nor U8464 (N_8464,N_6400,N_7464);
and U8465 (N_8465,N_7334,N_6902);
or U8466 (N_8466,N_7459,N_6094);
and U8467 (N_8467,N_6585,N_6695);
nand U8468 (N_8468,N_6331,N_7066);
or U8469 (N_8469,N_6907,N_7325);
nor U8470 (N_8470,N_7194,N_6316);
or U8471 (N_8471,N_6455,N_6889);
and U8472 (N_8472,N_6677,N_7311);
or U8473 (N_8473,N_7384,N_7293);
nand U8474 (N_8474,N_7147,N_7046);
nand U8475 (N_8475,N_7397,N_7400);
or U8476 (N_8476,N_6337,N_6854);
nand U8477 (N_8477,N_6352,N_6412);
and U8478 (N_8478,N_7404,N_7458);
and U8479 (N_8479,N_7334,N_7221);
nor U8480 (N_8480,N_6485,N_6656);
or U8481 (N_8481,N_7494,N_6233);
and U8482 (N_8482,N_7279,N_6703);
and U8483 (N_8483,N_6540,N_6916);
and U8484 (N_8484,N_6592,N_6590);
nand U8485 (N_8485,N_6253,N_6920);
or U8486 (N_8486,N_6201,N_6983);
nand U8487 (N_8487,N_6951,N_6783);
nor U8488 (N_8488,N_6944,N_7104);
and U8489 (N_8489,N_6656,N_6675);
nand U8490 (N_8490,N_7061,N_6340);
xnor U8491 (N_8491,N_6663,N_7399);
nor U8492 (N_8492,N_6247,N_6012);
nor U8493 (N_8493,N_6252,N_7413);
and U8494 (N_8494,N_7096,N_6728);
nor U8495 (N_8495,N_6432,N_6996);
nor U8496 (N_8496,N_6634,N_7271);
and U8497 (N_8497,N_7062,N_7087);
and U8498 (N_8498,N_7105,N_6531);
or U8499 (N_8499,N_7287,N_6073);
or U8500 (N_8500,N_6020,N_7450);
nor U8501 (N_8501,N_7404,N_6674);
nand U8502 (N_8502,N_6899,N_6851);
and U8503 (N_8503,N_6338,N_6421);
nand U8504 (N_8504,N_6806,N_7104);
nand U8505 (N_8505,N_7263,N_7149);
nor U8506 (N_8506,N_6244,N_6536);
nand U8507 (N_8507,N_6671,N_7219);
nor U8508 (N_8508,N_6807,N_6224);
and U8509 (N_8509,N_6323,N_7341);
nand U8510 (N_8510,N_6958,N_6438);
and U8511 (N_8511,N_6409,N_6462);
and U8512 (N_8512,N_7062,N_6479);
and U8513 (N_8513,N_6655,N_6359);
or U8514 (N_8514,N_7499,N_6415);
nor U8515 (N_8515,N_6917,N_7229);
or U8516 (N_8516,N_7382,N_6686);
nand U8517 (N_8517,N_6401,N_7186);
nor U8518 (N_8518,N_6559,N_6603);
and U8519 (N_8519,N_7312,N_6788);
and U8520 (N_8520,N_6872,N_7166);
and U8521 (N_8521,N_6284,N_7199);
or U8522 (N_8522,N_6477,N_6695);
and U8523 (N_8523,N_7320,N_6348);
and U8524 (N_8524,N_6889,N_6413);
or U8525 (N_8525,N_6597,N_7136);
nand U8526 (N_8526,N_7224,N_6245);
or U8527 (N_8527,N_6729,N_6092);
nand U8528 (N_8528,N_6648,N_6781);
nor U8529 (N_8529,N_6771,N_6242);
nor U8530 (N_8530,N_6952,N_7084);
or U8531 (N_8531,N_6665,N_6051);
nand U8532 (N_8532,N_7280,N_6030);
or U8533 (N_8533,N_7220,N_7385);
nor U8534 (N_8534,N_6636,N_6490);
or U8535 (N_8535,N_6351,N_6720);
or U8536 (N_8536,N_7122,N_6575);
nand U8537 (N_8537,N_6475,N_6744);
or U8538 (N_8538,N_7495,N_6864);
nand U8539 (N_8539,N_6721,N_6674);
and U8540 (N_8540,N_7200,N_7260);
nor U8541 (N_8541,N_7427,N_7385);
nor U8542 (N_8542,N_7007,N_6120);
nor U8543 (N_8543,N_6994,N_6055);
nor U8544 (N_8544,N_7387,N_6701);
and U8545 (N_8545,N_7295,N_7019);
nand U8546 (N_8546,N_6411,N_6799);
nand U8547 (N_8547,N_7242,N_6463);
and U8548 (N_8548,N_7065,N_7292);
nand U8549 (N_8549,N_7308,N_6689);
nor U8550 (N_8550,N_7046,N_6022);
or U8551 (N_8551,N_6929,N_6430);
nand U8552 (N_8552,N_6376,N_7369);
or U8553 (N_8553,N_6482,N_7459);
and U8554 (N_8554,N_6665,N_6045);
nand U8555 (N_8555,N_6534,N_7211);
or U8556 (N_8556,N_6998,N_7471);
nand U8557 (N_8557,N_7086,N_7465);
and U8558 (N_8558,N_7345,N_7321);
nand U8559 (N_8559,N_6666,N_7101);
and U8560 (N_8560,N_6725,N_6026);
or U8561 (N_8561,N_6090,N_6719);
or U8562 (N_8562,N_7131,N_6497);
nor U8563 (N_8563,N_7049,N_7109);
or U8564 (N_8564,N_7076,N_6851);
and U8565 (N_8565,N_6402,N_6317);
nor U8566 (N_8566,N_6081,N_6894);
nand U8567 (N_8567,N_6645,N_6385);
or U8568 (N_8568,N_6645,N_7411);
nand U8569 (N_8569,N_6290,N_7102);
xor U8570 (N_8570,N_6766,N_6742);
or U8571 (N_8571,N_6389,N_7025);
and U8572 (N_8572,N_7112,N_7428);
or U8573 (N_8573,N_6742,N_7217);
nor U8574 (N_8574,N_6496,N_7351);
nand U8575 (N_8575,N_6009,N_6693);
nor U8576 (N_8576,N_6935,N_6445);
nor U8577 (N_8577,N_6839,N_7005);
xnor U8578 (N_8578,N_7044,N_6667);
nor U8579 (N_8579,N_6636,N_6572);
or U8580 (N_8580,N_7057,N_6319);
nand U8581 (N_8581,N_7356,N_7393);
nor U8582 (N_8582,N_7120,N_6341);
or U8583 (N_8583,N_6483,N_7471);
and U8584 (N_8584,N_7028,N_6690);
nor U8585 (N_8585,N_6814,N_6422);
and U8586 (N_8586,N_6642,N_6831);
nand U8587 (N_8587,N_6086,N_6958);
nor U8588 (N_8588,N_6121,N_6555);
nand U8589 (N_8589,N_6978,N_7494);
and U8590 (N_8590,N_7490,N_6658);
and U8591 (N_8591,N_7363,N_6362);
or U8592 (N_8592,N_7128,N_6566);
and U8593 (N_8593,N_7004,N_7166);
nand U8594 (N_8594,N_7241,N_6108);
or U8595 (N_8595,N_6024,N_6182);
nor U8596 (N_8596,N_6655,N_6990);
and U8597 (N_8597,N_7004,N_6213);
nand U8598 (N_8598,N_7412,N_7122);
or U8599 (N_8599,N_6383,N_7297);
and U8600 (N_8600,N_6630,N_7107);
and U8601 (N_8601,N_7344,N_6754);
nand U8602 (N_8602,N_6919,N_7326);
xor U8603 (N_8603,N_6286,N_6229);
nand U8604 (N_8604,N_7084,N_6940);
nor U8605 (N_8605,N_6231,N_6089);
nand U8606 (N_8606,N_7155,N_6613);
nor U8607 (N_8607,N_6820,N_7040);
or U8608 (N_8608,N_6445,N_7252);
and U8609 (N_8609,N_7331,N_6226);
and U8610 (N_8610,N_6741,N_7336);
nor U8611 (N_8611,N_6352,N_6101);
or U8612 (N_8612,N_7351,N_6602);
nand U8613 (N_8613,N_6690,N_6176);
nand U8614 (N_8614,N_6379,N_6191);
nand U8615 (N_8615,N_6157,N_6658);
nor U8616 (N_8616,N_6171,N_6956);
nor U8617 (N_8617,N_6214,N_7439);
nand U8618 (N_8618,N_7034,N_7015);
and U8619 (N_8619,N_6946,N_7207);
nor U8620 (N_8620,N_6569,N_6885);
nand U8621 (N_8621,N_6941,N_6464);
or U8622 (N_8622,N_6703,N_6005);
nor U8623 (N_8623,N_6613,N_7016);
nor U8624 (N_8624,N_7094,N_6088);
xnor U8625 (N_8625,N_7377,N_7014);
nor U8626 (N_8626,N_7490,N_6653);
nor U8627 (N_8627,N_7408,N_6393);
and U8628 (N_8628,N_6982,N_7340);
or U8629 (N_8629,N_7119,N_7126);
and U8630 (N_8630,N_7451,N_6317);
nor U8631 (N_8631,N_6522,N_7357);
and U8632 (N_8632,N_6258,N_6405);
and U8633 (N_8633,N_6398,N_6908);
and U8634 (N_8634,N_7076,N_6100);
or U8635 (N_8635,N_6626,N_6036);
nor U8636 (N_8636,N_7004,N_7277);
xor U8637 (N_8637,N_6308,N_7007);
nand U8638 (N_8638,N_7469,N_6611);
nand U8639 (N_8639,N_6278,N_6606);
nand U8640 (N_8640,N_6604,N_7332);
and U8641 (N_8641,N_7131,N_6950);
and U8642 (N_8642,N_6470,N_7213);
nand U8643 (N_8643,N_6488,N_7456);
nor U8644 (N_8644,N_7033,N_7017);
and U8645 (N_8645,N_6830,N_6606);
or U8646 (N_8646,N_7302,N_6970);
and U8647 (N_8647,N_6108,N_6868);
or U8648 (N_8648,N_6669,N_7104);
nand U8649 (N_8649,N_6932,N_6632);
and U8650 (N_8650,N_6331,N_6080);
or U8651 (N_8651,N_7020,N_7383);
nor U8652 (N_8652,N_7345,N_6484);
nand U8653 (N_8653,N_7066,N_7443);
or U8654 (N_8654,N_6272,N_6315);
and U8655 (N_8655,N_6532,N_6588);
xnor U8656 (N_8656,N_6830,N_6788);
or U8657 (N_8657,N_6795,N_6442);
nor U8658 (N_8658,N_7374,N_6387);
nand U8659 (N_8659,N_6983,N_6217);
or U8660 (N_8660,N_6599,N_7452);
nor U8661 (N_8661,N_6333,N_7428);
and U8662 (N_8662,N_7394,N_7320);
nor U8663 (N_8663,N_7110,N_6668);
or U8664 (N_8664,N_7141,N_7388);
and U8665 (N_8665,N_6087,N_7362);
and U8666 (N_8666,N_6306,N_7044);
nor U8667 (N_8667,N_6050,N_6980);
or U8668 (N_8668,N_6245,N_7397);
nand U8669 (N_8669,N_7216,N_6205);
xnor U8670 (N_8670,N_6635,N_6809);
or U8671 (N_8671,N_7093,N_6615);
nor U8672 (N_8672,N_6456,N_6078);
nor U8673 (N_8673,N_6484,N_6098);
and U8674 (N_8674,N_7346,N_6109);
nor U8675 (N_8675,N_6440,N_7172);
nand U8676 (N_8676,N_7366,N_7479);
nor U8677 (N_8677,N_6061,N_6387);
and U8678 (N_8678,N_7007,N_6456);
nor U8679 (N_8679,N_6732,N_6526);
or U8680 (N_8680,N_7311,N_6216);
nor U8681 (N_8681,N_7015,N_7127);
nor U8682 (N_8682,N_6645,N_7355);
and U8683 (N_8683,N_7179,N_6996);
nor U8684 (N_8684,N_6403,N_7275);
and U8685 (N_8685,N_7297,N_6624);
nor U8686 (N_8686,N_6878,N_7461);
nor U8687 (N_8687,N_6212,N_6124);
and U8688 (N_8688,N_7070,N_7476);
and U8689 (N_8689,N_6556,N_6913);
nand U8690 (N_8690,N_6444,N_6819);
nand U8691 (N_8691,N_6995,N_7135);
xor U8692 (N_8692,N_6955,N_7176);
and U8693 (N_8693,N_7000,N_7275);
xor U8694 (N_8694,N_6631,N_7344);
or U8695 (N_8695,N_7108,N_7204);
and U8696 (N_8696,N_6757,N_6667);
nor U8697 (N_8697,N_6260,N_7118);
and U8698 (N_8698,N_6144,N_6170);
nor U8699 (N_8699,N_6878,N_7159);
and U8700 (N_8700,N_6449,N_6076);
nand U8701 (N_8701,N_6860,N_7263);
nand U8702 (N_8702,N_6379,N_6387);
or U8703 (N_8703,N_7201,N_7156);
nor U8704 (N_8704,N_7318,N_6747);
nor U8705 (N_8705,N_6338,N_6780);
or U8706 (N_8706,N_6153,N_6516);
or U8707 (N_8707,N_6198,N_6692);
and U8708 (N_8708,N_6650,N_6495);
nand U8709 (N_8709,N_6063,N_6118);
and U8710 (N_8710,N_6556,N_6016);
or U8711 (N_8711,N_6128,N_6375);
and U8712 (N_8712,N_7278,N_7301);
or U8713 (N_8713,N_6497,N_6676);
and U8714 (N_8714,N_6596,N_6440);
and U8715 (N_8715,N_6983,N_6255);
and U8716 (N_8716,N_6547,N_7317);
or U8717 (N_8717,N_6667,N_6765);
or U8718 (N_8718,N_6308,N_7206);
xor U8719 (N_8719,N_6584,N_6907);
nor U8720 (N_8720,N_7263,N_7055);
or U8721 (N_8721,N_7010,N_6725);
and U8722 (N_8722,N_6441,N_6996);
nand U8723 (N_8723,N_6951,N_7139);
or U8724 (N_8724,N_6380,N_6751);
nor U8725 (N_8725,N_6245,N_7496);
nand U8726 (N_8726,N_6149,N_7366);
and U8727 (N_8727,N_7445,N_7471);
nor U8728 (N_8728,N_6564,N_6685);
nand U8729 (N_8729,N_6319,N_6768);
or U8730 (N_8730,N_6313,N_7037);
and U8731 (N_8731,N_6304,N_7364);
and U8732 (N_8732,N_6543,N_6915);
or U8733 (N_8733,N_6970,N_6684);
nor U8734 (N_8734,N_6491,N_6196);
nand U8735 (N_8735,N_6266,N_6717);
or U8736 (N_8736,N_6873,N_6583);
xor U8737 (N_8737,N_6656,N_7347);
nand U8738 (N_8738,N_7131,N_6434);
or U8739 (N_8739,N_6070,N_6693);
nor U8740 (N_8740,N_7253,N_6117);
nor U8741 (N_8741,N_7274,N_6515);
and U8742 (N_8742,N_6681,N_6504);
or U8743 (N_8743,N_7493,N_6067);
or U8744 (N_8744,N_6718,N_7088);
nand U8745 (N_8745,N_7411,N_6957);
or U8746 (N_8746,N_7210,N_7160);
or U8747 (N_8747,N_7485,N_7365);
nor U8748 (N_8748,N_6922,N_7047);
nor U8749 (N_8749,N_6065,N_6538);
nand U8750 (N_8750,N_6295,N_6101);
nand U8751 (N_8751,N_6797,N_6776);
nor U8752 (N_8752,N_6260,N_6873);
and U8753 (N_8753,N_6365,N_6070);
or U8754 (N_8754,N_6963,N_7152);
and U8755 (N_8755,N_6525,N_6051);
and U8756 (N_8756,N_6236,N_6069);
and U8757 (N_8757,N_6820,N_6215);
nand U8758 (N_8758,N_6130,N_7042);
nor U8759 (N_8759,N_7406,N_6652);
or U8760 (N_8760,N_7077,N_7004);
and U8761 (N_8761,N_6891,N_7479);
nor U8762 (N_8762,N_6596,N_7467);
or U8763 (N_8763,N_6191,N_6905);
or U8764 (N_8764,N_7115,N_7060);
nor U8765 (N_8765,N_7248,N_6305);
nand U8766 (N_8766,N_6208,N_6548);
and U8767 (N_8767,N_6958,N_6421);
nand U8768 (N_8768,N_7165,N_7248);
xor U8769 (N_8769,N_6977,N_6412);
nor U8770 (N_8770,N_6576,N_6827);
or U8771 (N_8771,N_7487,N_7381);
nor U8772 (N_8772,N_7375,N_6148);
nor U8773 (N_8773,N_6461,N_6437);
nor U8774 (N_8774,N_6411,N_6335);
xor U8775 (N_8775,N_7243,N_6674);
nor U8776 (N_8776,N_6713,N_6834);
nor U8777 (N_8777,N_6242,N_7046);
nand U8778 (N_8778,N_7148,N_6522);
nand U8779 (N_8779,N_6749,N_6571);
or U8780 (N_8780,N_6456,N_6392);
nor U8781 (N_8781,N_6879,N_6242);
nor U8782 (N_8782,N_7301,N_7274);
nand U8783 (N_8783,N_6548,N_6188);
nand U8784 (N_8784,N_6819,N_6730);
and U8785 (N_8785,N_6727,N_7477);
nand U8786 (N_8786,N_6381,N_6403);
nand U8787 (N_8787,N_6794,N_6503);
and U8788 (N_8788,N_6436,N_6794);
and U8789 (N_8789,N_6936,N_6699);
and U8790 (N_8790,N_6971,N_6297);
and U8791 (N_8791,N_6903,N_7211);
nand U8792 (N_8792,N_6686,N_7170);
nand U8793 (N_8793,N_6887,N_6471);
nand U8794 (N_8794,N_6146,N_6281);
and U8795 (N_8795,N_6274,N_6259);
and U8796 (N_8796,N_7307,N_6961);
or U8797 (N_8797,N_6317,N_7034);
nor U8798 (N_8798,N_6245,N_6672);
or U8799 (N_8799,N_6052,N_6791);
nor U8800 (N_8800,N_6938,N_7188);
nor U8801 (N_8801,N_6653,N_6364);
and U8802 (N_8802,N_6465,N_7272);
nand U8803 (N_8803,N_7348,N_7376);
or U8804 (N_8804,N_6751,N_6302);
or U8805 (N_8805,N_6383,N_6658);
nor U8806 (N_8806,N_6613,N_6830);
nor U8807 (N_8807,N_7280,N_7046);
nor U8808 (N_8808,N_6824,N_6454);
and U8809 (N_8809,N_6570,N_6054);
nor U8810 (N_8810,N_7431,N_6196);
or U8811 (N_8811,N_7174,N_6733);
nand U8812 (N_8812,N_6191,N_6025);
or U8813 (N_8813,N_7178,N_6519);
and U8814 (N_8814,N_6794,N_7369);
or U8815 (N_8815,N_6872,N_6115);
nand U8816 (N_8816,N_7315,N_7220);
nor U8817 (N_8817,N_6040,N_6498);
nand U8818 (N_8818,N_6948,N_6709);
and U8819 (N_8819,N_7285,N_7480);
or U8820 (N_8820,N_6399,N_6099);
or U8821 (N_8821,N_6786,N_7487);
nand U8822 (N_8822,N_6399,N_6757);
nor U8823 (N_8823,N_6779,N_7450);
nor U8824 (N_8824,N_7009,N_6755);
or U8825 (N_8825,N_6347,N_6537);
nor U8826 (N_8826,N_7475,N_6253);
or U8827 (N_8827,N_6062,N_7256);
nor U8828 (N_8828,N_7009,N_6614);
nor U8829 (N_8829,N_6029,N_6536);
nand U8830 (N_8830,N_7416,N_6235);
nand U8831 (N_8831,N_7050,N_6248);
nor U8832 (N_8832,N_7294,N_6986);
nand U8833 (N_8833,N_7362,N_7218);
and U8834 (N_8834,N_6122,N_6565);
nand U8835 (N_8835,N_6341,N_7086);
nand U8836 (N_8836,N_7426,N_6341);
and U8837 (N_8837,N_6479,N_6463);
and U8838 (N_8838,N_6502,N_7161);
or U8839 (N_8839,N_7234,N_7276);
and U8840 (N_8840,N_6807,N_7011);
nand U8841 (N_8841,N_6846,N_6328);
or U8842 (N_8842,N_6637,N_7400);
nand U8843 (N_8843,N_6026,N_6659);
or U8844 (N_8844,N_6300,N_6917);
nand U8845 (N_8845,N_7206,N_6506);
nor U8846 (N_8846,N_6620,N_6758);
or U8847 (N_8847,N_6663,N_7346);
or U8848 (N_8848,N_6977,N_6621);
nand U8849 (N_8849,N_6463,N_7015);
nand U8850 (N_8850,N_7262,N_6060);
and U8851 (N_8851,N_6507,N_6708);
and U8852 (N_8852,N_6209,N_6817);
and U8853 (N_8853,N_6688,N_7160);
nor U8854 (N_8854,N_6156,N_6989);
and U8855 (N_8855,N_7202,N_7424);
and U8856 (N_8856,N_6831,N_6024);
or U8857 (N_8857,N_7242,N_7343);
nor U8858 (N_8858,N_6865,N_6964);
or U8859 (N_8859,N_7250,N_6770);
and U8860 (N_8860,N_6029,N_6073);
or U8861 (N_8861,N_6646,N_6863);
or U8862 (N_8862,N_7210,N_7088);
nor U8863 (N_8863,N_6692,N_6664);
nand U8864 (N_8864,N_7371,N_6938);
or U8865 (N_8865,N_6825,N_7224);
or U8866 (N_8866,N_6498,N_7312);
nor U8867 (N_8867,N_6912,N_6465);
nand U8868 (N_8868,N_6206,N_6376);
and U8869 (N_8869,N_6931,N_6755);
nor U8870 (N_8870,N_6322,N_6129);
or U8871 (N_8871,N_7443,N_6920);
nor U8872 (N_8872,N_6426,N_7277);
or U8873 (N_8873,N_6969,N_6009);
nand U8874 (N_8874,N_6722,N_6001);
or U8875 (N_8875,N_6802,N_6070);
or U8876 (N_8876,N_6367,N_6183);
and U8877 (N_8877,N_6726,N_6853);
and U8878 (N_8878,N_6332,N_6165);
or U8879 (N_8879,N_7038,N_6679);
or U8880 (N_8880,N_6686,N_6642);
nor U8881 (N_8881,N_6783,N_6899);
and U8882 (N_8882,N_6887,N_6350);
or U8883 (N_8883,N_6660,N_6014);
nand U8884 (N_8884,N_6841,N_6104);
nand U8885 (N_8885,N_6643,N_7163);
nor U8886 (N_8886,N_7176,N_6210);
or U8887 (N_8887,N_6715,N_6432);
nor U8888 (N_8888,N_7315,N_7076);
nand U8889 (N_8889,N_7249,N_7000);
and U8890 (N_8890,N_7134,N_7146);
nand U8891 (N_8891,N_6309,N_7012);
or U8892 (N_8892,N_6399,N_6176);
xor U8893 (N_8893,N_6394,N_6102);
and U8894 (N_8894,N_7141,N_6585);
or U8895 (N_8895,N_6546,N_7215);
nor U8896 (N_8896,N_7043,N_6123);
nor U8897 (N_8897,N_7235,N_7486);
nand U8898 (N_8898,N_6703,N_6952);
xor U8899 (N_8899,N_7339,N_6454);
and U8900 (N_8900,N_6464,N_6540);
nand U8901 (N_8901,N_6407,N_7132);
or U8902 (N_8902,N_6530,N_6723);
nor U8903 (N_8903,N_6731,N_7298);
nor U8904 (N_8904,N_7105,N_7085);
and U8905 (N_8905,N_6133,N_6337);
nand U8906 (N_8906,N_6100,N_6306);
nor U8907 (N_8907,N_6207,N_7129);
or U8908 (N_8908,N_6766,N_7302);
nand U8909 (N_8909,N_6739,N_6629);
nand U8910 (N_8910,N_6273,N_6695);
nand U8911 (N_8911,N_7425,N_6031);
nand U8912 (N_8912,N_6618,N_6540);
or U8913 (N_8913,N_7282,N_6532);
or U8914 (N_8914,N_7454,N_6504);
nor U8915 (N_8915,N_6082,N_6736);
and U8916 (N_8916,N_6048,N_6357);
and U8917 (N_8917,N_6087,N_6545);
nor U8918 (N_8918,N_7326,N_7421);
and U8919 (N_8919,N_6726,N_6183);
nor U8920 (N_8920,N_6866,N_6090);
nor U8921 (N_8921,N_7460,N_6621);
or U8922 (N_8922,N_6121,N_6943);
nand U8923 (N_8923,N_7371,N_6093);
and U8924 (N_8924,N_6013,N_6660);
nand U8925 (N_8925,N_7467,N_6569);
and U8926 (N_8926,N_6134,N_6794);
nand U8927 (N_8927,N_6833,N_7420);
nand U8928 (N_8928,N_6456,N_6471);
nand U8929 (N_8929,N_6233,N_6278);
nand U8930 (N_8930,N_6403,N_6412);
or U8931 (N_8931,N_6911,N_7160);
or U8932 (N_8932,N_6122,N_7371);
or U8933 (N_8933,N_7446,N_6967);
nor U8934 (N_8934,N_6344,N_6194);
or U8935 (N_8935,N_7353,N_7114);
and U8936 (N_8936,N_7087,N_6342);
or U8937 (N_8937,N_6126,N_7318);
or U8938 (N_8938,N_7019,N_6331);
nor U8939 (N_8939,N_6007,N_6324);
nand U8940 (N_8940,N_6626,N_6324);
nand U8941 (N_8941,N_6419,N_6046);
nor U8942 (N_8942,N_6671,N_6641);
and U8943 (N_8943,N_6199,N_6773);
or U8944 (N_8944,N_6725,N_7443);
or U8945 (N_8945,N_6936,N_6527);
nand U8946 (N_8946,N_6382,N_7353);
nand U8947 (N_8947,N_7049,N_6922);
or U8948 (N_8948,N_7255,N_7137);
xnor U8949 (N_8949,N_7185,N_7316);
or U8950 (N_8950,N_6993,N_7170);
nand U8951 (N_8951,N_6944,N_6101);
or U8952 (N_8952,N_6688,N_6639);
xnor U8953 (N_8953,N_7174,N_6225);
nor U8954 (N_8954,N_7435,N_6801);
nand U8955 (N_8955,N_6582,N_6493);
nor U8956 (N_8956,N_7418,N_6840);
nand U8957 (N_8957,N_6797,N_7082);
or U8958 (N_8958,N_6284,N_7200);
nand U8959 (N_8959,N_7473,N_6888);
and U8960 (N_8960,N_6933,N_7454);
xor U8961 (N_8961,N_7159,N_6506);
or U8962 (N_8962,N_6000,N_6120);
and U8963 (N_8963,N_7473,N_6034);
nand U8964 (N_8964,N_7462,N_7036);
and U8965 (N_8965,N_6626,N_6897);
nor U8966 (N_8966,N_6738,N_6097);
and U8967 (N_8967,N_6620,N_6814);
nand U8968 (N_8968,N_6324,N_7188);
nor U8969 (N_8969,N_6322,N_6851);
xnor U8970 (N_8970,N_6602,N_6952);
nor U8971 (N_8971,N_6438,N_7091);
nand U8972 (N_8972,N_6966,N_6357);
nand U8973 (N_8973,N_6072,N_6668);
nand U8974 (N_8974,N_7188,N_6129);
nand U8975 (N_8975,N_6823,N_7413);
nand U8976 (N_8976,N_7359,N_6718);
nand U8977 (N_8977,N_7335,N_6462);
and U8978 (N_8978,N_7290,N_6115);
nand U8979 (N_8979,N_6186,N_6578);
nand U8980 (N_8980,N_7098,N_6091);
or U8981 (N_8981,N_6288,N_6231);
nand U8982 (N_8982,N_7166,N_7020);
or U8983 (N_8983,N_6875,N_7482);
nand U8984 (N_8984,N_6493,N_6484);
or U8985 (N_8985,N_6376,N_7097);
nand U8986 (N_8986,N_7174,N_7113);
nor U8987 (N_8987,N_6227,N_7204);
or U8988 (N_8988,N_7251,N_6144);
nand U8989 (N_8989,N_7138,N_7372);
or U8990 (N_8990,N_7286,N_6961);
or U8991 (N_8991,N_6364,N_7118);
or U8992 (N_8992,N_7499,N_6490);
or U8993 (N_8993,N_6502,N_6507);
and U8994 (N_8994,N_6747,N_6400);
or U8995 (N_8995,N_6393,N_7396);
or U8996 (N_8996,N_7240,N_6510);
nand U8997 (N_8997,N_6454,N_7335);
or U8998 (N_8998,N_7138,N_6787);
or U8999 (N_8999,N_6577,N_7247);
nand U9000 (N_9000,N_7723,N_7798);
or U9001 (N_9001,N_7910,N_8554);
nand U9002 (N_9002,N_7847,N_8058);
or U9003 (N_9003,N_7650,N_7884);
nand U9004 (N_9004,N_8812,N_7516);
or U9005 (N_9005,N_8498,N_8491);
nand U9006 (N_9006,N_8199,N_7523);
nand U9007 (N_9007,N_7637,N_8042);
or U9008 (N_9008,N_7857,N_8173);
nor U9009 (N_9009,N_7975,N_8292);
nand U9010 (N_9010,N_8783,N_8793);
and U9011 (N_9011,N_8557,N_8249);
and U9012 (N_9012,N_8466,N_8123);
nor U9013 (N_9013,N_8006,N_8914);
nor U9014 (N_9014,N_8564,N_8116);
nor U9015 (N_9015,N_7564,N_7712);
and U9016 (N_9016,N_8069,N_7687);
nand U9017 (N_9017,N_8830,N_8332);
or U9018 (N_9018,N_8258,N_8220);
xnor U9019 (N_9019,N_8854,N_7554);
and U9020 (N_9020,N_8159,N_8255);
xor U9021 (N_9021,N_7827,N_7621);
nand U9022 (N_9022,N_7691,N_8031);
or U9023 (N_9023,N_7515,N_7826);
nand U9024 (N_9024,N_8716,N_8918);
or U9025 (N_9025,N_8883,N_7577);
or U9026 (N_9026,N_7856,N_8707);
nor U9027 (N_9027,N_8115,N_8270);
and U9028 (N_9028,N_7700,N_7665);
nand U9029 (N_9029,N_7941,N_8556);
or U9030 (N_9030,N_8448,N_8935);
or U9031 (N_9031,N_8364,N_7732);
or U9032 (N_9032,N_8369,N_8517);
or U9033 (N_9033,N_8382,N_8794);
or U9034 (N_9034,N_8765,N_8522);
and U9035 (N_9035,N_7570,N_8316);
nand U9036 (N_9036,N_8577,N_8379);
nor U9037 (N_9037,N_7654,N_7681);
nor U9038 (N_9038,N_8814,N_8322);
xor U9039 (N_9039,N_8462,N_7529);
and U9040 (N_9040,N_8790,N_8548);
or U9041 (N_9041,N_8430,N_8238);
or U9042 (N_9042,N_8455,N_7814);
and U9043 (N_9043,N_7722,N_7950);
and U9044 (N_9044,N_8032,N_8505);
nand U9045 (N_9045,N_8200,N_8020);
nand U9046 (N_9046,N_8097,N_7559);
or U9047 (N_9047,N_7573,N_8186);
or U9048 (N_9048,N_8131,N_8162);
and U9049 (N_9049,N_7824,N_8699);
nand U9050 (N_9050,N_8863,N_7728);
nor U9051 (N_9051,N_8834,N_8202);
nand U9052 (N_9052,N_8022,N_7575);
nor U9053 (N_9053,N_8867,N_8212);
nand U9054 (N_9054,N_8683,N_8372);
or U9055 (N_9055,N_8296,N_8756);
and U9056 (N_9056,N_7678,N_8282);
nand U9057 (N_9057,N_8074,N_8128);
or U9058 (N_9058,N_8518,N_8230);
nand U9059 (N_9059,N_8050,N_8968);
nor U9060 (N_9060,N_8330,N_8938);
nor U9061 (N_9061,N_7822,N_7789);
nor U9062 (N_9062,N_8616,N_7942);
nor U9063 (N_9063,N_8109,N_8713);
and U9064 (N_9064,N_8860,N_7737);
or U9065 (N_9065,N_8519,N_8954);
nor U9066 (N_9066,N_7717,N_8187);
nand U9067 (N_9067,N_8464,N_8908);
and U9068 (N_9068,N_8946,N_8797);
nand U9069 (N_9069,N_8171,N_8653);
and U9070 (N_9070,N_7679,N_8471);
or U9071 (N_9071,N_8185,N_8429);
nand U9072 (N_9072,N_8759,N_8383);
or U9073 (N_9073,N_8512,N_8996);
or U9074 (N_9074,N_8389,N_8843);
and U9075 (N_9075,N_8966,N_8664);
nor U9076 (N_9076,N_7749,N_7916);
nor U9077 (N_9077,N_8009,N_8126);
nand U9078 (N_9078,N_8813,N_8091);
and U9079 (N_9079,N_7602,N_8559);
nand U9080 (N_9080,N_7846,N_8514);
nor U9081 (N_9081,N_8399,N_8374);
nand U9082 (N_9082,N_8944,N_7599);
and U9083 (N_9083,N_8076,N_8825);
or U9084 (N_9084,N_8041,N_8142);
nor U9085 (N_9085,N_7859,N_7763);
and U9086 (N_9086,N_8301,N_8375);
nor U9087 (N_9087,N_8649,N_8335);
and U9088 (N_9088,N_7592,N_7802);
nor U9089 (N_9089,N_8515,N_8879);
nor U9090 (N_9090,N_8194,N_7956);
and U9091 (N_9091,N_8388,N_8085);
or U9092 (N_9092,N_8855,N_8082);
nand U9093 (N_9093,N_8392,N_8808);
and U9094 (N_9094,N_8784,N_8071);
or U9095 (N_9095,N_8774,N_8681);
xor U9096 (N_9096,N_7695,N_8799);
nand U9097 (N_9097,N_7897,N_8624);
and U9098 (N_9098,N_8838,N_8899);
and U9099 (N_9099,N_8546,N_8955);
nand U9100 (N_9100,N_8807,N_7873);
and U9101 (N_9101,N_8079,N_8357);
or U9102 (N_9102,N_8796,N_7848);
nor U9103 (N_9103,N_8562,N_8304);
and U9104 (N_9104,N_8333,N_8578);
nor U9105 (N_9105,N_8481,N_8534);
nand U9106 (N_9106,N_8129,N_8178);
nand U9107 (N_9107,N_7840,N_8198);
nand U9108 (N_9108,N_8362,N_7819);
nand U9109 (N_9109,N_7981,N_8054);
or U9110 (N_9110,N_8767,N_7553);
nor U9111 (N_9111,N_8605,N_8916);
or U9112 (N_9112,N_8975,N_8474);
nand U9113 (N_9113,N_7755,N_8581);
nand U9114 (N_9114,N_8601,N_7539);
or U9115 (N_9115,N_8727,N_7626);
or U9116 (N_9116,N_8911,N_8252);
nand U9117 (N_9117,N_7780,N_7607);
and U9118 (N_9118,N_7880,N_8422);
nor U9119 (N_9119,N_8469,N_8277);
and U9120 (N_9120,N_8510,N_7630);
xor U9121 (N_9121,N_8486,N_8254);
nand U9122 (N_9122,N_8211,N_8720);
nand U9123 (N_9123,N_8340,N_8743);
or U9124 (N_9124,N_8218,N_8444);
and U9125 (N_9125,N_8468,N_8235);
nor U9126 (N_9126,N_8351,N_8647);
or U9127 (N_9127,N_8603,N_7534);
nand U9128 (N_9128,N_8037,N_7514);
and U9129 (N_9129,N_8237,N_8673);
or U9130 (N_9130,N_8885,N_8105);
nand U9131 (N_9131,N_8490,N_8910);
nand U9132 (N_9132,N_8411,N_8046);
and U9133 (N_9133,N_8922,N_7508);
or U9134 (N_9134,N_8950,N_8284);
and U9135 (N_9135,N_7563,N_8421);
nand U9136 (N_9136,N_7813,N_7644);
nor U9137 (N_9137,N_7851,N_7904);
nor U9138 (N_9138,N_8192,N_7836);
or U9139 (N_9139,N_8070,N_7733);
nor U9140 (N_9140,N_8567,N_8053);
and U9141 (N_9141,N_7886,N_7697);
and U9142 (N_9142,N_7866,N_8524);
nor U9143 (N_9143,N_8775,N_8158);
nor U9144 (N_9144,N_7590,N_7993);
nor U9145 (N_9145,N_7593,N_8299);
or U9146 (N_9146,N_8163,N_8160);
nor U9147 (N_9147,N_7560,N_8538);
nor U9148 (N_9148,N_7582,N_7929);
and U9149 (N_9149,N_8589,N_8811);
nor U9150 (N_9150,N_8580,N_8485);
or U9151 (N_9151,N_7696,N_8182);
nand U9152 (N_9152,N_8776,N_7513);
or U9153 (N_9153,N_8225,N_8835);
nor U9154 (N_9154,N_8452,N_8312);
nor U9155 (N_9155,N_7624,N_7527);
nand U9156 (N_9156,N_8543,N_8446);
and U9157 (N_9157,N_8598,N_8663);
or U9158 (N_9158,N_7597,N_8532);
nor U9159 (N_9159,N_8431,N_8995);
or U9160 (N_9160,N_8615,N_7642);
and U9161 (N_9161,N_8810,N_8643);
nor U9162 (N_9162,N_8437,N_7990);
and U9163 (N_9163,N_8149,N_8994);
and U9164 (N_9164,N_8343,N_7883);
nand U9165 (N_9165,N_8461,N_8177);
nor U9166 (N_9166,N_8387,N_7812);
or U9167 (N_9167,N_8919,N_8831);
nand U9168 (N_9168,N_8253,N_8868);
or U9169 (N_9169,N_8926,N_8401);
or U9170 (N_9170,N_8426,N_7980);
nand U9171 (N_9171,N_8297,N_7953);
and U9172 (N_9172,N_8949,N_8859);
nor U9173 (N_9173,N_7730,N_8127);
or U9174 (N_9174,N_8658,N_7633);
or U9175 (N_9175,N_8817,N_8584);
xor U9176 (N_9176,N_7537,N_8685);
nor U9177 (N_9177,N_7977,N_7754);
and U9178 (N_9178,N_7815,N_7896);
and U9179 (N_9179,N_7984,N_8962);
or U9180 (N_9180,N_8690,N_8771);
and U9181 (N_9181,N_8875,N_8094);
and U9182 (N_9182,N_8132,N_7522);
or U9183 (N_9183,N_7585,N_8118);
or U9184 (N_9184,N_8969,N_8089);
nand U9185 (N_9185,N_8752,N_7881);
or U9186 (N_9186,N_8325,N_7799);
nor U9187 (N_9187,N_8978,N_7605);
or U9188 (N_9188,N_7647,N_8096);
and U9189 (N_9189,N_8721,N_8724);
nor U9190 (N_9190,N_8757,N_8956);
nand U9191 (N_9191,N_8582,N_8404);
nand U9192 (N_9192,N_8675,N_8599);
nand U9193 (N_9193,N_7578,N_7940);
or U9194 (N_9194,N_8030,N_8438);
nand U9195 (N_9195,N_8110,N_8820);
or U9196 (N_9196,N_7738,N_7546);
or U9197 (N_9197,N_7757,N_8206);
and U9198 (N_9198,N_8583,N_8674);
nor U9199 (N_9199,N_8066,N_8909);
and U9200 (N_9200,N_8953,N_8355);
and U9201 (N_9201,N_7907,N_7806);
and U9202 (N_9202,N_7962,N_8499);
or U9203 (N_9203,N_7507,N_8959);
nor U9204 (N_9204,N_8190,N_8529);
nand U9205 (N_9205,N_8288,N_8210);
xnor U9206 (N_9206,N_7983,N_7775);
or U9207 (N_9207,N_8666,N_8373);
nor U9208 (N_9208,N_8839,N_7862);
and U9209 (N_9209,N_8869,N_8081);
nand U9210 (N_9210,N_7876,N_8380);
or U9211 (N_9211,N_7782,N_7818);
nand U9212 (N_9212,N_7676,N_8723);
nand U9213 (N_9213,N_8465,N_8864);
nor U9214 (N_9214,N_8365,N_8413);
nand U9215 (N_9215,N_8648,N_8712);
and U9216 (N_9216,N_8736,N_8141);
and U9217 (N_9217,N_8795,N_7677);
and U9218 (N_9218,N_8528,N_7966);
or U9219 (N_9219,N_8751,N_8671);
or U9220 (N_9220,N_8596,N_8323);
or U9221 (N_9221,N_8439,N_8276);
or U9222 (N_9222,N_8023,N_7949);
or U9223 (N_9223,N_7622,N_7964);
or U9224 (N_9224,N_8530,N_7770);
nor U9225 (N_9225,N_7648,N_8568);
nor U9226 (N_9226,N_8882,N_7504);
and U9227 (N_9227,N_8035,N_8627);
nand U9228 (N_9228,N_8579,N_7552);
or U9229 (N_9229,N_8047,N_8733);
nor U9230 (N_9230,N_7837,N_7845);
nor U9231 (N_9231,N_8921,N_8272);
nand U9232 (N_9232,N_7863,N_8398);
or U9233 (N_9233,N_7868,N_8107);
nand U9234 (N_9234,N_8189,N_7903);
or U9235 (N_9235,N_8406,N_7569);
nor U9236 (N_9236,N_8878,N_8232);
nor U9237 (N_9237,N_8930,N_8961);
nand U9238 (N_9238,N_8114,N_8487);
nand U9239 (N_9239,N_8203,N_8130);
nand U9240 (N_9240,N_8670,N_7509);
nand U9241 (N_9241,N_7664,N_8083);
or U9242 (N_9242,N_7998,N_8872);
or U9243 (N_9243,N_8693,N_8507);
and U9244 (N_9244,N_8963,N_7611);
and U9245 (N_9245,N_8896,N_7609);
or U9246 (N_9246,N_8350,N_8136);
and U9247 (N_9247,N_8590,N_8493);
nand U9248 (N_9248,N_7973,N_8986);
and U9249 (N_9249,N_7744,N_8196);
nor U9250 (N_9250,N_8287,N_8488);
nand U9251 (N_9251,N_8034,N_7718);
nand U9252 (N_9252,N_7997,N_7976);
nand U9253 (N_9253,N_8201,N_7821);
nor U9254 (N_9254,N_7809,N_8473);
and U9255 (N_9255,N_7760,N_8367);
nor U9256 (N_9256,N_8958,N_7801);
nor U9257 (N_9257,N_7729,N_8092);
or U9258 (N_9258,N_8760,N_8659);
nor U9259 (N_9259,N_8656,N_8251);
and U9260 (N_9260,N_8880,N_8145);
and U9261 (N_9261,N_7703,N_7758);
or U9262 (N_9262,N_8895,N_7616);
nor U9263 (N_9263,N_8932,N_8993);
nor U9264 (N_9264,N_8527,N_8687);
or U9265 (N_9265,N_7957,N_8453);
and U9266 (N_9266,N_8551,N_7551);
nor U9267 (N_9267,N_7795,N_7685);
nand U9268 (N_9268,N_8140,N_8412);
nor U9269 (N_9269,N_7500,N_8040);
nand U9270 (N_9270,N_7538,N_8467);
or U9271 (N_9271,N_7882,N_8676);
and U9272 (N_9272,N_7714,N_7925);
and U9273 (N_9273,N_8423,N_8052);
nand U9274 (N_9274,N_8525,N_8463);
xor U9275 (N_9275,N_7943,N_7901);
or U9276 (N_9276,N_8798,N_7879);
or U9277 (N_9277,N_7740,N_7645);
nor U9278 (N_9278,N_8180,N_8940);
nor U9279 (N_9279,N_7946,N_7713);
and U9280 (N_9280,N_8894,N_7680);
nor U9281 (N_9281,N_8595,N_7536);
or U9282 (N_9282,N_7603,N_8492);
and U9283 (N_9283,N_7810,N_7939);
nand U9284 (N_9284,N_8824,N_8770);
nor U9285 (N_9285,N_8007,N_7584);
nor U9286 (N_9286,N_7833,N_8029);
or U9287 (N_9287,N_7594,N_8112);
or U9288 (N_9288,N_8732,N_7908);
nand U9289 (N_9289,N_8657,N_8851);
nor U9290 (N_9290,N_7888,N_7719);
xor U9291 (N_9291,N_8574,N_8336);
nand U9292 (N_9292,N_8078,N_7601);
and U9293 (N_9293,N_8572,N_8902);
nand U9294 (N_9294,N_8987,N_8747);
nand U9295 (N_9295,N_8191,N_8445);
xor U9296 (N_9296,N_8672,N_7731);
and U9297 (N_9297,N_8051,N_8036);
nor U9298 (N_9298,N_7699,N_8856);
nand U9299 (N_9299,N_8334,N_8165);
or U9300 (N_9300,N_8998,N_8804);
or U9301 (N_9301,N_7927,N_7853);
and U9302 (N_9302,N_8802,N_8964);
and U9303 (N_9303,N_8099,N_8791);
nand U9304 (N_9304,N_7978,N_8117);
or U9305 (N_9305,N_7938,N_8873);
or U9306 (N_9306,N_7777,N_8500);
or U9307 (N_9307,N_7985,N_8749);
or U9308 (N_9308,N_8447,N_8294);
or U9309 (N_9309,N_8702,N_8597);
or U9310 (N_9310,N_8630,N_8631);
nand U9311 (N_9311,N_8661,N_8424);
nand U9312 (N_9312,N_8652,N_7589);
and U9313 (N_9313,N_7869,N_8501);
or U9314 (N_9314,N_8618,N_8840);
nand U9315 (N_9315,N_8227,N_8945);
and U9316 (N_9316,N_8256,N_8848);
and U9317 (N_9317,N_8303,N_8719);
or U9318 (N_9318,N_7746,N_8061);
or U9319 (N_9319,N_7961,N_8917);
or U9320 (N_9320,N_8729,N_8637);
nor U9321 (N_9321,N_7674,N_7576);
nand U9322 (N_9322,N_8269,N_7670);
nand U9323 (N_9323,N_8612,N_8805);
or U9324 (N_9324,N_8260,N_7861);
and U9325 (N_9325,N_8460,N_8489);
nand U9326 (N_9326,N_8965,N_7671);
or U9327 (N_9327,N_8989,N_7568);
and U9328 (N_9328,N_8833,N_8806);
nor U9329 (N_9329,N_7924,N_8418);
nor U9330 (N_9330,N_8010,N_8542);
or U9331 (N_9331,N_8511,N_8347);
or U9332 (N_9332,N_8234,N_8067);
nor U9333 (N_9333,N_8495,N_8298);
nand U9334 (N_9334,N_7887,N_7711);
nand U9335 (N_9335,N_7581,N_7988);
nor U9336 (N_9336,N_8970,N_8090);
nor U9337 (N_9337,N_7690,N_8240);
xor U9338 (N_9338,N_8262,N_8435);
nor U9339 (N_9339,N_8148,N_7636);
or U9340 (N_9340,N_7811,N_8846);
or U9341 (N_9341,N_7535,N_8417);
or U9342 (N_9342,N_7741,N_7725);
nand U9343 (N_9343,N_7994,N_8892);
nand U9344 (N_9344,N_7528,N_7771);
nand U9345 (N_9345,N_7524,N_8513);
xnor U9346 (N_9346,N_8984,N_8957);
or U9347 (N_9347,N_8766,N_8651);
nand U9348 (N_9348,N_8261,N_8273);
nor U9349 (N_9349,N_7658,N_7951);
nor U9350 (N_9350,N_8170,N_8575);
or U9351 (N_9351,N_7686,N_8850);
xnor U9352 (N_9352,N_8742,N_8936);
nand U9353 (N_9353,N_8539,N_7540);
nor U9354 (N_9354,N_8329,N_8573);
nand U9355 (N_9355,N_8169,N_7517);
and U9356 (N_9356,N_8295,N_8345);
nor U9357 (N_9357,N_8718,N_7683);
or U9358 (N_9358,N_8000,N_7547);
nor U9359 (N_9359,N_7781,N_8646);
nor U9360 (N_9360,N_7505,N_8003);
and U9361 (N_9361,N_8988,N_8370);
and U9362 (N_9362,N_8062,N_7900);
nor U9363 (N_9363,N_7986,N_8701);
or U9364 (N_9364,N_8055,N_8059);
or U9365 (N_9365,N_8339,N_7992);
nand U9366 (N_9366,N_7914,N_8585);
or U9367 (N_9367,N_7835,N_7716);
and U9368 (N_9368,N_8363,N_8769);
nand U9369 (N_9369,N_7893,N_8346);
xor U9370 (N_9370,N_8890,N_8827);
nor U9371 (N_9371,N_7854,N_8545);
nor U9372 (N_9372,N_7767,N_7651);
and U9373 (N_9373,N_8915,N_8122);
nand U9374 (N_9374,N_8972,N_8537);
and U9375 (N_9375,N_8952,N_7608);
nand U9376 (N_9376,N_7971,N_7906);
nand U9377 (N_9377,N_7672,N_8617);
xnor U9378 (N_9378,N_7639,N_8451);
or U9379 (N_9379,N_7727,N_8569);
nand U9380 (N_9380,N_8809,N_8381);
nor U9381 (N_9381,N_8819,N_8600);
nor U9382 (N_9382,N_8432,N_8048);
nor U9383 (N_9383,N_8520,N_8320);
nor U9384 (N_9384,N_7788,N_8143);
or U9385 (N_9385,N_7944,N_8973);
nand U9386 (N_9386,N_8259,N_7586);
nor U9387 (N_9387,N_7501,N_8308);
nor U9388 (N_9388,N_7735,N_8610);
nand U9389 (N_9389,N_8475,N_8402);
nor U9390 (N_9390,N_7619,N_8606);
or U9391 (N_9391,N_7933,N_7792);
and U9392 (N_9392,N_8706,N_7743);
or U9393 (N_9393,N_8215,N_7702);
and U9394 (N_9394,N_8772,N_8385);
nor U9395 (N_9395,N_8102,N_8064);
and U9396 (N_9396,N_8309,N_8857);
xnor U9397 (N_9397,N_7894,N_8741);
nor U9398 (N_9398,N_7787,N_8265);
and U9399 (N_9399,N_7922,N_7634);
xor U9400 (N_9400,N_8591,N_8153);
and U9401 (N_9401,N_7928,N_8816);
nand U9402 (N_9402,N_8002,N_7673);
and U9403 (N_9403,N_8508,N_8847);
and U9404 (N_9404,N_7867,N_8934);
nor U9405 (N_9405,N_7600,N_8360);
nand U9406 (N_9406,N_8645,N_8845);
nor U9407 (N_9407,N_8366,N_8523);
nand U9408 (N_9408,N_8164,N_8119);
nor U9409 (N_9409,N_8400,N_8700);
nor U9410 (N_9410,N_8901,N_8726);
nand U9411 (N_9411,N_7595,N_8361);
or U9412 (N_9412,N_8516,N_7669);
nor U9413 (N_9413,N_8778,N_8941);
nor U9414 (N_9414,N_8877,N_7800);
nand U9415 (N_9415,N_8080,N_7808);
nand U9416 (N_9416,N_8302,N_8576);
xnor U9417 (N_9417,N_7963,N_7999);
nand U9418 (N_9418,N_8134,N_7917);
or U9419 (N_9419,N_8352,N_8120);
nand U9420 (N_9420,N_8415,N_8786);
and U9421 (N_9421,N_8744,N_8985);
nand U9422 (N_9422,N_8632,N_7521);
nand U9423 (N_9423,N_7969,N_8541);
nand U9424 (N_9424,N_7588,N_8450);
nand U9425 (N_9425,N_7783,N_8176);
nor U9426 (N_9426,N_8341,N_7545);
nand U9427 (N_9427,N_8920,N_8753);
nor U9428 (N_9428,N_8315,N_8665);
and U9429 (N_9429,N_8305,N_7682);
and U9430 (N_9430,N_7739,N_8205);
nand U9431 (N_9431,N_8750,N_8748);
nor U9432 (N_9432,N_8739,N_8818);
nand U9433 (N_9433,N_7874,N_7561);
nor U9434 (N_9434,N_8503,N_7709);
and U9435 (N_9435,N_7967,N_8371);
and U9436 (N_9436,N_8087,N_8391);
nor U9437 (N_9437,N_7526,N_7839);
and U9438 (N_9438,N_7706,N_7661);
and U9439 (N_9439,N_8084,N_8124);
nor U9440 (N_9440,N_8992,N_7979);
and U9441 (N_9441,N_8655,N_8146);
nor U9442 (N_9442,N_7587,N_8436);
nor U9443 (N_9443,N_8695,N_8161);
and U9444 (N_9444,N_8592,N_7913);
and U9445 (N_9445,N_7512,N_7959);
and U9446 (N_9446,N_8133,N_8561);
nand U9447 (N_9447,N_8267,N_7556);
nor U9448 (N_9448,N_7937,N_7708);
nand U9449 (N_9449,N_8593,N_8100);
or U9450 (N_9450,N_8484,N_7919);
nand U9451 (N_9451,N_8420,N_8318);
nor U9452 (N_9452,N_7583,N_7667);
nand U9453 (N_9453,N_8565,N_8121);
and U9454 (N_9454,N_7580,N_7656);
and U9455 (N_9455,N_8544,N_8506);
nor U9456 (N_9456,N_8937,N_8560);
or U9457 (N_9457,N_7668,N_7533);
and U9458 (N_9458,N_7653,N_8884);
or U9459 (N_9459,N_7871,N_8907);
and U9460 (N_9460,N_8641,N_8195);
nand U9461 (N_9461,N_7663,N_8927);
nor U9462 (N_9462,N_7518,N_8231);
or U9463 (N_9463,N_8095,N_8841);
and U9464 (N_9464,N_8478,N_8730);
and U9465 (N_9465,N_7555,N_8960);
or U9466 (N_9466,N_8980,N_7849);
nand U9467 (N_9467,N_7558,N_7797);
nand U9468 (N_9468,N_8947,N_8086);
nor U9469 (N_9469,N_8621,N_8540);
nand U9470 (N_9470,N_7794,N_7572);
nand U9471 (N_9471,N_8354,N_8224);
or U9472 (N_9472,N_8001,N_8497);
nand U9473 (N_9473,N_7649,N_8113);
and U9474 (N_9474,N_7571,N_8472);
nand U9475 (N_9475,N_7761,N_8217);
and U9476 (N_9476,N_7764,N_8773);
and U9477 (N_9477,N_8181,N_7707);
nand U9478 (N_9478,N_8063,N_8623);
or U9479 (N_9479,N_7694,N_8150);
nor U9480 (N_9480,N_7617,N_8682);
or U9481 (N_9481,N_8039,N_8628);
nor U9482 (N_9482,N_8625,N_8395);
nand U9483 (N_9483,N_8013,N_7503);
nand U9484 (N_9484,N_8755,N_7816);
and U9485 (N_9485,N_8982,N_7926);
nor U9486 (N_9486,N_8887,N_8416);
or U9487 (N_9487,N_8521,N_8016);
nor U9488 (N_9488,N_7548,N_8870);
and U9489 (N_9489,N_8045,N_8650);
nand U9490 (N_9490,N_8019,N_8990);
or U9491 (N_9491,N_7520,N_7885);
nand U9492 (N_9492,N_8533,N_8286);
or U9493 (N_9493,N_7784,N_8725);
nand U9494 (N_9494,N_7930,N_7629);
nor U9495 (N_9495,N_7724,N_8662);
nor U9496 (N_9496,N_7643,N_8979);
nor U9497 (N_9497,N_8397,N_8933);
and U9498 (N_9498,N_8931,N_8098);
or U9499 (N_9499,N_8571,N_8912);
nor U9500 (N_9500,N_8837,N_8680);
nand U9501 (N_9501,N_7541,N_7710);
xnor U9502 (N_9502,N_8057,N_8852);
and U9503 (N_9503,N_8629,N_8219);
or U9504 (N_9504,N_7972,N_8991);
nand U9505 (N_9505,N_8043,N_8155);
nand U9506 (N_9506,N_8138,N_8393);
nor U9507 (N_9507,N_7752,N_7768);
or U9508 (N_9508,N_8904,N_8075);
nor U9509 (N_9509,N_8550,N_8425);
nor U9510 (N_9510,N_8761,N_8326);
nand U9511 (N_9511,N_8874,N_8558);
nor U9512 (N_9512,N_8342,N_7895);
nor U9513 (N_9513,N_7898,N_8889);
or U9514 (N_9514,N_8028,N_8728);
nand U9515 (N_9515,N_8974,N_8531);
nor U9516 (N_9516,N_7870,N_8216);
and U9517 (N_9517,N_7773,N_8636);
nand U9518 (N_9518,N_8317,N_7796);
nor U9519 (N_9519,N_8587,N_7834);
or U9520 (N_9520,N_8324,N_8293);
nand U9521 (N_9521,N_8250,N_8633);
and U9522 (N_9522,N_7841,N_7909);
nand U9523 (N_9523,N_8640,N_7832);
or U9524 (N_9524,N_8939,N_8327);
xor U9525 (N_9525,N_7769,N_8456);
or U9526 (N_9526,N_7689,N_8768);
or U9527 (N_9527,N_8314,N_8871);
or U9528 (N_9528,N_7726,N_8686);
nor U9529 (N_9529,N_8913,N_8443);
nor U9530 (N_9530,N_7948,N_7542);
and U9531 (N_9531,N_8696,N_7579);
or U9532 (N_9532,N_7635,N_8971);
or U9533 (N_9533,N_8167,N_8792);
and U9534 (N_9534,N_7566,N_7778);
nand U9535 (N_9535,N_8072,N_8842);
or U9536 (N_9536,N_8106,N_8359);
or U9537 (N_9537,N_8236,N_8619);
or U9538 (N_9538,N_8614,N_8821);
and U9539 (N_9539,N_8356,N_7991);
or U9540 (N_9540,N_8745,N_8386);
nor U9541 (N_9541,N_7734,N_7899);
or U9542 (N_9542,N_8038,N_8535);
xnor U9543 (N_9543,N_8376,N_8483);
and U9544 (N_9544,N_7610,N_8570);
or U9545 (N_9545,N_8223,N_8454);
or U9546 (N_9546,N_8166,N_7550);
and U9547 (N_9547,N_7655,N_8348);
nor U9548 (N_9548,N_7952,N_8862);
nor U9549 (N_9549,N_7618,N_8073);
nor U9550 (N_9550,N_8710,N_7549);
nand U9551 (N_9551,N_8881,N_8017);
nor U9552 (N_9552,N_8943,N_7684);
and U9553 (N_9553,N_8609,N_7865);
nand U9554 (N_9554,N_8049,N_8248);
nor U9555 (N_9555,N_8103,N_8644);
nand U9556 (N_9556,N_8654,N_8801);
nor U9557 (N_9557,N_8144,N_8368);
and U9558 (N_9558,N_8479,N_8754);
and U9559 (N_9559,N_8734,N_8135);
and U9560 (N_9560,N_8209,N_8758);
or U9561 (N_9561,N_8278,N_7641);
nand U9562 (N_9562,N_8174,N_7831);
nand U9563 (N_9563,N_8983,N_8844);
nor U9564 (N_9564,N_8977,N_8300);
or U9565 (N_9565,N_7830,N_8781);
and U9566 (N_9566,N_8898,N_8151);
nand U9567 (N_9567,N_7779,N_8639);
nor U9568 (N_9568,N_8274,N_8997);
nand U9569 (N_9569,N_7531,N_7598);
and U9570 (N_9570,N_7850,N_7889);
nor U9571 (N_9571,N_8604,N_8291);
nand U9572 (N_9572,N_8708,N_7823);
and U9573 (N_9573,N_7666,N_7742);
or U9574 (N_9574,N_8433,N_7955);
and U9575 (N_9575,N_7704,N_8552);
nor U9576 (N_9576,N_7662,N_8154);
or U9577 (N_9577,N_7817,N_8214);
nand U9578 (N_9578,N_8929,N_8951);
nor U9579 (N_9579,N_8024,N_8731);
and U9580 (N_9580,N_8044,N_8183);
or U9581 (N_9581,N_7891,N_7632);
nand U9582 (N_9582,N_8635,N_8482);
nor U9583 (N_9583,N_7974,N_8509);
nand U9584 (N_9584,N_8782,N_8025);
and U9585 (N_9585,N_8613,N_8188);
nand U9586 (N_9586,N_8353,N_7688);
nor U9587 (N_9587,N_8068,N_8832);
or U9588 (N_9588,N_8763,N_8246);
nand U9589 (N_9589,N_7574,N_7519);
and U9590 (N_9590,N_7530,N_8139);
and U9591 (N_9591,N_8403,N_8384);
or U9592 (N_9592,N_7567,N_7628);
and U9593 (N_9593,N_7805,N_8321);
or U9594 (N_9594,N_8547,N_7892);
nor U9595 (N_9595,N_8476,N_7786);
nor U9596 (N_9596,N_8459,N_8328);
or U9597 (N_9597,N_7936,N_8407);
nor U9598 (N_9598,N_7872,N_7912);
and U9599 (N_9599,N_8319,N_8642);
nor U9600 (N_9600,N_8306,N_8800);
nor U9601 (N_9601,N_8976,N_7776);
or U9602 (N_9602,N_8689,N_8828);
or U9603 (N_9603,N_7506,N_8626);
nor U9604 (N_9604,N_7890,N_8213);
nor U9605 (N_9605,N_7511,N_8555);
nor U9606 (N_9606,N_7759,N_8245);
nor U9607 (N_9607,N_8396,N_8703);
nor U9608 (N_9608,N_8679,N_8012);
nand U9609 (N_9609,N_7502,N_7791);
nor U9610 (N_9610,N_7675,N_8408);
or U9611 (N_9611,N_7748,N_8942);
or U9612 (N_9612,N_8338,N_7947);
and U9613 (N_9613,N_8496,N_8803);
and U9614 (N_9614,N_7931,N_8088);
and U9615 (N_9615,N_8266,N_8263);
nor U9616 (N_9616,N_8221,N_7838);
nor U9617 (N_9617,N_8549,N_8660);
and U9618 (N_9618,N_8787,N_8536);
nor U9619 (N_9619,N_8428,N_8026);
nor U9620 (N_9620,N_8697,N_7921);
or U9621 (N_9621,N_7765,N_8243);
nand U9622 (N_9622,N_8108,N_7615);
nor U9623 (N_9623,N_8027,N_8257);
and U9624 (N_9624,N_8893,N_7750);
or U9625 (N_9625,N_8638,N_7844);
or U9626 (N_9626,N_8622,N_7987);
and U9627 (N_9627,N_7842,N_8865);
nor U9628 (N_9628,N_7920,N_8740);
nand U9629 (N_9629,N_8008,N_8668);
nand U9630 (N_9630,N_7596,N_8077);
nor U9631 (N_9631,N_8193,N_8409);
nor U9632 (N_9632,N_7638,N_8594);
or U9633 (N_9633,N_8715,N_8093);
and U9634 (N_9634,N_8866,N_8241);
and U9635 (N_9635,N_8586,N_8853);
nand U9636 (N_9636,N_8310,N_8358);
or U9637 (N_9637,N_7659,N_8711);
nand U9638 (N_9638,N_7934,N_8014);
nor U9639 (N_9639,N_8275,N_8829);
nand U9640 (N_9640,N_7557,N_8390);
and U9641 (N_9641,N_7762,N_8156);
nor U9642 (N_9642,N_7627,N_7970);
or U9643 (N_9643,N_8405,N_8111);
nand U9644 (N_9644,N_7945,N_7932);
nand U9645 (N_9645,N_7715,N_8888);
nand U9646 (N_9646,N_7923,N_8694);
nand U9647 (N_9647,N_8789,N_7625);
or U9648 (N_9648,N_8242,N_7774);
and U9649 (N_9649,N_8222,N_8905);
nand U9650 (N_9650,N_7623,N_8349);
nand U9651 (N_9651,N_8244,N_8999);
nand U9652 (N_9652,N_8788,N_7606);
or U9653 (N_9653,N_8207,N_7807);
or U9654 (N_9654,N_8313,N_8018);
and U9655 (N_9655,N_8184,N_8822);
or U9656 (N_9656,N_8228,N_8247);
and U9657 (N_9657,N_8204,N_8457);
nor U9658 (N_9658,N_7646,N_8152);
nand U9659 (N_9659,N_7829,N_7989);
and U9660 (N_9660,N_8285,N_8168);
nor U9661 (N_9661,N_8678,N_8738);
or U9662 (N_9662,N_7562,N_7877);
and U9663 (N_9663,N_8764,N_8229);
nor U9664 (N_9664,N_7543,N_7858);
and U9665 (N_9665,N_7745,N_8494);
nor U9666 (N_9666,N_7918,N_7860);
and U9667 (N_9667,N_8608,N_7701);
nand U9668 (N_9668,N_8634,N_8900);
nor U9669 (N_9669,N_8563,N_8667);
nand U9670 (N_9670,N_7828,N_8709);
nand U9671 (N_9671,N_8427,N_8137);
nand U9672 (N_9672,N_8271,N_8344);
or U9673 (N_9673,N_8377,N_8780);
or U9674 (N_9674,N_7804,N_8005);
nor U9675 (N_9675,N_8705,N_7911);
nor U9676 (N_9676,N_7525,N_8823);
and U9677 (N_9677,N_7996,N_8208);
and U9678 (N_9678,N_8836,N_8268);
nand U9679 (N_9679,N_8378,N_7954);
nand U9680 (N_9680,N_8858,N_8691);
nand U9681 (N_9681,N_8442,N_8688);
nor U9682 (N_9682,N_8331,N_7995);
or U9683 (N_9683,N_8440,N_8441);
or U9684 (N_9684,N_8722,N_7878);
xnor U9685 (N_9685,N_8504,N_8410);
or U9686 (N_9686,N_8897,N_8175);
xor U9687 (N_9687,N_7803,N_8414);
nor U9688 (N_9688,N_8826,N_7614);
nand U9689 (N_9689,N_8737,N_7721);
nor U9690 (N_9690,N_8011,N_8449);
and U9691 (N_9691,N_7693,N_8502);
or U9692 (N_9692,N_7652,N_8692);
and U9693 (N_9693,N_7785,N_7698);
nand U9694 (N_9694,N_7660,N_8861);
nor U9695 (N_9695,N_7875,N_7532);
or U9696 (N_9696,N_7631,N_8981);
and U9697 (N_9697,N_8279,N_7965);
or U9698 (N_9698,N_8226,N_8434);
nor U9699 (N_9699,N_7902,N_8620);
nor U9700 (N_9700,N_8553,N_8233);
nor U9701 (N_9701,N_8588,N_8698);
and U9702 (N_9702,N_8394,N_7510);
and U9703 (N_9703,N_8602,N_8876);
nor U9704 (N_9704,N_8056,N_8172);
nor U9705 (N_9705,N_8925,N_7747);
nand U9706 (N_9706,N_7720,N_8290);
nand U9707 (N_9707,N_8104,N_7692);
and U9708 (N_9708,N_8419,N_8891);
nor U9709 (N_9709,N_8015,N_7751);
or U9710 (N_9710,N_8611,N_7756);
and U9711 (N_9711,N_7982,N_8004);
nand U9712 (N_9712,N_8281,N_8924);
nor U9713 (N_9713,N_8280,N_8458);
or U9714 (N_9714,N_7820,N_7612);
xor U9715 (N_9715,N_7852,N_8886);
nor U9716 (N_9716,N_8526,N_8785);
or U9717 (N_9717,N_7960,N_8477);
nand U9718 (N_9718,N_8777,N_8283);
nand U9719 (N_9719,N_8179,N_8684);
and U9720 (N_9720,N_7640,N_8762);
nand U9721 (N_9721,N_8607,N_8307);
nor U9722 (N_9722,N_8815,N_7935);
and U9723 (N_9723,N_7604,N_7620);
or U9724 (N_9724,N_8033,N_8903);
nand U9725 (N_9725,N_7864,N_8928);
and U9726 (N_9726,N_7705,N_8677);
nand U9727 (N_9727,N_7753,N_8779);
or U9728 (N_9728,N_7565,N_7772);
nor U9729 (N_9729,N_8923,N_8264);
or U9730 (N_9730,N_7905,N_8746);
and U9731 (N_9731,N_7915,N_8566);
or U9732 (N_9732,N_8849,N_7657);
and U9733 (N_9733,N_7544,N_8337);
nand U9734 (N_9734,N_8906,N_7591);
or U9735 (N_9735,N_7825,N_8157);
nor U9736 (N_9736,N_8470,N_8065);
nand U9737 (N_9737,N_7855,N_8735);
nand U9738 (N_9738,N_8239,N_8060);
nand U9739 (N_9739,N_7958,N_7736);
nor U9740 (N_9740,N_7793,N_8101);
nand U9741 (N_9741,N_8704,N_7766);
or U9742 (N_9742,N_8289,N_7613);
nor U9743 (N_9743,N_8480,N_8714);
or U9744 (N_9744,N_7790,N_8948);
nor U9745 (N_9745,N_8147,N_8669);
and U9746 (N_9746,N_8021,N_8717);
and U9747 (N_9747,N_7968,N_8125);
and U9748 (N_9748,N_8311,N_7843);
nand U9749 (N_9749,N_8197,N_8967);
or U9750 (N_9750,N_7696,N_8360);
nor U9751 (N_9751,N_8916,N_7965);
or U9752 (N_9752,N_8998,N_8929);
nor U9753 (N_9753,N_8608,N_7531);
and U9754 (N_9754,N_8124,N_7984);
nor U9755 (N_9755,N_7689,N_7538);
or U9756 (N_9756,N_8207,N_7655);
nand U9757 (N_9757,N_8961,N_8906);
or U9758 (N_9758,N_8753,N_8506);
nand U9759 (N_9759,N_8635,N_7961);
nor U9760 (N_9760,N_8488,N_7710);
nand U9761 (N_9761,N_8297,N_8184);
nor U9762 (N_9762,N_8285,N_8121);
nand U9763 (N_9763,N_8825,N_7770);
and U9764 (N_9764,N_8879,N_8154);
nand U9765 (N_9765,N_8114,N_8833);
nor U9766 (N_9766,N_7747,N_7764);
nor U9767 (N_9767,N_7664,N_7558);
or U9768 (N_9768,N_7583,N_7570);
nand U9769 (N_9769,N_8239,N_8434);
xor U9770 (N_9770,N_8079,N_7504);
or U9771 (N_9771,N_8466,N_8357);
and U9772 (N_9772,N_8785,N_8515);
or U9773 (N_9773,N_8386,N_8738);
or U9774 (N_9774,N_7939,N_8450);
or U9775 (N_9775,N_8717,N_8755);
nor U9776 (N_9776,N_7917,N_8225);
or U9777 (N_9777,N_8126,N_8724);
nand U9778 (N_9778,N_7745,N_8808);
and U9779 (N_9779,N_8972,N_8062);
nor U9780 (N_9780,N_8877,N_8974);
xnor U9781 (N_9781,N_7540,N_8443);
and U9782 (N_9782,N_7705,N_8754);
nand U9783 (N_9783,N_8252,N_8830);
nand U9784 (N_9784,N_8879,N_7548);
nor U9785 (N_9785,N_8217,N_7523);
nand U9786 (N_9786,N_8907,N_8112);
and U9787 (N_9787,N_8205,N_8102);
nor U9788 (N_9788,N_8492,N_7643);
nor U9789 (N_9789,N_8956,N_7537);
or U9790 (N_9790,N_8165,N_8785);
or U9791 (N_9791,N_7504,N_7995);
nand U9792 (N_9792,N_7993,N_8074);
nor U9793 (N_9793,N_8819,N_7561);
nor U9794 (N_9794,N_8283,N_8613);
nor U9795 (N_9795,N_8090,N_8231);
and U9796 (N_9796,N_7631,N_7791);
and U9797 (N_9797,N_7616,N_7966);
or U9798 (N_9798,N_8525,N_7881);
nor U9799 (N_9799,N_8352,N_8597);
nand U9800 (N_9800,N_8722,N_8981);
and U9801 (N_9801,N_8209,N_7691);
nand U9802 (N_9802,N_7904,N_7925);
or U9803 (N_9803,N_7794,N_8110);
nand U9804 (N_9804,N_7781,N_8799);
nand U9805 (N_9805,N_8841,N_7880);
and U9806 (N_9806,N_8209,N_7575);
nand U9807 (N_9807,N_8007,N_7653);
or U9808 (N_9808,N_8090,N_8963);
nand U9809 (N_9809,N_7930,N_7745);
or U9810 (N_9810,N_7584,N_8241);
and U9811 (N_9811,N_7758,N_7787);
nor U9812 (N_9812,N_8445,N_8294);
nand U9813 (N_9813,N_8582,N_8767);
nand U9814 (N_9814,N_8785,N_8978);
or U9815 (N_9815,N_8241,N_8228);
nand U9816 (N_9816,N_8956,N_8423);
and U9817 (N_9817,N_8392,N_7899);
nand U9818 (N_9818,N_8301,N_8800);
nand U9819 (N_9819,N_8498,N_8205);
and U9820 (N_9820,N_7722,N_8649);
or U9821 (N_9821,N_8635,N_8905);
nand U9822 (N_9822,N_8334,N_8293);
or U9823 (N_9823,N_7533,N_7652);
nor U9824 (N_9824,N_8600,N_8394);
and U9825 (N_9825,N_8841,N_8654);
nand U9826 (N_9826,N_7543,N_8479);
nor U9827 (N_9827,N_7884,N_7971);
and U9828 (N_9828,N_8803,N_8661);
nand U9829 (N_9829,N_7868,N_8710);
nand U9830 (N_9830,N_7721,N_7734);
or U9831 (N_9831,N_8615,N_8467);
and U9832 (N_9832,N_8575,N_8295);
nor U9833 (N_9833,N_8758,N_7740);
and U9834 (N_9834,N_8576,N_7632);
or U9835 (N_9835,N_7649,N_8800);
and U9836 (N_9836,N_7978,N_8037);
and U9837 (N_9837,N_8985,N_8704);
nor U9838 (N_9838,N_8820,N_8688);
nor U9839 (N_9839,N_7792,N_7898);
nand U9840 (N_9840,N_8815,N_8989);
or U9841 (N_9841,N_8236,N_7898);
nand U9842 (N_9842,N_8997,N_8804);
and U9843 (N_9843,N_8994,N_7931);
or U9844 (N_9844,N_7808,N_7828);
and U9845 (N_9845,N_8004,N_7543);
nor U9846 (N_9846,N_8056,N_7745);
or U9847 (N_9847,N_8551,N_8460);
or U9848 (N_9848,N_8399,N_7803);
nor U9849 (N_9849,N_8149,N_8659);
nor U9850 (N_9850,N_8670,N_8260);
and U9851 (N_9851,N_8611,N_7504);
nand U9852 (N_9852,N_8232,N_8602);
xnor U9853 (N_9853,N_8782,N_7988);
and U9854 (N_9854,N_8117,N_8075);
nor U9855 (N_9855,N_8380,N_7909);
nor U9856 (N_9856,N_7709,N_8530);
and U9857 (N_9857,N_8009,N_8457);
nand U9858 (N_9858,N_8433,N_8599);
or U9859 (N_9859,N_8185,N_8933);
nor U9860 (N_9860,N_7697,N_8863);
nand U9861 (N_9861,N_8384,N_8837);
nand U9862 (N_9862,N_8106,N_8083);
or U9863 (N_9863,N_8666,N_8015);
nor U9864 (N_9864,N_7888,N_8445);
or U9865 (N_9865,N_7607,N_7828);
and U9866 (N_9866,N_7683,N_7999);
and U9867 (N_9867,N_7989,N_7796);
and U9868 (N_9868,N_8921,N_8007);
nand U9869 (N_9869,N_8628,N_7845);
xnor U9870 (N_9870,N_7705,N_8691);
nand U9871 (N_9871,N_8267,N_8182);
or U9872 (N_9872,N_8916,N_7512);
or U9873 (N_9873,N_8112,N_8461);
nor U9874 (N_9874,N_8576,N_7867);
or U9875 (N_9875,N_8302,N_7654);
or U9876 (N_9876,N_8181,N_8454);
nand U9877 (N_9877,N_8442,N_7636);
nor U9878 (N_9878,N_7821,N_7928);
nor U9879 (N_9879,N_7939,N_8593);
or U9880 (N_9880,N_8228,N_7526);
nand U9881 (N_9881,N_7541,N_8214);
or U9882 (N_9882,N_8663,N_7703);
or U9883 (N_9883,N_8047,N_8623);
or U9884 (N_9884,N_8920,N_8386);
nor U9885 (N_9885,N_8132,N_8824);
or U9886 (N_9886,N_7885,N_7617);
nor U9887 (N_9887,N_8869,N_7595);
or U9888 (N_9888,N_8173,N_8986);
and U9889 (N_9889,N_8858,N_7611);
and U9890 (N_9890,N_7518,N_8621);
nand U9891 (N_9891,N_8766,N_8577);
and U9892 (N_9892,N_8007,N_7716);
or U9893 (N_9893,N_8998,N_7638);
and U9894 (N_9894,N_8446,N_7748);
or U9895 (N_9895,N_8596,N_8679);
nor U9896 (N_9896,N_8970,N_8140);
nor U9897 (N_9897,N_8971,N_8789);
and U9898 (N_9898,N_7584,N_7867);
xnor U9899 (N_9899,N_7517,N_8194);
and U9900 (N_9900,N_7727,N_8029);
nor U9901 (N_9901,N_8440,N_8782);
or U9902 (N_9902,N_8065,N_8916);
nand U9903 (N_9903,N_8543,N_8638);
nor U9904 (N_9904,N_8381,N_8378);
and U9905 (N_9905,N_7917,N_8676);
or U9906 (N_9906,N_8728,N_8965);
or U9907 (N_9907,N_8514,N_7751);
nor U9908 (N_9908,N_7549,N_7767);
or U9909 (N_9909,N_7638,N_7997);
and U9910 (N_9910,N_8564,N_7560);
or U9911 (N_9911,N_7688,N_7526);
nor U9912 (N_9912,N_8307,N_8334);
and U9913 (N_9913,N_7764,N_8830);
or U9914 (N_9914,N_8007,N_8468);
xnor U9915 (N_9915,N_8555,N_7636);
or U9916 (N_9916,N_7954,N_8666);
and U9917 (N_9917,N_8229,N_7730);
or U9918 (N_9918,N_8335,N_7764);
and U9919 (N_9919,N_7613,N_7959);
or U9920 (N_9920,N_8410,N_8616);
nor U9921 (N_9921,N_7839,N_8943);
or U9922 (N_9922,N_8289,N_7928);
or U9923 (N_9923,N_8526,N_7925);
nor U9924 (N_9924,N_8663,N_8649);
and U9925 (N_9925,N_7971,N_7907);
nor U9926 (N_9926,N_8932,N_7721);
and U9927 (N_9927,N_7817,N_7940);
or U9928 (N_9928,N_7689,N_8432);
and U9929 (N_9929,N_7805,N_7801);
nor U9930 (N_9930,N_8682,N_7988);
nor U9931 (N_9931,N_8223,N_8424);
nand U9932 (N_9932,N_8633,N_8348);
nor U9933 (N_9933,N_8783,N_8990);
nand U9934 (N_9934,N_8298,N_7907);
nor U9935 (N_9935,N_8994,N_8748);
nand U9936 (N_9936,N_8995,N_8883);
or U9937 (N_9937,N_8638,N_7977);
nand U9938 (N_9938,N_7732,N_7826);
nand U9939 (N_9939,N_8763,N_7987);
nor U9940 (N_9940,N_8956,N_7638);
and U9941 (N_9941,N_7880,N_8677);
nor U9942 (N_9942,N_8223,N_8146);
nor U9943 (N_9943,N_7714,N_8354);
and U9944 (N_9944,N_8288,N_7905);
or U9945 (N_9945,N_8948,N_7729);
xnor U9946 (N_9946,N_7941,N_8619);
and U9947 (N_9947,N_8645,N_8576);
nor U9948 (N_9948,N_8516,N_8095);
or U9949 (N_9949,N_8360,N_7932);
and U9950 (N_9950,N_8792,N_7567);
or U9951 (N_9951,N_8894,N_8313);
nor U9952 (N_9952,N_7626,N_7892);
and U9953 (N_9953,N_8538,N_8962);
or U9954 (N_9954,N_8858,N_8348);
or U9955 (N_9955,N_8368,N_8097);
and U9956 (N_9956,N_8918,N_7625);
or U9957 (N_9957,N_8178,N_8989);
nor U9958 (N_9958,N_7504,N_8626);
nand U9959 (N_9959,N_7780,N_7582);
nor U9960 (N_9960,N_7926,N_8664);
and U9961 (N_9961,N_7877,N_8478);
or U9962 (N_9962,N_8094,N_8976);
nor U9963 (N_9963,N_8221,N_8232);
nor U9964 (N_9964,N_7932,N_8996);
or U9965 (N_9965,N_8155,N_7826);
nor U9966 (N_9966,N_7631,N_7832);
and U9967 (N_9967,N_7556,N_8277);
or U9968 (N_9968,N_7768,N_7823);
or U9969 (N_9969,N_8304,N_7724);
or U9970 (N_9970,N_8006,N_8726);
and U9971 (N_9971,N_8402,N_8120);
and U9972 (N_9972,N_8395,N_8443);
and U9973 (N_9973,N_8909,N_8593);
or U9974 (N_9974,N_7823,N_8504);
or U9975 (N_9975,N_8648,N_8070);
xor U9976 (N_9976,N_7713,N_8413);
nor U9977 (N_9977,N_8220,N_8612);
and U9978 (N_9978,N_7952,N_8564);
nand U9979 (N_9979,N_8090,N_7798);
or U9980 (N_9980,N_8303,N_8885);
nor U9981 (N_9981,N_7550,N_8032);
or U9982 (N_9982,N_8354,N_7734);
or U9983 (N_9983,N_8362,N_7870);
and U9984 (N_9984,N_7690,N_8266);
nor U9985 (N_9985,N_7627,N_8932);
or U9986 (N_9986,N_8935,N_8137);
nand U9987 (N_9987,N_7925,N_8192);
nor U9988 (N_9988,N_7790,N_8463);
nor U9989 (N_9989,N_8989,N_7666);
or U9990 (N_9990,N_8793,N_8570);
or U9991 (N_9991,N_8154,N_8240);
nand U9992 (N_9992,N_8951,N_7970);
or U9993 (N_9993,N_8691,N_8481);
and U9994 (N_9994,N_7970,N_7777);
and U9995 (N_9995,N_8922,N_8697);
and U9996 (N_9996,N_7628,N_8334);
and U9997 (N_9997,N_7971,N_8789);
nor U9998 (N_9998,N_8432,N_8993);
nor U9999 (N_9999,N_8932,N_8972);
nor U10000 (N_10000,N_8904,N_7955);
nand U10001 (N_10001,N_7573,N_7963);
nor U10002 (N_10002,N_7883,N_8679);
nor U10003 (N_10003,N_8413,N_8468);
nand U10004 (N_10004,N_8437,N_8358);
xnor U10005 (N_10005,N_8223,N_8195);
or U10006 (N_10006,N_8437,N_8945);
nand U10007 (N_10007,N_7700,N_8056);
nor U10008 (N_10008,N_7983,N_7629);
nand U10009 (N_10009,N_8615,N_8892);
nor U10010 (N_10010,N_8402,N_7887);
nand U10011 (N_10011,N_7982,N_8965);
or U10012 (N_10012,N_8780,N_7997);
or U10013 (N_10013,N_8289,N_8306);
and U10014 (N_10014,N_8394,N_8483);
or U10015 (N_10015,N_8118,N_7984);
or U10016 (N_10016,N_8934,N_8567);
or U10017 (N_10017,N_8873,N_8628);
and U10018 (N_10018,N_8371,N_7505);
or U10019 (N_10019,N_7612,N_7788);
nor U10020 (N_10020,N_8445,N_8093);
or U10021 (N_10021,N_8316,N_8949);
nand U10022 (N_10022,N_7501,N_7723);
nor U10023 (N_10023,N_8114,N_7746);
or U10024 (N_10024,N_8035,N_7846);
nand U10025 (N_10025,N_8968,N_7613);
and U10026 (N_10026,N_8493,N_8380);
or U10027 (N_10027,N_7907,N_8378);
and U10028 (N_10028,N_8134,N_8152);
nor U10029 (N_10029,N_8434,N_7660);
and U10030 (N_10030,N_7635,N_8164);
nor U10031 (N_10031,N_8692,N_7900);
xor U10032 (N_10032,N_8004,N_8390);
nand U10033 (N_10033,N_8683,N_8214);
or U10034 (N_10034,N_8444,N_8755);
nand U10035 (N_10035,N_8629,N_8796);
or U10036 (N_10036,N_8094,N_8240);
nand U10037 (N_10037,N_8060,N_7597);
nand U10038 (N_10038,N_8263,N_7758);
nor U10039 (N_10039,N_8425,N_7893);
or U10040 (N_10040,N_8392,N_7650);
or U10041 (N_10041,N_7593,N_7921);
nand U10042 (N_10042,N_7972,N_8745);
nand U10043 (N_10043,N_7765,N_7786);
nor U10044 (N_10044,N_8001,N_7940);
xnor U10045 (N_10045,N_8649,N_8817);
or U10046 (N_10046,N_8250,N_7597);
or U10047 (N_10047,N_7945,N_7521);
and U10048 (N_10048,N_7778,N_8938);
or U10049 (N_10049,N_7667,N_7759);
xnor U10050 (N_10050,N_8685,N_7729);
nand U10051 (N_10051,N_8170,N_7931);
nand U10052 (N_10052,N_8306,N_7847);
and U10053 (N_10053,N_8186,N_8968);
and U10054 (N_10054,N_8183,N_7840);
nand U10055 (N_10055,N_7509,N_8385);
nor U10056 (N_10056,N_8605,N_8761);
or U10057 (N_10057,N_8782,N_7716);
or U10058 (N_10058,N_8028,N_7680);
nand U10059 (N_10059,N_8740,N_7853);
nor U10060 (N_10060,N_8689,N_8192);
nor U10061 (N_10061,N_8434,N_8066);
and U10062 (N_10062,N_8653,N_7810);
or U10063 (N_10063,N_8051,N_7980);
nor U10064 (N_10064,N_8382,N_8030);
nand U10065 (N_10065,N_7668,N_8327);
nor U10066 (N_10066,N_7554,N_8762);
nand U10067 (N_10067,N_8118,N_8134);
or U10068 (N_10068,N_8443,N_8588);
nor U10069 (N_10069,N_8425,N_7693);
and U10070 (N_10070,N_8851,N_7857);
nand U10071 (N_10071,N_8144,N_8737);
or U10072 (N_10072,N_8308,N_7744);
or U10073 (N_10073,N_8943,N_7626);
nor U10074 (N_10074,N_8841,N_8908);
or U10075 (N_10075,N_7806,N_8955);
or U10076 (N_10076,N_7846,N_7629);
nor U10077 (N_10077,N_8722,N_8400);
nand U10078 (N_10078,N_8819,N_8337);
nor U10079 (N_10079,N_8097,N_7803);
nand U10080 (N_10080,N_8472,N_7798);
nor U10081 (N_10081,N_8447,N_8206);
or U10082 (N_10082,N_8381,N_8032);
and U10083 (N_10083,N_8981,N_8516);
or U10084 (N_10084,N_8270,N_8085);
and U10085 (N_10085,N_8941,N_7530);
nand U10086 (N_10086,N_8057,N_8961);
and U10087 (N_10087,N_7743,N_7647);
nor U10088 (N_10088,N_8050,N_7666);
nand U10089 (N_10089,N_8448,N_8292);
or U10090 (N_10090,N_8242,N_8683);
nor U10091 (N_10091,N_8043,N_7673);
xnor U10092 (N_10092,N_7538,N_7579);
nor U10093 (N_10093,N_8037,N_7685);
and U10094 (N_10094,N_8241,N_8309);
or U10095 (N_10095,N_8319,N_8334);
and U10096 (N_10096,N_8058,N_7767);
nor U10097 (N_10097,N_8475,N_8567);
or U10098 (N_10098,N_8111,N_7604);
and U10099 (N_10099,N_8243,N_8329);
and U10100 (N_10100,N_7551,N_8734);
and U10101 (N_10101,N_8997,N_8448);
nand U10102 (N_10102,N_8649,N_7985);
nor U10103 (N_10103,N_8919,N_8098);
nand U10104 (N_10104,N_8921,N_8047);
or U10105 (N_10105,N_7867,N_8932);
nor U10106 (N_10106,N_7841,N_8545);
and U10107 (N_10107,N_8376,N_8029);
nand U10108 (N_10108,N_7824,N_8207);
nor U10109 (N_10109,N_8891,N_8170);
or U10110 (N_10110,N_7704,N_8204);
or U10111 (N_10111,N_8899,N_8798);
or U10112 (N_10112,N_8231,N_7940);
nor U10113 (N_10113,N_8224,N_8556);
nand U10114 (N_10114,N_8908,N_8726);
nand U10115 (N_10115,N_7920,N_8741);
nor U10116 (N_10116,N_7612,N_8657);
nor U10117 (N_10117,N_7622,N_7888);
nor U10118 (N_10118,N_7596,N_7909);
xnor U10119 (N_10119,N_8553,N_8431);
nor U10120 (N_10120,N_8623,N_8657);
nor U10121 (N_10121,N_7635,N_7632);
and U10122 (N_10122,N_7752,N_8845);
and U10123 (N_10123,N_7975,N_7890);
nand U10124 (N_10124,N_8077,N_8293);
nand U10125 (N_10125,N_8389,N_8565);
and U10126 (N_10126,N_7865,N_8737);
or U10127 (N_10127,N_8042,N_8593);
nand U10128 (N_10128,N_8444,N_7731);
nand U10129 (N_10129,N_7853,N_8875);
or U10130 (N_10130,N_8787,N_8797);
and U10131 (N_10131,N_7977,N_8066);
nand U10132 (N_10132,N_7561,N_8952);
nand U10133 (N_10133,N_7545,N_8381);
or U10134 (N_10134,N_7917,N_8604);
nand U10135 (N_10135,N_7813,N_8707);
and U10136 (N_10136,N_7966,N_8017);
nand U10137 (N_10137,N_7923,N_8254);
or U10138 (N_10138,N_8807,N_8265);
or U10139 (N_10139,N_7880,N_8312);
nor U10140 (N_10140,N_7701,N_7598);
nand U10141 (N_10141,N_7759,N_8170);
nor U10142 (N_10142,N_7866,N_8251);
nand U10143 (N_10143,N_8206,N_7727);
and U10144 (N_10144,N_7770,N_8931);
nand U10145 (N_10145,N_8679,N_8201);
and U10146 (N_10146,N_8506,N_7661);
or U10147 (N_10147,N_7645,N_7982);
or U10148 (N_10148,N_7637,N_8471);
nand U10149 (N_10149,N_7827,N_7784);
nand U10150 (N_10150,N_8823,N_8240);
xnor U10151 (N_10151,N_8440,N_7709);
or U10152 (N_10152,N_8544,N_8686);
or U10153 (N_10153,N_8964,N_8430);
nand U10154 (N_10154,N_8318,N_7566);
nor U10155 (N_10155,N_8792,N_7911);
nand U10156 (N_10156,N_8470,N_8485);
or U10157 (N_10157,N_8116,N_8786);
and U10158 (N_10158,N_8784,N_7804);
nand U10159 (N_10159,N_8099,N_8529);
or U10160 (N_10160,N_8622,N_8954);
or U10161 (N_10161,N_8775,N_8818);
nand U10162 (N_10162,N_8116,N_8602);
and U10163 (N_10163,N_8895,N_8222);
nor U10164 (N_10164,N_8491,N_7835);
nor U10165 (N_10165,N_8674,N_8439);
nand U10166 (N_10166,N_8187,N_8715);
xnor U10167 (N_10167,N_8074,N_8457);
nand U10168 (N_10168,N_8488,N_8373);
xnor U10169 (N_10169,N_7721,N_7983);
and U10170 (N_10170,N_8736,N_7886);
nand U10171 (N_10171,N_8096,N_8700);
nor U10172 (N_10172,N_7513,N_7677);
and U10173 (N_10173,N_8544,N_8646);
nand U10174 (N_10174,N_8121,N_7785);
or U10175 (N_10175,N_8527,N_8794);
or U10176 (N_10176,N_8030,N_7515);
and U10177 (N_10177,N_7541,N_8597);
and U10178 (N_10178,N_7697,N_8580);
nand U10179 (N_10179,N_8857,N_8039);
and U10180 (N_10180,N_8790,N_8605);
and U10181 (N_10181,N_7908,N_8993);
nand U10182 (N_10182,N_8707,N_7774);
or U10183 (N_10183,N_8948,N_8423);
nand U10184 (N_10184,N_8326,N_8874);
or U10185 (N_10185,N_8847,N_8410);
and U10186 (N_10186,N_7900,N_8472);
or U10187 (N_10187,N_8600,N_8249);
and U10188 (N_10188,N_8261,N_8481);
nor U10189 (N_10189,N_8443,N_8382);
nand U10190 (N_10190,N_8884,N_8705);
nand U10191 (N_10191,N_7701,N_7794);
xor U10192 (N_10192,N_8674,N_8955);
and U10193 (N_10193,N_8594,N_7573);
and U10194 (N_10194,N_7576,N_7766);
nor U10195 (N_10195,N_8037,N_7537);
or U10196 (N_10196,N_7756,N_7543);
nand U10197 (N_10197,N_7936,N_8622);
and U10198 (N_10198,N_7618,N_8158);
nand U10199 (N_10199,N_8488,N_8515);
or U10200 (N_10200,N_8581,N_8119);
nand U10201 (N_10201,N_7925,N_8928);
or U10202 (N_10202,N_8197,N_8393);
or U10203 (N_10203,N_8455,N_8521);
or U10204 (N_10204,N_8136,N_7538);
and U10205 (N_10205,N_8202,N_7704);
or U10206 (N_10206,N_8972,N_8231);
nor U10207 (N_10207,N_8453,N_7810);
nor U10208 (N_10208,N_7897,N_8762);
nand U10209 (N_10209,N_8711,N_7620);
or U10210 (N_10210,N_8047,N_7574);
or U10211 (N_10211,N_8818,N_8040);
or U10212 (N_10212,N_8967,N_8729);
and U10213 (N_10213,N_8175,N_7749);
nor U10214 (N_10214,N_8028,N_8628);
and U10215 (N_10215,N_7677,N_7888);
nor U10216 (N_10216,N_8103,N_8353);
or U10217 (N_10217,N_8784,N_8845);
xor U10218 (N_10218,N_8222,N_7698);
or U10219 (N_10219,N_7979,N_8962);
or U10220 (N_10220,N_7638,N_8250);
or U10221 (N_10221,N_7966,N_7776);
and U10222 (N_10222,N_8771,N_8431);
nand U10223 (N_10223,N_7504,N_7698);
and U10224 (N_10224,N_8462,N_7779);
nand U10225 (N_10225,N_8979,N_7668);
nand U10226 (N_10226,N_8174,N_8340);
nand U10227 (N_10227,N_8490,N_8734);
xnor U10228 (N_10228,N_8048,N_8103);
or U10229 (N_10229,N_8553,N_8833);
and U10230 (N_10230,N_8697,N_7549);
nor U10231 (N_10231,N_8868,N_8344);
nand U10232 (N_10232,N_8010,N_8231);
or U10233 (N_10233,N_8860,N_7702);
nand U10234 (N_10234,N_8708,N_8351);
or U10235 (N_10235,N_7868,N_8624);
nor U10236 (N_10236,N_8247,N_8676);
nor U10237 (N_10237,N_8718,N_7875);
and U10238 (N_10238,N_8629,N_8030);
or U10239 (N_10239,N_8243,N_8874);
or U10240 (N_10240,N_7763,N_7824);
nor U10241 (N_10241,N_8213,N_7548);
or U10242 (N_10242,N_7812,N_7873);
nand U10243 (N_10243,N_7505,N_8976);
nand U10244 (N_10244,N_8395,N_8984);
and U10245 (N_10245,N_8350,N_8875);
or U10246 (N_10246,N_7514,N_8257);
or U10247 (N_10247,N_8128,N_8340);
and U10248 (N_10248,N_7506,N_7727);
nor U10249 (N_10249,N_8246,N_8148);
or U10250 (N_10250,N_8012,N_8973);
nor U10251 (N_10251,N_8131,N_8549);
nand U10252 (N_10252,N_7639,N_8631);
nor U10253 (N_10253,N_8761,N_8183);
and U10254 (N_10254,N_8529,N_8898);
and U10255 (N_10255,N_8315,N_8951);
xnor U10256 (N_10256,N_8238,N_8423);
nor U10257 (N_10257,N_8096,N_8637);
or U10258 (N_10258,N_8191,N_8883);
nor U10259 (N_10259,N_7952,N_8541);
nor U10260 (N_10260,N_8437,N_7982);
and U10261 (N_10261,N_8917,N_8884);
nor U10262 (N_10262,N_8260,N_8953);
nand U10263 (N_10263,N_7978,N_8987);
nand U10264 (N_10264,N_7794,N_8165);
nand U10265 (N_10265,N_7839,N_8243);
and U10266 (N_10266,N_8723,N_8235);
nand U10267 (N_10267,N_8475,N_8066);
or U10268 (N_10268,N_7985,N_8909);
nand U10269 (N_10269,N_8419,N_8108);
or U10270 (N_10270,N_8352,N_8917);
nand U10271 (N_10271,N_8773,N_7507);
nand U10272 (N_10272,N_8873,N_8203);
nand U10273 (N_10273,N_7550,N_8415);
and U10274 (N_10274,N_8611,N_8842);
nand U10275 (N_10275,N_7928,N_7818);
nor U10276 (N_10276,N_8265,N_8648);
nor U10277 (N_10277,N_8448,N_8894);
nor U10278 (N_10278,N_8247,N_7508);
nor U10279 (N_10279,N_7584,N_8872);
or U10280 (N_10280,N_7841,N_7623);
and U10281 (N_10281,N_7679,N_7754);
xnor U10282 (N_10282,N_7501,N_7803);
and U10283 (N_10283,N_7776,N_7995);
and U10284 (N_10284,N_8483,N_8410);
nor U10285 (N_10285,N_8142,N_8336);
nor U10286 (N_10286,N_8649,N_7655);
nor U10287 (N_10287,N_7813,N_8967);
nand U10288 (N_10288,N_8634,N_7630);
nand U10289 (N_10289,N_8609,N_8705);
nand U10290 (N_10290,N_8448,N_8721);
nand U10291 (N_10291,N_7873,N_8250);
nand U10292 (N_10292,N_7765,N_7944);
and U10293 (N_10293,N_8591,N_8143);
nor U10294 (N_10294,N_8621,N_8096);
and U10295 (N_10295,N_8613,N_8256);
nand U10296 (N_10296,N_8200,N_8613);
or U10297 (N_10297,N_8752,N_7670);
and U10298 (N_10298,N_7670,N_8617);
and U10299 (N_10299,N_8441,N_8470);
and U10300 (N_10300,N_8922,N_8490);
nor U10301 (N_10301,N_8251,N_7850);
nor U10302 (N_10302,N_7793,N_7589);
nor U10303 (N_10303,N_8970,N_7689);
nor U10304 (N_10304,N_8628,N_7963);
nand U10305 (N_10305,N_7695,N_8215);
or U10306 (N_10306,N_8225,N_8720);
nand U10307 (N_10307,N_8535,N_8004);
or U10308 (N_10308,N_8227,N_8359);
and U10309 (N_10309,N_8614,N_7847);
nand U10310 (N_10310,N_8029,N_7901);
and U10311 (N_10311,N_7950,N_8847);
or U10312 (N_10312,N_8672,N_7514);
and U10313 (N_10313,N_7896,N_8347);
or U10314 (N_10314,N_8751,N_8134);
and U10315 (N_10315,N_8452,N_7724);
and U10316 (N_10316,N_8245,N_8406);
nand U10317 (N_10317,N_7762,N_8311);
or U10318 (N_10318,N_8920,N_8620);
nand U10319 (N_10319,N_8090,N_8621);
nor U10320 (N_10320,N_7992,N_7932);
or U10321 (N_10321,N_8994,N_7785);
and U10322 (N_10322,N_7760,N_8264);
or U10323 (N_10323,N_8649,N_8400);
or U10324 (N_10324,N_7517,N_8262);
nand U10325 (N_10325,N_7950,N_8145);
xor U10326 (N_10326,N_7668,N_7915);
nor U10327 (N_10327,N_7857,N_8103);
or U10328 (N_10328,N_7649,N_8643);
nand U10329 (N_10329,N_8607,N_7744);
and U10330 (N_10330,N_7897,N_8704);
and U10331 (N_10331,N_8088,N_8586);
nor U10332 (N_10332,N_7687,N_8709);
nor U10333 (N_10333,N_7544,N_8530);
or U10334 (N_10334,N_7762,N_8936);
nand U10335 (N_10335,N_8849,N_8846);
nand U10336 (N_10336,N_8034,N_7771);
nand U10337 (N_10337,N_8298,N_7583);
nand U10338 (N_10338,N_7658,N_8443);
nor U10339 (N_10339,N_7526,N_7845);
and U10340 (N_10340,N_8717,N_8692);
nand U10341 (N_10341,N_7647,N_8415);
nand U10342 (N_10342,N_8124,N_8671);
xnor U10343 (N_10343,N_8820,N_7917);
nand U10344 (N_10344,N_8543,N_7765);
nor U10345 (N_10345,N_8385,N_8312);
nand U10346 (N_10346,N_7706,N_8350);
nor U10347 (N_10347,N_8889,N_8351);
nor U10348 (N_10348,N_8785,N_8479);
or U10349 (N_10349,N_7884,N_8441);
nand U10350 (N_10350,N_7523,N_7544);
nor U10351 (N_10351,N_8320,N_8875);
or U10352 (N_10352,N_7665,N_8637);
or U10353 (N_10353,N_7935,N_8059);
nor U10354 (N_10354,N_8292,N_7900);
or U10355 (N_10355,N_8335,N_8745);
or U10356 (N_10356,N_7681,N_7910);
nor U10357 (N_10357,N_8201,N_8884);
or U10358 (N_10358,N_7747,N_7816);
or U10359 (N_10359,N_7722,N_8431);
nor U10360 (N_10360,N_8921,N_8034);
nor U10361 (N_10361,N_8017,N_7747);
or U10362 (N_10362,N_8044,N_7856);
nor U10363 (N_10363,N_7597,N_8324);
and U10364 (N_10364,N_7568,N_8342);
nand U10365 (N_10365,N_7748,N_7943);
and U10366 (N_10366,N_7519,N_8494);
or U10367 (N_10367,N_7789,N_8456);
nor U10368 (N_10368,N_8782,N_7658);
and U10369 (N_10369,N_7865,N_8702);
or U10370 (N_10370,N_8842,N_8091);
nand U10371 (N_10371,N_8176,N_8648);
or U10372 (N_10372,N_8169,N_8279);
nand U10373 (N_10373,N_7807,N_8246);
nand U10374 (N_10374,N_7504,N_7776);
or U10375 (N_10375,N_8844,N_7933);
or U10376 (N_10376,N_7796,N_7662);
nand U10377 (N_10377,N_8899,N_8747);
and U10378 (N_10378,N_8866,N_8566);
nand U10379 (N_10379,N_7754,N_8169);
nor U10380 (N_10380,N_8236,N_8112);
nand U10381 (N_10381,N_8805,N_8121);
nand U10382 (N_10382,N_8247,N_8600);
nand U10383 (N_10383,N_7746,N_8675);
nand U10384 (N_10384,N_8038,N_8103);
nand U10385 (N_10385,N_8092,N_8656);
nor U10386 (N_10386,N_8830,N_8099);
and U10387 (N_10387,N_8256,N_7602);
or U10388 (N_10388,N_7680,N_8689);
and U10389 (N_10389,N_8138,N_7546);
or U10390 (N_10390,N_8912,N_8117);
and U10391 (N_10391,N_8477,N_7620);
nor U10392 (N_10392,N_8094,N_8649);
nand U10393 (N_10393,N_7703,N_8931);
nand U10394 (N_10394,N_7895,N_7607);
and U10395 (N_10395,N_7850,N_8841);
or U10396 (N_10396,N_8858,N_7734);
xnor U10397 (N_10397,N_7652,N_8850);
or U10398 (N_10398,N_8797,N_8467);
nand U10399 (N_10399,N_7575,N_7893);
and U10400 (N_10400,N_8529,N_8405);
and U10401 (N_10401,N_8147,N_7716);
nor U10402 (N_10402,N_8903,N_8606);
nor U10403 (N_10403,N_8363,N_8390);
or U10404 (N_10404,N_8620,N_8633);
or U10405 (N_10405,N_8462,N_8672);
or U10406 (N_10406,N_7824,N_8144);
nor U10407 (N_10407,N_7782,N_8624);
or U10408 (N_10408,N_8055,N_8252);
nor U10409 (N_10409,N_7807,N_8196);
and U10410 (N_10410,N_8693,N_7864);
or U10411 (N_10411,N_8620,N_8322);
nor U10412 (N_10412,N_8074,N_8034);
or U10413 (N_10413,N_7931,N_7713);
nor U10414 (N_10414,N_7821,N_8603);
nor U10415 (N_10415,N_8592,N_7922);
and U10416 (N_10416,N_8392,N_8883);
nand U10417 (N_10417,N_8487,N_8784);
or U10418 (N_10418,N_7523,N_7594);
or U10419 (N_10419,N_8454,N_8400);
or U10420 (N_10420,N_7872,N_8777);
and U10421 (N_10421,N_8546,N_8490);
and U10422 (N_10422,N_8539,N_7584);
nor U10423 (N_10423,N_8993,N_7873);
nand U10424 (N_10424,N_8843,N_8953);
or U10425 (N_10425,N_7574,N_8018);
nor U10426 (N_10426,N_8855,N_8229);
nor U10427 (N_10427,N_7748,N_7650);
nor U10428 (N_10428,N_8766,N_7503);
or U10429 (N_10429,N_8450,N_8274);
and U10430 (N_10430,N_8946,N_8706);
nor U10431 (N_10431,N_8978,N_8593);
and U10432 (N_10432,N_8393,N_8110);
and U10433 (N_10433,N_8007,N_8355);
or U10434 (N_10434,N_8954,N_8318);
or U10435 (N_10435,N_8389,N_8818);
nor U10436 (N_10436,N_7904,N_8587);
and U10437 (N_10437,N_8734,N_7513);
or U10438 (N_10438,N_7536,N_7757);
nor U10439 (N_10439,N_8728,N_8245);
nand U10440 (N_10440,N_7694,N_7671);
or U10441 (N_10441,N_7652,N_7641);
nor U10442 (N_10442,N_7943,N_7843);
nand U10443 (N_10443,N_8641,N_7544);
or U10444 (N_10444,N_7670,N_8594);
xnor U10445 (N_10445,N_8324,N_7707);
and U10446 (N_10446,N_8825,N_8397);
and U10447 (N_10447,N_8308,N_8674);
and U10448 (N_10448,N_8119,N_8663);
nand U10449 (N_10449,N_8623,N_7944);
nor U10450 (N_10450,N_8720,N_7916);
and U10451 (N_10451,N_7644,N_8211);
nand U10452 (N_10452,N_8623,N_8163);
or U10453 (N_10453,N_7693,N_8910);
or U10454 (N_10454,N_7565,N_7774);
or U10455 (N_10455,N_7692,N_7635);
nor U10456 (N_10456,N_8430,N_8959);
or U10457 (N_10457,N_7765,N_8317);
nand U10458 (N_10458,N_8272,N_8293);
or U10459 (N_10459,N_8141,N_8564);
nand U10460 (N_10460,N_8206,N_8032);
nor U10461 (N_10461,N_7884,N_8824);
nor U10462 (N_10462,N_8543,N_8951);
or U10463 (N_10463,N_8705,N_8479);
nor U10464 (N_10464,N_8159,N_8167);
or U10465 (N_10465,N_8939,N_7644);
or U10466 (N_10466,N_8954,N_8468);
and U10467 (N_10467,N_8149,N_8045);
xor U10468 (N_10468,N_8549,N_7807);
nor U10469 (N_10469,N_8858,N_8658);
nor U10470 (N_10470,N_8725,N_8569);
nand U10471 (N_10471,N_8276,N_7848);
nor U10472 (N_10472,N_8771,N_8415);
nand U10473 (N_10473,N_8381,N_8324);
nor U10474 (N_10474,N_7797,N_8197);
nor U10475 (N_10475,N_8660,N_8929);
nand U10476 (N_10476,N_8050,N_8609);
and U10477 (N_10477,N_8825,N_8361);
nand U10478 (N_10478,N_8859,N_8975);
nor U10479 (N_10479,N_8983,N_8155);
nand U10480 (N_10480,N_8617,N_8456);
and U10481 (N_10481,N_8920,N_8722);
nor U10482 (N_10482,N_7676,N_7605);
and U10483 (N_10483,N_8748,N_8295);
or U10484 (N_10484,N_7510,N_8609);
and U10485 (N_10485,N_8176,N_8758);
and U10486 (N_10486,N_8915,N_8335);
and U10487 (N_10487,N_8822,N_7680);
nor U10488 (N_10488,N_8653,N_7947);
nor U10489 (N_10489,N_7721,N_7836);
nand U10490 (N_10490,N_8702,N_8045);
or U10491 (N_10491,N_8543,N_8539);
and U10492 (N_10492,N_8703,N_7859);
nor U10493 (N_10493,N_8365,N_7523);
nor U10494 (N_10494,N_8578,N_8663);
and U10495 (N_10495,N_8876,N_8733);
nor U10496 (N_10496,N_8875,N_7722);
xnor U10497 (N_10497,N_7762,N_8640);
or U10498 (N_10498,N_8899,N_8801);
or U10499 (N_10499,N_8849,N_8206);
nor U10500 (N_10500,N_9756,N_9677);
nand U10501 (N_10501,N_9325,N_9049);
or U10502 (N_10502,N_10392,N_10009);
xnor U10503 (N_10503,N_9273,N_9088);
or U10504 (N_10504,N_9211,N_9656);
nand U10505 (N_10505,N_10338,N_9402);
and U10506 (N_10506,N_9743,N_9221);
nand U10507 (N_10507,N_9702,N_9499);
nand U10508 (N_10508,N_9801,N_10391);
or U10509 (N_10509,N_10289,N_9246);
or U10510 (N_10510,N_9632,N_10141);
nand U10511 (N_10511,N_9000,N_9306);
or U10512 (N_10512,N_10277,N_10308);
nor U10513 (N_10513,N_9114,N_9324);
nand U10514 (N_10514,N_10484,N_9422);
and U10515 (N_10515,N_9643,N_10068);
nor U10516 (N_10516,N_9960,N_9400);
nor U10517 (N_10517,N_9660,N_9909);
nand U10518 (N_10518,N_10489,N_10447);
or U10519 (N_10519,N_10359,N_10232);
nor U10520 (N_10520,N_9526,N_9045);
and U10521 (N_10521,N_9321,N_9963);
and U10522 (N_10522,N_9369,N_9782);
nand U10523 (N_10523,N_9089,N_9223);
nor U10524 (N_10524,N_9747,N_9760);
nor U10525 (N_10525,N_9816,N_10167);
nor U10526 (N_10526,N_9435,N_9812);
or U10527 (N_10527,N_9887,N_10438);
and U10528 (N_10528,N_9787,N_9992);
nor U10529 (N_10529,N_10081,N_9419);
nand U10530 (N_10530,N_9824,N_9018);
nor U10531 (N_10531,N_9978,N_9692);
nand U10532 (N_10532,N_10299,N_10098);
or U10533 (N_10533,N_9279,N_9733);
or U10534 (N_10534,N_10417,N_9872);
or U10535 (N_10535,N_9942,N_9574);
nor U10536 (N_10536,N_10314,N_9235);
nand U10537 (N_10537,N_9074,N_9858);
nor U10538 (N_10538,N_10468,N_10346);
or U10539 (N_10539,N_9388,N_10432);
nor U10540 (N_10540,N_10161,N_9976);
nand U10541 (N_10541,N_9258,N_9350);
and U10542 (N_10542,N_9688,N_9448);
nor U10543 (N_10543,N_9224,N_10353);
or U10544 (N_10544,N_9810,N_10347);
nor U10545 (N_10545,N_9030,N_10216);
nor U10546 (N_10546,N_10485,N_9160);
nand U10547 (N_10547,N_9763,N_9930);
nor U10548 (N_10548,N_9794,N_9167);
nand U10549 (N_10549,N_10085,N_9550);
and U10550 (N_10550,N_9594,N_9637);
and U10551 (N_10551,N_9043,N_9515);
nand U10552 (N_10552,N_9806,N_9482);
nor U10553 (N_10553,N_10117,N_9840);
or U10554 (N_10554,N_9520,N_9480);
nand U10555 (N_10555,N_9151,N_9944);
or U10556 (N_10556,N_10178,N_9393);
nand U10557 (N_10557,N_9729,N_10386);
or U10558 (N_10558,N_9013,N_9943);
nand U10559 (N_10559,N_10249,N_10415);
nor U10560 (N_10560,N_9502,N_9905);
or U10561 (N_10561,N_9430,N_10390);
nor U10562 (N_10562,N_10186,N_9778);
nand U10563 (N_10563,N_9041,N_9478);
and U10564 (N_10564,N_10193,N_9335);
or U10565 (N_10565,N_9161,N_10145);
nand U10566 (N_10566,N_10394,N_10477);
or U10567 (N_10567,N_10240,N_9257);
or U10568 (N_10568,N_10451,N_10144);
nand U10569 (N_10569,N_9039,N_10088);
nand U10570 (N_10570,N_9189,N_9069);
or U10571 (N_10571,N_9395,N_10032);
nor U10572 (N_10572,N_9183,N_9843);
and U10573 (N_10573,N_10062,N_10022);
and U10574 (N_10574,N_10310,N_9815);
nand U10575 (N_10575,N_9484,N_9655);
nor U10576 (N_10576,N_9300,N_9710);
and U10577 (N_10577,N_10472,N_10475);
nor U10578 (N_10578,N_9033,N_10031);
nor U10579 (N_10579,N_9761,N_9740);
nor U10580 (N_10580,N_9025,N_9052);
nand U10581 (N_10581,N_9627,N_9294);
and U10582 (N_10582,N_9922,N_9842);
and U10583 (N_10583,N_10054,N_10076);
or U10584 (N_10584,N_9267,N_10125);
nand U10585 (N_10585,N_10162,N_10056);
and U10586 (N_10586,N_10266,N_9899);
or U10587 (N_10587,N_9586,N_9973);
and U10588 (N_10588,N_9295,N_9204);
or U10589 (N_10589,N_9219,N_9690);
or U10590 (N_10590,N_9636,N_10011);
nand U10591 (N_10591,N_9653,N_9083);
nand U10592 (N_10592,N_9471,N_10225);
and U10593 (N_10593,N_9617,N_9714);
nor U10594 (N_10594,N_9738,N_10416);
and U10595 (N_10595,N_9330,N_9141);
and U10596 (N_10596,N_10187,N_9622);
or U10597 (N_10597,N_10066,N_9648);
or U10598 (N_10598,N_9540,N_9110);
and U10599 (N_10599,N_9260,N_9012);
nand U10600 (N_10600,N_9621,N_10356);
nand U10601 (N_10601,N_9265,N_9570);
and U10602 (N_10602,N_9460,N_9486);
xor U10603 (N_10603,N_10093,N_9202);
and U10604 (N_10604,N_9477,N_10109);
xor U10605 (N_10605,N_9831,N_9796);
or U10606 (N_10606,N_9387,N_10008);
or U10607 (N_10607,N_10307,N_9382);
xnor U10608 (N_10608,N_9775,N_9463);
nand U10609 (N_10609,N_9323,N_9607);
or U10610 (N_10610,N_9370,N_9972);
nor U10611 (N_10611,N_10280,N_10173);
and U10612 (N_10612,N_10378,N_9085);
nand U10613 (N_10613,N_10092,N_9708);
nor U10614 (N_10614,N_10369,N_9524);
nor U10615 (N_10615,N_10483,N_10450);
nor U10616 (N_10616,N_9491,N_9150);
and U10617 (N_10617,N_10150,N_9634);
and U10618 (N_10618,N_9061,N_10149);
or U10619 (N_10619,N_9820,N_10445);
and U10620 (N_10620,N_9935,N_9554);
nand U10621 (N_10621,N_10016,N_9615);
or U10622 (N_10622,N_10146,N_9493);
nor U10623 (N_10623,N_9641,N_9340);
or U10624 (N_10624,N_10034,N_9937);
nor U10625 (N_10625,N_10351,N_9344);
or U10626 (N_10626,N_9606,N_10360);
nor U10627 (N_10627,N_9585,N_9666);
nand U10628 (N_10628,N_9543,N_9414);
nor U10629 (N_10629,N_10033,N_9754);
or U10630 (N_10630,N_9256,N_10278);
or U10631 (N_10631,N_9099,N_9307);
nand U10632 (N_10632,N_9910,N_9312);
nor U10633 (N_10633,N_9758,N_10184);
nor U10634 (N_10634,N_10449,N_9195);
nand U10635 (N_10635,N_9216,N_9588);
nand U10636 (N_10636,N_9440,N_10212);
nand U10637 (N_10637,N_10252,N_9091);
nor U10638 (N_10638,N_9277,N_9599);
nor U10639 (N_10639,N_9557,N_9838);
or U10640 (N_10640,N_9113,N_10486);
and U10641 (N_10641,N_9956,N_9188);
nor U10642 (N_10642,N_9203,N_9427);
and U10643 (N_10643,N_10015,N_9149);
nor U10644 (N_10644,N_9144,N_9252);
or U10645 (N_10645,N_9987,N_9605);
or U10646 (N_10646,N_9248,N_9210);
nand U10647 (N_10647,N_9379,N_9239);
and U10648 (N_10648,N_9732,N_9962);
nor U10649 (N_10649,N_9559,N_9693);
nand U10650 (N_10650,N_10474,N_10222);
nand U10651 (N_10651,N_9527,N_10463);
nor U10652 (N_10652,N_9062,N_9583);
nand U10653 (N_10653,N_9871,N_10430);
nand U10654 (N_10654,N_9337,N_9122);
or U10655 (N_10655,N_9187,N_10330);
and U10656 (N_10656,N_9124,N_9462);
nor U10657 (N_10657,N_9951,N_9888);
or U10658 (N_10658,N_9560,N_10148);
nor U10659 (N_10659,N_9251,N_9284);
nor U10660 (N_10660,N_9105,N_9695);
xor U10661 (N_10661,N_9548,N_9867);
and U10662 (N_10662,N_9713,N_10448);
and U10663 (N_10663,N_10132,N_9184);
nand U10664 (N_10664,N_10423,N_9050);
nand U10665 (N_10665,N_9022,N_9054);
nor U10666 (N_10666,N_9006,N_9142);
nor U10667 (N_10667,N_9642,N_9949);
or U10668 (N_10668,N_10379,N_9722);
nand U10669 (N_10669,N_9551,N_9556);
nand U10670 (N_10670,N_9681,N_10136);
nand U10671 (N_10671,N_9862,N_9800);
nor U10672 (N_10672,N_10418,N_9261);
and U10673 (N_10673,N_10482,N_9539);
or U10674 (N_10674,N_9880,N_9115);
and U10675 (N_10675,N_9023,N_9181);
nor U10676 (N_10676,N_10110,N_9117);
nand U10677 (N_10677,N_9029,N_9886);
nor U10678 (N_10678,N_9581,N_10010);
nor U10679 (N_10679,N_9669,N_9194);
xnor U10680 (N_10680,N_10261,N_9250);
nand U10681 (N_10681,N_9673,N_9241);
nand U10682 (N_10682,N_9966,N_10272);
and U10683 (N_10683,N_10365,N_9936);
nand U10684 (N_10684,N_9523,N_10368);
nand U10685 (N_10685,N_9229,N_9109);
nor U10686 (N_10686,N_9870,N_10460);
nand U10687 (N_10687,N_10080,N_10035);
nor U10688 (N_10688,N_9839,N_9620);
nand U10689 (N_10689,N_10082,N_10334);
or U10690 (N_10690,N_9496,N_9865);
nor U10691 (N_10691,N_10456,N_10180);
or U10692 (N_10692,N_10052,N_10270);
or U10693 (N_10693,N_10013,N_10227);
and U10694 (N_10694,N_10263,N_10287);
nor U10695 (N_10695,N_9542,N_10172);
nand U10696 (N_10696,N_10409,N_10407);
and U10697 (N_10697,N_9811,N_9734);
and U10698 (N_10698,N_9222,N_10376);
and U10699 (N_10699,N_9670,N_9952);
xnor U10700 (N_10700,N_10290,N_9508);
and U10701 (N_10701,N_9311,N_9741);
nor U10702 (N_10702,N_9968,N_10211);
and U10703 (N_10703,N_9107,N_9852);
and U10704 (N_10704,N_9674,N_10064);
or U10705 (N_10705,N_10246,N_9441);
nor U10706 (N_10706,N_10103,N_9644);
or U10707 (N_10707,N_10118,N_9595);
nor U10708 (N_10708,N_9932,N_9657);
and U10709 (N_10709,N_10251,N_9073);
nor U10710 (N_10710,N_9771,N_10166);
nor U10711 (N_10711,N_9197,N_9361);
nand U10712 (N_10712,N_10079,N_9007);
nand U10713 (N_10713,N_9940,N_9730);
nand U10714 (N_10714,N_9234,N_9918);
nand U10715 (N_10715,N_9333,N_9928);
nand U10716 (N_10716,N_9240,N_9631);
and U10717 (N_10717,N_10399,N_9404);
nand U10718 (N_10718,N_9549,N_9565);
nand U10719 (N_10719,N_9903,N_9360);
nand U10720 (N_10720,N_9139,N_9822);
nor U10721 (N_10721,N_9895,N_9879);
or U10722 (N_10722,N_9517,N_9809);
or U10723 (N_10723,N_9534,N_10428);
or U10724 (N_10724,N_9112,N_10095);
nand U10725 (N_10725,N_9345,N_10333);
nand U10726 (N_10726,N_9390,N_9072);
and U10727 (N_10727,N_9485,N_9442);
nand U10728 (N_10728,N_9797,N_9953);
nand U10729 (N_10729,N_9916,N_9803);
or U10730 (N_10730,N_9920,N_9532);
nor U10731 (N_10731,N_9985,N_10454);
nor U10732 (N_10732,N_9925,N_9134);
or U10733 (N_10733,N_9443,N_10275);
or U10734 (N_10734,N_10320,N_10182);
and U10735 (N_10735,N_9476,N_9076);
xor U10736 (N_10736,N_10041,N_10181);
nand U10737 (N_10737,N_10191,N_9707);
and U10738 (N_10738,N_10493,N_9140);
or U10739 (N_10739,N_9717,N_9979);
or U10740 (N_10740,N_9037,N_9026);
and U10741 (N_10741,N_10206,N_9900);
and U10742 (N_10742,N_10140,N_10316);
and U10743 (N_10743,N_9721,N_9123);
nor U10744 (N_10744,N_9452,N_10265);
nor U10745 (N_10745,N_9504,N_10366);
and U10746 (N_10746,N_10143,N_10214);
and U10747 (N_10747,N_10242,N_9954);
or U10748 (N_10748,N_10377,N_10237);
nand U10749 (N_10749,N_9431,N_10005);
nand U10750 (N_10750,N_9845,N_9065);
xor U10751 (N_10751,N_9343,N_10337);
nor U10752 (N_10752,N_9682,N_9165);
or U10753 (N_10753,N_9399,N_9613);
nand U10754 (N_10754,N_10241,N_9982);
and U10755 (N_10755,N_9084,N_9612);
or U10756 (N_10756,N_9371,N_9401);
xnor U10757 (N_10757,N_9863,N_10481);
or U10758 (N_10758,N_9469,N_9193);
nor U10759 (N_10759,N_10344,N_9719);
and U10760 (N_10760,N_10464,N_9948);
nand U10761 (N_10761,N_9227,N_9226);
or U10762 (N_10762,N_10458,N_9813);
nand U10763 (N_10763,N_10127,N_9587);
nor U10764 (N_10764,N_9757,N_10048);
nand U10765 (N_10765,N_9933,N_9603);
nor U10766 (N_10766,N_9190,N_10205);
nand U10767 (N_10767,N_9971,N_10324);
nand U10768 (N_10768,N_10163,N_9047);
nand U10769 (N_10769,N_9433,N_10147);
nor U10770 (N_10770,N_9159,N_9731);
or U10771 (N_10771,N_9292,N_10404);
nand U10772 (N_10772,N_9638,N_10023);
and U10773 (N_10773,N_9341,N_9266);
or U10774 (N_10774,N_10123,N_9132);
and U10775 (N_10775,N_9403,N_10453);
nor U10776 (N_10776,N_10340,N_10350);
nand U10777 (N_10777,N_9964,N_9411);
xor U10778 (N_10778,N_9339,N_9322);
nand U10779 (N_10779,N_10139,N_9255);
nand U10780 (N_10780,N_9991,N_10304);
or U10781 (N_10781,N_9623,N_9199);
and U10782 (N_10782,N_9684,N_9817);
and U10783 (N_10783,N_9882,N_9749);
and U10784 (N_10784,N_9002,N_9215);
nor U10785 (N_10785,N_10020,N_9133);
and U10786 (N_10786,N_9506,N_9793);
and U10787 (N_10787,N_9700,N_10306);
nand U10788 (N_10788,N_9108,N_10395);
and U10789 (N_10789,N_9897,N_9040);
or U10790 (N_10790,N_9200,N_10188);
nand U10791 (N_10791,N_9214,N_10107);
or U10792 (N_10792,N_9590,N_9051);
xor U10793 (N_10793,N_9889,N_9630);
nor U10794 (N_10794,N_10003,N_9823);
nor U10795 (N_10795,N_10221,N_9434);
nor U10796 (N_10796,N_10159,N_9497);
nand U10797 (N_10797,N_10497,N_9179);
and U10798 (N_10798,N_9629,N_10440);
or U10799 (N_10799,N_9773,N_9474);
and U10800 (N_10800,N_9358,N_9170);
and U10801 (N_10801,N_10298,N_9596);
or U10802 (N_10802,N_10325,N_9699);
nor U10803 (N_10803,N_9444,N_9297);
or U10804 (N_10804,N_9659,N_9009);
nor U10805 (N_10805,N_10437,N_9394);
nand U10806 (N_10806,N_9173,N_9171);
nor U10807 (N_10807,N_9698,N_9407);
nor U10808 (N_10808,N_10490,N_10012);
nand U10809 (N_10809,N_9281,N_9847);
nand U10810 (N_10810,N_10154,N_10429);
nand U10811 (N_10811,N_9753,N_10248);
nand U10812 (N_10812,N_9553,N_9172);
nand U10813 (N_10813,N_9475,N_10345);
nor U10814 (N_10814,N_9016,N_10367);
and U10815 (N_10815,N_9011,N_10393);
nand U10816 (N_10816,N_10315,N_9042);
and U10817 (N_10817,N_9230,N_10348);
nand U10818 (N_10818,N_9946,N_9131);
nor U10819 (N_10819,N_9286,N_9704);
nor U10820 (N_10820,N_10327,N_9327);
nor U10821 (N_10821,N_9875,N_9676);
nor U10822 (N_10822,N_9153,N_9280);
or U10823 (N_10823,N_9737,N_9687);
nand U10824 (N_10824,N_10371,N_9004);
or U10825 (N_10825,N_9896,N_9119);
or U10826 (N_10826,N_9299,N_10074);
or U10827 (N_10827,N_9950,N_9336);
and U10828 (N_10828,N_9201,N_9449);
or U10829 (N_10829,N_9850,N_9518);
or U10830 (N_10830,N_9313,N_9432);
nor U10831 (N_10831,N_10274,N_9316);
and U10832 (N_10832,N_10219,N_9262);
or U10833 (N_10833,N_9137,N_9728);
nor U10834 (N_10834,N_9245,N_9175);
nor U10835 (N_10835,N_9331,N_9828);
nand U10836 (N_10836,N_9367,N_9198);
and U10837 (N_10837,N_9868,N_10115);
or U10838 (N_10838,N_9683,N_9102);
or U10839 (N_10839,N_10235,N_10383);
nand U10840 (N_10840,N_10382,N_9777);
or U10841 (N_10841,N_10075,N_9055);
and U10842 (N_10842,N_10065,N_10256);
and U10843 (N_10843,N_9989,N_10017);
or U10844 (N_10844,N_10268,N_9254);
or U10845 (N_10845,N_10467,N_9329);
xor U10846 (N_10846,N_9466,N_10250);
or U10847 (N_10847,N_10189,N_10491);
or U10848 (N_10848,N_10309,N_9079);
or U10849 (N_10849,N_9685,N_9374);
or U10850 (N_10850,N_9618,N_9456);
or U10851 (N_10851,N_9884,N_9802);
and U10852 (N_10852,N_9287,N_9075);
nor U10853 (N_10853,N_9036,N_10087);
and U10854 (N_10854,N_10312,N_9652);
nor U10855 (N_10855,N_9939,N_9785);
xnor U10856 (N_10856,N_9278,N_9436);
and U10857 (N_10857,N_10183,N_9536);
and U10858 (N_10858,N_9326,N_9237);
or U10859 (N_10859,N_9912,N_10398);
nand U10860 (N_10860,N_9437,N_9513);
nand U10861 (N_10861,N_10119,N_10069);
and U10862 (N_10862,N_9579,N_9375);
and U10863 (N_10863,N_10282,N_10201);
nand U10864 (N_10864,N_10461,N_10202);
nand U10865 (N_10865,N_9592,N_9694);
and U10866 (N_10866,N_9014,N_9097);
nand U10867 (N_10867,N_9063,N_10495);
and U10868 (N_10868,N_9604,N_9064);
nor U10869 (N_10869,N_9851,N_9856);
nand U10870 (N_10870,N_10155,N_9247);
and U10871 (N_10871,N_9853,N_10037);
or U10872 (N_10872,N_9945,N_10257);
or U10873 (N_10873,N_9472,N_9242);
or U10874 (N_10874,N_9155,N_9470);
and U10875 (N_10875,N_9993,N_9176);
or U10876 (N_10876,N_9885,N_10028);
nor U10877 (N_10877,N_10479,N_9791);
or U10878 (N_10878,N_9667,N_9894);
nor U10879 (N_10879,N_10083,N_9917);
nand U10880 (N_10880,N_9464,N_9019);
nor U10881 (N_10881,N_9755,N_10311);
or U10882 (N_10882,N_10019,N_9135);
nand U10883 (N_10883,N_9034,N_10165);
or U10884 (N_10884,N_10247,N_9145);
nand U10885 (N_10885,N_9650,N_9528);
and U10886 (N_10886,N_9712,N_9389);
nor U10887 (N_10887,N_9908,N_9772);
or U10888 (N_10888,N_10412,N_9696);
or U10889 (N_10889,N_9829,N_9348);
nand U10890 (N_10890,N_9154,N_10478);
and U10891 (N_10891,N_9104,N_10317);
and U10892 (N_10892,N_9383,N_9697);
or U10893 (N_10893,N_9111,N_9031);
nand U10894 (N_10894,N_10496,N_10025);
nand U10895 (N_10895,N_10018,N_9639);
and U10896 (N_10896,N_9156,N_10046);
or U10897 (N_10897,N_10444,N_10462);
nor U10898 (N_10898,N_9409,N_10396);
or U10899 (N_10899,N_9931,N_10070);
and U10900 (N_10900,N_9762,N_9315);
nand U10901 (N_10901,N_9275,N_9391);
or U10902 (N_10902,N_10194,N_10370);
and U10903 (N_10903,N_10465,N_9303);
nor U10904 (N_10904,N_9904,N_10318);
and U10905 (N_10905,N_10476,N_9938);
and U10906 (N_10906,N_10057,N_9582);
nor U10907 (N_10907,N_10158,N_9724);
nand U10908 (N_10908,N_10199,N_9274);
and U10909 (N_10909,N_9148,N_9308);
and U10910 (N_10910,N_10264,N_10285);
nand U10911 (N_10911,N_10197,N_10343);
nor U10912 (N_10912,N_9561,N_9832);
nor U10913 (N_10913,N_9378,N_9799);
nand U10914 (N_10914,N_9774,N_9934);
and U10915 (N_10915,N_9790,N_9525);
nor U10916 (N_10916,N_9208,N_10133);
or U10917 (N_10917,N_9866,N_9723);
nor U10918 (N_10918,N_9901,N_9347);
nand U10919 (N_10919,N_9413,N_10058);
or U10920 (N_10920,N_9205,N_9218);
nor U10921 (N_10921,N_9467,N_9024);
nand U10922 (N_10922,N_9529,N_10209);
or U10923 (N_10923,N_9876,N_10000);
nand U10924 (N_10924,N_9368,N_9298);
and U10925 (N_10925,N_9487,N_9332);
nor U10926 (N_10926,N_9573,N_9302);
nor U10927 (N_10927,N_10466,N_10038);
nor U10928 (N_10928,N_9418,N_10039);
or U10929 (N_10929,N_10230,N_9609);
nor U10930 (N_10930,N_9010,N_10036);
or U10931 (N_10931,N_10494,N_9021);
and U10932 (N_10932,N_9309,N_9874);
and U10933 (N_10933,N_10200,N_9649);
or U10934 (N_10934,N_10294,N_10323);
nor U10935 (N_10935,N_9709,N_9098);
and U10936 (N_10936,N_9269,N_10223);
and U10937 (N_10937,N_10196,N_10279);
and U10938 (N_10938,N_10099,N_10402);
nand U10939 (N_10939,N_9398,N_9983);
or U10940 (N_10940,N_9301,N_9317);
and U10941 (N_10941,N_9027,N_9384);
nor U10942 (N_10942,N_9352,N_9001);
nand U10943 (N_10943,N_9781,N_9998);
nor U10944 (N_10944,N_10130,N_9869);
or U10945 (N_10945,N_10419,N_9959);
nor U10946 (N_10946,N_9505,N_9633);
nand U10947 (N_10947,N_9805,N_9366);
nand U10948 (N_10948,N_9584,N_9967);
or U10949 (N_10949,N_9078,N_9451);
or U10950 (N_10950,N_10339,N_10029);
nand U10951 (N_10951,N_9503,N_10372);
or U10952 (N_10952,N_9490,N_9571);
nand U10953 (N_10953,N_10300,N_9718);
nand U10954 (N_10954,N_9380,N_9293);
or U10955 (N_10955,N_9921,N_9096);
nor U10956 (N_10956,N_9835,N_9498);
nand U10957 (N_10957,N_9680,N_10385);
nand U10958 (N_10958,N_9126,N_9819);
or U10959 (N_10959,N_9365,N_9779);
and U10960 (N_10960,N_10185,N_9645);
or U10961 (N_10961,N_9898,N_9555);
and U10962 (N_10962,N_9915,N_9489);
and U10963 (N_10963,N_9459,N_9070);
nor U10964 (N_10964,N_10096,N_9020);
and U10965 (N_10965,N_10434,N_10425);
or U10966 (N_10966,N_9077,N_9958);
and U10967 (N_10967,N_10061,N_9977);
nor U10968 (N_10968,N_9535,N_9169);
nor U10969 (N_10969,N_9726,N_9919);
nor U10970 (N_10970,N_10168,N_9665);
or U10971 (N_10971,N_9186,N_10441);
and U10972 (N_10972,N_9715,N_10255);
and U10973 (N_10973,N_10195,N_9093);
nor U10974 (N_10974,N_9562,N_10030);
nor U10975 (N_10975,N_9635,N_9878);
nand U10976 (N_10976,N_10326,N_10470);
or U10977 (N_10977,N_10374,N_10260);
nand U10978 (N_10978,N_9357,N_9338);
nor U10979 (N_10979,N_10271,N_9415);
and U10980 (N_10980,N_9530,N_9028);
nand U10981 (N_10981,N_10153,N_10480);
or U10982 (N_10982,N_9209,N_9746);
and U10983 (N_10983,N_10105,N_9182);
nand U10984 (N_10984,N_10269,N_10455);
nor U10985 (N_10985,N_9397,N_9924);
and U10986 (N_10986,N_9121,N_9577);
and U10987 (N_10987,N_9501,N_9318);
nor U10988 (N_10988,N_9305,N_9957);
nor U10989 (N_10989,N_9748,N_9668);
xnor U10990 (N_10990,N_9488,N_10234);
nand U10991 (N_10991,N_9883,N_9844);
nand U10992 (N_10992,N_9727,N_10375);
and U10993 (N_10993,N_9969,N_9481);
nand U10994 (N_10994,N_9406,N_9744);
and U10995 (N_10995,N_9351,N_10090);
or U10996 (N_10996,N_10111,N_9103);
or U10997 (N_10997,N_10142,N_10175);
and U10998 (N_10998,N_9626,N_10388);
or U10999 (N_10999,N_10335,N_9507);
nand U11000 (N_11000,N_10498,N_9911);
nor U11001 (N_11001,N_10435,N_10421);
nor U11002 (N_11002,N_9848,N_9243);
nand U11003 (N_11003,N_10457,N_10492);
and U11004 (N_11004,N_9362,N_9511);
and U11005 (N_11005,N_9664,N_9453);
and U11006 (N_11006,N_9980,N_10204);
nor U11007 (N_11007,N_9999,N_10439);
and U11008 (N_11008,N_9941,N_10152);
nand U11009 (N_11009,N_9058,N_10443);
or U11010 (N_11010,N_9759,N_9568);
nor U11011 (N_11011,N_10413,N_10245);
nand U11012 (N_11012,N_9833,N_9483);
nor U11013 (N_11013,N_10384,N_9233);
or U11014 (N_11014,N_9236,N_9616);
and U11015 (N_11015,N_10156,N_9408);
xnor U11016 (N_11016,N_10488,N_10129);
nor U11017 (N_11017,N_9547,N_9742);
or U11018 (N_11018,N_9125,N_10253);
and U11019 (N_11019,N_9720,N_10342);
and U11020 (N_11020,N_9138,N_10420);
nand U11021 (N_11021,N_9057,N_9786);
nand U11022 (N_11022,N_10177,N_9814);
nor U11023 (N_11023,N_9446,N_9576);
and U11024 (N_11024,N_9625,N_9975);
nand U11025 (N_11025,N_10389,N_10414);
or U11026 (N_11026,N_9457,N_9567);
or U11027 (N_11027,N_9191,N_10084);
and U11028 (N_11028,N_9906,N_10471);
or U11029 (N_11029,N_9213,N_9038);
and U11030 (N_11030,N_9751,N_9776);
or U11031 (N_11031,N_10276,N_10094);
nand U11032 (N_11032,N_10291,N_9291);
or U11033 (N_11033,N_9996,N_10410);
nor U11034 (N_11034,N_9087,N_9468);
nor U11035 (N_11035,N_9118,N_9647);
and U11036 (N_11036,N_9807,N_9129);
nand U11037 (N_11037,N_9304,N_9531);
nor U11038 (N_11038,N_10352,N_9624);
or U11039 (N_11039,N_9271,N_9522);
nor U11040 (N_11040,N_9166,N_10302);
nor U11041 (N_11041,N_9372,N_9168);
and U11042 (N_11042,N_10361,N_9003);
and U11043 (N_11043,N_10469,N_9902);
xnor U11044 (N_11044,N_10258,N_9745);
nor U11045 (N_11045,N_9359,N_9283);
or U11046 (N_11046,N_9289,N_10364);
and U11047 (N_11047,N_9355,N_9185);
nor U11048 (N_11048,N_9591,N_9981);
nand U11049 (N_11049,N_9225,N_9066);
nand U11050 (N_11050,N_9947,N_9310);
nor U11051 (N_11051,N_9412,N_9558);
nor U11052 (N_11052,N_10121,N_10051);
nor U11053 (N_11053,N_10243,N_10024);
nor U11054 (N_11054,N_10100,N_9736);
and U11055 (N_11055,N_9207,N_9494);
and U11056 (N_11056,N_9857,N_10071);
nand U11057 (N_11057,N_10236,N_9552);
or U11058 (N_11058,N_10305,N_9827);
nand U11059 (N_11059,N_10192,N_10297);
nor U11060 (N_11060,N_10336,N_9739);
and U11061 (N_11061,N_9846,N_10215);
or U11062 (N_11062,N_9675,N_9164);
nor U11063 (N_11063,N_9923,N_9147);
and U11064 (N_11064,N_9986,N_10401);
and U11065 (N_11065,N_9231,N_10007);
and U11066 (N_11066,N_10040,N_10358);
and U11067 (N_11067,N_10286,N_10120);
or U11068 (N_11068,N_10400,N_9479);
nor U11069 (N_11069,N_10403,N_9662);
or U11070 (N_11070,N_9593,N_10239);
nor U11071 (N_11071,N_9619,N_9798);
or U11072 (N_11072,N_10231,N_10208);
nand U11073 (N_11073,N_10473,N_9891);
and U11074 (N_11074,N_10433,N_9363);
and U11075 (N_11075,N_10176,N_9082);
nor U11076 (N_11076,N_9837,N_9127);
nor U11077 (N_11077,N_10026,N_9101);
xor U11078 (N_11078,N_10203,N_10170);
nor U11079 (N_11079,N_9015,N_10053);
and U11080 (N_11080,N_10408,N_10108);
nor U11081 (N_11081,N_9601,N_10499);
or U11082 (N_11082,N_9546,N_10171);
and U11083 (N_11083,N_9927,N_10134);
or U11084 (N_11084,N_9410,N_9081);
nor U11085 (N_11085,N_9495,N_9244);
nor U11086 (N_11086,N_9238,N_10355);
or U11087 (N_11087,N_9438,N_9864);
nor U11088 (N_11088,N_9961,N_9572);
or U11089 (N_11089,N_9752,N_10288);
or U11090 (N_11090,N_9672,N_9420);
or U11091 (N_11091,N_9705,N_9580);
or U11092 (N_11092,N_9276,N_10233);
nor U11093 (N_11093,N_9095,N_9545);
and U11094 (N_11094,N_10045,N_9764);
nor U11095 (N_11095,N_9792,N_9509);
nor U11096 (N_11096,N_10313,N_9855);
xor U11097 (N_11097,N_9830,N_9997);
nand U11098 (N_11098,N_9533,N_9514);
xor U11099 (N_11099,N_9272,N_10422);
nand U11100 (N_11100,N_9766,N_9067);
or U11101 (N_11101,N_9228,N_9881);
nor U11102 (N_11102,N_10089,N_9860);
nor U11103 (N_11103,N_9100,N_9725);
or U11104 (N_11104,N_10331,N_9120);
or U11105 (N_11105,N_10228,N_9068);
or U11106 (N_11106,N_9610,N_10073);
and U11107 (N_11107,N_10292,N_10044);
nand U11108 (N_11108,N_9319,N_10332);
nand U11109 (N_11109,N_10397,N_9821);
and U11110 (N_11110,N_9735,N_9465);
and U11111 (N_11111,N_9473,N_9841);
nand U11112 (N_11112,N_9396,N_9686);
nor U11113 (N_11113,N_9264,N_10104);
nor U11114 (N_11114,N_10328,N_10060);
and U11115 (N_11115,N_9059,N_9263);
nor U11116 (N_11116,N_9206,N_9854);
nand U11117 (N_11117,N_9516,N_10487);
nor U11118 (N_11118,N_9417,N_9017);
or U11119 (N_11119,N_9174,N_9146);
and U11120 (N_11120,N_9455,N_10067);
and U11121 (N_11121,N_9035,N_9290);
and U11122 (N_11122,N_10213,N_10244);
or U11123 (N_11123,N_9541,N_9614);
and U11124 (N_11124,N_10321,N_9320);
nor U11125 (N_11125,N_9519,N_9538);
or U11126 (N_11126,N_10091,N_10021);
or U11127 (N_11127,N_9965,N_10284);
nor U11128 (N_11128,N_9701,N_9056);
and U11129 (N_11129,N_9769,N_10226);
nand U11130 (N_11130,N_10112,N_9178);
or U11131 (N_11131,N_10319,N_9439);
nor U11132 (N_11132,N_10424,N_9767);
nor U11133 (N_11133,N_9544,N_9890);
or U11134 (N_11134,N_9768,N_9086);
and U11135 (N_11135,N_10113,N_9640);
nand U11136 (N_11136,N_10293,N_9354);
nand U11137 (N_11137,N_10116,N_9285);
nand U11138 (N_11138,N_10072,N_9575);
nor U11139 (N_11139,N_10262,N_10436);
and U11140 (N_11140,N_9196,N_10097);
and U11141 (N_11141,N_9770,N_9849);
and U11142 (N_11142,N_9611,N_9994);
and U11143 (N_11143,N_10063,N_10137);
and U11144 (N_11144,N_9044,N_9716);
or U11145 (N_11145,N_10281,N_9405);
and U11146 (N_11146,N_9249,N_9988);
or U11147 (N_11147,N_10106,N_9376);
or U11148 (N_11148,N_10411,N_9808);
or U11149 (N_11149,N_10102,N_9492);
and U11150 (N_11150,N_9157,N_9445);
or U11151 (N_11151,N_9600,N_9220);
and U11152 (N_11152,N_10002,N_9349);
nand U11153 (N_11153,N_9663,N_9342);
nand U11154 (N_11154,N_9356,N_9053);
nor U11155 (N_11155,N_9654,N_10381);
nor U11156 (N_11156,N_9232,N_10362);
and U11157 (N_11157,N_10190,N_9162);
nor U11158 (N_11158,N_9566,N_9907);
and U11159 (N_11159,N_10055,N_9500);
and U11160 (N_11160,N_10047,N_9461);
and U11161 (N_11161,N_9929,N_9458);
and U11162 (N_11162,N_9424,N_9282);
nor U11163 (N_11163,N_9130,N_10014);
nor U11164 (N_11164,N_10220,N_10101);
nor U11165 (N_11165,N_10164,N_9447);
nor U11166 (N_11166,N_10001,N_9537);
and U11167 (N_11167,N_9217,N_9646);
and U11168 (N_11168,N_9046,N_10049);
nor U11169 (N_11169,N_9578,N_9795);
xnor U11170 (N_11170,N_9804,N_9974);
xnor U11171 (N_11171,N_9106,N_9914);
nand U11172 (N_11172,N_9288,N_9008);
and U11173 (N_11173,N_10259,N_9836);
nor U11174 (N_11174,N_9689,N_10452);
nor U11175 (N_11175,N_10405,N_9454);
nand U11176 (N_11176,N_9268,N_9679);
nor U11177 (N_11177,N_9892,N_10431);
or U11178 (N_11178,N_9589,N_9955);
nor U11179 (N_11179,N_9080,N_10301);
or U11180 (N_11180,N_9598,N_10198);
nor U11181 (N_11181,N_9877,N_9094);
or U11182 (N_11182,N_9296,N_10283);
or U11183 (N_11183,N_10218,N_10354);
and U11184 (N_11184,N_10160,N_10169);
xnor U11185 (N_11185,N_9783,N_9116);
nand U11186 (N_11186,N_10267,N_10427);
nor U11187 (N_11187,N_9421,N_9661);
and U11188 (N_11188,N_9060,N_9180);
or U11189 (N_11189,N_9428,N_10131);
nand U11190 (N_11190,N_9628,N_10349);
nor U11191 (N_11191,N_9152,N_9995);
or U11192 (N_11192,N_9970,N_10124);
nand U11193 (N_11193,N_9564,N_9386);
nor U11194 (N_11194,N_9678,N_10446);
nand U11195 (N_11195,N_10179,N_10042);
nor U11196 (N_11196,N_9861,N_9788);
nor U11197 (N_11197,N_9177,N_9859);
nor U11198 (N_11198,N_10122,N_9429);
and U11199 (N_11199,N_10135,N_9158);
nand U11200 (N_11200,N_9090,N_9784);
and U11201 (N_11201,N_9608,N_10426);
nor U11202 (N_11202,N_9913,N_10254);
or U11203 (N_11203,N_10174,N_9253);
nor U11204 (N_11204,N_9377,N_9789);
or U11205 (N_11205,N_10128,N_9048);
and U11206 (N_11206,N_9423,N_9512);
nand U11207 (N_11207,N_10086,N_9658);
nor U11208 (N_11208,N_9373,N_10273);
nor U11209 (N_11209,N_9510,N_9334);
nor U11210 (N_11210,N_9143,N_9385);
or U11211 (N_11211,N_9873,N_9765);
and U11212 (N_11212,N_9328,N_10217);
and U11213 (N_11213,N_9834,N_9826);
or U11214 (N_11214,N_9780,N_10363);
or U11215 (N_11215,N_9259,N_10224);
nor U11216 (N_11216,N_9314,N_9671);
nand U11217 (N_11217,N_9893,N_9703);
and U11218 (N_11218,N_9990,N_9426);
or U11219 (N_11219,N_10077,N_9926);
and U11220 (N_11220,N_10373,N_10114);
and U11221 (N_11221,N_10406,N_10229);
nor U11222 (N_11222,N_10059,N_10329);
or U11223 (N_11223,N_9691,N_9192);
nor U11224 (N_11224,N_9071,N_10238);
and U11225 (N_11225,N_10151,N_9984);
and U11226 (N_11226,N_9163,N_10322);
nand U11227 (N_11227,N_10210,N_9128);
nor U11228 (N_11228,N_10138,N_9450);
or U11229 (N_11229,N_9032,N_9602);
nand U11230 (N_11230,N_9353,N_10341);
nand U11231 (N_11231,N_10303,N_9392);
nor U11232 (N_11232,N_9092,N_10078);
nand U11233 (N_11233,N_9569,N_10442);
and U11234 (N_11234,N_9521,N_9563);
and U11235 (N_11235,N_9825,N_10207);
or U11236 (N_11236,N_9212,N_10027);
or U11237 (N_11237,N_10126,N_10357);
nor U11238 (N_11238,N_10050,N_9136);
nor U11239 (N_11239,N_9425,N_9005);
nor U11240 (N_11240,N_9416,N_10006);
nand U11241 (N_11241,N_10380,N_10459);
or U11242 (N_11242,N_9651,N_10295);
and U11243 (N_11243,N_9711,N_9270);
nor U11244 (N_11244,N_9364,N_9381);
nor U11245 (N_11245,N_10387,N_10296);
and U11246 (N_11246,N_10157,N_9818);
nor U11247 (N_11247,N_10004,N_9750);
xnor U11248 (N_11248,N_9706,N_9346);
or U11249 (N_11249,N_10043,N_9597);
nand U11250 (N_11250,N_9782,N_9914);
and U11251 (N_11251,N_9684,N_10076);
and U11252 (N_11252,N_9570,N_10014);
or U11253 (N_11253,N_9194,N_9697);
or U11254 (N_11254,N_9730,N_9273);
nand U11255 (N_11255,N_10166,N_9197);
nand U11256 (N_11256,N_9387,N_9763);
nand U11257 (N_11257,N_10435,N_9379);
or U11258 (N_11258,N_9786,N_9212);
nor U11259 (N_11259,N_9057,N_9098);
and U11260 (N_11260,N_9874,N_9851);
or U11261 (N_11261,N_9213,N_9414);
xnor U11262 (N_11262,N_9313,N_9881);
or U11263 (N_11263,N_10209,N_9697);
xnor U11264 (N_11264,N_9843,N_10322);
and U11265 (N_11265,N_10105,N_9265);
nand U11266 (N_11266,N_10481,N_9291);
or U11267 (N_11267,N_9159,N_10118);
or U11268 (N_11268,N_9506,N_9769);
nor U11269 (N_11269,N_9156,N_9693);
nand U11270 (N_11270,N_9442,N_9529);
nor U11271 (N_11271,N_9020,N_10044);
and U11272 (N_11272,N_10094,N_9203);
xor U11273 (N_11273,N_9720,N_9358);
and U11274 (N_11274,N_9302,N_10263);
nand U11275 (N_11275,N_10180,N_9365);
and U11276 (N_11276,N_9312,N_10391);
or U11277 (N_11277,N_9796,N_10117);
nor U11278 (N_11278,N_9350,N_9574);
nor U11279 (N_11279,N_9240,N_9549);
or U11280 (N_11280,N_9824,N_9173);
and U11281 (N_11281,N_9199,N_9061);
and U11282 (N_11282,N_9971,N_9859);
nand U11283 (N_11283,N_9406,N_10195);
or U11284 (N_11284,N_10050,N_9858);
nor U11285 (N_11285,N_10002,N_10054);
nor U11286 (N_11286,N_9991,N_10129);
or U11287 (N_11287,N_9146,N_9319);
and U11288 (N_11288,N_9785,N_9053);
and U11289 (N_11289,N_9415,N_9797);
and U11290 (N_11290,N_9705,N_10108);
or U11291 (N_11291,N_9675,N_9132);
nand U11292 (N_11292,N_10162,N_9730);
and U11293 (N_11293,N_9486,N_9237);
nor U11294 (N_11294,N_10190,N_10015);
or U11295 (N_11295,N_9031,N_9651);
nand U11296 (N_11296,N_10164,N_10012);
and U11297 (N_11297,N_9306,N_9199);
xor U11298 (N_11298,N_9501,N_9821);
and U11299 (N_11299,N_10260,N_9244);
and U11300 (N_11300,N_9189,N_10118);
and U11301 (N_11301,N_9895,N_9275);
nor U11302 (N_11302,N_9031,N_9015);
or U11303 (N_11303,N_9597,N_9176);
or U11304 (N_11304,N_10153,N_9074);
and U11305 (N_11305,N_10067,N_9957);
nor U11306 (N_11306,N_9989,N_9784);
nand U11307 (N_11307,N_10390,N_9005);
or U11308 (N_11308,N_9515,N_10100);
and U11309 (N_11309,N_9520,N_9780);
nand U11310 (N_11310,N_10348,N_9108);
nor U11311 (N_11311,N_10060,N_10131);
or U11312 (N_11312,N_10356,N_9677);
or U11313 (N_11313,N_9045,N_9274);
xor U11314 (N_11314,N_9186,N_9308);
and U11315 (N_11315,N_10144,N_9121);
and U11316 (N_11316,N_9445,N_10297);
nand U11317 (N_11317,N_10218,N_10397);
or U11318 (N_11318,N_9186,N_9325);
or U11319 (N_11319,N_10486,N_9710);
and U11320 (N_11320,N_10065,N_10276);
xor U11321 (N_11321,N_9752,N_9033);
or U11322 (N_11322,N_9313,N_9500);
or U11323 (N_11323,N_10365,N_9805);
nor U11324 (N_11324,N_9143,N_9827);
and U11325 (N_11325,N_9008,N_10446);
nand U11326 (N_11326,N_9479,N_9580);
or U11327 (N_11327,N_9194,N_9284);
nand U11328 (N_11328,N_9561,N_9214);
nor U11329 (N_11329,N_9066,N_10336);
nor U11330 (N_11330,N_10091,N_9171);
nand U11331 (N_11331,N_9153,N_10025);
nor U11332 (N_11332,N_9485,N_9643);
xor U11333 (N_11333,N_9785,N_10490);
nor U11334 (N_11334,N_9355,N_10130);
and U11335 (N_11335,N_10276,N_10139);
or U11336 (N_11336,N_9661,N_9255);
nand U11337 (N_11337,N_9503,N_9131);
nor U11338 (N_11338,N_10121,N_10434);
or U11339 (N_11339,N_10341,N_10046);
nand U11340 (N_11340,N_10109,N_9474);
nor U11341 (N_11341,N_9165,N_10486);
or U11342 (N_11342,N_9655,N_10415);
and U11343 (N_11343,N_10482,N_9777);
xnor U11344 (N_11344,N_9998,N_9295);
nor U11345 (N_11345,N_10329,N_10314);
nor U11346 (N_11346,N_9828,N_10464);
or U11347 (N_11347,N_10324,N_9077);
and U11348 (N_11348,N_9744,N_10091);
nand U11349 (N_11349,N_10463,N_9619);
or U11350 (N_11350,N_9482,N_10145);
nor U11351 (N_11351,N_9912,N_9019);
and U11352 (N_11352,N_10492,N_9820);
and U11353 (N_11353,N_9445,N_9001);
nor U11354 (N_11354,N_9040,N_9076);
nor U11355 (N_11355,N_10391,N_9818);
nand U11356 (N_11356,N_9416,N_9878);
nor U11357 (N_11357,N_9757,N_10406);
nand U11358 (N_11358,N_9708,N_10420);
and U11359 (N_11359,N_9689,N_9928);
or U11360 (N_11360,N_9338,N_9174);
or U11361 (N_11361,N_9131,N_9095);
and U11362 (N_11362,N_9642,N_9615);
or U11363 (N_11363,N_9978,N_9835);
nor U11364 (N_11364,N_9652,N_10276);
or U11365 (N_11365,N_9297,N_10451);
nor U11366 (N_11366,N_9095,N_10449);
xor U11367 (N_11367,N_10452,N_10364);
or U11368 (N_11368,N_10396,N_10024);
or U11369 (N_11369,N_9814,N_10068);
nor U11370 (N_11370,N_10380,N_9791);
nor U11371 (N_11371,N_9718,N_9226);
nor U11372 (N_11372,N_9379,N_9492);
or U11373 (N_11373,N_9846,N_9686);
nand U11374 (N_11374,N_9790,N_10191);
nor U11375 (N_11375,N_9626,N_10357);
and U11376 (N_11376,N_9780,N_9393);
nand U11377 (N_11377,N_10282,N_10162);
and U11378 (N_11378,N_9988,N_9104);
or U11379 (N_11379,N_10167,N_9242);
and U11380 (N_11380,N_9838,N_9433);
nand U11381 (N_11381,N_10381,N_9619);
nor U11382 (N_11382,N_9928,N_9835);
nor U11383 (N_11383,N_10026,N_9567);
and U11384 (N_11384,N_9778,N_10247);
nand U11385 (N_11385,N_10301,N_9247);
nand U11386 (N_11386,N_9112,N_9675);
nor U11387 (N_11387,N_10201,N_9236);
or U11388 (N_11388,N_9909,N_9010);
nand U11389 (N_11389,N_10274,N_9478);
or U11390 (N_11390,N_9392,N_10107);
nor U11391 (N_11391,N_9549,N_10405);
and U11392 (N_11392,N_9234,N_10118);
nor U11393 (N_11393,N_9994,N_10367);
nor U11394 (N_11394,N_10470,N_9974);
nand U11395 (N_11395,N_9323,N_9463);
or U11396 (N_11396,N_9903,N_10147);
nor U11397 (N_11397,N_9706,N_9154);
nand U11398 (N_11398,N_9772,N_9291);
and U11399 (N_11399,N_9411,N_9464);
and U11400 (N_11400,N_9347,N_9187);
or U11401 (N_11401,N_10283,N_10217);
or U11402 (N_11402,N_9522,N_10024);
nand U11403 (N_11403,N_9113,N_10056);
and U11404 (N_11404,N_9682,N_10400);
nor U11405 (N_11405,N_9428,N_9868);
and U11406 (N_11406,N_9874,N_9237);
nand U11407 (N_11407,N_9020,N_10280);
or U11408 (N_11408,N_10206,N_9699);
or U11409 (N_11409,N_9112,N_9418);
nor U11410 (N_11410,N_9722,N_9262);
or U11411 (N_11411,N_9821,N_9631);
nor U11412 (N_11412,N_9309,N_9947);
nand U11413 (N_11413,N_10328,N_10103);
nand U11414 (N_11414,N_9805,N_9132);
or U11415 (N_11415,N_9040,N_9936);
and U11416 (N_11416,N_10172,N_9844);
nand U11417 (N_11417,N_9118,N_9038);
nor U11418 (N_11418,N_9139,N_9929);
and U11419 (N_11419,N_9729,N_10246);
nand U11420 (N_11420,N_9004,N_9673);
nor U11421 (N_11421,N_10322,N_10418);
or U11422 (N_11422,N_9134,N_9721);
and U11423 (N_11423,N_10254,N_9953);
and U11424 (N_11424,N_9913,N_9809);
nor U11425 (N_11425,N_9512,N_9201);
nor U11426 (N_11426,N_10114,N_10379);
or U11427 (N_11427,N_10323,N_10158);
nand U11428 (N_11428,N_9861,N_10194);
nor U11429 (N_11429,N_9855,N_9917);
and U11430 (N_11430,N_9960,N_10002);
or U11431 (N_11431,N_10068,N_10037);
nand U11432 (N_11432,N_9513,N_9129);
nand U11433 (N_11433,N_10279,N_10153);
nand U11434 (N_11434,N_9595,N_10252);
or U11435 (N_11435,N_9931,N_9143);
nand U11436 (N_11436,N_9239,N_9339);
nand U11437 (N_11437,N_9257,N_9674);
or U11438 (N_11438,N_10253,N_9442);
nand U11439 (N_11439,N_9659,N_9418);
xnor U11440 (N_11440,N_9293,N_9460);
nor U11441 (N_11441,N_9025,N_9894);
or U11442 (N_11442,N_9346,N_10079);
and U11443 (N_11443,N_9831,N_9136);
nor U11444 (N_11444,N_9234,N_10302);
and U11445 (N_11445,N_10062,N_9783);
or U11446 (N_11446,N_9451,N_9755);
nand U11447 (N_11447,N_10281,N_9161);
and U11448 (N_11448,N_9359,N_9083);
or U11449 (N_11449,N_9467,N_10111);
or U11450 (N_11450,N_9340,N_10490);
nand U11451 (N_11451,N_9812,N_9451);
or U11452 (N_11452,N_9441,N_10158);
nor U11453 (N_11453,N_9405,N_10303);
nor U11454 (N_11454,N_9099,N_9432);
nand U11455 (N_11455,N_9299,N_9833);
or U11456 (N_11456,N_10181,N_9509);
nor U11457 (N_11457,N_9201,N_9434);
and U11458 (N_11458,N_9342,N_9878);
or U11459 (N_11459,N_10483,N_9290);
nand U11460 (N_11460,N_9611,N_9794);
or U11461 (N_11461,N_9462,N_10018);
nor U11462 (N_11462,N_9491,N_9533);
and U11463 (N_11463,N_9619,N_10435);
nor U11464 (N_11464,N_10167,N_9448);
nand U11465 (N_11465,N_10212,N_9060);
or U11466 (N_11466,N_9577,N_9546);
nand U11467 (N_11467,N_10271,N_10471);
or U11468 (N_11468,N_10136,N_9710);
and U11469 (N_11469,N_9331,N_9847);
nor U11470 (N_11470,N_9361,N_9998);
and U11471 (N_11471,N_9702,N_9712);
and U11472 (N_11472,N_9232,N_9735);
nor U11473 (N_11473,N_9430,N_10314);
nor U11474 (N_11474,N_10279,N_9024);
nand U11475 (N_11475,N_9091,N_10326);
or U11476 (N_11476,N_9774,N_9303);
and U11477 (N_11477,N_9578,N_9463);
and U11478 (N_11478,N_10397,N_9029);
nand U11479 (N_11479,N_10420,N_9896);
and U11480 (N_11480,N_9101,N_9149);
nor U11481 (N_11481,N_10241,N_10345);
or U11482 (N_11482,N_9621,N_10309);
nand U11483 (N_11483,N_9147,N_9128);
or U11484 (N_11484,N_9157,N_9647);
nand U11485 (N_11485,N_9642,N_9461);
or U11486 (N_11486,N_9519,N_9550);
xor U11487 (N_11487,N_10149,N_9073);
nor U11488 (N_11488,N_10280,N_10176);
or U11489 (N_11489,N_9395,N_9852);
xor U11490 (N_11490,N_9486,N_10148);
and U11491 (N_11491,N_9677,N_9753);
nor U11492 (N_11492,N_9841,N_9906);
and U11493 (N_11493,N_9872,N_9212);
and U11494 (N_11494,N_9295,N_9061);
nor U11495 (N_11495,N_9660,N_10445);
or U11496 (N_11496,N_9541,N_9013);
or U11497 (N_11497,N_9625,N_9796);
or U11498 (N_11498,N_9268,N_9843);
or U11499 (N_11499,N_9333,N_9962);
and U11500 (N_11500,N_9206,N_9318);
nor U11501 (N_11501,N_9719,N_10245);
and U11502 (N_11502,N_9732,N_9594);
nor U11503 (N_11503,N_9257,N_10321);
and U11504 (N_11504,N_9651,N_9389);
nor U11505 (N_11505,N_9489,N_9211);
nor U11506 (N_11506,N_9958,N_10497);
and U11507 (N_11507,N_9197,N_10369);
or U11508 (N_11508,N_10012,N_9222);
xnor U11509 (N_11509,N_9183,N_9481);
nand U11510 (N_11510,N_9810,N_9107);
nor U11511 (N_11511,N_9705,N_9831);
nor U11512 (N_11512,N_9275,N_9554);
nor U11513 (N_11513,N_10439,N_10469);
or U11514 (N_11514,N_10400,N_10019);
and U11515 (N_11515,N_10283,N_9508);
nor U11516 (N_11516,N_10071,N_9371);
nor U11517 (N_11517,N_10084,N_9385);
nor U11518 (N_11518,N_9490,N_10323);
and U11519 (N_11519,N_9642,N_10444);
nand U11520 (N_11520,N_9496,N_10408);
nor U11521 (N_11521,N_9318,N_9419);
and U11522 (N_11522,N_9459,N_10156);
or U11523 (N_11523,N_9227,N_10249);
and U11524 (N_11524,N_10090,N_9369);
nor U11525 (N_11525,N_10121,N_9430);
nor U11526 (N_11526,N_9594,N_10419);
and U11527 (N_11527,N_9852,N_10051);
nand U11528 (N_11528,N_10257,N_9176);
or U11529 (N_11529,N_9317,N_10198);
nand U11530 (N_11530,N_10177,N_10365);
nor U11531 (N_11531,N_9882,N_9942);
or U11532 (N_11532,N_10387,N_9598);
and U11533 (N_11533,N_9889,N_10055);
nor U11534 (N_11534,N_10068,N_9029);
and U11535 (N_11535,N_9794,N_9987);
xor U11536 (N_11536,N_9124,N_9237);
or U11537 (N_11537,N_10072,N_9258);
or U11538 (N_11538,N_9855,N_9051);
nor U11539 (N_11539,N_10330,N_9985);
nor U11540 (N_11540,N_9965,N_9367);
nand U11541 (N_11541,N_9779,N_9738);
and U11542 (N_11542,N_9426,N_9613);
or U11543 (N_11543,N_10310,N_10401);
nand U11544 (N_11544,N_9835,N_9862);
or U11545 (N_11545,N_9243,N_9705);
and U11546 (N_11546,N_9093,N_10079);
or U11547 (N_11547,N_9448,N_9834);
nor U11548 (N_11548,N_9325,N_9934);
xor U11549 (N_11549,N_10180,N_9789);
nor U11550 (N_11550,N_9587,N_9760);
and U11551 (N_11551,N_10065,N_9806);
nand U11552 (N_11552,N_10184,N_9383);
or U11553 (N_11553,N_9369,N_10472);
nor U11554 (N_11554,N_9398,N_9166);
or U11555 (N_11555,N_9416,N_9082);
nand U11556 (N_11556,N_9847,N_9023);
and U11557 (N_11557,N_9637,N_9034);
nand U11558 (N_11558,N_9598,N_9506);
nand U11559 (N_11559,N_9757,N_10294);
nand U11560 (N_11560,N_9354,N_9727);
and U11561 (N_11561,N_9316,N_9105);
and U11562 (N_11562,N_9291,N_9430);
and U11563 (N_11563,N_9779,N_10430);
or U11564 (N_11564,N_9977,N_9295);
nand U11565 (N_11565,N_9272,N_9108);
or U11566 (N_11566,N_9667,N_9699);
and U11567 (N_11567,N_9839,N_10439);
nand U11568 (N_11568,N_10008,N_10198);
nand U11569 (N_11569,N_9375,N_9954);
nor U11570 (N_11570,N_9980,N_9770);
or U11571 (N_11571,N_9561,N_10046);
nand U11572 (N_11572,N_10003,N_9508);
and U11573 (N_11573,N_10479,N_9065);
nand U11574 (N_11574,N_10209,N_9112);
nand U11575 (N_11575,N_9009,N_9448);
and U11576 (N_11576,N_10340,N_9878);
and U11577 (N_11577,N_9395,N_10046);
nor U11578 (N_11578,N_10123,N_9939);
nor U11579 (N_11579,N_10069,N_9399);
xnor U11580 (N_11580,N_10300,N_9302);
or U11581 (N_11581,N_9904,N_9124);
and U11582 (N_11582,N_9270,N_9293);
nor U11583 (N_11583,N_9994,N_9766);
or U11584 (N_11584,N_9670,N_10121);
and U11585 (N_11585,N_10179,N_9742);
nor U11586 (N_11586,N_10233,N_9038);
or U11587 (N_11587,N_9443,N_9301);
and U11588 (N_11588,N_9389,N_9747);
and U11589 (N_11589,N_9215,N_10073);
or U11590 (N_11590,N_9915,N_9546);
and U11591 (N_11591,N_9044,N_10108);
nand U11592 (N_11592,N_9773,N_10375);
or U11593 (N_11593,N_10098,N_9325);
nor U11594 (N_11594,N_9887,N_9509);
and U11595 (N_11595,N_9087,N_9794);
or U11596 (N_11596,N_9226,N_10439);
or U11597 (N_11597,N_9929,N_9716);
nand U11598 (N_11598,N_9195,N_9567);
and U11599 (N_11599,N_10131,N_9777);
nand U11600 (N_11600,N_9901,N_9655);
nand U11601 (N_11601,N_9870,N_9528);
or U11602 (N_11602,N_9778,N_10326);
nand U11603 (N_11603,N_9138,N_9055);
or U11604 (N_11604,N_10336,N_10113);
nand U11605 (N_11605,N_9580,N_9954);
or U11606 (N_11606,N_10212,N_9822);
or U11607 (N_11607,N_9935,N_9934);
xor U11608 (N_11608,N_9220,N_10405);
or U11609 (N_11609,N_9914,N_9857);
or U11610 (N_11610,N_9748,N_9020);
or U11611 (N_11611,N_9319,N_9685);
nand U11612 (N_11612,N_10217,N_9705);
nor U11613 (N_11613,N_9240,N_9736);
and U11614 (N_11614,N_10260,N_9522);
and U11615 (N_11615,N_10266,N_9704);
or U11616 (N_11616,N_10394,N_10311);
or U11617 (N_11617,N_9304,N_9034);
nor U11618 (N_11618,N_9674,N_9101);
nor U11619 (N_11619,N_10401,N_10159);
or U11620 (N_11620,N_10414,N_9771);
and U11621 (N_11621,N_9661,N_9720);
or U11622 (N_11622,N_10163,N_9375);
xor U11623 (N_11623,N_9292,N_10045);
or U11624 (N_11624,N_9158,N_9604);
or U11625 (N_11625,N_10246,N_9698);
or U11626 (N_11626,N_9620,N_10058);
and U11627 (N_11627,N_9893,N_10068);
nor U11628 (N_11628,N_10184,N_10259);
nand U11629 (N_11629,N_9780,N_10367);
nand U11630 (N_11630,N_9774,N_9341);
nor U11631 (N_11631,N_10326,N_9732);
nand U11632 (N_11632,N_9322,N_9328);
nor U11633 (N_11633,N_9079,N_9857);
nor U11634 (N_11634,N_9941,N_10148);
nand U11635 (N_11635,N_10090,N_9371);
or U11636 (N_11636,N_9361,N_9418);
and U11637 (N_11637,N_9552,N_9989);
and U11638 (N_11638,N_9806,N_10452);
nor U11639 (N_11639,N_9212,N_9298);
and U11640 (N_11640,N_9093,N_10311);
and U11641 (N_11641,N_9820,N_9742);
or U11642 (N_11642,N_9586,N_9205);
or U11643 (N_11643,N_10166,N_10347);
nor U11644 (N_11644,N_9119,N_9250);
nor U11645 (N_11645,N_9872,N_9676);
nand U11646 (N_11646,N_9452,N_10028);
and U11647 (N_11647,N_10376,N_10369);
nor U11648 (N_11648,N_9463,N_9003);
and U11649 (N_11649,N_10145,N_10384);
and U11650 (N_11650,N_9641,N_10235);
nand U11651 (N_11651,N_9538,N_9530);
nor U11652 (N_11652,N_10446,N_10087);
nand U11653 (N_11653,N_9137,N_9380);
nand U11654 (N_11654,N_9321,N_9000);
or U11655 (N_11655,N_10221,N_9928);
nor U11656 (N_11656,N_10101,N_9716);
nor U11657 (N_11657,N_9160,N_9780);
xnor U11658 (N_11658,N_9794,N_9763);
and U11659 (N_11659,N_9573,N_9138);
or U11660 (N_11660,N_9769,N_9603);
nand U11661 (N_11661,N_9444,N_10341);
nor U11662 (N_11662,N_9045,N_10125);
nand U11663 (N_11663,N_9110,N_9045);
or U11664 (N_11664,N_9388,N_9047);
and U11665 (N_11665,N_9309,N_9786);
and U11666 (N_11666,N_10340,N_9575);
nor U11667 (N_11667,N_9633,N_10014);
or U11668 (N_11668,N_10460,N_9481);
nor U11669 (N_11669,N_10160,N_10212);
nand U11670 (N_11670,N_9717,N_9138);
nand U11671 (N_11671,N_9881,N_9042);
and U11672 (N_11672,N_9385,N_9630);
and U11673 (N_11673,N_9597,N_9787);
and U11674 (N_11674,N_9948,N_9346);
and U11675 (N_11675,N_9694,N_9722);
or U11676 (N_11676,N_10301,N_9541);
nor U11677 (N_11677,N_9229,N_10170);
and U11678 (N_11678,N_9977,N_9208);
and U11679 (N_11679,N_10076,N_10077);
or U11680 (N_11680,N_9110,N_9030);
and U11681 (N_11681,N_9947,N_9286);
or U11682 (N_11682,N_10306,N_9197);
nand U11683 (N_11683,N_9658,N_9774);
nand U11684 (N_11684,N_9907,N_9048);
nor U11685 (N_11685,N_9017,N_9455);
or U11686 (N_11686,N_9414,N_9694);
nand U11687 (N_11687,N_10475,N_10328);
nand U11688 (N_11688,N_9966,N_10113);
nor U11689 (N_11689,N_10339,N_9199);
or U11690 (N_11690,N_9782,N_10115);
nor U11691 (N_11691,N_9655,N_9473);
nor U11692 (N_11692,N_9607,N_10017);
nand U11693 (N_11693,N_9476,N_9062);
or U11694 (N_11694,N_9210,N_10042);
xor U11695 (N_11695,N_10393,N_10271);
and U11696 (N_11696,N_10287,N_9472);
nand U11697 (N_11697,N_10421,N_10067);
or U11698 (N_11698,N_9466,N_9183);
and U11699 (N_11699,N_10143,N_9005);
and U11700 (N_11700,N_9236,N_9526);
nor U11701 (N_11701,N_9854,N_9552);
and U11702 (N_11702,N_9376,N_9110);
and U11703 (N_11703,N_10305,N_10009);
or U11704 (N_11704,N_10247,N_10225);
nor U11705 (N_11705,N_9100,N_9728);
nand U11706 (N_11706,N_9019,N_9536);
and U11707 (N_11707,N_10476,N_10238);
or U11708 (N_11708,N_10238,N_9562);
nor U11709 (N_11709,N_9832,N_9192);
nand U11710 (N_11710,N_9993,N_9991);
and U11711 (N_11711,N_9104,N_10187);
nand U11712 (N_11712,N_9598,N_9549);
nand U11713 (N_11713,N_9279,N_9176);
nor U11714 (N_11714,N_10254,N_9483);
nand U11715 (N_11715,N_9319,N_9642);
nor U11716 (N_11716,N_9623,N_9277);
xor U11717 (N_11717,N_10225,N_9129);
nor U11718 (N_11718,N_9310,N_10030);
or U11719 (N_11719,N_9313,N_10414);
nor U11720 (N_11720,N_9867,N_10102);
nor U11721 (N_11721,N_9154,N_9148);
and U11722 (N_11722,N_9381,N_10290);
or U11723 (N_11723,N_10201,N_10449);
or U11724 (N_11724,N_10394,N_10383);
and U11725 (N_11725,N_9429,N_9940);
xnor U11726 (N_11726,N_9850,N_9958);
nand U11727 (N_11727,N_9873,N_10133);
nor U11728 (N_11728,N_9089,N_9693);
nand U11729 (N_11729,N_9613,N_9842);
or U11730 (N_11730,N_10108,N_10413);
or U11731 (N_11731,N_10411,N_9728);
nand U11732 (N_11732,N_9968,N_9243);
nand U11733 (N_11733,N_9315,N_9651);
nor U11734 (N_11734,N_10065,N_9140);
nand U11735 (N_11735,N_9509,N_9653);
and U11736 (N_11736,N_10443,N_9443);
nor U11737 (N_11737,N_9244,N_9928);
and U11738 (N_11738,N_9415,N_10287);
nor U11739 (N_11739,N_9082,N_9705);
xnor U11740 (N_11740,N_9407,N_9475);
or U11741 (N_11741,N_9165,N_9302);
and U11742 (N_11742,N_10024,N_9283);
nor U11743 (N_11743,N_9226,N_9780);
nor U11744 (N_11744,N_10471,N_9124);
nor U11745 (N_11745,N_9675,N_9594);
nor U11746 (N_11746,N_9077,N_9949);
nand U11747 (N_11747,N_10083,N_10216);
nor U11748 (N_11748,N_10137,N_9683);
nor U11749 (N_11749,N_9058,N_9123);
or U11750 (N_11750,N_9469,N_10024);
and U11751 (N_11751,N_9316,N_9811);
xnor U11752 (N_11752,N_10001,N_9830);
nand U11753 (N_11753,N_9419,N_10396);
or U11754 (N_11754,N_9878,N_10468);
xor U11755 (N_11755,N_10411,N_10376);
nor U11756 (N_11756,N_9232,N_9008);
nor U11757 (N_11757,N_10107,N_10366);
nor U11758 (N_11758,N_9590,N_9064);
nand U11759 (N_11759,N_9935,N_9411);
nand U11760 (N_11760,N_9652,N_9350);
or U11761 (N_11761,N_9089,N_10468);
nand U11762 (N_11762,N_10251,N_10160);
or U11763 (N_11763,N_9496,N_10335);
xnor U11764 (N_11764,N_9092,N_9659);
nand U11765 (N_11765,N_10275,N_10281);
or U11766 (N_11766,N_10481,N_9779);
nor U11767 (N_11767,N_9052,N_9238);
nor U11768 (N_11768,N_9959,N_10218);
or U11769 (N_11769,N_9422,N_9800);
and U11770 (N_11770,N_9232,N_9663);
or U11771 (N_11771,N_9627,N_9499);
and U11772 (N_11772,N_9519,N_9399);
or U11773 (N_11773,N_9122,N_9113);
nor U11774 (N_11774,N_9564,N_9634);
nor U11775 (N_11775,N_9991,N_9589);
nand U11776 (N_11776,N_9299,N_10236);
xnor U11777 (N_11777,N_9493,N_9594);
and U11778 (N_11778,N_10470,N_9093);
nor U11779 (N_11779,N_9652,N_9044);
or U11780 (N_11780,N_10297,N_9292);
and U11781 (N_11781,N_9048,N_9618);
nor U11782 (N_11782,N_10491,N_9010);
nor U11783 (N_11783,N_9644,N_10344);
or U11784 (N_11784,N_9562,N_9303);
nor U11785 (N_11785,N_10422,N_10031);
nand U11786 (N_11786,N_9253,N_9514);
nand U11787 (N_11787,N_9363,N_9782);
nand U11788 (N_11788,N_9601,N_9897);
or U11789 (N_11789,N_9549,N_10013);
and U11790 (N_11790,N_9270,N_9948);
nor U11791 (N_11791,N_10308,N_9657);
and U11792 (N_11792,N_9763,N_10076);
nand U11793 (N_11793,N_9384,N_9714);
nor U11794 (N_11794,N_10148,N_9715);
nor U11795 (N_11795,N_9890,N_9010);
xnor U11796 (N_11796,N_9907,N_9547);
and U11797 (N_11797,N_9974,N_9839);
nand U11798 (N_11798,N_9947,N_9962);
nor U11799 (N_11799,N_9592,N_9776);
or U11800 (N_11800,N_10324,N_9700);
and U11801 (N_11801,N_9175,N_9816);
xnor U11802 (N_11802,N_10035,N_10190);
nor U11803 (N_11803,N_10051,N_10011);
and U11804 (N_11804,N_9442,N_10409);
or U11805 (N_11805,N_9666,N_9069);
or U11806 (N_11806,N_10383,N_9640);
nor U11807 (N_11807,N_10175,N_10268);
nand U11808 (N_11808,N_9856,N_9470);
xnor U11809 (N_11809,N_10190,N_9663);
and U11810 (N_11810,N_9554,N_9667);
nand U11811 (N_11811,N_9702,N_9337);
nor U11812 (N_11812,N_9111,N_10145);
nand U11813 (N_11813,N_9141,N_9626);
or U11814 (N_11814,N_10461,N_10002);
nor U11815 (N_11815,N_9756,N_9451);
and U11816 (N_11816,N_10162,N_10183);
nand U11817 (N_11817,N_10204,N_10008);
nor U11818 (N_11818,N_9917,N_9115);
and U11819 (N_11819,N_10461,N_10419);
nand U11820 (N_11820,N_9850,N_10099);
or U11821 (N_11821,N_9555,N_9803);
nand U11822 (N_11822,N_9272,N_9380);
nor U11823 (N_11823,N_9869,N_9683);
or U11824 (N_11824,N_10075,N_9624);
or U11825 (N_11825,N_10440,N_10029);
nor U11826 (N_11826,N_9011,N_9882);
nor U11827 (N_11827,N_9866,N_9913);
and U11828 (N_11828,N_9278,N_9484);
and U11829 (N_11829,N_9428,N_9418);
nand U11830 (N_11830,N_10096,N_10370);
or U11831 (N_11831,N_10263,N_10152);
nand U11832 (N_11832,N_10147,N_9275);
and U11833 (N_11833,N_9602,N_9572);
or U11834 (N_11834,N_9098,N_9028);
and U11835 (N_11835,N_9843,N_9158);
or U11836 (N_11836,N_9536,N_10045);
and U11837 (N_11837,N_9169,N_9332);
and U11838 (N_11838,N_9838,N_9459);
or U11839 (N_11839,N_9198,N_9979);
nor U11840 (N_11840,N_10301,N_9206);
nand U11841 (N_11841,N_9501,N_9926);
nand U11842 (N_11842,N_10095,N_9217);
or U11843 (N_11843,N_9526,N_10129);
nand U11844 (N_11844,N_10422,N_10093);
nand U11845 (N_11845,N_9450,N_9711);
nand U11846 (N_11846,N_10334,N_10285);
nor U11847 (N_11847,N_10097,N_9682);
nand U11848 (N_11848,N_10030,N_9877);
nor U11849 (N_11849,N_10492,N_9837);
nand U11850 (N_11850,N_9599,N_9474);
and U11851 (N_11851,N_9067,N_10140);
nor U11852 (N_11852,N_10350,N_9673);
nand U11853 (N_11853,N_10075,N_9350);
and U11854 (N_11854,N_9017,N_10126);
nor U11855 (N_11855,N_9025,N_9635);
and U11856 (N_11856,N_10460,N_9284);
nand U11857 (N_11857,N_9739,N_9582);
and U11858 (N_11858,N_9132,N_9753);
nor U11859 (N_11859,N_9068,N_10131);
and U11860 (N_11860,N_10309,N_10150);
nand U11861 (N_11861,N_10015,N_9860);
xor U11862 (N_11862,N_9575,N_9660);
nand U11863 (N_11863,N_10105,N_9347);
and U11864 (N_11864,N_9505,N_10089);
and U11865 (N_11865,N_9667,N_9774);
or U11866 (N_11866,N_9102,N_10306);
nor U11867 (N_11867,N_10250,N_9477);
or U11868 (N_11868,N_9927,N_9112);
and U11869 (N_11869,N_10124,N_9492);
or U11870 (N_11870,N_9221,N_10013);
and U11871 (N_11871,N_10437,N_9335);
or U11872 (N_11872,N_9164,N_9023);
and U11873 (N_11873,N_10203,N_10208);
or U11874 (N_11874,N_10183,N_9710);
nor U11875 (N_11875,N_10075,N_9203);
and U11876 (N_11876,N_10439,N_9125);
or U11877 (N_11877,N_10409,N_10232);
and U11878 (N_11878,N_9317,N_9011);
and U11879 (N_11879,N_9737,N_9639);
nand U11880 (N_11880,N_9373,N_9021);
nand U11881 (N_11881,N_9923,N_10472);
and U11882 (N_11882,N_9671,N_9722);
or U11883 (N_11883,N_9699,N_9802);
or U11884 (N_11884,N_10297,N_9755);
or U11885 (N_11885,N_9839,N_9536);
and U11886 (N_11886,N_10351,N_10440);
xor U11887 (N_11887,N_9400,N_10465);
or U11888 (N_11888,N_9630,N_9773);
or U11889 (N_11889,N_9328,N_9064);
or U11890 (N_11890,N_9555,N_9676);
and U11891 (N_11891,N_9665,N_9766);
nand U11892 (N_11892,N_9331,N_9997);
or U11893 (N_11893,N_9824,N_9904);
nor U11894 (N_11894,N_9748,N_9106);
or U11895 (N_11895,N_9504,N_9841);
nand U11896 (N_11896,N_10206,N_10147);
and U11897 (N_11897,N_9839,N_10231);
xnor U11898 (N_11898,N_9113,N_9428);
nor U11899 (N_11899,N_9821,N_9355);
and U11900 (N_11900,N_10167,N_10425);
nor U11901 (N_11901,N_9840,N_10471);
nand U11902 (N_11902,N_9584,N_9353);
and U11903 (N_11903,N_10017,N_9295);
and U11904 (N_11904,N_9415,N_10161);
nor U11905 (N_11905,N_10433,N_10408);
nor U11906 (N_11906,N_9832,N_10439);
nand U11907 (N_11907,N_9846,N_10242);
and U11908 (N_11908,N_9024,N_9414);
and U11909 (N_11909,N_10213,N_9420);
nand U11910 (N_11910,N_10272,N_10082);
and U11911 (N_11911,N_9151,N_10361);
nand U11912 (N_11912,N_10498,N_9192);
nand U11913 (N_11913,N_10406,N_9566);
nor U11914 (N_11914,N_9070,N_9127);
and U11915 (N_11915,N_9539,N_9608);
nand U11916 (N_11916,N_9917,N_9018);
nor U11917 (N_11917,N_10436,N_9581);
nand U11918 (N_11918,N_9461,N_10387);
nor U11919 (N_11919,N_9176,N_9949);
xor U11920 (N_11920,N_10119,N_10200);
nor U11921 (N_11921,N_9133,N_9892);
nor U11922 (N_11922,N_9090,N_10202);
and U11923 (N_11923,N_10040,N_9202);
and U11924 (N_11924,N_10042,N_9594);
nor U11925 (N_11925,N_10218,N_10310);
nor U11926 (N_11926,N_10378,N_9800);
nand U11927 (N_11927,N_9373,N_9659);
nand U11928 (N_11928,N_9469,N_10091);
and U11929 (N_11929,N_9371,N_10308);
or U11930 (N_11930,N_9352,N_9743);
nand U11931 (N_11931,N_10177,N_10443);
and U11932 (N_11932,N_10307,N_9340);
nand U11933 (N_11933,N_9616,N_9916);
nand U11934 (N_11934,N_10194,N_9268);
nand U11935 (N_11935,N_9576,N_10454);
or U11936 (N_11936,N_9430,N_9247);
or U11937 (N_11937,N_9385,N_9030);
nand U11938 (N_11938,N_9036,N_9880);
nand U11939 (N_11939,N_9925,N_10490);
nor U11940 (N_11940,N_10438,N_9749);
or U11941 (N_11941,N_9249,N_10289);
or U11942 (N_11942,N_9004,N_9202);
nand U11943 (N_11943,N_10120,N_10307);
nor U11944 (N_11944,N_10420,N_9965);
nor U11945 (N_11945,N_9977,N_10134);
and U11946 (N_11946,N_10391,N_10045);
and U11947 (N_11947,N_9592,N_9188);
and U11948 (N_11948,N_10448,N_9710);
and U11949 (N_11949,N_9743,N_10154);
and U11950 (N_11950,N_9661,N_10077);
or U11951 (N_11951,N_9356,N_9786);
or U11952 (N_11952,N_9748,N_9656);
nor U11953 (N_11953,N_9057,N_9327);
nor U11954 (N_11954,N_10326,N_10480);
nor U11955 (N_11955,N_10081,N_10061);
and U11956 (N_11956,N_9468,N_9862);
and U11957 (N_11957,N_9796,N_10340);
and U11958 (N_11958,N_9254,N_9478);
or U11959 (N_11959,N_9397,N_9334);
or U11960 (N_11960,N_10067,N_9345);
nand U11961 (N_11961,N_9695,N_9879);
nor U11962 (N_11962,N_9132,N_10096);
nor U11963 (N_11963,N_10263,N_9560);
nand U11964 (N_11964,N_9474,N_9552);
nand U11965 (N_11965,N_9866,N_9529);
nor U11966 (N_11966,N_9878,N_9758);
nand U11967 (N_11967,N_9549,N_9238);
and U11968 (N_11968,N_9487,N_9519);
nor U11969 (N_11969,N_9458,N_10200);
or U11970 (N_11970,N_9497,N_9891);
and U11971 (N_11971,N_9520,N_9270);
and U11972 (N_11972,N_9984,N_9396);
nand U11973 (N_11973,N_10365,N_10170);
or U11974 (N_11974,N_9958,N_9484);
nor U11975 (N_11975,N_10097,N_9539);
nand U11976 (N_11976,N_10272,N_10410);
and U11977 (N_11977,N_10037,N_9137);
nand U11978 (N_11978,N_10338,N_9969);
and U11979 (N_11979,N_9096,N_9153);
and U11980 (N_11980,N_9860,N_9256);
nand U11981 (N_11981,N_9488,N_9410);
or U11982 (N_11982,N_9959,N_10386);
nand U11983 (N_11983,N_9971,N_9972);
nand U11984 (N_11984,N_10147,N_10256);
or U11985 (N_11985,N_9245,N_9138);
nand U11986 (N_11986,N_10363,N_9169);
nand U11987 (N_11987,N_10251,N_9782);
or U11988 (N_11988,N_9862,N_10280);
and U11989 (N_11989,N_9449,N_10256);
nand U11990 (N_11990,N_10308,N_10047);
and U11991 (N_11991,N_10056,N_9823);
nand U11992 (N_11992,N_9606,N_9294);
or U11993 (N_11993,N_9193,N_9361);
nand U11994 (N_11994,N_9386,N_9767);
and U11995 (N_11995,N_9278,N_10394);
nand U11996 (N_11996,N_10332,N_9805);
nand U11997 (N_11997,N_10447,N_9712);
nand U11998 (N_11998,N_9797,N_9441);
nor U11999 (N_11999,N_9128,N_9780);
and U12000 (N_12000,N_11224,N_10519);
and U12001 (N_12001,N_11532,N_11801);
xnor U12002 (N_12002,N_11995,N_11614);
nand U12003 (N_12003,N_11952,N_11325);
nor U12004 (N_12004,N_10564,N_11146);
and U12005 (N_12005,N_11354,N_11135);
nor U12006 (N_12006,N_11658,N_10523);
nor U12007 (N_12007,N_10711,N_11333);
nor U12008 (N_12008,N_11774,N_11517);
nand U12009 (N_12009,N_11545,N_11964);
or U12010 (N_12010,N_11133,N_10816);
nor U12011 (N_12011,N_11698,N_11652);
and U12012 (N_12012,N_11846,N_11375);
or U12013 (N_12013,N_10797,N_11611);
or U12014 (N_12014,N_10759,N_10725);
xnor U12015 (N_12015,N_10817,N_11295);
and U12016 (N_12016,N_10669,N_11009);
and U12017 (N_12017,N_10729,N_11579);
and U12018 (N_12018,N_11370,N_11398);
nor U12019 (N_12019,N_11866,N_11853);
or U12020 (N_12020,N_11882,N_11881);
nor U12021 (N_12021,N_11759,N_11033);
or U12022 (N_12022,N_11353,N_11606);
nand U12023 (N_12023,N_11576,N_11613);
and U12024 (N_12024,N_11128,N_11645);
or U12025 (N_12025,N_10902,N_11512);
nand U12026 (N_12026,N_11176,N_11998);
and U12027 (N_12027,N_11025,N_10624);
or U12028 (N_12028,N_11102,N_11364);
nor U12029 (N_12029,N_10779,N_11720);
nor U12030 (N_12030,N_10893,N_11931);
or U12031 (N_12031,N_11967,N_11197);
or U12032 (N_12032,N_10806,N_10527);
nand U12033 (N_12033,N_10610,N_10608);
or U12034 (N_12034,N_11923,N_11466);
nor U12035 (N_12035,N_10538,N_11175);
nand U12036 (N_12036,N_10672,N_10855);
nand U12037 (N_12037,N_10613,N_10941);
nor U12038 (N_12038,N_11419,N_11994);
and U12039 (N_12039,N_11660,N_10567);
nor U12040 (N_12040,N_11805,N_11118);
nor U12041 (N_12041,N_11913,N_11654);
nand U12042 (N_12042,N_11607,N_10542);
and U12043 (N_12043,N_11343,N_10598);
and U12044 (N_12044,N_11477,N_11429);
and U12045 (N_12045,N_11799,N_11657);
or U12046 (N_12046,N_11493,N_10753);
nor U12047 (N_12047,N_10928,N_10627);
or U12048 (N_12048,N_10699,N_11121);
or U12049 (N_12049,N_11484,N_11717);
and U12050 (N_12050,N_11089,N_10754);
or U12051 (N_12051,N_10801,N_11473);
xnor U12052 (N_12052,N_11861,N_11815);
and U12053 (N_12053,N_11879,N_11685);
nand U12054 (N_12054,N_11854,N_10728);
or U12055 (N_12055,N_11891,N_11249);
and U12056 (N_12056,N_11075,N_11986);
nand U12057 (N_12057,N_10548,N_11294);
or U12058 (N_12058,N_11303,N_11851);
nor U12059 (N_12059,N_10999,N_11661);
or U12060 (N_12060,N_11961,N_11792);
nor U12061 (N_12061,N_10529,N_11402);
or U12062 (N_12062,N_10926,N_10674);
or U12063 (N_12063,N_10705,N_11305);
nand U12064 (N_12064,N_10968,N_11350);
nand U12065 (N_12065,N_11060,N_11829);
and U12066 (N_12066,N_11908,N_11085);
nor U12067 (N_12067,N_11320,N_10813);
nand U12068 (N_12068,N_10736,N_11349);
and U12069 (N_12069,N_10951,N_11708);
nand U12070 (N_12070,N_10819,N_11744);
nor U12071 (N_12071,N_11684,N_11006);
nand U12072 (N_12072,N_11090,N_11471);
and U12073 (N_12073,N_10706,N_11003);
nand U12074 (N_12074,N_11676,N_11245);
and U12075 (N_12075,N_11702,N_11083);
or U12076 (N_12076,N_11713,N_11005);
nand U12077 (N_12077,N_10774,N_10919);
nand U12078 (N_12078,N_11629,N_10569);
and U12079 (N_12079,N_11459,N_11818);
nor U12080 (N_12080,N_11288,N_11730);
nor U12081 (N_12081,N_10916,N_10515);
and U12082 (N_12082,N_11105,N_10534);
or U12083 (N_12083,N_11926,N_11895);
and U12084 (N_12084,N_11640,N_10782);
and U12085 (N_12085,N_11662,N_10937);
nand U12086 (N_12086,N_11583,N_11737);
nor U12087 (N_12087,N_10865,N_11220);
and U12088 (N_12088,N_11946,N_10825);
nand U12089 (N_12089,N_11235,N_11951);
and U12090 (N_12090,N_10740,N_11763);
or U12091 (N_12091,N_11700,N_11503);
or U12092 (N_12092,N_11059,N_10884);
and U12093 (N_12093,N_11689,N_11502);
nor U12094 (N_12094,N_11174,N_10522);
nand U12095 (N_12095,N_10899,N_11841);
nor U12096 (N_12096,N_11810,N_11740);
and U12097 (N_12097,N_11768,N_11780);
nor U12098 (N_12098,N_11647,N_11515);
nor U12099 (N_12099,N_10526,N_10546);
or U12100 (N_12100,N_10953,N_11575);
nor U12101 (N_12101,N_11947,N_11577);
and U12102 (N_12102,N_10986,N_10554);
and U12103 (N_12103,N_11803,N_11871);
or U12104 (N_12104,N_10805,N_11050);
or U12105 (N_12105,N_11560,N_10908);
and U12106 (N_12106,N_11488,N_10808);
and U12107 (N_12107,N_11725,N_11394);
and U12108 (N_12108,N_11734,N_11157);
nor U12109 (N_12109,N_11439,N_10799);
nand U12110 (N_12110,N_11748,N_11848);
and U12111 (N_12111,N_11336,N_10861);
nand U12112 (N_12112,N_11564,N_10576);
nor U12113 (N_12113,N_11230,N_11642);
nand U12114 (N_12114,N_11639,N_11314);
or U12115 (N_12115,N_11738,N_11587);
or U12116 (N_12116,N_11234,N_10536);
nand U12117 (N_12117,N_11046,N_11599);
or U12118 (N_12118,N_11032,N_10551);
or U12119 (N_12119,N_11806,N_10579);
nand U12120 (N_12120,N_10667,N_11911);
and U12121 (N_12121,N_10880,N_11378);
nand U12122 (N_12122,N_10824,N_11476);
and U12123 (N_12123,N_11001,N_10688);
and U12124 (N_12124,N_10602,N_11754);
nand U12125 (N_12125,N_11022,N_10676);
or U12126 (N_12126,N_10900,N_11411);
nand U12127 (N_12127,N_11044,N_11558);
and U12128 (N_12128,N_10601,N_11572);
nor U12129 (N_12129,N_11980,N_11705);
nand U12130 (N_12130,N_11387,N_10849);
nor U12131 (N_12131,N_10850,N_10914);
nor U12132 (N_12132,N_10639,N_11600);
nor U12133 (N_12133,N_11603,N_11489);
or U12134 (N_12134,N_11819,N_11412);
nand U12135 (N_12135,N_10925,N_11096);
or U12136 (N_12136,N_10609,N_10524);
and U12137 (N_12137,N_10691,N_11139);
or U12138 (N_12138,N_11296,N_11218);
nand U12139 (N_12139,N_10581,N_11581);
nand U12140 (N_12140,N_11427,N_11772);
or U12141 (N_12141,N_10794,N_11876);
nor U12142 (N_12142,N_10943,N_10786);
or U12143 (N_12143,N_11597,N_11322);
or U12144 (N_12144,N_10870,N_10503);
or U12145 (N_12145,N_10989,N_11458);
nand U12146 (N_12146,N_11445,N_10773);
nand U12147 (N_12147,N_11274,N_10731);
and U12148 (N_12148,N_11268,N_11306);
nor U12149 (N_12149,N_10510,N_11329);
and U12150 (N_12150,N_10556,N_11750);
or U12151 (N_12151,N_11399,N_11987);
nand U12152 (N_12152,N_11878,N_11867);
and U12153 (N_12153,N_11531,N_11932);
nand U12154 (N_12154,N_11852,N_11307);
nand U12155 (N_12155,N_11182,N_11401);
nand U12156 (N_12156,N_11634,N_10513);
and U12157 (N_12157,N_11783,N_10678);
or U12158 (N_12158,N_10845,N_10985);
nor U12159 (N_12159,N_10836,N_10839);
and U12160 (N_12160,N_11834,N_10783);
nand U12161 (N_12161,N_11478,N_10878);
nor U12162 (N_12162,N_11368,N_11650);
and U12163 (N_12163,N_11860,N_11051);
nor U12164 (N_12164,N_11021,N_10858);
nand U12165 (N_12165,N_11875,N_10826);
nor U12166 (N_12166,N_10781,N_11984);
or U12167 (N_12167,N_11087,N_11537);
or U12168 (N_12168,N_11345,N_11800);
nor U12169 (N_12169,N_10734,N_10887);
or U12170 (N_12170,N_11462,N_11376);
nand U12171 (N_12171,N_11062,N_11252);
nand U12172 (N_12172,N_11019,N_10501);
nor U12173 (N_12173,N_10988,N_10637);
or U12174 (N_12174,N_11070,N_11226);
or U12175 (N_12175,N_11934,N_11066);
nor U12176 (N_12176,N_11865,N_11390);
or U12177 (N_12177,N_11656,N_11108);
and U12178 (N_12178,N_10516,N_11842);
xnor U12179 (N_12179,N_11273,N_11681);
nor U12180 (N_12180,N_10938,N_10785);
or U12181 (N_12181,N_10612,N_10715);
nand U12182 (N_12182,N_11110,N_11340);
or U12183 (N_12183,N_10507,N_10505);
and U12184 (N_12184,N_10979,N_11648);
or U12185 (N_12185,N_11208,N_11735);
nor U12186 (N_12186,N_11098,N_10620);
and U12187 (N_12187,N_11004,N_11683);
nor U12188 (N_12188,N_10772,N_10795);
nor U12189 (N_12189,N_11200,N_11877);
and U12190 (N_12190,N_11739,N_11279);
or U12191 (N_12191,N_10964,N_10952);
nor U12192 (N_12192,N_10578,N_11454);
or U12193 (N_12193,N_11147,N_11906);
or U12194 (N_12194,N_10570,N_11250);
xnor U12195 (N_12195,N_11836,N_10657);
or U12196 (N_12196,N_11557,N_11358);
nor U12197 (N_12197,N_11468,N_11384);
and U12198 (N_12198,N_11982,N_11610);
nor U12199 (N_12199,N_11627,N_10718);
nor U12200 (N_12200,N_11873,N_11366);
or U12201 (N_12201,N_11337,N_11113);
xnor U12202 (N_12202,N_11541,N_11292);
nor U12203 (N_12203,N_11686,N_11706);
nor U12204 (N_12204,N_11495,N_11511);
nand U12205 (N_12205,N_10838,N_10793);
or U12206 (N_12206,N_11981,N_10622);
xnor U12207 (N_12207,N_11859,N_11828);
nor U12208 (N_12208,N_10588,N_11921);
or U12209 (N_12209,N_10568,N_11518);
nand U12210 (N_12210,N_10934,N_11138);
nor U12211 (N_12211,N_11433,N_11030);
nor U12212 (N_12212,N_11764,N_11898);
and U12213 (N_12213,N_10746,N_11552);
nand U12214 (N_12214,N_10654,N_11100);
or U12215 (N_12215,N_11775,N_11688);
nor U12216 (N_12216,N_11669,N_10972);
or U12217 (N_12217,N_10790,N_10763);
nand U12218 (N_12218,N_11101,N_11410);
and U12219 (N_12219,N_11886,N_11616);
and U12220 (N_12220,N_10573,N_10980);
or U12221 (N_12221,N_11054,N_11598);
nand U12222 (N_12222,N_10502,N_11535);
nand U12223 (N_12223,N_11036,N_10692);
nand U12224 (N_12224,N_11826,N_10896);
or U12225 (N_12225,N_10566,N_11975);
and U12226 (N_12226,N_10589,N_11530);
nor U12227 (N_12227,N_11088,N_11862);
or U12228 (N_12228,N_10702,N_11544);
or U12229 (N_12229,N_10704,N_11240);
nand U12230 (N_12230,N_10686,N_10831);
or U12231 (N_12231,N_10971,N_11726);
and U12232 (N_12232,N_11093,N_11620);
and U12233 (N_12233,N_11324,N_11363);
nor U12234 (N_12234,N_11793,N_11263);
xnor U12235 (N_12235,N_11171,N_11731);
nand U12236 (N_12236,N_10851,N_11017);
nand U12237 (N_12237,N_11525,N_11381);
nor U12238 (N_12238,N_11048,N_11483);
or U12239 (N_12239,N_11203,N_11703);
nand U12240 (N_12240,N_11816,N_10606);
nand U12241 (N_12241,N_11628,N_11413);
nor U12242 (N_12242,N_10636,N_11486);
nand U12243 (N_12243,N_11475,N_11902);
nor U12244 (N_12244,N_11786,N_11892);
and U12245 (N_12245,N_11528,N_11812);
or U12246 (N_12246,N_11672,N_10684);
nand U12247 (N_12247,N_10881,N_10963);
and U12248 (N_12248,N_11126,N_10830);
and U12249 (N_12249,N_10973,N_11061);
or U12250 (N_12250,N_11408,N_10967);
or U12251 (N_12251,N_10827,N_11920);
or U12252 (N_12252,N_11523,N_11519);
nor U12253 (N_12253,N_11903,N_11141);
nand U12254 (N_12254,N_10743,N_11896);
nor U12255 (N_12255,N_10658,N_10644);
and U12256 (N_12256,N_11199,N_10628);
or U12257 (N_12257,N_11238,N_11665);
and U12258 (N_12258,N_11936,N_11561);
or U12259 (N_12259,N_11960,N_11396);
and U12260 (N_12260,N_10592,N_11372);
xnor U12261 (N_12261,N_10742,N_11534);
or U12262 (N_12262,N_11418,N_11996);
or U12263 (N_12263,N_11181,N_11073);
nand U12264 (N_12264,N_10539,N_10804);
nor U12265 (N_12265,N_11715,N_11359);
nand U12266 (N_12266,N_11326,N_10891);
or U12267 (N_12267,N_11290,N_11521);
or U12268 (N_12268,N_10532,N_10769);
and U12269 (N_12269,N_11777,N_10927);
and U12270 (N_12270,N_10681,N_11659);
nor U12271 (N_12271,N_11010,N_10531);
and U12272 (N_12272,N_10732,N_11778);
or U12273 (N_12273,N_10605,N_11928);
nand U12274 (N_12274,N_11441,N_11312);
nand U12275 (N_12275,N_10648,N_11971);
and U12276 (N_12276,N_10521,N_11106);
nor U12277 (N_12277,N_11420,N_11527);
and U12278 (N_12278,N_11666,N_11491);
and U12279 (N_12279,N_11474,N_11404);
or U12280 (N_12280,N_10511,N_11553);
nor U12281 (N_12281,N_11130,N_11506);
or U12282 (N_12282,N_10617,N_10885);
nand U12283 (N_12283,N_11855,N_11280);
or U12284 (N_12284,N_11894,N_11885);
nand U12285 (N_12285,N_10848,N_10557);
nand U12286 (N_12286,N_11131,N_10660);
or U12287 (N_12287,N_10575,N_11955);
and U12288 (N_12288,N_11283,N_11916);
nand U12289 (N_12289,N_11566,N_10915);
nand U12290 (N_12290,N_11546,N_10664);
nand U12291 (N_12291,N_10528,N_11569);
and U12292 (N_12292,N_11028,N_10700);
nor U12293 (N_12293,N_11516,N_10882);
or U12294 (N_12294,N_10898,N_10626);
or U12295 (N_12295,N_11257,N_11596);
or U12296 (N_12296,N_10955,N_11567);
and U12297 (N_12297,N_11189,N_10550);
or U12298 (N_12298,N_10707,N_11136);
or U12299 (N_12299,N_11453,N_11785);
and U12300 (N_12300,N_11940,N_11284);
or U12301 (N_12301,N_10832,N_11173);
or U12302 (N_12302,N_10871,N_11456);
nand U12303 (N_12303,N_11119,N_11554);
nand U12304 (N_12304,N_10944,N_11663);
and U12305 (N_12305,N_11052,N_10597);
or U12306 (N_12306,N_10932,N_11893);
nand U12307 (N_12307,N_11559,N_11346);
and U12308 (N_12308,N_11198,N_11624);
and U12309 (N_12309,N_11985,N_11278);
nand U12310 (N_12310,N_10721,N_11031);
or U12311 (N_12311,N_11332,N_11573);
nand U12312 (N_12312,N_11183,N_11943);
or U12313 (N_12313,N_11887,N_11724);
nor U12314 (N_12314,N_11945,N_11766);
nor U12315 (N_12315,N_11547,N_10812);
nand U12316 (N_12316,N_11978,N_11543);
nand U12317 (N_12317,N_11501,N_11428);
nor U12318 (N_12318,N_11115,N_10975);
nor U12319 (N_12319,N_10543,N_11991);
xnor U12320 (N_12320,N_11677,N_11927);
nand U12321 (N_12321,N_10745,N_11425);
or U12322 (N_12322,N_11190,N_10907);
or U12323 (N_12323,N_11049,N_11762);
nand U12324 (N_12324,N_11297,N_11221);
and U12325 (N_12325,N_11905,N_11505);
nor U12326 (N_12326,N_11837,N_11064);
and U12327 (N_12327,N_10947,N_11237);
or U12328 (N_12328,N_11298,N_11435);
or U12329 (N_12329,N_11563,N_11802);
nand U12330 (N_12330,N_11243,N_11968);
xor U12331 (N_12331,N_11365,N_10533);
or U12332 (N_12332,N_11154,N_11275);
nor U12333 (N_12333,N_11151,N_10994);
nand U12334 (N_12334,N_11712,N_10993);
nand U12335 (N_12335,N_10571,N_11919);
nor U12336 (N_12336,N_10872,N_11356);
nand U12337 (N_12337,N_11219,N_11619);
and U12338 (N_12338,N_10580,N_10894);
nor U12339 (N_12339,N_10561,N_10641);
or U12340 (N_12340,N_10913,N_11371);
and U12341 (N_12341,N_11522,N_11948);
nor U12342 (N_12342,N_11348,N_11770);
nor U12343 (N_12343,N_11057,N_11170);
or U12344 (N_12344,N_11161,N_11788);
or U12345 (N_12345,N_11626,N_10811);
and U12346 (N_12346,N_11016,N_10775);
nand U12347 (N_12347,N_11351,N_10633);
nor U12348 (N_12348,N_11122,N_11310);
or U12349 (N_12349,N_11416,N_10559);
or U12350 (N_12350,N_10879,N_11589);
and U12351 (N_12351,N_10835,N_11701);
or U12352 (N_12352,N_11123,N_10991);
xor U12353 (N_12353,N_11227,N_10623);
or U12354 (N_12354,N_11069,N_10866);
nor U12355 (N_12355,N_10792,N_11782);
nand U12356 (N_12356,N_11962,N_11186);
or U12357 (N_12357,N_10696,N_11668);
or U12358 (N_12358,N_10766,N_10869);
and U12359 (N_12359,N_11153,N_11167);
and U12360 (N_12360,N_11236,N_11117);
nor U12361 (N_12361,N_11432,N_11630);
nand U12362 (N_12362,N_10512,N_11008);
and U12363 (N_12363,N_10594,N_11301);
nand U12364 (N_12364,N_11449,N_11957);
nand U12365 (N_12365,N_11849,N_11617);
or U12366 (N_12366,N_11260,N_11749);
nand U12367 (N_12367,N_11144,N_11431);
nand U12368 (N_12368,N_11205,N_11385);
nor U12369 (N_12369,N_10757,N_10738);
and U12370 (N_12370,N_11727,N_11832);
or U12371 (N_12371,N_10862,N_10917);
nand U12372 (N_12372,N_11922,N_11386);
and U12373 (N_12373,N_11092,N_11584);
or U12374 (N_12374,N_11452,N_10517);
nand U12375 (N_12375,N_10749,N_11958);
or U12376 (N_12376,N_11265,N_11209);
nand U12377 (N_12377,N_11556,N_11675);
nor U12378 (N_12378,N_10614,N_11231);
or U12379 (N_12379,N_11974,N_10504);
nand U12380 (N_12380,N_11592,N_10535);
nand U12381 (N_12381,N_11438,N_11339);
or U12382 (N_12382,N_11213,N_11674);
xor U12383 (N_12383,N_10823,N_10841);
nor U12384 (N_12384,N_11124,N_10655);
xor U12385 (N_12385,N_10921,N_11870);
nor U12386 (N_12386,N_10547,N_11787);
xnor U12387 (N_12387,N_11637,N_11953);
nand U12388 (N_12388,N_11733,N_11211);
and U12389 (N_12389,N_10922,N_10920);
or U12390 (N_12390,N_11910,N_10712);
or U12391 (N_12391,N_10671,N_10990);
nand U12392 (N_12392,N_10936,N_11697);
or U12393 (N_12393,N_11935,N_11142);
and U12394 (N_12394,N_10663,N_11426);
and U12395 (N_12395,N_11999,N_10695);
and U12396 (N_12396,N_10710,N_10611);
and U12397 (N_12397,N_10549,N_10895);
or U12398 (N_12398,N_11448,N_11538);
and U12399 (N_12399,N_11890,N_10800);
nand U12400 (N_12400,N_11670,N_11825);
nand U12401 (N_12401,N_11470,N_10810);
nand U12402 (N_12402,N_10860,N_10905);
or U12403 (N_12403,N_11074,N_11973);
and U12404 (N_12404,N_11415,N_10514);
or U12405 (N_12405,N_10868,N_11682);
nor U12406 (N_12406,N_11299,N_10616);
nor U12407 (N_12407,N_10596,N_10587);
nor U12408 (N_12408,N_11261,N_10815);
nand U12409 (N_12409,N_10603,N_10809);
nand U12410 (N_12410,N_11929,N_11369);
and U12411 (N_12411,N_11664,N_11414);
or U12412 (N_12412,N_11289,N_11382);
nor U12413 (N_12413,N_11103,N_11747);
nor U12414 (N_12414,N_10645,N_11977);
nor U12415 (N_12415,N_11990,N_11490);
and U12416 (N_12416,N_10778,N_11160);
nor U12417 (N_12417,N_10600,N_11077);
or U12418 (N_12418,N_10733,N_10789);
or U12419 (N_12419,N_10708,N_11678);
nand U12420 (N_12420,N_11868,N_10981);
and U12421 (N_12421,N_11736,N_11496);
nor U12422 (N_12422,N_11604,N_10552);
and U12423 (N_12423,N_11026,N_11918);
nand U12424 (N_12424,N_10918,N_11796);
nand U12425 (N_12425,N_11889,N_11817);
or U12426 (N_12426,N_11824,N_10525);
nand U12427 (N_12427,N_10814,N_10650);
or U12428 (N_12428,N_11821,N_11360);
nor U12429 (N_12429,N_10701,N_11018);
or U12430 (N_12430,N_11976,N_10888);
nor U12431 (N_12431,N_11344,N_11091);
nand U12432 (N_12432,N_10520,N_11756);
and U12433 (N_12433,N_10714,N_11149);
nor U12434 (N_12434,N_11309,N_11330);
and U12435 (N_12435,N_10776,N_11482);
and U12436 (N_12436,N_10768,N_11671);
nor U12437 (N_12437,N_10719,N_10730);
nor U12438 (N_12438,N_11814,N_11063);
nor U12439 (N_12439,N_11162,N_11513);
nand U12440 (N_12440,N_10724,N_10662);
and U12441 (N_12441,N_11751,N_10970);
nor U12442 (N_12442,N_11043,N_10807);
nor U12443 (N_12443,N_11168,N_11317);
and U12444 (N_12444,N_10987,N_11965);
nor U12445 (N_12445,N_11056,N_10901);
nand U12446 (N_12446,N_11111,N_10969);
or U12447 (N_12447,N_11443,N_11781);
nor U12448 (N_12448,N_11950,N_11225);
or U12449 (N_12449,N_10682,N_11313);
and U12450 (N_12450,N_10558,N_11758);
nand U12451 (N_12451,N_10574,N_11421);
nand U12452 (N_12452,N_11692,N_10942);
nand U12453 (N_12453,N_11076,N_11323);
nor U12454 (N_12454,N_11695,N_10646);
nand U12455 (N_12455,N_11807,N_10995);
xnor U12456 (N_12456,N_10931,N_10966);
and U12457 (N_12457,N_11362,N_11210);
and U12458 (N_12458,N_11746,N_11196);
nor U12459 (N_12459,N_11972,N_11742);
or U12460 (N_12460,N_10828,N_11334);
and U12461 (N_12461,N_11042,N_11992);
or U12462 (N_12462,N_11704,N_11403);
nor U12463 (N_12463,N_11029,N_11040);
nor U12464 (N_12464,N_10744,N_10717);
nor U12465 (N_12465,N_10630,N_11514);
or U12466 (N_12466,N_11388,N_10634);
nand U12467 (N_12467,N_10974,N_11794);
nand U12468 (N_12468,N_11500,N_10666);
nand U12469 (N_12469,N_11188,N_11784);
nand U12470 (N_12470,N_10933,N_11444);
nor U12471 (N_12471,N_11393,N_11460);
and U12472 (N_12472,N_10840,N_11520);
nor U12473 (N_12473,N_11690,N_10877);
xor U12474 (N_12474,N_11983,N_10764);
nand U12475 (N_12475,N_11694,N_11229);
or U12476 (N_12476,N_11481,N_11869);
and U12477 (N_12477,N_11673,N_10619);
or U12478 (N_12478,N_11389,N_11638);
or U12479 (N_12479,N_10679,N_10685);
and U12480 (N_12480,N_11367,N_10565);
and U12481 (N_12481,N_11395,N_11507);
nand U12482 (N_12482,N_11752,N_11888);
nand U12483 (N_12483,N_11494,N_11707);
and U12484 (N_12484,N_11055,N_11693);
nand U12485 (N_12485,N_11079,N_10929);
or U12486 (N_12486,N_11068,N_11207);
nor U12487 (N_12487,N_11321,N_11741);
and U12488 (N_12488,N_11158,N_10847);
and U12489 (N_12489,N_10962,N_11020);
nor U12490 (N_12490,N_11863,N_11548);
or U12491 (N_12491,N_10788,N_11844);
nor U12492 (N_12492,N_10798,N_11266);
nand U12493 (N_12493,N_11201,N_11461);
xnor U12494 (N_12494,N_11467,N_11156);
nor U12495 (N_12495,N_11422,N_11549);
nor U12496 (N_12496,N_11843,N_11612);
or U12497 (N_12497,N_10852,N_11437);
and U12498 (N_12498,N_11463,N_10912);
and U12499 (N_12499,N_10687,N_10640);
or U12500 (N_12500,N_11191,N_11080);
nand U12501 (N_12501,N_11760,N_11858);
or U12502 (N_12502,N_10583,N_11721);
and U12503 (N_12503,N_11820,N_11850);
and U12504 (N_12504,N_11058,N_10883);
nand U12505 (N_12505,N_11551,N_10903);
nand U12506 (N_12506,N_10954,N_10618);
nor U12507 (N_12507,N_11510,N_10604);
nand U12508 (N_12508,N_11838,N_10846);
nor U12509 (N_12509,N_10818,N_10737);
and U12510 (N_12510,N_11912,N_10750);
and U12511 (N_12511,N_11311,N_11574);
nor U12512 (N_12512,N_11267,N_11722);
or U12513 (N_12513,N_11969,N_11570);
nor U12514 (N_12514,N_11621,N_11811);
xnor U12515 (N_12515,N_10727,N_11251);
nor U12516 (N_12516,N_11595,N_11622);
and U12517 (N_12517,N_10820,N_11907);
or U12518 (N_12518,N_11338,N_10632);
nor U12519 (N_12519,N_10857,N_10940);
nand U12520 (N_12520,N_10585,N_10906);
nand U12521 (N_12521,N_11540,N_11643);
nand U12522 (N_12522,N_11696,N_11272);
or U12523 (N_12523,N_10822,N_10876);
nor U12524 (N_12524,N_11202,N_10791);
nor U12525 (N_12525,N_11152,N_11757);
or U12526 (N_12526,N_11014,N_10690);
or U12527 (N_12527,N_11729,N_11711);
nor U12528 (N_12528,N_11641,N_10544);
nor U12529 (N_12529,N_11644,N_11765);
nand U12530 (N_12530,N_11710,N_10939);
nand U12531 (N_12531,N_10923,N_10500);
nor U12532 (N_12532,N_11623,N_11901);
xnor U12533 (N_12533,N_11880,N_11479);
or U12534 (N_12534,N_11586,N_11216);
nor U12535 (N_12535,N_11352,N_11839);
or U12536 (N_12536,N_11631,N_10765);
and U12537 (N_12537,N_10837,N_11127);
nand U12538 (N_12538,N_11125,N_11094);
nand U12539 (N_12539,N_11791,N_11159);
and U12540 (N_12540,N_11457,N_11104);
nand U12541 (N_12541,N_10961,N_11129);
or U12542 (N_12542,N_10697,N_10977);
nand U12543 (N_12543,N_11716,N_10615);
and U12544 (N_12544,N_11508,N_11608);
and U12545 (N_12545,N_11909,N_10863);
xnor U12546 (N_12546,N_11653,N_11047);
and U12547 (N_12547,N_10665,N_11071);
nand U12548 (N_12548,N_11120,N_10892);
nor U12549 (N_12549,N_11723,N_10625);
nand U12550 (N_12550,N_10873,N_10950);
or U12551 (N_12551,N_11809,N_10586);
or U12552 (N_12552,N_11469,N_11864);
and U12553 (N_12553,N_10960,N_11590);
and U12554 (N_12554,N_11347,N_11937);
nor U12555 (N_12555,N_11165,N_11699);
and U12556 (N_12556,N_10506,N_11446);
nor U12557 (N_12557,N_11178,N_11591);
nor U12558 (N_12558,N_10752,N_10998);
nand U12559 (N_12559,N_10910,N_11959);
and U12560 (N_12560,N_10756,N_10540);
nand U12561 (N_12561,N_10996,N_10693);
or U12562 (N_12562,N_11308,N_11897);
and U12563 (N_12563,N_11097,N_11035);
nand U12564 (N_12564,N_11779,N_11011);
nand U12565 (N_12565,N_11155,N_11112);
nor U12566 (N_12566,N_11039,N_11602);
nor U12567 (N_12567,N_10844,N_11193);
and U12568 (N_12568,N_11542,N_11078);
or U12569 (N_12569,N_10735,N_11023);
or U12570 (N_12570,N_11822,N_11790);
and U12571 (N_12571,N_11072,N_11609);
or U12572 (N_12572,N_10957,N_10959);
and U12573 (N_12573,N_10741,N_11392);
or U12574 (N_12574,N_11813,N_11761);
and U12575 (N_12575,N_11134,N_11732);
nand U12576 (N_12576,N_10935,N_11571);
or U12577 (N_12577,N_11450,N_11374);
nor U12578 (N_12578,N_10948,N_10859);
and U12579 (N_12579,N_11293,N_11857);
or U12580 (N_12580,N_11373,N_11254);
or U12581 (N_12581,N_10760,N_11084);
or U12582 (N_12582,N_11745,N_10949);
nand U12583 (N_12583,N_11938,N_11804);
nor U12584 (N_12584,N_11436,N_10787);
and U12585 (N_12585,N_11169,N_10997);
or U12586 (N_12586,N_10590,N_10629);
nor U12587 (N_12587,N_11434,N_11555);
and U12588 (N_12588,N_10647,N_11835);
and U12589 (N_12589,N_11038,N_11409);
and U12590 (N_12590,N_11899,N_11989);
or U12591 (N_12591,N_11593,N_11979);
nor U12592 (N_12592,N_11424,N_11045);
nand U12593 (N_12593,N_10677,N_11259);
nor U12594 (N_12594,N_10802,N_10751);
and U12595 (N_12595,N_11148,N_11255);
and U12596 (N_12596,N_11588,N_11002);
and U12597 (N_12597,N_11914,N_11529);
nor U12598 (N_12598,N_10541,N_10572);
or U12599 (N_12599,N_11256,N_11081);
and U12600 (N_12600,N_11150,N_11405);
nand U12601 (N_12601,N_11568,N_10621);
or U12602 (N_12602,N_10982,N_11651);
nand U12603 (N_12603,N_10761,N_11132);
or U12604 (N_12604,N_11954,N_11797);
and U12605 (N_12605,N_11380,N_11194);
nor U12606 (N_12606,N_10723,N_11397);
or U12607 (N_12607,N_11550,N_11798);
and U12608 (N_12608,N_11430,N_11248);
or U12609 (N_12609,N_11107,N_10582);
and U12610 (N_12610,N_10518,N_10748);
or U12611 (N_12611,N_10976,N_11172);
and U12612 (N_12612,N_11988,N_11993);
and U12613 (N_12613,N_11872,N_11487);
nor U12614 (N_12614,N_11539,N_10703);
nor U12615 (N_12615,N_11253,N_11884);
and U12616 (N_12616,N_11709,N_11109);
nand U12617 (N_12617,N_11632,N_10689);
or U12618 (N_12618,N_11847,N_10875);
nand U12619 (N_12619,N_11391,N_11166);
nand U12620 (N_12620,N_10758,N_11318);
and U12621 (N_12621,N_10930,N_11246);
nor U12622 (N_12622,N_10545,N_10978);
or U12623 (N_12623,N_11966,N_11217);
nand U12624 (N_12624,N_11264,N_11963);
and U12625 (N_12625,N_11095,N_11625);
nand U12626 (N_12626,N_11179,N_11455);
nor U12627 (N_12627,N_10833,N_10638);
and U12628 (N_12628,N_10595,N_10683);
nand U12629 (N_12629,N_10747,N_11192);
and U12630 (N_12630,N_11222,N_11184);
nand U12631 (N_12631,N_10656,N_11315);
xnor U12632 (N_12632,N_11041,N_10842);
or U12633 (N_12633,N_11615,N_11714);
nand U12634 (N_12634,N_10653,N_10694);
nor U12635 (N_12635,N_11565,N_11180);
or U12636 (N_12636,N_11417,N_10509);
nand U12637 (N_12637,N_10983,N_11485);
nor U12638 (N_12638,N_11185,N_11383);
and U12639 (N_12639,N_11719,N_11291);
nand U12640 (N_12640,N_10853,N_11667);
or U12641 (N_12641,N_11177,N_11140);
and U12642 (N_12642,N_10673,N_11524);
and U12643 (N_12643,N_11239,N_11065);
nand U12644 (N_12644,N_11845,N_10909);
nand U12645 (N_12645,N_11823,N_11451);
nand U12646 (N_12646,N_11440,N_11223);
nand U12647 (N_12647,N_11582,N_10867);
or U12648 (N_12648,N_11000,N_10651);
and U12649 (N_12649,N_11163,N_11406);
and U12650 (N_12650,N_11808,N_11578);
and U12651 (N_12651,N_11942,N_11789);
and U12652 (N_12652,N_11327,N_11944);
xor U12653 (N_12653,N_11776,N_11442);
or U12654 (N_12654,N_11633,N_11526);
nor U12655 (N_12655,N_10767,N_11605);
and U12656 (N_12656,N_11655,N_11755);
nand U12657 (N_12657,N_11465,N_11232);
and U12658 (N_12658,N_11636,N_11504);
nand U12659 (N_12659,N_10796,N_10668);
nor U12660 (N_12660,N_11316,N_11024);
and U12661 (N_12661,N_11361,N_10599);
nor U12662 (N_12662,N_11939,N_10553);
nand U12663 (N_12663,N_11244,N_10675);
nand U12664 (N_12664,N_10631,N_11585);
nor U12665 (N_12665,N_11771,N_11856);
nor U12666 (N_12666,N_10555,N_10886);
nand U12667 (N_12667,N_11013,N_11228);
or U12668 (N_12668,N_10924,N_11498);
and U12669 (N_12669,N_11407,N_11915);
nor U12670 (N_12670,N_11480,N_11562);
and U12671 (N_12671,N_11833,N_11304);
or U12672 (N_12672,N_11241,N_11830);
or U12673 (N_12673,N_10890,N_10856);
nand U12674 (N_12674,N_10635,N_11116);
nand U12675 (N_12675,N_11286,N_10698);
nor U12676 (N_12676,N_11377,N_10593);
nor U12677 (N_12677,N_11447,N_11649);
nor U12678 (N_12678,N_11114,N_11342);
or U12679 (N_12679,N_11580,N_11956);
or U12680 (N_12680,N_10670,N_11718);
nand U12681 (N_12681,N_11287,N_11341);
and U12682 (N_12682,N_11214,N_11464);
nand U12683 (N_12683,N_11357,N_10563);
or U12684 (N_12684,N_11099,N_11933);
nor U12685 (N_12685,N_11282,N_10770);
nand U12686 (N_12686,N_10984,N_11242);
and U12687 (N_12687,N_11067,N_10661);
xnor U12688 (N_12688,N_10722,N_10562);
and U12689 (N_12689,N_10874,N_10843);
and U12690 (N_12690,N_11027,N_11007);
and U12691 (N_12691,N_10508,N_11949);
or U12692 (N_12692,N_10803,N_11400);
and U12693 (N_12693,N_11997,N_11281);
or U12694 (N_12694,N_11379,N_11053);
nand U12695 (N_12695,N_11883,N_11499);
or U12696 (N_12696,N_11195,N_11840);
nand U12697 (N_12697,N_11355,N_11970);
or U12698 (N_12698,N_10643,N_11924);
nor U12699 (N_12699,N_11769,N_11874);
and U12700 (N_12700,N_11533,N_11204);
and U12701 (N_12701,N_11034,N_11917);
or U12702 (N_12702,N_11302,N_11618);
or U12703 (N_12703,N_11497,N_11037);
and U12704 (N_12704,N_11276,N_11328);
or U12705 (N_12705,N_10992,N_10854);
nand U12706 (N_12706,N_11472,N_11687);
nor U12707 (N_12707,N_10537,N_11212);
and U12708 (N_12708,N_11145,N_11164);
and U12709 (N_12709,N_11319,N_10829);
or U12710 (N_12710,N_10945,N_11635);
and U12711 (N_12711,N_11753,N_11187);
nor U12712 (N_12712,N_11137,N_10762);
nand U12713 (N_12713,N_10771,N_11277);
nor U12714 (N_12714,N_10821,N_10864);
nand U12715 (N_12715,N_11900,N_10784);
nor U12716 (N_12716,N_11646,N_11492);
nor U12717 (N_12717,N_11206,N_10720);
nor U12718 (N_12718,N_10649,N_10897);
xnor U12719 (N_12719,N_11335,N_11285);
and U12720 (N_12720,N_10680,N_10642);
nor U12721 (N_12721,N_10591,N_11795);
xnor U12722 (N_12722,N_10904,N_10652);
nor U12723 (N_12723,N_10577,N_10739);
or U12724 (N_12724,N_10607,N_10834);
and U12725 (N_12725,N_11925,N_11215);
and U12726 (N_12726,N_11082,N_10584);
nand U12727 (N_12727,N_10659,N_11300);
nor U12728 (N_12728,N_10530,N_10777);
or U12729 (N_12729,N_10726,N_11269);
or U12730 (N_12730,N_11827,N_11767);
nand U12731 (N_12731,N_11262,N_10911);
nor U12732 (N_12732,N_10780,N_10946);
nand U12733 (N_12733,N_11258,N_11143);
nor U12734 (N_12734,N_10965,N_10560);
nand U12735 (N_12735,N_10956,N_11679);
and U12736 (N_12736,N_11270,N_11247);
or U12737 (N_12737,N_11594,N_10755);
nand U12738 (N_12738,N_11831,N_10713);
nor U12739 (N_12739,N_11012,N_10716);
nor U12740 (N_12740,N_11233,N_11601);
nand U12741 (N_12741,N_11904,N_10709);
nand U12742 (N_12742,N_11773,N_11509);
or U12743 (N_12743,N_11015,N_11536);
nor U12744 (N_12744,N_11680,N_10958);
nand U12745 (N_12745,N_11728,N_11423);
nand U12746 (N_12746,N_11743,N_11930);
nand U12747 (N_12747,N_11691,N_10889);
and U12748 (N_12748,N_11271,N_11941);
nand U12749 (N_12749,N_11331,N_11086);
nor U12750 (N_12750,N_11134,N_11873);
and U12751 (N_12751,N_10785,N_11482);
or U12752 (N_12752,N_11305,N_11472);
nand U12753 (N_12753,N_11064,N_11329);
and U12754 (N_12754,N_10898,N_10642);
nor U12755 (N_12755,N_11272,N_11058);
xnor U12756 (N_12756,N_11234,N_10520);
or U12757 (N_12757,N_10965,N_11896);
nand U12758 (N_12758,N_11136,N_11405);
nand U12759 (N_12759,N_10512,N_11893);
nand U12760 (N_12760,N_11452,N_10685);
or U12761 (N_12761,N_11852,N_11560);
nor U12762 (N_12762,N_11549,N_11673);
nor U12763 (N_12763,N_11864,N_11751);
nor U12764 (N_12764,N_11983,N_11925);
and U12765 (N_12765,N_11302,N_11985);
nor U12766 (N_12766,N_11341,N_10980);
nand U12767 (N_12767,N_11983,N_11954);
or U12768 (N_12768,N_11455,N_10707);
nor U12769 (N_12769,N_11264,N_11322);
nand U12770 (N_12770,N_11981,N_11324);
nor U12771 (N_12771,N_11321,N_11766);
nor U12772 (N_12772,N_11247,N_10633);
and U12773 (N_12773,N_11131,N_11213);
or U12774 (N_12774,N_10629,N_11884);
nand U12775 (N_12775,N_11836,N_11725);
nor U12776 (N_12776,N_11990,N_10715);
nor U12777 (N_12777,N_11899,N_11737);
nor U12778 (N_12778,N_10760,N_11145);
nor U12779 (N_12779,N_11537,N_11074);
or U12780 (N_12780,N_11736,N_10792);
nor U12781 (N_12781,N_10837,N_10713);
nor U12782 (N_12782,N_11832,N_11557);
nand U12783 (N_12783,N_11181,N_11133);
or U12784 (N_12784,N_10507,N_11677);
or U12785 (N_12785,N_11468,N_10601);
and U12786 (N_12786,N_10532,N_10947);
or U12787 (N_12787,N_10790,N_11067);
nand U12788 (N_12788,N_10595,N_10870);
nand U12789 (N_12789,N_10626,N_11097);
or U12790 (N_12790,N_10679,N_11685);
and U12791 (N_12791,N_10621,N_10758);
and U12792 (N_12792,N_11293,N_11533);
and U12793 (N_12793,N_11770,N_11538);
and U12794 (N_12794,N_11184,N_10517);
nand U12795 (N_12795,N_11478,N_10681);
and U12796 (N_12796,N_11696,N_11127);
and U12797 (N_12797,N_10992,N_11445);
and U12798 (N_12798,N_10699,N_11879);
xnor U12799 (N_12799,N_10635,N_11295);
or U12800 (N_12800,N_10774,N_10894);
nand U12801 (N_12801,N_10951,N_10638);
nand U12802 (N_12802,N_10891,N_11068);
or U12803 (N_12803,N_10523,N_11813);
or U12804 (N_12804,N_10655,N_10971);
nand U12805 (N_12805,N_10887,N_11900);
nor U12806 (N_12806,N_10789,N_11046);
or U12807 (N_12807,N_11714,N_11490);
or U12808 (N_12808,N_11999,N_10970);
nand U12809 (N_12809,N_11820,N_11444);
and U12810 (N_12810,N_11194,N_11376);
nand U12811 (N_12811,N_10507,N_11500);
nor U12812 (N_12812,N_10810,N_10619);
or U12813 (N_12813,N_11131,N_10861);
or U12814 (N_12814,N_11906,N_10605);
nand U12815 (N_12815,N_10598,N_11947);
nand U12816 (N_12816,N_10652,N_11507);
nor U12817 (N_12817,N_11942,N_10588);
nor U12818 (N_12818,N_10599,N_10632);
and U12819 (N_12819,N_11528,N_11322);
or U12820 (N_12820,N_11801,N_11920);
and U12821 (N_12821,N_10618,N_11359);
and U12822 (N_12822,N_10963,N_11627);
nand U12823 (N_12823,N_11322,N_10728);
or U12824 (N_12824,N_11031,N_11039);
nand U12825 (N_12825,N_11742,N_10829);
and U12826 (N_12826,N_11149,N_11679);
nor U12827 (N_12827,N_10979,N_11870);
or U12828 (N_12828,N_11366,N_10917);
nand U12829 (N_12829,N_11140,N_11147);
and U12830 (N_12830,N_11920,N_11936);
or U12831 (N_12831,N_11340,N_11999);
and U12832 (N_12832,N_10840,N_10764);
or U12833 (N_12833,N_11209,N_10741);
and U12834 (N_12834,N_11427,N_10982);
nor U12835 (N_12835,N_10905,N_10810);
or U12836 (N_12836,N_11070,N_11158);
nor U12837 (N_12837,N_10665,N_11519);
nand U12838 (N_12838,N_11797,N_11419);
nor U12839 (N_12839,N_11128,N_10531);
or U12840 (N_12840,N_11460,N_11579);
nand U12841 (N_12841,N_10755,N_10655);
nand U12842 (N_12842,N_11589,N_11976);
nor U12843 (N_12843,N_11447,N_11999);
nor U12844 (N_12844,N_11136,N_11904);
nand U12845 (N_12845,N_11091,N_10726);
or U12846 (N_12846,N_10820,N_11404);
nand U12847 (N_12847,N_11117,N_11567);
or U12848 (N_12848,N_11105,N_11856);
and U12849 (N_12849,N_11737,N_11023);
and U12850 (N_12850,N_10769,N_11273);
nor U12851 (N_12851,N_11623,N_11591);
and U12852 (N_12852,N_11190,N_11911);
or U12853 (N_12853,N_10592,N_11311);
nor U12854 (N_12854,N_10683,N_11914);
nor U12855 (N_12855,N_11680,N_11410);
or U12856 (N_12856,N_11357,N_11117);
and U12857 (N_12857,N_11802,N_10578);
and U12858 (N_12858,N_10968,N_11733);
or U12859 (N_12859,N_11348,N_10625);
or U12860 (N_12860,N_11862,N_10924);
nor U12861 (N_12861,N_11613,N_11298);
and U12862 (N_12862,N_11918,N_10816);
and U12863 (N_12863,N_11753,N_11704);
nor U12864 (N_12864,N_11211,N_10751);
or U12865 (N_12865,N_10955,N_11514);
nor U12866 (N_12866,N_11103,N_11177);
and U12867 (N_12867,N_11166,N_11565);
and U12868 (N_12868,N_11135,N_10765);
nand U12869 (N_12869,N_10995,N_11870);
and U12870 (N_12870,N_11273,N_10836);
nand U12871 (N_12871,N_11678,N_11035);
nor U12872 (N_12872,N_11387,N_11028);
and U12873 (N_12873,N_11122,N_11289);
nand U12874 (N_12874,N_11321,N_10804);
nand U12875 (N_12875,N_11096,N_11452);
nor U12876 (N_12876,N_11348,N_10631);
or U12877 (N_12877,N_10815,N_11940);
and U12878 (N_12878,N_11574,N_11161);
and U12879 (N_12879,N_11609,N_10705);
nand U12880 (N_12880,N_11591,N_10906);
nand U12881 (N_12881,N_11564,N_11010);
nor U12882 (N_12882,N_11278,N_11129);
or U12883 (N_12883,N_11102,N_11916);
and U12884 (N_12884,N_11703,N_11442);
and U12885 (N_12885,N_11511,N_10572);
or U12886 (N_12886,N_10975,N_11531);
or U12887 (N_12887,N_11070,N_11270);
or U12888 (N_12888,N_11277,N_11474);
nand U12889 (N_12889,N_11291,N_10983);
nor U12890 (N_12890,N_11038,N_11551);
and U12891 (N_12891,N_11618,N_11290);
xor U12892 (N_12892,N_10728,N_10643);
or U12893 (N_12893,N_10561,N_11669);
or U12894 (N_12894,N_10511,N_11269);
and U12895 (N_12895,N_11588,N_11549);
or U12896 (N_12896,N_11517,N_10717);
nor U12897 (N_12897,N_11572,N_11730);
and U12898 (N_12898,N_11349,N_11655);
nand U12899 (N_12899,N_11989,N_11235);
or U12900 (N_12900,N_10996,N_10753);
nand U12901 (N_12901,N_10603,N_11289);
or U12902 (N_12902,N_11180,N_11641);
nor U12903 (N_12903,N_11566,N_11916);
or U12904 (N_12904,N_10819,N_11972);
nor U12905 (N_12905,N_10699,N_10763);
or U12906 (N_12906,N_11318,N_11861);
nor U12907 (N_12907,N_11670,N_11891);
nor U12908 (N_12908,N_11553,N_11104);
nand U12909 (N_12909,N_11316,N_11374);
or U12910 (N_12910,N_11294,N_11744);
and U12911 (N_12911,N_10986,N_11539);
or U12912 (N_12912,N_10963,N_10741);
nor U12913 (N_12913,N_11387,N_10900);
or U12914 (N_12914,N_10713,N_11770);
xor U12915 (N_12915,N_11077,N_11125);
nand U12916 (N_12916,N_11097,N_11385);
and U12917 (N_12917,N_11194,N_10936);
nor U12918 (N_12918,N_11540,N_11573);
nor U12919 (N_12919,N_10960,N_11874);
or U12920 (N_12920,N_11344,N_10750);
or U12921 (N_12921,N_10806,N_11138);
nand U12922 (N_12922,N_11658,N_11789);
and U12923 (N_12923,N_11942,N_11053);
and U12924 (N_12924,N_11115,N_11574);
and U12925 (N_12925,N_10714,N_11120);
nand U12926 (N_12926,N_11418,N_11935);
or U12927 (N_12927,N_10697,N_10892);
nand U12928 (N_12928,N_11679,N_11123);
or U12929 (N_12929,N_11356,N_11649);
nor U12930 (N_12930,N_11208,N_11163);
or U12931 (N_12931,N_11951,N_11048);
nor U12932 (N_12932,N_11779,N_11565);
nand U12933 (N_12933,N_11827,N_10898);
nand U12934 (N_12934,N_11579,N_11555);
nor U12935 (N_12935,N_11637,N_11809);
or U12936 (N_12936,N_11663,N_10816);
and U12937 (N_12937,N_10674,N_11512);
and U12938 (N_12938,N_10624,N_11853);
and U12939 (N_12939,N_11438,N_10761);
nand U12940 (N_12940,N_10926,N_10960);
xor U12941 (N_12941,N_11262,N_11414);
and U12942 (N_12942,N_11301,N_10802);
nor U12943 (N_12943,N_10786,N_10658);
nor U12944 (N_12944,N_11305,N_11540);
and U12945 (N_12945,N_11314,N_10980);
nand U12946 (N_12946,N_11164,N_11165);
nand U12947 (N_12947,N_10526,N_11921);
nor U12948 (N_12948,N_10849,N_10970);
or U12949 (N_12949,N_11674,N_11777);
xnor U12950 (N_12950,N_10804,N_10897);
nand U12951 (N_12951,N_10808,N_11553);
and U12952 (N_12952,N_11658,N_11624);
or U12953 (N_12953,N_10783,N_10976);
nand U12954 (N_12954,N_11659,N_11813);
and U12955 (N_12955,N_11454,N_11047);
xor U12956 (N_12956,N_11608,N_11281);
and U12957 (N_12957,N_10985,N_10601);
nor U12958 (N_12958,N_10995,N_11349);
and U12959 (N_12959,N_10832,N_11285);
or U12960 (N_12960,N_10754,N_11597);
xnor U12961 (N_12961,N_11433,N_11838);
and U12962 (N_12962,N_10890,N_11301);
nor U12963 (N_12963,N_10936,N_11601);
nand U12964 (N_12964,N_10695,N_11877);
and U12965 (N_12965,N_11850,N_11097);
and U12966 (N_12966,N_10868,N_11069);
or U12967 (N_12967,N_10642,N_11865);
nor U12968 (N_12968,N_11527,N_11223);
and U12969 (N_12969,N_11526,N_11449);
and U12970 (N_12970,N_11943,N_11300);
or U12971 (N_12971,N_11982,N_10666);
and U12972 (N_12972,N_11964,N_10579);
nor U12973 (N_12973,N_11910,N_11659);
and U12974 (N_12974,N_11230,N_11211);
nand U12975 (N_12975,N_11061,N_11106);
or U12976 (N_12976,N_11060,N_11930);
nand U12977 (N_12977,N_10992,N_11407);
nand U12978 (N_12978,N_10756,N_10686);
nand U12979 (N_12979,N_11688,N_11615);
or U12980 (N_12980,N_11797,N_10719);
xor U12981 (N_12981,N_11669,N_11583);
and U12982 (N_12982,N_11473,N_11769);
or U12983 (N_12983,N_10798,N_11481);
nor U12984 (N_12984,N_11543,N_11950);
nor U12985 (N_12985,N_11921,N_11011);
and U12986 (N_12986,N_11305,N_11340);
nor U12987 (N_12987,N_11077,N_10784);
and U12988 (N_12988,N_11969,N_11039);
and U12989 (N_12989,N_11721,N_11966);
nand U12990 (N_12990,N_11921,N_11181);
nor U12991 (N_12991,N_10961,N_11905);
and U12992 (N_12992,N_11368,N_10649);
and U12993 (N_12993,N_11670,N_11316);
nor U12994 (N_12994,N_11575,N_11019);
or U12995 (N_12995,N_11652,N_11618);
and U12996 (N_12996,N_10702,N_10917);
xor U12997 (N_12997,N_11822,N_11978);
nand U12998 (N_12998,N_10787,N_11508);
nand U12999 (N_12999,N_11457,N_10801);
xor U13000 (N_13000,N_10943,N_11853);
and U13001 (N_13001,N_11211,N_10937);
nand U13002 (N_13002,N_11817,N_11720);
or U13003 (N_13003,N_11270,N_10688);
nor U13004 (N_13004,N_10802,N_11873);
and U13005 (N_13005,N_11272,N_11371);
nand U13006 (N_13006,N_10706,N_11911);
or U13007 (N_13007,N_11244,N_11666);
or U13008 (N_13008,N_10980,N_11117);
nand U13009 (N_13009,N_10795,N_11961);
nand U13010 (N_13010,N_11704,N_11404);
or U13011 (N_13011,N_11801,N_11322);
nor U13012 (N_13012,N_11490,N_11428);
or U13013 (N_13013,N_10802,N_11840);
nor U13014 (N_13014,N_10525,N_11879);
nor U13015 (N_13015,N_11551,N_11062);
nand U13016 (N_13016,N_10613,N_11288);
and U13017 (N_13017,N_11209,N_10825);
nand U13018 (N_13018,N_10677,N_10584);
and U13019 (N_13019,N_11863,N_11366);
or U13020 (N_13020,N_11300,N_11620);
nand U13021 (N_13021,N_10823,N_11712);
nand U13022 (N_13022,N_10768,N_10553);
nand U13023 (N_13023,N_10948,N_11512);
or U13024 (N_13024,N_11065,N_10570);
and U13025 (N_13025,N_10614,N_11179);
nor U13026 (N_13026,N_11029,N_11168);
or U13027 (N_13027,N_10854,N_10838);
nor U13028 (N_13028,N_11908,N_11415);
nor U13029 (N_13029,N_10607,N_11441);
or U13030 (N_13030,N_11699,N_10983);
and U13031 (N_13031,N_10662,N_11996);
nand U13032 (N_13032,N_10861,N_11901);
and U13033 (N_13033,N_11264,N_11169);
or U13034 (N_13034,N_10931,N_10589);
and U13035 (N_13035,N_11052,N_11132);
nor U13036 (N_13036,N_11739,N_11161);
and U13037 (N_13037,N_11749,N_11504);
nand U13038 (N_13038,N_11233,N_11340);
nor U13039 (N_13039,N_11247,N_10971);
nor U13040 (N_13040,N_11024,N_11243);
nand U13041 (N_13041,N_11647,N_11347);
and U13042 (N_13042,N_11755,N_11749);
or U13043 (N_13043,N_10758,N_11912);
and U13044 (N_13044,N_11762,N_10546);
nand U13045 (N_13045,N_10523,N_11921);
and U13046 (N_13046,N_11058,N_11742);
nand U13047 (N_13047,N_11903,N_11219);
and U13048 (N_13048,N_11082,N_10572);
nand U13049 (N_13049,N_11174,N_11510);
and U13050 (N_13050,N_10727,N_11319);
nand U13051 (N_13051,N_11267,N_10748);
or U13052 (N_13052,N_11058,N_11990);
nor U13053 (N_13053,N_11710,N_11502);
nand U13054 (N_13054,N_11350,N_10956);
nor U13055 (N_13055,N_11615,N_11285);
nand U13056 (N_13056,N_11610,N_11618);
or U13057 (N_13057,N_10941,N_10698);
and U13058 (N_13058,N_11039,N_11398);
nand U13059 (N_13059,N_11751,N_11863);
or U13060 (N_13060,N_11270,N_10817);
and U13061 (N_13061,N_11732,N_10566);
nor U13062 (N_13062,N_10828,N_10902);
nor U13063 (N_13063,N_10986,N_10968);
and U13064 (N_13064,N_10591,N_11545);
nor U13065 (N_13065,N_11365,N_10749);
nand U13066 (N_13066,N_11421,N_11376);
or U13067 (N_13067,N_11078,N_11930);
nand U13068 (N_13068,N_10967,N_11043);
nor U13069 (N_13069,N_11588,N_11097);
or U13070 (N_13070,N_10771,N_11480);
nand U13071 (N_13071,N_11797,N_10504);
and U13072 (N_13072,N_11704,N_10860);
xnor U13073 (N_13073,N_11710,N_11891);
nor U13074 (N_13074,N_10911,N_10554);
and U13075 (N_13075,N_10561,N_10960);
or U13076 (N_13076,N_10717,N_10792);
and U13077 (N_13077,N_10553,N_11173);
and U13078 (N_13078,N_11115,N_11662);
and U13079 (N_13079,N_10690,N_10550);
nand U13080 (N_13080,N_11502,N_10519);
and U13081 (N_13081,N_11988,N_10623);
xor U13082 (N_13082,N_11943,N_11824);
xnor U13083 (N_13083,N_10614,N_11977);
or U13084 (N_13084,N_11176,N_10727);
nor U13085 (N_13085,N_11754,N_11932);
or U13086 (N_13086,N_11399,N_11196);
nand U13087 (N_13087,N_11708,N_11451);
and U13088 (N_13088,N_10973,N_11870);
or U13089 (N_13089,N_11217,N_11481);
and U13090 (N_13090,N_11778,N_10579);
nor U13091 (N_13091,N_10834,N_11225);
and U13092 (N_13092,N_11367,N_11519);
or U13093 (N_13093,N_10745,N_11102);
and U13094 (N_13094,N_10805,N_11708);
or U13095 (N_13095,N_11329,N_10914);
and U13096 (N_13096,N_11111,N_11974);
and U13097 (N_13097,N_11520,N_10855);
and U13098 (N_13098,N_11499,N_11135);
or U13099 (N_13099,N_11023,N_10861);
nand U13100 (N_13100,N_11437,N_10583);
nand U13101 (N_13101,N_10922,N_10911);
xor U13102 (N_13102,N_10611,N_11710);
and U13103 (N_13103,N_11803,N_11927);
xor U13104 (N_13104,N_11604,N_11447);
nand U13105 (N_13105,N_10772,N_10822);
or U13106 (N_13106,N_10980,N_11151);
and U13107 (N_13107,N_11967,N_11923);
nand U13108 (N_13108,N_11577,N_10719);
nor U13109 (N_13109,N_10916,N_11796);
or U13110 (N_13110,N_11353,N_11684);
or U13111 (N_13111,N_10843,N_10680);
or U13112 (N_13112,N_10856,N_10507);
nand U13113 (N_13113,N_11340,N_11174);
nand U13114 (N_13114,N_11669,N_10799);
nor U13115 (N_13115,N_11443,N_10964);
nor U13116 (N_13116,N_11862,N_10543);
nand U13117 (N_13117,N_10900,N_10874);
and U13118 (N_13118,N_11807,N_11342);
or U13119 (N_13119,N_10930,N_11696);
xor U13120 (N_13120,N_11266,N_11022);
and U13121 (N_13121,N_11042,N_11648);
or U13122 (N_13122,N_11596,N_11744);
or U13123 (N_13123,N_11407,N_11220);
and U13124 (N_13124,N_10773,N_10847);
or U13125 (N_13125,N_10662,N_10832);
nand U13126 (N_13126,N_10954,N_11201);
and U13127 (N_13127,N_10523,N_10819);
nand U13128 (N_13128,N_11330,N_11824);
or U13129 (N_13129,N_10592,N_10910);
or U13130 (N_13130,N_10798,N_11646);
and U13131 (N_13131,N_11063,N_11557);
nand U13132 (N_13132,N_11745,N_10706);
and U13133 (N_13133,N_11830,N_10636);
nor U13134 (N_13134,N_10530,N_10558);
nand U13135 (N_13135,N_10854,N_10656);
nor U13136 (N_13136,N_11020,N_11950);
or U13137 (N_13137,N_11075,N_11330);
nand U13138 (N_13138,N_11456,N_11513);
and U13139 (N_13139,N_11602,N_10591);
or U13140 (N_13140,N_10841,N_11676);
nand U13141 (N_13141,N_10808,N_11964);
and U13142 (N_13142,N_11489,N_11007);
and U13143 (N_13143,N_11153,N_11321);
nand U13144 (N_13144,N_11041,N_10727);
or U13145 (N_13145,N_10690,N_11741);
and U13146 (N_13146,N_11735,N_10517);
or U13147 (N_13147,N_11603,N_10935);
or U13148 (N_13148,N_11711,N_10797);
nand U13149 (N_13149,N_11380,N_11665);
or U13150 (N_13150,N_10914,N_11664);
or U13151 (N_13151,N_10705,N_11308);
and U13152 (N_13152,N_10633,N_11386);
nor U13153 (N_13153,N_11733,N_11920);
and U13154 (N_13154,N_11150,N_11662);
nand U13155 (N_13155,N_10913,N_11180);
nand U13156 (N_13156,N_11550,N_11274);
or U13157 (N_13157,N_11519,N_11804);
nand U13158 (N_13158,N_11214,N_10791);
or U13159 (N_13159,N_10849,N_11819);
or U13160 (N_13160,N_10789,N_11029);
and U13161 (N_13161,N_11885,N_11851);
or U13162 (N_13162,N_11068,N_10726);
and U13163 (N_13163,N_11544,N_10881);
nor U13164 (N_13164,N_11536,N_11615);
nand U13165 (N_13165,N_10559,N_10986);
nor U13166 (N_13166,N_11647,N_11014);
and U13167 (N_13167,N_11401,N_11468);
nand U13168 (N_13168,N_10732,N_10826);
nand U13169 (N_13169,N_11413,N_11726);
and U13170 (N_13170,N_11479,N_11220);
and U13171 (N_13171,N_10590,N_11315);
and U13172 (N_13172,N_11858,N_11027);
nor U13173 (N_13173,N_10992,N_11223);
nor U13174 (N_13174,N_11465,N_11055);
nor U13175 (N_13175,N_10564,N_11446);
xor U13176 (N_13176,N_11154,N_10898);
and U13177 (N_13177,N_11281,N_11158);
or U13178 (N_13178,N_10854,N_10901);
nand U13179 (N_13179,N_11916,N_11096);
nand U13180 (N_13180,N_10768,N_10973);
xnor U13181 (N_13181,N_11940,N_10686);
nor U13182 (N_13182,N_10934,N_11967);
and U13183 (N_13183,N_11451,N_10779);
or U13184 (N_13184,N_11721,N_11712);
xor U13185 (N_13185,N_11848,N_11333);
nand U13186 (N_13186,N_11862,N_11159);
or U13187 (N_13187,N_10983,N_11039);
nor U13188 (N_13188,N_10695,N_10822);
nand U13189 (N_13189,N_11204,N_11714);
nor U13190 (N_13190,N_11813,N_11997);
or U13191 (N_13191,N_10777,N_10599);
nand U13192 (N_13192,N_10718,N_11674);
nor U13193 (N_13193,N_10714,N_11584);
nor U13194 (N_13194,N_11110,N_10971);
nor U13195 (N_13195,N_10505,N_10929);
and U13196 (N_13196,N_10615,N_11820);
and U13197 (N_13197,N_11990,N_11826);
and U13198 (N_13198,N_11957,N_11256);
nor U13199 (N_13199,N_11096,N_10953);
nand U13200 (N_13200,N_10866,N_11807);
or U13201 (N_13201,N_11981,N_11665);
nor U13202 (N_13202,N_11342,N_11920);
nand U13203 (N_13203,N_11719,N_10850);
nor U13204 (N_13204,N_11003,N_11840);
nand U13205 (N_13205,N_11322,N_11518);
or U13206 (N_13206,N_10564,N_11874);
nand U13207 (N_13207,N_11102,N_11988);
and U13208 (N_13208,N_11050,N_11487);
and U13209 (N_13209,N_11867,N_11514);
nor U13210 (N_13210,N_10602,N_11972);
nand U13211 (N_13211,N_11779,N_11312);
and U13212 (N_13212,N_11087,N_11775);
nor U13213 (N_13213,N_11271,N_11924);
or U13214 (N_13214,N_11556,N_11790);
or U13215 (N_13215,N_11609,N_10994);
and U13216 (N_13216,N_11043,N_11467);
nor U13217 (N_13217,N_10855,N_11955);
or U13218 (N_13218,N_11368,N_11280);
nand U13219 (N_13219,N_11377,N_11094);
nor U13220 (N_13220,N_10774,N_11082);
or U13221 (N_13221,N_10562,N_10809);
nor U13222 (N_13222,N_11745,N_11839);
and U13223 (N_13223,N_11399,N_10658);
and U13224 (N_13224,N_11233,N_10541);
nor U13225 (N_13225,N_11158,N_10764);
or U13226 (N_13226,N_11059,N_11452);
and U13227 (N_13227,N_11392,N_10657);
and U13228 (N_13228,N_11667,N_10661);
nor U13229 (N_13229,N_11403,N_11078);
nand U13230 (N_13230,N_11243,N_11727);
nor U13231 (N_13231,N_11457,N_11875);
nor U13232 (N_13232,N_11915,N_10942);
or U13233 (N_13233,N_11285,N_11518);
or U13234 (N_13234,N_11333,N_10546);
nor U13235 (N_13235,N_10943,N_11303);
and U13236 (N_13236,N_11193,N_11236);
nand U13237 (N_13237,N_11973,N_11306);
nand U13238 (N_13238,N_11727,N_11630);
nand U13239 (N_13239,N_11432,N_11880);
or U13240 (N_13240,N_11972,N_11029);
or U13241 (N_13241,N_11221,N_11119);
nor U13242 (N_13242,N_10694,N_10608);
nor U13243 (N_13243,N_10574,N_11474);
or U13244 (N_13244,N_11749,N_11175);
nor U13245 (N_13245,N_11426,N_10626);
nand U13246 (N_13246,N_11246,N_11957);
nand U13247 (N_13247,N_11347,N_10711);
nand U13248 (N_13248,N_11161,N_11051);
and U13249 (N_13249,N_11104,N_10534);
or U13250 (N_13250,N_11871,N_11227);
and U13251 (N_13251,N_11162,N_10520);
and U13252 (N_13252,N_11295,N_11902);
and U13253 (N_13253,N_11642,N_11997);
nor U13254 (N_13254,N_10761,N_10967);
and U13255 (N_13255,N_11798,N_10583);
or U13256 (N_13256,N_11031,N_11991);
and U13257 (N_13257,N_10742,N_11910);
nand U13258 (N_13258,N_10900,N_11042);
nor U13259 (N_13259,N_10552,N_11998);
nand U13260 (N_13260,N_11353,N_11084);
and U13261 (N_13261,N_10548,N_10910);
or U13262 (N_13262,N_11449,N_11285);
and U13263 (N_13263,N_10599,N_10710);
and U13264 (N_13264,N_11780,N_11214);
or U13265 (N_13265,N_10573,N_10882);
or U13266 (N_13266,N_11121,N_11035);
nor U13267 (N_13267,N_10635,N_11774);
nor U13268 (N_13268,N_11973,N_10959);
and U13269 (N_13269,N_11212,N_11386);
nand U13270 (N_13270,N_10825,N_10766);
nand U13271 (N_13271,N_11662,N_11518);
nand U13272 (N_13272,N_10557,N_11097);
and U13273 (N_13273,N_11553,N_10764);
and U13274 (N_13274,N_11254,N_10783);
xor U13275 (N_13275,N_11968,N_10571);
nand U13276 (N_13276,N_11844,N_11493);
nand U13277 (N_13277,N_11518,N_11175);
and U13278 (N_13278,N_10781,N_11933);
nor U13279 (N_13279,N_11981,N_11506);
nand U13280 (N_13280,N_10778,N_11435);
or U13281 (N_13281,N_10618,N_10545);
nand U13282 (N_13282,N_11217,N_11223);
nor U13283 (N_13283,N_11461,N_11172);
and U13284 (N_13284,N_11435,N_11116);
or U13285 (N_13285,N_10697,N_11193);
xor U13286 (N_13286,N_10821,N_11044);
nor U13287 (N_13287,N_11208,N_11874);
or U13288 (N_13288,N_11466,N_11135);
nand U13289 (N_13289,N_11478,N_11017);
or U13290 (N_13290,N_11559,N_11747);
nor U13291 (N_13291,N_11773,N_11273);
nand U13292 (N_13292,N_11915,N_10745);
and U13293 (N_13293,N_11879,N_10587);
nor U13294 (N_13294,N_10639,N_11448);
nor U13295 (N_13295,N_10801,N_11249);
nor U13296 (N_13296,N_11071,N_11542);
and U13297 (N_13297,N_10840,N_11279);
and U13298 (N_13298,N_10740,N_11931);
and U13299 (N_13299,N_11565,N_11559);
or U13300 (N_13300,N_10854,N_11748);
nor U13301 (N_13301,N_11302,N_11367);
nand U13302 (N_13302,N_10860,N_11529);
nor U13303 (N_13303,N_11175,N_11954);
and U13304 (N_13304,N_11558,N_11298);
or U13305 (N_13305,N_11224,N_10756);
or U13306 (N_13306,N_10615,N_11543);
nor U13307 (N_13307,N_11829,N_11414);
or U13308 (N_13308,N_11143,N_11632);
nand U13309 (N_13309,N_10831,N_11182);
nand U13310 (N_13310,N_11013,N_11583);
nor U13311 (N_13311,N_10525,N_11538);
or U13312 (N_13312,N_11320,N_10739);
nor U13313 (N_13313,N_11655,N_11076);
and U13314 (N_13314,N_11394,N_10781);
and U13315 (N_13315,N_10554,N_11269);
nor U13316 (N_13316,N_10935,N_11509);
or U13317 (N_13317,N_10993,N_10845);
nor U13318 (N_13318,N_10887,N_11172);
and U13319 (N_13319,N_11911,N_11015);
and U13320 (N_13320,N_11473,N_11841);
xnor U13321 (N_13321,N_11984,N_11556);
nand U13322 (N_13322,N_10856,N_11443);
nand U13323 (N_13323,N_10620,N_11315);
or U13324 (N_13324,N_11582,N_11937);
and U13325 (N_13325,N_11851,N_11237);
and U13326 (N_13326,N_11872,N_11827);
nand U13327 (N_13327,N_10796,N_11879);
nand U13328 (N_13328,N_11145,N_11167);
or U13329 (N_13329,N_10918,N_11347);
nor U13330 (N_13330,N_11853,N_11322);
nand U13331 (N_13331,N_11391,N_11412);
xnor U13332 (N_13332,N_11951,N_11558);
nor U13333 (N_13333,N_10775,N_11131);
nor U13334 (N_13334,N_11734,N_10757);
nor U13335 (N_13335,N_11814,N_11229);
nor U13336 (N_13336,N_11444,N_11595);
or U13337 (N_13337,N_11304,N_10898);
nand U13338 (N_13338,N_10876,N_10664);
nor U13339 (N_13339,N_11001,N_11226);
or U13340 (N_13340,N_11465,N_10883);
nor U13341 (N_13341,N_11013,N_11387);
nor U13342 (N_13342,N_10662,N_10983);
or U13343 (N_13343,N_11248,N_11189);
nand U13344 (N_13344,N_11933,N_11615);
nor U13345 (N_13345,N_11573,N_11665);
nor U13346 (N_13346,N_11301,N_10881);
nand U13347 (N_13347,N_11586,N_10982);
nand U13348 (N_13348,N_11132,N_11479);
nand U13349 (N_13349,N_11872,N_11813);
nor U13350 (N_13350,N_10501,N_10688);
or U13351 (N_13351,N_11121,N_11957);
or U13352 (N_13352,N_11166,N_11992);
or U13353 (N_13353,N_11569,N_11787);
nor U13354 (N_13354,N_10505,N_10965);
or U13355 (N_13355,N_10583,N_11851);
nand U13356 (N_13356,N_11614,N_11647);
nand U13357 (N_13357,N_10948,N_11161);
nor U13358 (N_13358,N_11499,N_10944);
and U13359 (N_13359,N_11824,N_10649);
and U13360 (N_13360,N_11148,N_11693);
or U13361 (N_13361,N_11013,N_11727);
or U13362 (N_13362,N_11765,N_11278);
nor U13363 (N_13363,N_11878,N_10678);
or U13364 (N_13364,N_11902,N_11769);
nand U13365 (N_13365,N_11098,N_11437);
nor U13366 (N_13366,N_11058,N_11979);
and U13367 (N_13367,N_11878,N_11411);
or U13368 (N_13368,N_11117,N_11409);
nand U13369 (N_13369,N_11522,N_11277);
nor U13370 (N_13370,N_11030,N_10633);
xnor U13371 (N_13371,N_11251,N_11884);
or U13372 (N_13372,N_10594,N_11497);
and U13373 (N_13373,N_11400,N_11500);
or U13374 (N_13374,N_10842,N_11570);
and U13375 (N_13375,N_11019,N_11278);
nor U13376 (N_13376,N_11581,N_10795);
nor U13377 (N_13377,N_11335,N_10757);
or U13378 (N_13378,N_10643,N_11060);
nor U13379 (N_13379,N_10699,N_10839);
nor U13380 (N_13380,N_11499,N_10889);
and U13381 (N_13381,N_11020,N_11031);
nor U13382 (N_13382,N_11570,N_11849);
and U13383 (N_13383,N_11875,N_11470);
and U13384 (N_13384,N_11021,N_11071);
nand U13385 (N_13385,N_11162,N_11777);
nand U13386 (N_13386,N_11415,N_11698);
or U13387 (N_13387,N_11140,N_10977);
or U13388 (N_13388,N_11649,N_11759);
and U13389 (N_13389,N_11146,N_11967);
and U13390 (N_13390,N_11357,N_11413);
nand U13391 (N_13391,N_11598,N_11502);
and U13392 (N_13392,N_11809,N_11778);
nand U13393 (N_13393,N_11503,N_11839);
or U13394 (N_13394,N_11285,N_10576);
and U13395 (N_13395,N_11408,N_11246);
and U13396 (N_13396,N_11650,N_11032);
or U13397 (N_13397,N_11290,N_10953);
or U13398 (N_13398,N_10824,N_11737);
nor U13399 (N_13399,N_11659,N_11068);
or U13400 (N_13400,N_10894,N_11711);
nand U13401 (N_13401,N_10700,N_11973);
and U13402 (N_13402,N_10591,N_10850);
and U13403 (N_13403,N_10923,N_11603);
and U13404 (N_13404,N_11871,N_10905);
nand U13405 (N_13405,N_11417,N_11279);
or U13406 (N_13406,N_10554,N_11828);
and U13407 (N_13407,N_11958,N_11744);
nand U13408 (N_13408,N_10981,N_11602);
or U13409 (N_13409,N_11221,N_11427);
nand U13410 (N_13410,N_11329,N_11730);
and U13411 (N_13411,N_10658,N_11279);
or U13412 (N_13412,N_11693,N_11244);
or U13413 (N_13413,N_11900,N_11102);
and U13414 (N_13414,N_11233,N_10971);
and U13415 (N_13415,N_10866,N_11618);
or U13416 (N_13416,N_10892,N_10562);
nand U13417 (N_13417,N_11169,N_11542);
or U13418 (N_13418,N_11764,N_11327);
and U13419 (N_13419,N_11489,N_10785);
and U13420 (N_13420,N_11904,N_10750);
nor U13421 (N_13421,N_10975,N_11694);
nor U13422 (N_13422,N_11751,N_11853);
nor U13423 (N_13423,N_10688,N_11980);
nand U13424 (N_13424,N_11551,N_10685);
and U13425 (N_13425,N_10668,N_11491);
nor U13426 (N_13426,N_10714,N_11840);
nand U13427 (N_13427,N_10847,N_11773);
and U13428 (N_13428,N_11519,N_11368);
nor U13429 (N_13429,N_11092,N_10692);
nand U13430 (N_13430,N_10652,N_10959);
nor U13431 (N_13431,N_10864,N_10610);
or U13432 (N_13432,N_11096,N_10527);
or U13433 (N_13433,N_10594,N_11906);
or U13434 (N_13434,N_11990,N_11643);
and U13435 (N_13435,N_10807,N_10848);
or U13436 (N_13436,N_11434,N_11345);
or U13437 (N_13437,N_11745,N_11366);
nor U13438 (N_13438,N_10867,N_11687);
nand U13439 (N_13439,N_10711,N_10988);
xor U13440 (N_13440,N_11376,N_10611);
or U13441 (N_13441,N_11809,N_10891);
or U13442 (N_13442,N_11426,N_10644);
nand U13443 (N_13443,N_11217,N_11345);
and U13444 (N_13444,N_10553,N_11017);
and U13445 (N_13445,N_11151,N_10913);
and U13446 (N_13446,N_11897,N_10564);
nand U13447 (N_13447,N_11583,N_11086);
or U13448 (N_13448,N_11926,N_10855);
nor U13449 (N_13449,N_10858,N_10672);
or U13450 (N_13450,N_11748,N_11189);
nor U13451 (N_13451,N_11863,N_11479);
nor U13452 (N_13452,N_11866,N_11936);
or U13453 (N_13453,N_10573,N_11485);
nand U13454 (N_13454,N_11386,N_11688);
nor U13455 (N_13455,N_11661,N_10811);
and U13456 (N_13456,N_11944,N_11693);
and U13457 (N_13457,N_11576,N_11490);
nor U13458 (N_13458,N_11327,N_10827);
or U13459 (N_13459,N_11279,N_10861);
nand U13460 (N_13460,N_10718,N_11904);
and U13461 (N_13461,N_11255,N_11450);
and U13462 (N_13462,N_11366,N_10723);
xor U13463 (N_13463,N_11733,N_11275);
nand U13464 (N_13464,N_10561,N_11008);
and U13465 (N_13465,N_11009,N_11586);
and U13466 (N_13466,N_10712,N_11252);
or U13467 (N_13467,N_11660,N_11972);
nand U13468 (N_13468,N_10533,N_11019);
and U13469 (N_13469,N_11572,N_11289);
and U13470 (N_13470,N_10669,N_10578);
nand U13471 (N_13471,N_11675,N_10533);
nand U13472 (N_13472,N_11128,N_11030);
and U13473 (N_13473,N_11791,N_11360);
or U13474 (N_13474,N_11614,N_11227);
nand U13475 (N_13475,N_10966,N_11540);
or U13476 (N_13476,N_10665,N_11673);
nor U13477 (N_13477,N_11071,N_10817);
nor U13478 (N_13478,N_11080,N_11800);
or U13479 (N_13479,N_11161,N_11177);
nor U13480 (N_13480,N_11317,N_10612);
nor U13481 (N_13481,N_10854,N_11465);
nor U13482 (N_13482,N_11093,N_10869);
or U13483 (N_13483,N_10785,N_11693);
or U13484 (N_13484,N_11038,N_11214);
or U13485 (N_13485,N_11327,N_11414);
nand U13486 (N_13486,N_10883,N_11761);
and U13487 (N_13487,N_10620,N_11312);
nor U13488 (N_13488,N_11475,N_10746);
nor U13489 (N_13489,N_11643,N_11521);
and U13490 (N_13490,N_11330,N_11605);
nor U13491 (N_13491,N_11074,N_10768);
or U13492 (N_13492,N_10683,N_11513);
nand U13493 (N_13493,N_11802,N_10526);
and U13494 (N_13494,N_10649,N_11465);
or U13495 (N_13495,N_11922,N_11236);
nand U13496 (N_13496,N_11634,N_11240);
nor U13497 (N_13497,N_10698,N_11065);
or U13498 (N_13498,N_10997,N_11358);
and U13499 (N_13499,N_10682,N_10956);
xor U13500 (N_13500,N_12370,N_12036);
or U13501 (N_13501,N_12249,N_12324);
nor U13502 (N_13502,N_12379,N_12316);
or U13503 (N_13503,N_12609,N_13099);
and U13504 (N_13504,N_13299,N_12431);
nand U13505 (N_13505,N_12943,N_12646);
or U13506 (N_13506,N_12771,N_13138);
nand U13507 (N_13507,N_12950,N_12886);
or U13508 (N_13508,N_12260,N_12435);
and U13509 (N_13509,N_13376,N_12519);
nand U13510 (N_13510,N_13186,N_12509);
and U13511 (N_13511,N_12375,N_12376);
and U13512 (N_13512,N_12186,N_13198);
nor U13513 (N_13513,N_12098,N_12472);
nor U13514 (N_13514,N_12150,N_12183);
nand U13515 (N_13515,N_13481,N_12693);
or U13516 (N_13516,N_12785,N_12978);
xnor U13517 (N_13517,N_12939,N_12457);
nor U13518 (N_13518,N_12167,N_13109);
or U13519 (N_13519,N_12562,N_12440);
or U13520 (N_13520,N_13359,N_12443);
and U13521 (N_13521,N_13036,N_12746);
nand U13522 (N_13522,N_12603,N_12709);
nor U13523 (N_13523,N_12304,N_12147);
and U13524 (N_13524,N_13314,N_13363);
and U13525 (N_13525,N_13083,N_12121);
and U13526 (N_13526,N_12497,N_13132);
and U13527 (N_13527,N_12954,N_13051);
nor U13528 (N_13528,N_12348,N_13331);
and U13529 (N_13529,N_13303,N_12907);
nor U13530 (N_13530,N_13443,N_13453);
nand U13531 (N_13531,N_12952,N_12703);
or U13532 (N_13532,N_12054,N_12148);
nor U13533 (N_13533,N_12560,N_13330);
xnor U13534 (N_13534,N_12759,N_13284);
or U13535 (N_13535,N_12427,N_12206);
nand U13536 (N_13536,N_12994,N_12701);
or U13537 (N_13537,N_13412,N_12941);
and U13538 (N_13538,N_12488,N_12853);
and U13539 (N_13539,N_13302,N_12223);
nor U13540 (N_13540,N_13072,N_12586);
nand U13541 (N_13541,N_12113,N_12250);
xor U13542 (N_13542,N_13400,N_12708);
nand U13543 (N_13543,N_12066,N_12135);
and U13544 (N_13544,N_13043,N_12384);
or U13545 (N_13545,N_12373,N_12908);
nor U13546 (N_13546,N_12974,N_12474);
nor U13547 (N_13547,N_12489,N_12003);
or U13548 (N_13548,N_12395,N_13269);
nand U13549 (N_13549,N_12969,N_12116);
and U13550 (N_13550,N_13248,N_12213);
nand U13551 (N_13551,N_12485,N_13200);
nor U13552 (N_13552,N_12920,N_12254);
nand U13553 (N_13553,N_12060,N_12571);
nand U13554 (N_13554,N_13029,N_13432);
nor U13555 (N_13555,N_12778,N_13146);
nor U13556 (N_13556,N_13047,N_12508);
nor U13557 (N_13557,N_12847,N_13477);
and U13558 (N_13558,N_12180,N_12381);
or U13559 (N_13559,N_12181,N_12932);
nand U13560 (N_13560,N_13081,N_13354);
nor U13561 (N_13561,N_12720,N_13166);
xnor U13562 (N_13562,N_12937,N_12292);
nand U13563 (N_13563,N_12951,N_12346);
and U13564 (N_13564,N_13246,N_12545);
nand U13565 (N_13565,N_12033,N_12607);
nand U13566 (N_13566,N_12416,N_12735);
or U13567 (N_13567,N_12491,N_12215);
and U13568 (N_13568,N_12936,N_13430);
and U13569 (N_13569,N_12914,N_13387);
or U13570 (N_13570,N_12363,N_12288);
nor U13571 (N_13571,N_12385,N_13046);
and U13572 (N_13572,N_12097,N_12757);
nand U13573 (N_13573,N_13471,N_12927);
nor U13574 (N_13574,N_12817,N_12818);
nor U13575 (N_13575,N_12122,N_13320);
xnor U13576 (N_13576,N_12595,N_12336);
and U13577 (N_13577,N_12469,N_13384);
nand U13578 (N_13578,N_13064,N_12530);
and U13579 (N_13579,N_13071,N_12449);
nor U13580 (N_13580,N_13237,N_13195);
nor U13581 (N_13581,N_12411,N_12698);
nor U13582 (N_13582,N_12640,N_12128);
nand U13583 (N_13583,N_12333,N_12161);
nor U13584 (N_13584,N_12059,N_12547);
or U13585 (N_13585,N_13017,N_12825);
xnor U13586 (N_13586,N_13114,N_12776);
or U13587 (N_13587,N_13256,N_12524);
nor U13588 (N_13588,N_13209,N_13446);
or U13589 (N_13589,N_12794,N_12184);
or U13590 (N_13590,N_12768,N_12513);
nor U13591 (N_13591,N_12037,N_13052);
or U13592 (N_13592,N_13357,N_12362);
or U13593 (N_13593,N_12087,N_13457);
nor U13594 (N_13594,N_12231,N_12169);
and U13595 (N_13595,N_12715,N_12652);
nand U13596 (N_13596,N_12643,N_12834);
and U13597 (N_13597,N_12252,N_12714);
nor U13598 (N_13598,N_12806,N_13317);
or U13599 (N_13599,N_12748,N_13241);
and U13600 (N_13600,N_12117,N_12680);
nand U13601 (N_13601,N_13399,N_12134);
or U13602 (N_13602,N_12366,N_12456);
nor U13603 (N_13603,N_12775,N_12506);
and U13604 (N_13604,N_13203,N_12455);
and U13605 (N_13605,N_12168,N_13104);
nand U13606 (N_13606,N_12897,N_12368);
or U13607 (N_13607,N_13003,N_12217);
nor U13608 (N_13608,N_12599,N_12082);
nor U13609 (N_13609,N_12727,N_12964);
or U13610 (N_13610,N_13000,N_13042);
xnor U13611 (N_13611,N_13202,N_12017);
nor U13612 (N_13612,N_13461,N_12690);
and U13613 (N_13613,N_12833,N_12844);
and U13614 (N_13614,N_12975,N_12542);
and U13615 (N_13615,N_12582,N_13444);
or U13616 (N_13616,N_13434,N_12405);
nor U13617 (N_13617,N_13134,N_12888);
nor U13618 (N_13618,N_12535,N_12419);
nor U13619 (N_13619,N_12662,N_13379);
or U13620 (N_13620,N_13228,N_12481);
xnor U13621 (N_13621,N_12425,N_12073);
or U13622 (N_13622,N_12691,N_13226);
and U13623 (N_13623,N_12325,N_13011);
xnor U13624 (N_13624,N_13490,N_12555);
nor U13625 (N_13625,N_13067,N_13116);
nand U13626 (N_13626,N_12380,N_12983);
or U13627 (N_13627,N_12014,N_12156);
nor U13628 (N_13628,N_12482,N_13101);
and U13629 (N_13629,N_13021,N_13406);
nor U13630 (N_13630,N_13436,N_13037);
nor U13631 (N_13631,N_12523,N_13165);
and U13632 (N_13632,N_13267,N_12922);
nor U13633 (N_13633,N_13086,N_12256);
and U13634 (N_13634,N_12232,N_12928);
or U13635 (N_13635,N_12210,N_12350);
nor U13636 (N_13636,N_12917,N_12123);
and U13637 (N_13637,N_12633,N_12092);
or U13638 (N_13638,N_13061,N_12171);
nor U13639 (N_13639,N_12531,N_13442);
or U13640 (N_13640,N_12044,N_12202);
or U13641 (N_13641,N_12587,N_13440);
nand U13642 (N_13642,N_12575,N_12000);
nor U13643 (N_13643,N_12107,N_12742);
nand U13644 (N_13644,N_13343,N_12711);
nor U13645 (N_13645,N_12904,N_12397);
xnor U13646 (N_13646,N_12620,N_12734);
nor U13647 (N_13647,N_12654,N_12938);
or U13648 (N_13648,N_12876,N_13026);
xor U13649 (N_13649,N_12129,N_12919);
or U13650 (N_13650,N_12358,N_12793);
nor U13651 (N_13651,N_12747,N_12758);
nor U13652 (N_13652,N_12966,N_12548);
nor U13653 (N_13653,N_13445,N_12313);
nor U13654 (N_13654,N_12552,N_12110);
or U13655 (N_13655,N_13173,N_13274);
or U13656 (N_13656,N_12343,N_12371);
xor U13657 (N_13657,N_13245,N_12270);
nor U13658 (N_13658,N_12835,N_13048);
nor U13659 (N_13659,N_12792,N_13148);
nor U13660 (N_13660,N_12301,N_12702);
and U13661 (N_13661,N_13482,N_12877);
and U13662 (N_13662,N_12674,N_12899);
or U13663 (N_13663,N_12052,N_13325);
or U13664 (N_13664,N_12887,N_13233);
and U13665 (N_13665,N_13118,N_13008);
nor U13666 (N_13666,N_13153,N_13057);
and U13667 (N_13667,N_12131,N_12191);
nand U13668 (N_13668,N_13022,N_12067);
nand U13669 (N_13669,N_12903,N_13077);
or U13670 (N_13670,N_12549,N_12063);
nor U13671 (N_13671,N_12255,N_13106);
nor U13672 (N_13672,N_12621,N_12164);
nor U13673 (N_13673,N_12536,N_13313);
and U13674 (N_13674,N_12661,N_13161);
nand U13675 (N_13675,N_13335,N_12868);
or U13676 (N_13676,N_12179,N_12590);
and U13677 (N_13677,N_12880,N_12664);
nor U13678 (N_13678,N_13414,N_13030);
nor U13679 (N_13679,N_12174,N_13425);
or U13680 (N_13680,N_13316,N_12145);
nand U13681 (N_13681,N_13369,N_13049);
nor U13682 (N_13682,N_13403,N_12334);
xor U13683 (N_13683,N_13221,N_13110);
or U13684 (N_13684,N_13038,N_12239);
and U13685 (N_13685,N_12660,N_13291);
and U13686 (N_13686,N_12843,N_12525);
or U13687 (N_13687,N_12364,N_13385);
nor U13688 (N_13688,N_12803,N_13162);
or U13689 (N_13689,N_13091,N_12342);
or U13690 (N_13690,N_13377,N_12881);
nand U13691 (N_13691,N_13348,N_12677);
or U13692 (N_13692,N_13281,N_12671);
or U13693 (N_13693,N_13082,N_13183);
nand U13694 (N_13694,N_12650,N_12041);
nor U13695 (N_13695,N_12789,N_12009);
and U13696 (N_13696,N_12885,N_13147);
nor U13697 (N_13697,N_13454,N_13389);
or U13698 (N_13698,N_12724,N_12527);
nor U13699 (N_13699,N_12540,N_12352);
or U13700 (N_13700,N_13062,N_12185);
nor U13701 (N_13701,N_12743,N_13366);
or U13702 (N_13702,N_12824,N_13009);
or U13703 (N_13703,N_13392,N_12741);
nor U13704 (N_13704,N_12638,N_13260);
and U13705 (N_13705,N_13044,N_12763);
nor U13706 (N_13706,N_12815,N_13273);
nor U13707 (N_13707,N_12257,N_12241);
nor U13708 (N_13708,N_12570,N_12039);
or U13709 (N_13709,N_12011,N_13340);
nand U13710 (N_13710,N_13227,N_13383);
nand U13711 (N_13711,N_13250,N_12221);
and U13712 (N_13712,N_13327,N_13438);
or U13713 (N_13713,N_12996,N_12682);
nor U13714 (N_13714,N_12277,N_12421);
nor U13715 (N_13715,N_12811,N_12644);
and U13716 (N_13716,N_12767,N_12502);
nor U13717 (N_13717,N_12740,N_12068);
nor U13718 (N_13718,N_12813,N_13450);
nand U13719 (N_13719,N_12426,N_13492);
nand U13720 (N_13720,N_12420,N_12208);
or U13721 (N_13721,N_12948,N_12865);
and U13722 (N_13722,N_12476,N_13181);
or U13723 (N_13723,N_13361,N_12062);
or U13724 (N_13724,N_12049,N_13184);
xnor U13725 (N_13725,N_12389,N_13424);
nand U13726 (N_13726,N_13353,N_12687);
nor U13727 (N_13727,N_12152,N_12728);
or U13728 (N_13728,N_12988,N_13164);
nor U13729 (N_13729,N_13133,N_13012);
nand U13730 (N_13730,N_12490,N_13097);
nand U13731 (N_13731,N_12719,N_13229);
nand U13732 (N_13732,N_12556,N_13103);
nand U13733 (N_13733,N_12867,N_13130);
nand U13734 (N_13734,N_12308,N_12520);
and U13735 (N_13735,N_13411,N_12772);
or U13736 (N_13736,N_12568,N_12980);
nor U13737 (N_13737,N_13449,N_12335);
nor U13738 (N_13738,N_12807,N_12189);
and U13739 (N_13739,N_12705,N_13422);
or U13740 (N_13740,N_12819,N_13407);
nand U13741 (N_13741,N_12263,N_12925);
or U13742 (N_13742,N_12264,N_12534);
nor U13743 (N_13743,N_12851,N_12546);
or U13744 (N_13744,N_12790,N_12639);
xnor U13745 (N_13745,N_12329,N_12856);
or U13746 (N_13746,N_13096,N_12672);
or U13747 (N_13747,N_12697,N_13433);
and U13748 (N_13748,N_12158,N_13336);
nor U13749 (N_13749,N_13395,N_12173);
and U13750 (N_13750,N_12057,N_13123);
xnor U13751 (N_13751,N_12015,N_12132);
or U13752 (N_13752,N_13063,N_12207);
nand U13753 (N_13753,N_12801,N_13386);
or U13754 (N_13754,N_12648,N_12989);
nand U13755 (N_13755,N_12515,N_13367);
nor U13756 (N_13756,N_12561,N_12267);
nor U13757 (N_13757,N_13373,N_12203);
nand U13758 (N_13758,N_12753,N_12750);
and U13759 (N_13759,N_12918,N_13027);
or U13760 (N_13760,N_12657,N_12396);
and U13761 (N_13761,N_12955,N_12944);
or U13762 (N_13762,N_12172,N_13150);
or U13763 (N_13763,N_12940,N_13337);
and U13764 (N_13764,N_12528,N_12829);
or U13765 (N_13765,N_12372,N_12784);
and U13766 (N_13766,N_12023,N_12499);
nor U13767 (N_13767,N_12689,N_12896);
or U13768 (N_13768,N_13350,N_12088);
or U13769 (N_13769,N_12665,N_13290);
or U13770 (N_13770,N_12608,N_12659);
nand U13771 (N_13771,N_13194,N_12175);
nand U13772 (N_13772,N_13427,N_13002);
or U13773 (N_13773,N_12898,N_12971);
nor U13774 (N_13774,N_13120,N_13159);
or U13775 (N_13775,N_12494,N_12780);
nor U13776 (N_13776,N_13177,N_12788);
or U13777 (N_13777,N_12684,N_13447);
nand U13778 (N_13778,N_13388,N_12669);
nand U13779 (N_13779,N_13362,N_12018);
nand U13780 (N_13780,N_12816,N_12559);
nor U13781 (N_13781,N_13401,N_13416);
xor U13782 (N_13782,N_12606,N_13033);
and U13783 (N_13783,N_13470,N_12629);
nor U13784 (N_13784,N_12878,N_12394);
nor U13785 (N_13785,N_12448,N_12602);
and U13786 (N_13786,N_12500,N_12874);
nor U13787 (N_13787,N_13280,N_13451);
nand U13788 (N_13788,N_12997,N_12533);
and U13789 (N_13789,N_13121,N_12585);
or U13790 (N_13790,N_12762,N_12605);
and U13791 (N_13791,N_12451,N_12286);
nand U13792 (N_13792,N_12745,N_12473);
nor U13793 (N_13793,N_13251,N_13041);
or U13794 (N_13794,N_12276,N_12354);
and U13795 (N_13795,N_12809,N_13370);
nand U13796 (N_13796,N_12287,N_13201);
or U13797 (N_13797,N_13467,N_12635);
or U13798 (N_13798,N_12906,N_12096);
and U13799 (N_13799,N_12297,N_12246);
nor U13800 (N_13800,N_12934,N_12091);
or U13801 (N_13801,N_12826,N_12837);
and U13802 (N_13802,N_13190,N_12114);
nand U13803 (N_13803,N_12912,N_13418);
nand U13804 (N_13804,N_13468,N_12323);
nor U13805 (N_13805,N_13075,N_13485);
or U13806 (N_13806,N_12137,N_12351);
nand U13807 (N_13807,N_12730,N_12081);
and U13808 (N_13808,N_12507,N_12024);
or U13809 (N_13809,N_12306,N_13179);
or U13810 (N_13810,N_12594,N_13309);
nor U13811 (N_13811,N_13435,N_12356);
or U13812 (N_13812,N_12756,N_13452);
nand U13813 (N_13813,N_12170,N_12773);
or U13814 (N_13814,N_13344,N_12109);
nand U13815 (N_13815,N_13206,N_13489);
nand U13816 (N_13816,N_13020,N_12083);
nand U13817 (N_13817,N_12227,N_12331);
and U13818 (N_13818,N_12086,N_12320);
nand U13819 (N_13819,N_12958,N_13157);
nand U13820 (N_13820,N_13423,N_12557);
nand U13821 (N_13821,N_12162,N_12900);
or U13822 (N_13822,N_13483,N_12589);
nor U13823 (N_13823,N_12831,N_13259);
or U13824 (N_13824,N_12760,N_12864);
nor U13825 (N_13825,N_13170,N_12013);
nand U13826 (N_13826,N_13115,N_13225);
nor U13827 (N_13827,N_12694,N_13001);
or U13828 (N_13828,N_12972,N_13469);
nand U13829 (N_13829,N_12840,N_12273);
nor U13830 (N_13830,N_12349,N_12025);
nor U13831 (N_13831,N_12236,N_13408);
or U13832 (N_13832,N_12611,N_13019);
or U13833 (N_13833,N_13122,N_13287);
nand U13834 (N_13834,N_12862,N_12322);
nand U13835 (N_13835,N_12187,N_12787);
nand U13836 (N_13836,N_12295,N_13487);
nand U13837 (N_13837,N_13479,N_12251);
or U13838 (N_13838,N_12610,N_12402);
and U13839 (N_13839,N_13093,N_12987);
or U13840 (N_13840,N_12111,N_12892);
nor U13841 (N_13841,N_12642,N_13187);
or U13842 (N_13842,N_13092,N_13242);
nor U13843 (N_13843,N_12667,N_12721);
nand U13844 (N_13844,N_13142,N_12647);
nand U13845 (N_13845,N_12298,N_12883);
nor U13846 (N_13846,N_12468,N_12676);
and U13847 (N_13847,N_12075,N_13169);
nand U13848 (N_13848,N_12655,N_12957);
and U13849 (N_13849,N_13193,N_13235);
and U13850 (N_13850,N_13004,N_12563);
or U13851 (N_13851,N_12076,N_12022);
nor U13852 (N_13852,N_13239,N_12592);
and U13853 (N_13853,N_13283,N_13311);
nand U13854 (N_13854,N_13264,N_13334);
nor U13855 (N_13855,N_12583,N_12108);
nand U13856 (N_13856,N_13391,N_12890);
and U13857 (N_13857,N_12779,N_12504);
nor U13858 (N_13858,N_12299,N_12795);
nand U13859 (N_13859,N_12212,N_13419);
nand U13860 (N_13860,N_13382,N_12514);
nand U13861 (N_13861,N_13488,N_12543);
or U13862 (N_13862,N_12544,N_12942);
nand U13863 (N_13863,N_12205,N_13428);
and U13864 (N_13864,N_12751,N_12965);
xor U13865 (N_13865,N_12230,N_12112);
or U13866 (N_13866,N_13060,N_13378);
nand U13867 (N_13867,N_12099,N_13231);
or U13868 (N_13868,N_12237,N_12459);
and U13869 (N_13869,N_12142,N_12923);
nor U13870 (N_13870,N_12200,N_13217);
nor U13871 (N_13871,N_12700,N_12139);
nand U13872 (N_13872,N_13297,N_12492);
and U13873 (N_13873,N_12275,N_13272);
nor U13874 (N_13874,N_12242,N_12439);
nand U13875 (N_13875,N_12125,N_13080);
nor U13876 (N_13876,N_12028,N_12712);
nor U13877 (N_13877,N_12317,N_12050);
and U13878 (N_13878,N_12666,N_12077);
nor U13879 (N_13879,N_12812,N_12045);
or U13880 (N_13880,N_12115,N_13288);
nand U13881 (N_13881,N_12340,N_12319);
nand U13882 (N_13882,N_12302,N_12658);
and U13883 (N_13883,N_13265,N_13394);
and U13884 (N_13884,N_12103,N_12581);
and U13885 (N_13885,N_12962,N_12401);
xnor U13886 (N_13886,N_12947,N_13277);
nand U13887 (N_13887,N_12852,N_12194);
and U13888 (N_13888,N_12986,N_12861);
nor U13889 (N_13889,N_12085,N_13448);
and U13890 (N_13890,N_12102,N_12369);
xnor U13891 (N_13891,N_12569,N_13404);
and U13892 (N_13892,N_12631,N_12414);
and U13893 (N_13893,N_12328,N_12460);
nand U13894 (N_13894,N_12827,N_13455);
and U13895 (N_13895,N_12685,N_13050);
nand U13896 (N_13896,N_12889,N_13380);
nor U13897 (N_13897,N_12554,N_12977);
nand U13898 (N_13898,N_12056,N_13126);
xnor U13899 (N_13899,N_12193,N_12188);
and U13900 (N_13900,N_13405,N_13494);
or U13901 (N_13901,N_13255,N_12870);
nor U13902 (N_13902,N_12423,N_13285);
and U13903 (N_13903,N_12915,N_12461);
and U13904 (N_13904,N_12360,N_13480);
or U13905 (N_13905,N_12138,N_12437);
nand U13906 (N_13906,N_13293,N_13484);
and U13907 (N_13907,N_13295,N_12090);
nor U13908 (N_13908,N_12248,N_13028);
nand U13909 (N_13909,N_12995,N_12921);
or U13910 (N_13910,N_12752,N_12956);
nor U13911 (N_13911,N_12584,N_13497);
nand U13912 (N_13912,N_13420,N_13315);
and U13913 (N_13913,N_12529,N_12289);
or U13914 (N_13914,N_12632,N_13143);
nor U13915 (N_13915,N_12344,N_13466);
nand U13916 (N_13916,N_13107,N_12493);
and U13917 (N_13917,N_12550,N_13111);
and U13918 (N_13918,N_13182,N_12961);
nand U13919 (N_13919,N_12828,N_12444);
or U13920 (N_13920,N_12143,N_12731);
nor U13921 (N_13921,N_12296,N_12177);
and U13922 (N_13922,N_12151,N_12235);
or U13923 (N_13923,N_13349,N_12019);
and U13924 (N_13924,N_13084,N_12154);
or U13925 (N_13925,N_12769,N_13240);
nor U13926 (N_13926,N_12211,N_12126);
nand U13927 (N_13927,N_12749,N_13282);
nand U13928 (N_13928,N_13261,N_12696);
nor U13929 (N_13929,N_12484,N_12305);
nor U13930 (N_13930,N_13180,N_13223);
nor U13931 (N_13931,N_12532,N_12332);
nand U13932 (N_13932,N_12967,N_12007);
xnor U13933 (N_13933,N_13216,N_12120);
nor U13934 (N_13934,N_13465,N_13257);
nor U13935 (N_13935,N_12617,N_12035);
nor U13936 (N_13936,N_13141,N_12220);
and U13937 (N_13937,N_12798,N_12253);
nand U13938 (N_13938,N_12551,N_12681);
or U13939 (N_13939,N_13095,N_13006);
and U13940 (N_13940,N_12244,N_12797);
nand U13941 (N_13941,N_12409,N_12580);
or U13942 (N_13942,N_12093,N_12383);
and U13943 (N_13943,N_12510,N_12430);
nor U13944 (N_13944,N_12616,N_12872);
nor U13945 (N_13945,N_12879,N_13196);
and U13946 (N_13946,N_12136,N_12699);
nand U13947 (N_13947,N_13185,N_12641);
nand U13948 (N_13948,N_12567,N_13338);
nor U13949 (N_13949,N_12293,N_12467);
and U13950 (N_13950,N_13300,N_12192);
or U13951 (N_13951,N_13139,N_12623);
xor U13952 (N_13952,N_12258,N_12234);
and U13953 (N_13953,N_12214,N_13381);
and U13954 (N_13954,N_12020,N_13347);
and U13955 (N_13955,N_12001,N_13421);
and U13956 (N_13956,N_12404,N_12058);
nor U13957 (N_13957,N_12300,N_13458);
nor U13958 (N_13958,N_13332,N_13174);
nor U13959 (N_13959,N_13472,N_12432);
or U13960 (N_13960,N_12838,N_13224);
or U13961 (N_13961,N_12436,N_13253);
nand U13962 (N_13962,N_13154,N_12141);
nand U13963 (N_13963,N_12280,N_12931);
and U13964 (N_13964,N_13219,N_12021);
nor U13965 (N_13965,N_12291,N_12651);
nand U13966 (N_13966,N_12539,N_12338);
and U13967 (N_13967,N_13234,N_12558);
or U13968 (N_13968,N_12327,N_12008);
nand U13969 (N_13969,N_12290,N_12579);
or U13970 (N_13970,N_12754,N_12839);
and U13971 (N_13971,N_13499,N_12992);
and U13972 (N_13972,N_12814,N_12871);
and U13973 (N_13973,N_13131,N_12155);
or U13974 (N_13974,N_12245,N_12913);
nand U13975 (N_13975,N_13199,N_12630);
or U13976 (N_13976,N_13137,N_13270);
and U13977 (N_13977,N_12478,N_13306);
nor U13978 (N_13978,N_12854,N_13304);
or U13979 (N_13979,N_13136,N_12882);
nand U13980 (N_13980,N_12311,N_13476);
xor U13981 (N_13981,N_13417,N_13189);
and U13982 (N_13982,N_12269,N_12591);
or U13983 (N_13983,N_12279,N_12675);
and U13984 (N_13984,N_13214,N_12566);
nand U13985 (N_13985,N_13441,N_12774);
or U13986 (N_13986,N_13073,N_12688);
nor U13987 (N_13987,N_12284,N_12704);
nand U13988 (N_13988,N_12968,N_12808);
and U13989 (N_13989,N_12916,N_12588);
and U13990 (N_13990,N_12106,N_12417);
nand U13991 (N_13991,N_12755,N_12863);
nor U13992 (N_13992,N_13149,N_12737);
or U13993 (N_13993,N_12668,N_13212);
nor U13994 (N_13994,N_12518,N_13208);
or U13995 (N_13995,N_13346,N_12670);
or U13996 (N_13996,N_13085,N_13056);
nor U13997 (N_13997,N_12653,N_13220);
nor U13998 (N_13998,N_12893,N_12261);
or U13999 (N_13999,N_12166,N_12683);
nor U14000 (N_14000,N_12199,N_13125);
or U14001 (N_14001,N_13374,N_13058);
nor U14002 (N_14002,N_12692,N_12470);
or U14003 (N_14003,N_13390,N_13351);
nand U14004 (N_14004,N_13113,N_12447);
nand U14005 (N_14005,N_12307,N_12901);
nor U14006 (N_14006,N_12196,N_13054);
nor U14007 (N_14007,N_12910,N_12367);
and U14008 (N_14008,N_12377,N_13397);
and U14009 (N_14009,N_12209,N_12361);
and U14010 (N_14010,N_12832,N_12442);
nand U14011 (N_14011,N_12040,N_13218);
nand U14012 (N_14012,N_12226,N_13191);
or U14013 (N_14013,N_13031,N_12403);
and U14014 (N_14014,N_12802,N_13355);
nand U14015 (N_14015,N_12935,N_13319);
and U14016 (N_14016,N_12782,N_12454);
and U14017 (N_14017,N_13360,N_12118);
or U14018 (N_14018,N_13230,N_12875);
or U14019 (N_14019,N_12722,N_12615);
and U14020 (N_14020,N_12744,N_12198);
or U14021 (N_14021,N_12723,N_12391);
nor U14022 (N_14022,N_12218,N_12479);
and U14023 (N_14023,N_12718,N_12326);
nand U14024 (N_14024,N_13493,N_12153);
or U14025 (N_14025,N_12619,N_12963);
nand U14026 (N_14026,N_12949,N_13409);
and U14027 (N_14027,N_12222,N_12374);
nand U14028 (N_14028,N_13252,N_12716);
or U14029 (N_14029,N_13108,N_13135);
nand U14030 (N_14030,N_12388,N_12991);
or U14031 (N_14031,N_12842,N_12216);
nor U14032 (N_14032,N_12130,N_12841);
nand U14033 (N_14033,N_13339,N_13478);
nand U14034 (N_14034,N_12149,N_12030);
or U14035 (N_14035,N_12970,N_13496);
and U14036 (N_14036,N_12070,N_12031);
or U14037 (N_14037,N_12400,N_12578);
and U14038 (N_14038,N_13358,N_12710);
and U14039 (N_14039,N_12766,N_13068);
and U14040 (N_14040,N_12783,N_13247);
and U14041 (N_14041,N_12786,N_13464);
and U14042 (N_14042,N_12764,N_13266);
nand U14043 (N_14043,N_13323,N_13215);
and U14044 (N_14044,N_12176,N_12471);
or U14045 (N_14045,N_13079,N_12624);
and U14046 (N_14046,N_13329,N_12310);
nand U14047 (N_14047,N_13254,N_12341);
and U14048 (N_14048,N_12501,N_12100);
nand U14049 (N_14049,N_13151,N_13402);
or U14050 (N_14050,N_12503,N_12738);
nand U14051 (N_14051,N_13024,N_13356);
nand U14052 (N_14052,N_12359,N_12124);
and U14053 (N_14053,N_12998,N_12160);
xor U14054 (N_14054,N_13460,N_13167);
nand U14055 (N_14055,N_12016,N_12224);
nor U14056 (N_14056,N_12424,N_13474);
and U14057 (N_14057,N_13128,N_12593);
or U14058 (N_14058,N_12905,N_12706);
nand U14059 (N_14059,N_12281,N_12564);
nor U14060 (N_14060,N_12378,N_12604);
nor U14061 (N_14061,N_12574,N_13262);
nand U14062 (N_14062,N_12278,N_12739);
and U14063 (N_14063,N_13105,N_13426);
or U14064 (N_14064,N_12663,N_13495);
nor U14065 (N_14065,N_12673,N_12268);
nand U14066 (N_14066,N_12355,N_13053);
nand U14067 (N_14067,N_12428,N_12999);
nor U14068 (N_14068,N_13462,N_12190);
nand U14069 (N_14069,N_12055,N_12860);
nand U14070 (N_14070,N_12240,N_12197);
nor U14071 (N_14071,N_12993,N_12821);
and U14072 (N_14072,N_12144,N_13018);
nand U14073 (N_14073,N_13144,N_13439);
nor U14074 (N_14074,N_12713,N_12733);
xor U14075 (N_14075,N_12781,N_13168);
nand U14076 (N_14076,N_12976,N_12929);
nand U14077 (N_14077,N_12010,N_13039);
and U14078 (N_14078,N_12601,N_12765);
and U14079 (N_14079,N_12565,N_12483);
nor U14080 (N_14080,N_12101,N_13486);
or U14081 (N_14081,N_12365,N_12064);
or U14082 (N_14082,N_12095,N_13119);
nand U14083 (N_14083,N_13055,N_13013);
and U14084 (N_14084,N_12433,N_12429);
nand U14085 (N_14085,N_12283,N_12981);
or U14086 (N_14086,N_13310,N_12848);
nor U14087 (N_14087,N_13078,N_13396);
or U14088 (N_14088,N_12415,N_13301);
or U14089 (N_14089,N_12462,N_12229);
nand U14090 (N_14090,N_12859,N_13140);
nand U14091 (N_14091,N_12262,N_12475);
nand U14092 (N_14092,N_13232,N_12822);
or U14093 (N_14093,N_13238,N_12649);
and U14094 (N_14094,N_12163,N_12736);
nand U14095 (N_14095,N_12080,N_13365);
nor U14096 (N_14096,N_13088,N_12353);
and U14097 (N_14097,N_12127,N_13207);
nor U14098 (N_14098,N_12071,N_12791);
nand U14099 (N_14099,N_12512,N_12182);
and U14100 (N_14100,N_13278,N_13005);
nor U14101 (N_14101,N_12902,N_13307);
and U14102 (N_14102,N_12266,N_12707);
and U14103 (N_14103,N_12466,N_12272);
or U14104 (N_14104,N_12805,N_12732);
or U14105 (N_14105,N_12225,N_13098);
nor U14106 (N_14106,N_12480,N_13244);
nor U14107 (N_14107,N_12386,N_12393);
nand U14108 (N_14108,N_13393,N_12464);
nand U14109 (N_14109,N_13074,N_12634);
nand U14110 (N_14110,N_13090,N_13045);
nor U14111 (N_14111,N_12157,N_12104);
or U14112 (N_14112,N_13371,N_13263);
nor U14113 (N_14113,N_13286,N_12032);
nand U14114 (N_14114,N_12845,N_12004);
nand U14115 (N_14115,N_12855,N_12498);
and U14116 (N_14116,N_12576,N_13155);
nor U14117 (N_14117,N_13197,N_12625);
and U14118 (N_14118,N_12796,N_13279);
nand U14119 (N_14119,N_12398,N_13066);
nand U14120 (N_14120,N_12945,N_12487);
nand U14121 (N_14121,N_12382,N_12729);
nor U14122 (N_14122,N_12496,N_12303);
or U14123 (N_14123,N_13210,N_12990);
or U14124 (N_14124,N_12984,N_12979);
nor U14125 (N_14125,N_12146,N_12820);
or U14126 (N_14126,N_12959,N_13014);
or U14127 (N_14127,N_12985,N_13222);
or U14128 (N_14128,N_12982,N_12285);
or U14129 (N_14129,N_13459,N_12463);
and U14130 (N_14130,N_12051,N_13321);
nor U14131 (N_14131,N_12165,N_12521);
nand U14132 (N_14132,N_12895,N_13318);
and U14133 (N_14133,N_12598,N_13275);
nor U14134 (N_14134,N_12960,N_13035);
xnor U14135 (N_14135,N_12046,N_12777);
nor U14136 (N_14136,N_12247,N_12572);
or U14137 (N_14137,N_12836,N_13413);
nor U14138 (N_14138,N_13236,N_13429);
or U14139 (N_14139,N_12446,N_13178);
and U14140 (N_14140,N_13271,N_12330);
nand U14141 (N_14141,N_12597,N_13276);
nor U14142 (N_14142,N_12458,N_12034);
and U14143 (N_14143,N_12538,N_12347);
nand U14144 (N_14144,N_13160,N_13023);
or U14145 (N_14145,N_12627,N_12933);
nand U14146 (N_14146,N_12259,N_12517);
or U14147 (N_14147,N_13475,N_12695);
or U14148 (N_14148,N_12228,N_12407);
xnor U14149 (N_14149,N_12622,N_12069);
xnor U14150 (N_14150,N_13089,N_12159);
and U14151 (N_14151,N_12048,N_12679);
nor U14152 (N_14152,N_13156,N_13076);
or U14153 (N_14153,N_12511,N_13129);
nand U14154 (N_14154,N_12452,N_12686);
nor U14155 (N_14155,N_12445,N_12973);
and U14156 (N_14156,N_13268,N_12846);
or U14157 (N_14157,N_13213,N_12516);
and U14158 (N_14158,N_12884,N_13352);
nand U14159 (N_14159,N_13117,N_12315);
nor U14160 (N_14160,N_12412,N_12866);
or U14161 (N_14161,N_12636,N_12613);
nand U14162 (N_14162,N_13100,N_13473);
nand U14163 (N_14163,N_13158,N_12873);
nand U14164 (N_14164,N_12422,N_13112);
nor U14165 (N_14165,N_12645,N_12294);
nor U14166 (N_14166,N_12717,N_12318);
or U14167 (N_14167,N_12027,N_13059);
or U14168 (N_14168,N_12002,N_12823);
nand U14169 (N_14169,N_13152,N_13372);
nand U14170 (N_14170,N_13124,N_12526);
nand U14171 (N_14171,N_13491,N_12438);
nor U14172 (N_14172,N_12038,N_12006);
nor U14173 (N_14173,N_12858,N_12577);
nor U14174 (N_14174,N_13296,N_13040);
nor U14175 (N_14175,N_12105,N_12265);
nor U14176 (N_14176,N_13127,N_13289);
and U14177 (N_14177,N_12537,N_13410);
or U14178 (N_14178,N_12005,N_12849);
nand U14179 (N_14179,N_12233,N_12894);
nand U14180 (N_14180,N_12800,N_13211);
nand U14181 (N_14181,N_12450,N_12195);
and U14182 (N_14182,N_13069,N_13034);
or U14183 (N_14183,N_12612,N_13375);
and U14184 (N_14184,N_13010,N_12029);
nand U14185 (N_14185,N_12600,N_12770);
nor U14186 (N_14186,N_13204,N_12274);
and U14187 (N_14187,N_13415,N_12042);
nor U14188 (N_14188,N_13175,N_12465);
and U14189 (N_14189,N_12618,N_12094);
nor U14190 (N_14190,N_12357,N_13007);
nor U14191 (N_14191,N_12178,N_12477);
nand U14192 (N_14192,N_12891,N_12810);
and U14193 (N_14193,N_13171,N_12953);
nor U14194 (N_14194,N_12078,N_12930);
nand U14195 (N_14195,N_13342,N_12946);
and U14196 (N_14196,N_12119,N_13333);
and U14197 (N_14197,N_13065,N_12505);
and U14198 (N_14198,N_13298,N_13324);
or U14199 (N_14199,N_12026,N_12441);
nor U14200 (N_14200,N_13192,N_12628);
and U14201 (N_14201,N_12133,N_13456);
or U14202 (N_14202,N_12282,N_12924);
and U14203 (N_14203,N_12678,N_13016);
or U14204 (N_14204,N_12238,N_12410);
nor U14205 (N_14205,N_13205,N_12637);
nor U14206 (N_14206,N_13176,N_12656);
or U14207 (N_14207,N_12043,N_12626);
nand U14208 (N_14208,N_12553,N_12857);
nand U14209 (N_14209,N_13015,N_13498);
xor U14210 (N_14210,N_12541,N_12614);
and U14211 (N_14211,N_13463,N_13258);
nand U14212 (N_14212,N_12201,N_13188);
nor U14213 (N_14213,N_12850,N_12084);
or U14214 (N_14214,N_13341,N_13326);
nand U14215 (N_14215,N_13292,N_12314);
and U14216 (N_14216,N_13145,N_12406);
nor U14217 (N_14217,N_12053,N_13025);
or U14218 (N_14218,N_12345,N_13398);
xnor U14219 (N_14219,N_13368,N_12413);
nand U14220 (N_14220,N_12522,N_12869);
or U14221 (N_14221,N_12399,N_12392);
or U14222 (N_14222,N_12012,N_12761);
or U14223 (N_14223,N_13328,N_13094);
and U14224 (N_14224,N_12065,N_12061);
nor U14225 (N_14225,N_12079,N_12799);
nor U14226 (N_14226,N_12495,N_12596);
nand U14227 (N_14227,N_12926,N_12339);
nand U14228 (N_14228,N_12390,N_13172);
and U14229 (N_14229,N_13032,N_12830);
nor U14230 (N_14230,N_12387,N_13249);
nor U14231 (N_14231,N_12219,N_12725);
nand U14232 (N_14232,N_12337,N_12271);
and U14233 (N_14233,N_12309,N_12909);
or U14234 (N_14234,N_12312,N_12434);
nand U14235 (N_14235,N_12243,N_13102);
nor U14236 (N_14236,N_12418,N_13087);
nor U14237 (N_14237,N_12486,N_13437);
nand U14238 (N_14238,N_12321,N_13294);
nand U14239 (N_14239,N_13243,N_13308);
and U14240 (N_14240,N_12804,N_12047);
nand U14241 (N_14241,N_12453,N_12573);
and U14242 (N_14242,N_12726,N_12074);
or U14243 (N_14243,N_13163,N_13345);
nand U14244 (N_14244,N_13322,N_12204);
or U14245 (N_14245,N_12140,N_12911);
nand U14246 (N_14246,N_13431,N_12089);
nand U14247 (N_14247,N_13364,N_13070);
or U14248 (N_14248,N_13305,N_12408);
nand U14249 (N_14249,N_12072,N_13312);
and U14250 (N_14250,N_12466,N_13140);
nor U14251 (N_14251,N_12784,N_13097);
xor U14252 (N_14252,N_12543,N_12648);
or U14253 (N_14253,N_13119,N_13146);
or U14254 (N_14254,N_12613,N_13120);
or U14255 (N_14255,N_13354,N_13016);
and U14256 (N_14256,N_13067,N_13291);
and U14257 (N_14257,N_12742,N_12318);
or U14258 (N_14258,N_12467,N_12102);
nand U14259 (N_14259,N_13395,N_12560);
and U14260 (N_14260,N_12381,N_12069);
and U14261 (N_14261,N_12970,N_12095);
and U14262 (N_14262,N_12998,N_13430);
nand U14263 (N_14263,N_13372,N_13281);
or U14264 (N_14264,N_12062,N_13133);
or U14265 (N_14265,N_12776,N_12611);
or U14266 (N_14266,N_12804,N_13412);
nand U14267 (N_14267,N_12863,N_12281);
or U14268 (N_14268,N_12745,N_12361);
nand U14269 (N_14269,N_12851,N_13116);
or U14270 (N_14270,N_12575,N_12634);
nor U14271 (N_14271,N_12632,N_12845);
or U14272 (N_14272,N_12627,N_12818);
nand U14273 (N_14273,N_12179,N_12747);
and U14274 (N_14274,N_12224,N_12017);
nor U14275 (N_14275,N_12492,N_13237);
or U14276 (N_14276,N_12632,N_12318);
and U14277 (N_14277,N_12260,N_12204);
or U14278 (N_14278,N_12003,N_12706);
or U14279 (N_14279,N_12180,N_12844);
or U14280 (N_14280,N_12627,N_13261);
nor U14281 (N_14281,N_13499,N_13230);
nor U14282 (N_14282,N_12272,N_12779);
nor U14283 (N_14283,N_13057,N_13089);
nand U14284 (N_14284,N_13154,N_12724);
and U14285 (N_14285,N_12536,N_13219);
nand U14286 (N_14286,N_13277,N_12843);
nand U14287 (N_14287,N_12690,N_12110);
nor U14288 (N_14288,N_13068,N_12025);
or U14289 (N_14289,N_13029,N_13276);
nand U14290 (N_14290,N_13249,N_13177);
nand U14291 (N_14291,N_12637,N_12904);
nor U14292 (N_14292,N_12615,N_12244);
nand U14293 (N_14293,N_13176,N_12917);
or U14294 (N_14294,N_13112,N_13121);
nand U14295 (N_14295,N_12298,N_13375);
nor U14296 (N_14296,N_12969,N_13395);
and U14297 (N_14297,N_12929,N_12012);
and U14298 (N_14298,N_13323,N_13474);
nand U14299 (N_14299,N_12998,N_12676);
nand U14300 (N_14300,N_12420,N_13334);
nor U14301 (N_14301,N_12857,N_12422);
or U14302 (N_14302,N_13174,N_12072);
or U14303 (N_14303,N_12325,N_13335);
xor U14304 (N_14304,N_13321,N_12368);
nand U14305 (N_14305,N_12839,N_12999);
and U14306 (N_14306,N_13352,N_12995);
nor U14307 (N_14307,N_13348,N_12849);
nand U14308 (N_14308,N_13454,N_12397);
and U14309 (N_14309,N_12821,N_12254);
nor U14310 (N_14310,N_12148,N_12740);
nor U14311 (N_14311,N_12449,N_13204);
nand U14312 (N_14312,N_12028,N_12288);
or U14313 (N_14313,N_13033,N_13429);
and U14314 (N_14314,N_12686,N_12820);
nand U14315 (N_14315,N_12018,N_13276);
xor U14316 (N_14316,N_13431,N_12580);
nor U14317 (N_14317,N_12266,N_12051);
nand U14318 (N_14318,N_12924,N_13100);
nor U14319 (N_14319,N_13275,N_13103);
nand U14320 (N_14320,N_13329,N_12797);
nand U14321 (N_14321,N_13238,N_13338);
and U14322 (N_14322,N_12563,N_13477);
and U14323 (N_14323,N_12997,N_12650);
and U14324 (N_14324,N_13222,N_12072);
nand U14325 (N_14325,N_12055,N_12494);
or U14326 (N_14326,N_12534,N_13004);
nand U14327 (N_14327,N_12915,N_13384);
or U14328 (N_14328,N_13449,N_12393);
nor U14329 (N_14329,N_12812,N_12765);
or U14330 (N_14330,N_12670,N_12716);
xor U14331 (N_14331,N_12753,N_12051);
and U14332 (N_14332,N_12345,N_12351);
and U14333 (N_14333,N_12961,N_12411);
nand U14334 (N_14334,N_12476,N_12600);
nor U14335 (N_14335,N_13113,N_13397);
nand U14336 (N_14336,N_12295,N_12216);
and U14337 (N_14337,N_12687,N_12481);
or U14338 (N_14338,N_13198,N_12206);
nor U14339 (N_14339,N_13112,N_12744);
nand U14340 (N_14340,N_12574,N_12761);
or U14341 (N_14341,N_13090,N_12346);
nor U14342 (N_14342,N_13299,N_12042);
nor U14343 (N_14343,N_12521,N_12023);
and U14344 (N_14344,N_12011,N_13183);
nor U14345 (N_14345,N_12474,N_13087);
nor U14346 (N_14346,N_13187,N_13392);
or U14347 (N_14347,N_13086,N_12883);
nor U14348 (N_14348,N_13487,N_13155);
nand U14349 (N_14349,N_13040,N_12054);
nor U14350 (N_14350,N_12857,N_12279);
or U14351 (N_14351,N_12666,N_12689);
nor U14352 (N_14352,N_13353,N_13332);
nor U14353 (N_14353,N_13473,N_12682);
or U14354 (N_14354,N_12254,N_12685);
and U14355 (N_14355,N_12983,N_12228);
nand U14356 (N_14356,N_12566,N_13301);
nand U14357 (N_14357,N_12892,N_12301);
nand U14358 (N_14358,N_12985,N_13444);
and U14359 (N_14359,N_12572,N_13045);
or U14360 (N_14360,N_13238,N_13101);
nand U14361 (N_14361,N_12627,N_12633);
nor U14362 (N_14362,N_13483,N_12249);
nand U14363 (N_14363,N_12876,N_13318);
nand U14364 (N_14364,N_12717,N_12670);
or U14365 (N_14365,N_13261,N_13335);
nor U14366 (N_14366,N_12548,N_13404);
nand U14367 (N_14367,N_13206,N_12157);
and U14368 (N_14368,N_12362,N_13450);
and U14369 (N_14369,N_13070,N_12270);
nand U14370 (N_14370,N_12920,N_12598);
nand U14371 (N_14371,N_13196,N_13144);
nand U14372 (N_14372,N_13090,N_12759);
nand U14373 (N_14373,N_12944,N_13167);
or U14374 (N_14374,N_12847,N_12288);
nor U14375 (N_14375,N_12806,N_12188);
nor U14376 (N_14376,N_12993,N_12477);
or U14377 (N_14377,N_12542,N_12096);
and U14378 (N_14378,N_13069,N_13365);
nand U14379 (N_14379,N_13016,N_12721);
nand U14380 (N_14380,N_12685,N_12079);
nor U14381 (N_14381,N_12375,N_13175);
nor U14382 (N_14382,N_12942,N_13120);
or U14383 (N_14383,N_13376,N_12728);
nand U14384 (N_14384,N_13039,N_12609);
or U14385 (N_14385,N_12104,N_13266);
or U14386 (N_14386,N_12826,N_13471);
nand U14387 (N_14387,N_13097,N_12297);
and U14388 (N_14388,N_13399,N_13065);
nand U14389 (N_14389,N_12008,N_13220);
nor U14390 (N_14390,N_13034,N_13276);
and U14391 (N_14391,N_13111,N_13073);
or U14392 (N_14392,N_12288,N_12946);
nor U14393 (N_14393,N_13492,N_12527);
and U14394 (N_14394,N_12474,N_13306);
nand U14395 (N_14395,N_12442,N_12432);
nor U14396 (N_14396,N_12834,N_13079);
and U14397 (N_14397,N_13254,N_12458);
or U14398 (N_14398,N_12697,N_12468);
and U14399 (N_14399,N_12193,N_12555);
and U14400 (N_14400,N_13302,N_12809);
or U14401 (N_14401,N_13468,N_13237);
and U14402 (N_14402,N_12105,N_12895);
or U14403 (N_14403,N_13393,N_13178);
nand U14404 (N_14404,N_12626,N_12755);
nor U14405 (N_14405,N_13238,N_12947);
nor U14406 (N_14406,N_12848,N_12827);
or U14407 (N_14407,N_13017,N_13261);
and U14408 (N_14408,N_12404,N_12268);
nor U14409 (N_14409,N_12639,N_12111);
and U14410 (N_14410,N_12058,N_12816);
nor U14411 (N_14411,N_13396,N_12815);
nand U14412 (N_14412,N_12185,N_12837);
nand U14413 (N_14413,N_12510,N_12329);
and U14414 (N_14414,N_12275,N_12441);
or U14415 (N_14415,N_13141,N_12283);
and U14416 (N_14416,N_12264,N_12272);
and U14417 (N_14417,N_13436,N_12190);
and U14418 (N_14418,N_12372,N_13395);
and U14419 (N_14419,N_12535,N_13164);
and U14420 (N_14420,N_12932,N_12476);
and U14421 (N_14421,N_12420,N_12406);
nand U14422 (N_14422,N_13341,N_13346);
nand U14423 (N_14423,N_13126,N_13288);
nor U14424 (N_14424,N_12617,N_12538);
and U14425 (N_14425,N_13445,N_12744);
or U14426 (N_14426,N_12493,N_13434);
nor U14427 (N_14427,N_12824,N_12893);
and U14428 (N_14428,N_12414,N_13247);
and U14429 (N_14429,N_12293,N_12581);
nand U14430 (N_14430,N_13473,N_12522);
nand U14431 (N_14431,N_12624,N_12030);
nand U14432 (N_14432,N_12126,N_12075);
nand U14433 (N_14433,N_13265,N_13206);
or U14434 (N_14434,N_13447,N_13397);
or U14435 (N_14435,N_12351,N_12986);
xnor U14436 (N_14436,N_13005,N_12152);
and U14437 (N_14437,N_12663,N_12627);
nor U14438 (N_14438,N_13309,N_13057);
and U14439 (N_14439,N_12468,N_12091);
or U14440 (N_14440,N_12591,N_13468);
and U14441 (N_14441,N_13333,N_13101);
nor U14442 (N_14442,N_12527,N_12354);
nor U14443 (N_14443,N_13414,N_13368);
nor U14444 (N_14444,N_12739,N_13048);
and U14445 (N_14445,N_13434,N_13350);
xnor U14446 (N_14446,N_13064,N_12624);
nor U14447 (N_14447,N_12723,N_12306);
or U14448 (N_14448,N_13314,N_13017);
nand U14449 (N_14449,N_13094,N_13362);
or U14450 (N_14450,N_13235,N_12314);
nand U14451 (N_14451,N_13107,N_12933);
and U14452 (N_14452,N_12154,N_12676);
and U14453 (N_14453,N_13212,N_12781);
nor U14454 (N_14454,N_13114,N_13101);
and U14455 (N_14455,N_12129,N_12193);
and U14456 (N_14456,N_12672,N_12585);
or U14457 (N_14457,N_12406,N_12581);
nand U14458 (N_14458,N_13087,N_12063);
or U14459 (N_14459,N_13056,N_12655);
or U14460 (N_14460,N_12047,N_12338);
or U14461 (N_14461,N_12419,N_12183);
and U14462 (N_14462,N_12709,N_13499);
and U14463 (N_14463,N_12243,N_12414);
nor U14464 (N_14464,N_12719,N_12444);
and U14465 (N_14465,N_13342,N_13034);
nand U14466 (N_14466,N_12205,N_13316);
or U14467 (N_14467,N_12216,N_12118);
or U14468 (N_14468,N_12773,N_12895);
nor U14469 (N_14469,N_13431,N_13028);
nor U14470 (N_14470,N_13237,N_12529);
nor U14471 (N_14471,N_12642,N_13369);
nand U14472 (N_14472,N_13066,N_12512);
nor U14473 (N_14473,N_12304,N_12971);
nor U14474 (N_14474,N_12448,N_13067);
nor U14475 (N_14475,N_13349,N_12463);
and U14476 (N_14476,N_13264,N_12185);
nand U14477 (N_14477,N_13330,N_12494);
and U14478 (N_14478,N_12942,N_13261);
nand U14479 (N_14479,N_13019,N_12534);
or U14480 (N_14480,N_13186,N_13436);
nand U14481 (N_14481,N_12083,N_12840);
or U14482 (N_14482,N_12090,N_13089);
nor U14483 (N_14483,N_13491,N_12626);
nor U14484 (N_14484,N_12403,N_12871);
or U14485 (N_14485,N_12105,N_13478);
or U14486 (N_14486,N_13376,N_13035);
and U14487 (N_14487,N_13034,N_12371);
nor U14488 (N_14488,N_13015,N_12237);
xnor U14489 (N_14489,N_13317,N_13432);
or U14490 (N_14490,N_12833,N_12278);
or U14491 (N_14491,N_12838,N_13047);
or U14492 (N_14492,N_12712,N_12227);
and U14493 (N_14493,N_12418,N_13023);
or U14494 (N_14494,N_12420,N_12364);
and U14495 (N_14495,N_13103,N_13380);
or U14496 (N_14496,N_13291,N_12733);
nor U14497 (N_14497,N_13371,N_12272);
nor U14498 (N_14498,N_13334,N_12717);
nand U14499 (N_14499,N_12358,N_13422);
or U14500 (N_14500,N_13151,N_12569);
or U14501 (N_14501,N_13063,N_13269);
nand U14502 (N_14502,N_13386,N_12738);
nand U14503 (N_14503,N_12377,N_13016);
nor U14504 (N_14504,N_12815,N_12464);
nor U14505 (N_14505,N_12653,N_13125);
or U14506 (N_14506,N_12482,N_13383);
or U14507 (N_14507,N_12422,N_12340);
nand U14508 (N_14508,N_13332,N_12728);
nand U14509 (N_14509,N_13218,N_12053);
nor U14510 (N_14510,N_13143,N_13184);
and U14511 (N_14511,N_12948,N_12009);
nand U14512 (N_14512,N_12026,N_13241);
nor U14513 (N_14513,N_12679,N_12673);
or U14514 (N_14514,N_12576,N_13304);
nand U14515 (N_14515,N_12100,N_13419);
nand U14516 (N_14516,N_12194,N_12588);
and U14517 (N_14517,N_12491,N_12727);
or U14518 (N_14518,N_12303,N_13277);
or U14519 (N_14519,N_13381,N_13421);
and U14520 (N_14520,N_12340,N_13131);
nor U14521 (N_14521,N_12596,N_12309);
nor U14522 (N_14522,N_12207,N_12018);
nand U14523 (N_14523,N_13383,N_13167);
or U14524 (N_14524,N_12955,N_13176);
nor U14525 (N_14525,N_12978,N_12628);
nor U14526 (N_14526,N_12394,N_13224);
nand U14527 (N_14527,N_12339,N_12847);
xor U14528 (N_14528,N_12157,N_12549);
and U14529 (N_14529,N_12103,N_13320);
or U14530 (N_14530,N_12608,N_12938);
or U14531 (N_14531,N_12047,N_12254);
nor U14532 (N_14532,N_12015,N_13214);
or U14533 (N_14533,N_12991,N_12170);
nand U14534 (N_14534,N_13310,N_12078);
nand U14535 (N_14535,N_12629,N_12560);
nand U14536 (N_14536,N_13341,N_12264);
and U14537 (N_14537,N_12490,N_12130);
nand U14538 (N_14538,N_12647,N_12715);
or U14539 (N_14539,N_13097,N_13273);
nand U14540 (N_14540,N_13276,N_13097);
or U14541 (N_14541,N_12512,N_13305);
or U14542 (N_14542,N_12720,N_12339);
xor U14543 (N_14543,N_12175,N_12743);
nand U14544 (N_14544,N_12213,N_13375);
and U14545 (N_14545,N_12475,N_12203);
nor U14546 (N_14546,N_12307,N_12834);
nor U14547 (N_14547,N_12125,N_12216);
and U14548 (N_14548,N_13155,N_12593);
nand U14549 (N_14549,N_12212,N_12014);
nor U14550 (N_14550,N_12982,N_12172);
or U14551 (N_14551,N_12397,N_12015);
and U14552 (N_14552,N_12662,N_13079);
nand U14553 (N_14553,N_12460,N_12785);
and U14554 (N_14554,N_12991,N_12028);
and U14555 (N_14555,N_12496,N_12945);
and U14556 (N_14556,N_13004,N_12207);
or U14557 (N_14557,N_12239,N_12615);
xor U14558 (N_14558,N_12083,N_12751);
nor U14559 (N_14559,N_13300,N_12661);
nor U14560 (N_14560,N_13432,N_12134);
nand U14561 (N_14561,N_12712,N_13486);
nor U14562 (N_14562,N_12703,N_12202);
nand U14563 (N_14563,N_12813,N_12522);
nand U14564 (N_14564,N_12514,N_12759);
nor U14565 (N_14565,N_13425,N_12033);
or U14566 (N_14566,N_12890,N_13277);
or U14567 (N_14567,N_13319,N_12687);
or U14568 (N_14568,N_12413,N_12405);
nand U14569 (N_14569,N_12594,N_13144);
or U14570 (N_14570,N_12328,N_12189);
nor U14571 (N_14571,N_13042,N_12376);
nor U14572 (N_14572,N_13219,N_12202);
and U14573 (N_14573,N_12681,N_12095);
xor U14574 (N_14574,N_13118,N_13495);
and U14575 (N_14575,N_12265,N_12592);
nor U14576 (N_14576,N_12919,N_12041);
and U14577 (N_14577,N_12232,N_13277);
nand U14578 (N_14578,N_12673,N_12459);
or U14579 (N_14579,N_12229,N_12857);
nor U14580 (N_14580,N_12286,N_13086);
and U14581 (N_14581,N_12904,N_12677);
or U14582 (N_14582,N_12515,N_13466);
or U14583 (N_14583,N_12048,N_13409);
xor U14584 (N_14584,N_12979,N_13432);
nand U14585 (N_14585,N_12028,N_12051);
nand U14586 (N_14586,N_12994,N_12229);
and U14587 (N_14587,N_12783,N_12138);
nand U14588 (N_14588,N_13299,N_12813);
or U14589 (N_14589,N_12164,N_13341);
or U14590 (N_14590,N_12181,N_12216);
nor U14591 (N_14591,N_12629,N_12059);
or U14592 (N_14592,N_13384,N_12866);
nand U14593 (N_14593,N_12859,N_12603);
nor U14594 (N_14594,N_12898,N_12660);
nand U14595 (N_14595,N_12833,N_12941);
and U14596 (N_14596,N_12881,N_13330);
and U14597 (N_14597,N_12228,N_12636);
or U14598 (N_14598,N_12005,N_12685);
and U14599 (N_14599,N_13379,N_13261);
and U14600 (N_14600,N_12261,N_12671);
nand U14601 (N_14601,N_13390,N_12552);
or U14602 (N_14602,N_13206,N_13313);
nand U14603 (N_14603,N_12762,N_12032);
and U14604 (N_14604,N_13297,N_13155);
or U14605 (N_14605,N_13201,N_13069);
xnor U14606 (N_14606,N_13289,N_12595);
and U14607 (N_14607,N_13200,N_12543);
nand U14608 (N_14608,N_12589,N_12573);
or U14609 (N_14609,N_12357,N_12131);
nand U14610 (N_14610,N_12071,N_12497);
xor U14611 (N_14611,N_13332,N_12640);
nand U14612 (N_14612,N_12145,N_13033);
nand U14613 (N_14613,N_12865,N_13130);
nand U14614 (N_14614,N_13440,N_12595);
and U14615 (N_14615,N_12052,N_13376);
nor U14616 (N_14616,N_13135,N_12189);
nor U14617 (N_14617,N_12770,N_12613);
or U14618 (N_14618,N_12114,N_13208);
nor U14619 (N_14619,N_12443,N_12999);
or U14620 (N_14620,N_13499,N_12322);
and U14621 (N_14621,N_12710,N_12325);
or U14622 (N_14622,N_13152,N_13387);
and U14623 (N_14623,N_12239,N_12204);
nand U14624 (N_14624,N_13070,N_13394);
nor U14625 (N_14625,N_12611,N_13461);
or U14626 (N_14626,N_13286,N_12709);
nor U14627 (N_14627,N_13140,N_12639);
or U14628 (N_14628,N_12892,N_12428);
and U14629 (N_14629,N_12338,N_12922);
or U14630 (N_14630,N_13104,N_13092);
nand U14631 (N_14631,N_13295,N_13315);
nand U14632 (N_14632,N_12300,N_12806);
nor U14633 (N_14633,N_12311,N_13034);
or U14634 (N_14634,N_12710,N_12341);
nand U14635 (N_14635,N_12838,N_12776);
nand U14636 (N_14636,N_12746,N_13159);
nor U14637 (N_14637,N_12001,N_12375);
or U14638 (N_14638,N_13332,N_12105);
nor U14639 (N_14639,N_12554,N_12492);
nor U14640 (N_14640,N_12683,N_12565);
nor U14641 (N_14641,N_12291,N_12252);
and U14642 (N_14642,N_12239,N_13062);
nand U14643 (N_14643,N_12008,N_12126);
nor U14644 (N_14644,N_12906,N_12884);
nor U14645 (N_14645,N_13288,N_13435);
nand U14646 (N_14646,N_12289,N_12456);
nor U14647 (N_14647,N_13487,N_12222);
and U14648 (N_14648,N_13340,N_12335);
nand U14649 (N_14649,N_12301,N_12373);
nand U14650 (N_14650,N_12190,N_12501);
or U14651 (N_14651,N_13424,N_13449);
nand U14652 (N_14652,N_12904,N_12058);
and U14653 (N_14653,N_12510,N_13450);
nor U14654 (N_14654,N_12060,N_12833);
nand U14655 (N_14655,N_12564,N_12830);
and U14656 (N_14656,N_12970,N_12844);
nor U14657 (N_14657,N_12143,N_13203);
and U14658 (N_14658,N_13084,N_13337);
nand U14659 (N_14659,N_12300,N_12655);
nand U14660 (N_14660,N_12153,N_12183);
or U14661 (N_14661,N_12963,N_12820);
and U14662 (N_14662,N_12634,N_13106);
nor U14663 (N_14663,N_12345,N_13017);
nand U14664 (N_14664,N_13214,N_12271);
xor U14665 (N_14665,N_12154,N_13314);
or U14666 (N_14666,N_13375,N_12182);
nand U14667 (N_14667,N_12868,N_12411);
or U14668 (N_14668,N_12769,N_12742);
nand U14669 (N_14669,N_13262,N_12787);
and U14670 (N_14670,N_13066,N_12346);
nand U14671 (N_14671,N_12671,N_12041);
or U14672 (N_14672,N_13200,N_12079);
nor U14673 (N_14673,N_12716,N_12639);
or U14674 (N_14674,N_12089,N_13360);
and U14675 (N_14675,N_13056,N_12921);
nand U14676 (N_14676,N_12121,N_12748);
or U14677 (N_14677,N_12589,N_13149);
and U14678 (N_14678,N_13150,N_12664);
and U14679 (N_14679,N_12089,N_13464);
and U14680 (N_14680,N_13224,N_12923);
and U14681 (N_14681,N_13132,N_13030);
or U14682 (N_14682,N_13337,N_12889);
nand U14683 (N_14683,N_12736,N_12130);
and U14684 (N_14684,N_12315,N_12360);
nand U14685 (N_14685,N_12712,N_12763);
and U14686 (N_14686,N_13435,N_13049);
and U14687 (N_14687,N_12994,N_13091);
nor U14688 (N_14688,N_12532,N_13360);
and U14689 (N_14689,N_12514,N_13475);
and U14690 (N_14690,N_12789,N_12391);
or U14691 (N_14691,N_12348,N_12703);
and U14692 (N_14692,N_12540,N_12929);
nand U14693 (N_14693,N_12051,N_13186);
and U14694 (N_14694,N_13122,N_13111);
nand U14695 (N_14695,N_12919,N_12233);
and U14696 (N_14696,N_13460,N_13348);
nor U14697 (N_14697,N_12164,N_13113);
nand U14698 (N_14698,N_12751,N_12617);
or U14699 (N_14699,N_12893,N_13217);
nor U14700 (N_14700,N_13305,N_13154);
and U14701 (N_14701,N_12284,N_13399);
and U14702 (N_14702,N_13120,N_12000);
and U14703 (N_14703,N_12888,N_12022);
and U14704 (N_14704,N_12508,N_12612);
nor U14705 (N_14705,N_13270,N_12077);
and U14706 (N_14706,N_12513,N_12045);
or U14707 (N_14707,N_12322,N_13072);
nand U14708 (N_14708,N_13399,N_13266);
or U14709 (N_14709,N_12942,N_13415);
and U14710 (N_14710,N_12818,N_13496);
nor U14711 (N_14711,N_12726,N_12265);
nand U14712 (N_14712,N_12589,N_12423);
nor U14713 (N_14713,N_13436,N_13244);
nor U14714 (N_14714,N_12925,N_12876);
and U14715 (N_14715,N_13309,N_12080);
nand U14716 (N_14716,N_13058,N_13131);
and U14717 (N_14717,N_13482,N_12040);
or U14718 (N_14718,N_12395,N_12315);
or U14719 (N_14719,N_13066,N_12119);
or U14720 (N_14720,N_12158,N_13117);
or U14721 (N_14721,N_12409,N_13487);
nand U14722 (N_14722,N_13146,N_12012);
nor U14723 (N_14723,N_13485,N_12510);
or U14724 (N_14724,N_12839,N_13157);
nand U14725 (N_14725,N_12323,N_13221);
nand U14726 (N_14726,N_13439,N_12684);
nor U14727 (N_14727,N_13024,N_12162);
xnor U14728 (N_14728,N_12879,N_12895);
and U14729 (N_14729,N_12539,N_12463);
nor U14730 (N_14730,N_13141,N_12515);
nor U14731 (N_14731,N_12857,N_12514);
or U14732 (N_14732,N_12347,N_12578);
nor U14733 (N_14733,N_13467,N_12436);
or U14734 (N_14734,N_12293,N_12407);
and U14735 (N_14735,N_12035,N_12735);
or U14736 (N_14736,N_12199,N_12289);
nor U14737 (N_14737,N_12812,N_13373);
nand U14738 (N_14738,N_12979,N_12194);
nor U14739 (N_14739,N_12864,N_12948);
nor U14740 (N_14740,N_12753,N_12055);
nor U14741 (N_14741,N_12200,N_12713);
nand U14742 (N_14742,N_12343,N_13200);
nor U14743 (N_14743,N_12935,N_13291);
nand U14744 (N_14744,N_12490,N_12595);
or U14745 (N_14745,N_13347,N_12855);
and U14746 (N_14746,N_12251,N_13358);
and U14747 (N_14747,N_13123,N_12552);
nor U14748 (N_14748,N_13142,N_13187);
and U14749 (N_14749,N_12281,N_12413);
nand U14750 (N_14750,N_12112,N_12425);
or U14751 (N_14751,N_13267,N_13135);
xnor U14752 (N_14752,N_12147,N_12484);
and U14753 (N_14753,N_13167,N_12998);
nand U14754 (N_14754,N_13126,N_12266);
nand U14755 (N_14755,N_12183,N_12423);
nor U14756 (N_14756,N_12854,N_12202);
nor U14757 (N_14757,N_13412,N_13216);
nand U14758 (N_14758,N_13006,N_13204);
nor U14759 (N_14759,N_12842,N_13411);
and U14760 (N_14760,N_13482,N_12331);
nor U14761 (N_14761,N_13038,N_12890);
nand U14762 (N_14762,N_13407,N_12970);
nor U14763 (N_14763,N_12312,N_13336);
nor U14764 (N_14764,N_12491,N_13218);
and U14765 (N_14765,N_13416,N_12179);
and U14766 (N_14766,N_13304,N_13442);
xnor U14767 (N_14767,N_12962,N_12505);
or U14768 (N_14768,N_12498,N_12872);
nor U14769 (N_14769,N_12304,N_13248);
nor U14770 (N_14770,N_12331,N_12055);
and U14771 (N_14771,N_12384,N_12614);
nand U14772 (N_14772,N_12888,N_13451);
nor U14773 (N_14773,N_12337,N_13281);
nand U14774 (N_14774,N_12629,N_12053);
nor U14775 (N_14775,N_12026,N_12498);
or U14776 (N_14776,N_13447,N_12110);
or U14777 (N_14777,N_12785,N_13194);
nor U14778 (N_14778,N_12526,N_13006);
nor U14779 (N_14779,N_12993,N_12064);
or U14780 (N_14780,N_13431,N_12120);
nand U14781 (N_14781,N_13446,N_12236);
or U14782 (N_14782,N_13330,N_12804);
and U14783 (N_14783,N_13282,N_12823);
nand U14784 (N_14784,N_13342,N_13025);
or U14785 (N_14785,N_13056,N_13028);
nand U14786 (N_14786,N_12428,N_13423);
nor U14787 (N_14787,N_13056,N_12483);
and U14788 (N_14788,N_13357,N_12019);
and U14789 (N_14789,N_12142,N_12777);
or U14790 (N_14790,N_12046,N_13097);
nand U14791 (N_14791,N_13311,N_12713);
nor U14792 (N_14792,N_13058,N_12106);
or U14793 (N_14793,N_13433,N_13116);
and U14794 (N_14794,N_12389,N_13055);
xor U14795 (N_14795,N_12043,N_12673);
and U14796 (N_14796,N_12891,N_13432);
and U14797 (N_14797,N_12482,N_13352);
and U14798 (N_14798,N_12974,N_13264);
nor U14799 (N_14799,N_12284,N_12231);
and U14800 (N_14800,N_13281,N_12227);
nor U14801 (N_14801,N_13175,N_13247);
nand U14802 (N_14802,N_12982,N_13002);
or U14803 (N_14803,N_12677,N_13097);
and U14804 (N_14804,N_13072,N_13236);
nor U14805 (N_14805,N_13400,N_12275);
and U14806 (N_14806,N_12064,N_12457);
nor U14807 (N_14807,N_12146,N_12790);
nor U14808 (N_14808,N_12875,N_12252);
or U14809 (N_14809,N_12425,N_12689);
and U14810 (N_14810,N_12553,N_12945);
nor U14811 (N_14811,N_12926,N_13398);
or U14812 (N_14812,N_12610,N_13008);
nand U14813 (N_14813,N_13076,N_12882);
nand U14814 (N_14814,N_13019,N_12435);
nand U14815 (N_14815,N_12489,N_12770);
or U14816 (N_14816,N_13351,N_12276);
or U14817 (N_14817,N_12623,N_12675);
nand U14818 (N_14818,N_12920,N_12717);
or U14819 (N_14819,N_12610,N_12151);
nand U14820 (N_14820,N_12246,N_12452);
nor U14821 (N_14821,N_12506,N_13464);
nand U14822 (N_14822,N_13144,N_12657);
nand U14823 (N_14823,N_12983,N_12169);
and U14824 (N_14824,N_12915,N_13389);
nor U14825 (N_14825,N_12269,N_12342);
and U14826 (N_14826,N_12122,N_12030);
or U14827 (N_14827,N_13135,N_12957);
and U14828 (N_14828,N_13432,N_12432);
xnor U14829 (N_14829,N_12007,N_12586);
nor U14830 (N_14830,N_12895,N_13094);
or U14831 (N_14831,N_12688,N_12048);
or U14832 (N_14832,N_13271,N_12024);
and U14833 (N_14833,N_13081,N_13138);
and U14834 (N_14834,N_12911,N_13125);
nor U14835 (N_14835,N_12175,N_12345);
or U14836 (N_14836,N_12508,N_12860);
xnor U14837 (N_14837,N_12426,N_12256);
xor U14838 (N_14838,N_13311,N_13242);
nor U14839 (N_14839,N_13134,N_12674);
nor U14840 (N_14840,N_13208,N_12367);
and U14841 (N_14841,N_12798,N_12533);
nand U14842 (N_14842,N_13286,N_12100);
or U14843 (N_14843,N_12576,N_12415);
xor U14844 (N_14844,N_12197,N_12527);
and U14845 (N_14845,N_12781,N_12148);
or U14846 (N_14846,N_12155,N_12202);
nor U14847 (N_14847,N_13421,N_12207);
nand U14848 (N_14848,N_12982,N_12876);
nor U14849 (N_14849,N_12593,N_13006);
and U14850 (N_14850,N_13146,N_12568);
and U14851 (N_14851,N_12277,N_13285);
and U14852 (N_14852,N_12318,N_12719);
nor U14853 (N_14853,N_13439,N_12445);
nand U14854 (N_14854,N_13311,N_13251);
and U14855 (N_14855,N_12659,N_13462);
and U14856 (N_14856,N_13003,N_12791);
nor U14857 (N_14857,N_13431,N_12333);
nand U14858 (N_14858,N_12372,N_12727);
or U14859 (N_14859,N_13426,N_12700);
and U14860 (N_14860,N_12052,N_12214);
or U14861 (N_14861,N_12815,N_12064);
and U14862 (N_14862,N_12167,N_12914);
nor U14863 (N_14863,N_13346,N_13064);
and U14864 (N_14864,N_13079,N_13261);
or U14865 (N_14865,N_12186,N_12118);
or U14866 (N_14866,N_12454,N_12689);
and U14867 (N_14867,N_12452,N_13496);
nand U14868 (N_14868,N_13117,N_13265);
and U14869 (N_14869,N_12367,N_13173);
nand U14870 (N_14870,N_12284,N_13408);
and U14871 (N_14871,N_12267,N_13244);
or U14872 (N_14872,N_12812,N_13379);
nor U14873 (N_14873,N_12280,N_13402);
and U14874 (N_14874,N_13068,N_12277);
or U14875 (N_14875,N_12870,N_12396);
or U14876 (N_14876,N_12424,N_13380);
nand U14877 (N_14877,N_12640,N_13241);
or U14878 (N_14878,N_12267,N_12855);
nor U14879 (N_14879,N_13172,N_12585);
or U14880 (N_14880,N_12099,N_13128);
or U14881 (N_14881,N_12990,N_12100);
nor U14882 (N_14882,N_12203,N_12346);
nand U14883 (N_14883,N_13135,N_12667);
and U14884 (N_14884,N_12223,N_12667);
nand U14885 (N_14885,N_12038,N_12183);
nor U14886 (N_14886,N_12663,N_12470);
and U14887 (N_14887,N_12404,N_13468);
or U14888 (N_14888,N_12390,N_12591);
nor U14889 (N_14889,N_12946,N_13079);
or U14890 (N_14890,N_12450,N_12915);
nand U14891 (N_14891,N_12767,N_12640);
nand U14892 (N_14892,N_12911,N_12836);
or U14893 (N_14893,N_12162,N_13169);
or U14894 (N_14894,N_12831,N_12515);
or U14895 (N_14895,N_13244,N_12303);
or U14896 (N_14896,N_12132,N_13241);
nand U14897 (N_14897,N_12926,N_13125);
nand U14898 (N_14898,N_12088,N_12890);
nor U14899 (N_14899,N_13461,N_12195);
nor U14900 (N_14900,N_12379,N_13124);
nor U14901 (N_14901,N_12454,N_13398);
and U14902 (N_14902,N_12517,N_12941);
or U14903 (N_14903,N_12288,N_12145);
or U14904 (N_14904,N_12502,N_12946);
or U14905 (N_14905,N_12740,N_13417);
or U14906 (N_14906,N_12172,N_13034);
and U14907 (N_14907,N_13283,N_12829);
and U14908 (N_14908,N_12683,N_12046);
nand U14909 (N_14909,N_12304,N_12067);
nor U14910 (N_14910,N_12592,N_13337);
nor U14911 (N_14911,N_12084,N_12392);
nor U14912 (N_14912,N_12430,N_12594);
nor U14913 (N_14913,N_13220,N_13256);
or U14914 (N_14914,N_12838,N_12871);
nor U14915 (N_14915,N_12016,N_12260);
nand U14916 (N_14916,N_13365,N_13451);
or U14917 (N_14917,N_13337,N_12234);
and U14918 (N_14918,N_12414,N_12372);
or U14919 (N_14919,N_13434,N_12115);
nor U14920 (N_14920,N_13245,N_12170);
nor U14921 (N_14921,N_12038,N_13315);
nand U14922 (N_14922,N_13241,N_12793);
or U14923 (N_14923,N_12039,N_12498);
nor U14924 (N_14924,N_12664,N_13085);
xor U14925 (N_14925,N_13437,N_12817);
nor U14926 (N_14926,N_12935,N_12339);
nor U14927 (N_14927,N_13079,N_13085);
nand U14928 (N_14928,N_13401,N_12275);
nand U14929 (N_14929,N_12531,N_13329);
nand U14930 (N_14930,N_13442,N_12147);
or U14931 (N_14931,N_13089,N_12261);
and U14932 (N_14932,N_12715,N_13215);
or U14933 (N_14933,N_12057,N_12613);
or U14934 (N_14934,N_12569,N_12142);
nor U14935 (N_14935,N_12687,N_12997);
and U14936 (N_14936,N_12376,N_12286);
xor U14937 (N_14937,N_12169,N_13477);
or U14938 (N_14938,N_12117,N_13063);
nand U14939 (N_14939,N_13203,N_12741);
nand U14940 (N_14940,N_12452,N_12319);
or U14941 (N_14941,N_13036,N_12960);
and U14942 (N_14942,N_12553,N_13175);
and U14943 (N_14943,N_12340,N_12954);
nand U14944 (N_14944,N_13249,N_12254);
nor U14945 (N_14945,N_12903,N_13313);
and U14946 (N_14946,N_12975,N_13021);
nor U14947 (N_14947,N_13107,N_12843);
nor U14948 (N_14948,N_13151,N_13394);
nor U14949 (N_14949,N_12794,N_12062);
nand U14950 (N_14950,N_13281,N_12214);
or U14951 (N_14951,N_12577,N_12211);
nor U14952 (N_14952,N_13180,N_13358);
and U14953 (N_14953,N_12684,N_13122);
nor U14954 (N_14954,N_12703,N_13227);
nor U14955 (N_14955,N_12574,N_13458);
nor U14956 (N_14956,N_12516,N_13208);
nor U14957 (N_14957,N_12582,N_12064);
nor U14958 (N_14958,N_12431,N_12614);
and U14959 (N_14959,N_12234,N_13335);
and U14960 (N_14960,N_12440,N_12768);
and U14961 (N_14961,N_12702,N_12970);
nor U14962 (N_14962,N_13467,N_13249);
or U14963 (N_14963,N_12926,N_12760);
nand U14964 (N_14964,N_12841,N_13360);
or U14965 (N_14965,N_12334,N_12589);
nor U14966 (N_14966,N_12925,N_13414);
nor U14967 (N_14967,N_13380,N_13490);
nand U14968 (N_14968,N_12834,N_13186);
and U14969 (N_14969,N_12901,N_12645);
or U14970 (N_14970,N_13047,N_12197);
xor U14971 (N_14971,N_12197,N_13366);
nand U14972 (N_14972,N_12192,N_12669);
nor U14973 (N_14973,N_12183,N_13274);
xnor U14974 (N_14974,N_13176,N_13417);
nand U14975 (N_14975,N_12133,N_12725);
nand U14976 (N_14976,N_13168,N_12075);
nand U14977 (N_14977,N_13163,N_12761);
nand U14978 (N_14978,N_12251,N_12412);
nand U14979 (N_14979,N_12096,N_12829);
and U14980 (N_14980,N_13118,N_12256);
and U14981 (N_14981,N_12060,N_12416);
or U14982 (N_14982,N_12716,N_13288);
and U14983 (N_14983,N_13373,N_12052);
xor U14984 (N_14984,N_13228,N_12155);
nor U14985 (N_14985,N_12874,N_13354);
nor U14986 (N_14986,N_13290,N_12235);
nor U14987 (N_14987,N_12094,N_12351);
or U14988 (N_14988,N_12962,N_12383);
nand U14989 (N_14989,N_13190,N_12239);
or U14990 (N_14990,N_12613,N_13381);
nand U14991 (N_14991,N_12041,N_12092);
nor U14992 (N_14992,N_12720,N_12383);
nor U14993 (N_14993,N_12520,N_13095);
nor U14994 (N_14994,N_12331,N_13267);
nand U14995 (N_14995,N_13074,N_12452);
nand U14996 (N_14996,N_12329,N_12156);
xnor U14997 (N_14997,N_13173,N_13362);
nand U14998 (N_14998,N_12295,N_13240);
nor U14999 (N_14999,N_13393,N_13450);
nand UO_0 (O_0,N_14352,N_13755);
and UO_1 (O_1,N_14579,N_14702);
or UO_2 (O_2,N_14479,N_14822);
and UO_3 (O_3,N_14431,N_13991);
or UO_4 (O_4,N_14904,N_14168);
and UO_5 (O_5,N_14187,N_14972);
nor UO_6 (O_6,N_13556,N_14262);
or UO_7 (O_7,N_14940,N_13651);
nand UO_8 (O_8,N_13683,N_14632);
and UO_9 (O_9,N_14865,N_14199);
nor UO_10 (O_10,N_14722,N_14678);
or UO_11 (O_11,N_13828,N_13987);
nor UO_12 (O_12,N_14857,N_13719);
nand UO_13 (O_13,N_13580,N_14365);
nand UO_14 (O_14,N_14984,N_13525);
and UO_15 (O_15,N_14920,N_13748);
nor UO_16 (O_16,N_14967,N_14404);
nand UO_17 (O_17,N_14564,N_14921);
nand UO_18 (O_18,N_14995,N_14955);
and UO_19 (O_19,N_14536,N_13809);
nor UO_20 (O_20,N_13822,N_14739);
or UO_21 (O_21,N_13776,N_14061);
nor UO_22 (O_22,N_13887,N_13905);
nand UO_23 (O_23,N_14785,N_13502);
and UO_24 (O_24,N_14935,N_13765);
or UO_25 (O_25,N_13676,N_13554);
nand UO_26 (O_26,N_14477,N_14381);
nand UO_27 (O_27,N_13654,N_14795);
or UO_28 (O_28,N_13992,N_14213);
nand UO_29 (O_29,N_14566,N_13604);
or UO_30 (O_30,N_14613,N_14724);
or UO_31 (O_31,N_13871,N_14245);
or UO_32 (O_32,N_13607,N_14716);
nor UO_33 (O_33,N_14682,N_13996);
nor UO_34 (O_34,N_13590,N_14417);
nand UO_35 (O_35,N_14472,N_14660);
and UO_36 (O_36,N_14048,N_14686);
or UO_37 (O_37,N_14943,N_13908);
or UO_38 (O_38,N_14309,N_14058);
and UO_39 (O_39,N_14080,N_14898);
xnor UO_40 (O_40,N_13851,N_14528);
nand UO_41 (O_41,N_13726,N_13565);
nor UO_42 (O_42,N_14428,N_14993);
nand UO_43 (O_43,N_14205,N_14620);
nor UO_44 (O_44,N_14779,N_14126);
or UO_45 (O_45,N_13658,N_14375);
nor UO_46 (O_46,N_14176,N_14997);
or UO_47 (O_47,N_14831,N_14546);
or UO_48 (O_48,N_13969,N_14543);
and UO_49 (O_49,N_13513,N_14712);
and UO_50 (O_50,N_14941,N_14774);
and UO_51 (O_51,N_14582,N_14590);
or UO_52 (O_52,N_13617,N_14458);
nand UO_53 (O_53,N_14685,N_14446);
nor UO_54 (O_54,N_13558,N_13818);
or UO_55 (O_55,N_13699,N_13735);
and UO_56 (O_56,N_14122,N_14485);
and UO_57 (O_57,N_14344,N_13797);
and UO_58 (O_58,N_13618,N_13555);
and UO_59 (O_59,N_14082,N_14312);
and UO_60 (O_60,N_14196,N_14848);
nand UO_61 (O_61,N_14743,N_13531);
nor UO_62 (O_62,N_13646,N_14075);
nand UO_63 (O_63,N_14009,N_14515);
nor UO_64 (O_64,N_13904,N_14149);
xnor UO_65 (O_65,N_14958,N_14820);
and UO_66 (O_66,N_14229,N_13725);
nand UO_67 (O_67,N_14760,N_13701);
or UO_68 (O_68,N_14744,N_14527);
nand UO_69 (O_69,N_14944,N_14367);
nand UO_70 (O_70,N_13518,N_14456);
and UO_71 (O_71,N_14704,N_14191);
nand UO_72 (O_72,N_14714,N_14999);
nand UO_73 (O_73,N_13631,N_14088);
and UO_74 (O_74,N_14784,N_13762);
and UO_75 (O_75,N_13856,N_14690);
nor UO_76 (O_76,N_14637,N_14839);
nand UO_77 (O_77,N_13707,N_13613);
nand UO_78 (O_78,N_13913,N_14570);
or UO_79 (O_79,N_14805,N_13847);
nor UO_80 (O_80,N_14235,N_14490);
and UO_81 (O_81,N_14017,N_14541);
nor UO_82 (O_82,N_14110,N_14286);
nor UO_83 (O_83,N_14227,N_14128);
and UO_84 (O_84,N_13626,N_14910);
or UO_85 (O_85,N_14480,N_14254);
nand UO_86 (O_86,N_13655,N_14342);
or UO_87 (O_87,N_14538,N_14347);
or UO_88 (O_88,N_13619,N_14139);
nor UO_89 (O_89,N_13672,N_14019);
or UO_90 (O_90,N_13875,N_14797);
or UO_91 (O_91,N_13694,N_14876);
and UO_92 (O_92,N_14575,N_14137);
or UO_93 (O_93,N_14600,N_14841);
and UO_94 (O_94,N_14288,N_14589);
and UO_95 (O_95,N_13819,N_14932);
or UO_96 (O_96,N_14099,N_14155);
nand UO_97 (O_97,N_14648,N_14074);
or UO_98 (O_98,N_14775,N_14810);
nor UO_99 (O_99,N_14078,N_14809);
and UO_100 (O_100,N_14033,N_13849);
nor UO_101 (O_101,N_13878,N_13840);
xnor UO_102 (O_102,N_14291,N_14409);
nor UO_103 (O_103,N_14406,N_13572);
and UO_104 (O_104,N_13812,N_14355);
nor UO_105 (O_105,N_14946,N_14320);
or UO_106 (O_106,N_14974,N_14448);
nand UO_107 (O_107,N_14786,N_13890);
or UO_108 (O_108,N_14425,N_14952);
nor UO_109 (O_109,N_14497,N_14265);
and UO_110 (O_110,N_14851,N_14526);
or UO_111 (O_111,N_14182,N_13899);
and UO_112 (O_112,N_13528,N_14297);
nor UO_113 (O_113,N_13961,N_13622);
and UO_114 (O_114,N_14387,N_14246);
nor UO_115 (O_115,N_13730,N_14150);
nor UO_116 (O_116,N_14959,N_13564);
nand UO_117 (O_117,N_13820,N_14237);
xor UO_118 (O_118,N_14147,N_14195);
and UO_119 (O_119,N_14443,N_13915);
nor UO_120 (O_120,N_14407,N_13504);
and UO_121 (O_121,N_14811,N_14525);
or UO_122 (O_122,N_14378,N_14449);
nand UO_123 (O_123,N_14450,N_14891);
or UO_124 (O_124,N_14607,N_14234);
xor UO_125 (O_125,N_13743,N_14817);
or UO_126 (O_126,N_14437,N_14430);
and UO_127 (O_127,N_13586,N_14560);
and UO_128 (O_128,N_13722,N_13921);
nand UO_129 (O_129,N_14735,N_13811);
and UO_130 (O_130,N_13608,N_14558);
nand UO_131 (O_131,N_14323,N_14695);
and UO_132 (O_132,N_13951,N_13958);
or UO_133 (O_133,N_14177,N_14498);
and UO_134 (O_134,N_14394,N_13897);
or UO_135 (O_135,N_13581,N_13667);
and UO_136 (O_136,N_14701,N_13761);
or UO_137 (O_137,N_14152,N_13827);
and UO_138 (O_138,N_14516,N_14539);
or UO_139 (O_139,N_13882,N_14217);
or UO_140 (O_140,N_13903,N_14100);
and UO_141 (O_141,N_13954,N_14738);
nand UO_142 (O_142,N_13627,N_13829);
or UO_143 (O_143,N_14687,N_14734);
nand UO_144 (O_144,N_14405,N_13593);
nand UO_145 (O_145,N_14571,N_14872);
nand UO_146 (O_146,N_14986,N_14178);
or UO_147 (O_147,N_14639,N_14509);
nand UO_148 (O_148,N_14753,N_13671);
nor UO_149 (O_149,N_13584,N_14951);
and UO_150 (O_150,N_14064,N_13652);
and UO_151 (O_151,N_14051,N_14487);
or UO_152 (O_152,N_13955,N_14859);
nor UO_153 (O_153,N_14750,N_13937);
xor UO_154 (O_154,N_13749,N_14927);
and UO_155 (O_155,N_14556,N_14204);
nand UO_156 (O_156,N_14386,N_13548);
nand UO_157 (O_157,N_14219,N_13640);
or UO_158 (O_158,N_14518,N_14561);
or UO_159 (O_159,N_14520,N_13912);
nand UO_160 (O_160,N_14231,N_13988);
nor UO_161 (O_161,N_14803,N_14513);
and UO_162 (O_162,N_13984,N_14770);
or UO_163 (O_163,N_14745,N_14053);
and UO_164 (O_164,N_14296,N_13677);
nor UO_165 (O_165,N_14087,N_14138);
or UO_166 (O_166,N_14684,N_13744);
nand UO_167 (O_167,N_14573,N_14511);
nor UO_168 (O_168,N_13850,N_14752);
and UO_169 (O_169,N_14076,N_14843);
nor UO_170 (O_170,N_14190,N_14905);
or UO_171 (O_171,N_14718,N_14079);
nor UO_172 (O_172,N_14292,N_14025);
nand UO_173 (O_173,N_14036,N_14192);
nand UO_174 (O_174,N_13745,N_13509);
nor UO_175 (O_175,N_14090,N_13876);
nor UO_176 (O_176,N_14243,N_13968);
nand UO_177 (O_177,N_14433,N_14228);
nor UO_178 (O_178,N_13634,N_14798);
nor UO_179 (O_179,N_13536,N_13709);
nor UO_180 (O_180,N_14316,N_14978);
nand UO_181 (O_181,N_13643,N_14812);
nor UO_182 (O_182,N_14066,N_14141);
and UO_183 (O_183,N_14844,N_14041);
nand UO_184 (O_184,N_14277,N_14188);
and UO_185 (O_185,N_13893,N_13734);
or UO_186 (O_186,N_13663,N_14880);
nand UO_187 (O_187,N_14395,N_14358);
nor UO_188 (O_188,N_13886,N_14555);
and UO_189 (O_189,N_13546,N_14062);
or UO_190 (O_190,N_14635,N_14484);
nor UO_191 (O_191,N_14112,N_13834);
nand UO_192 (O_192,N_13680,N_14736);
nand UO_193 (O_193,N_13506,N_14623);
or UO_194 (O_194,N_14102,N_13629);
nand UO_195 (O_195,N_14045,N_13741);
and UO_196 (O_196,N_13610,N_14432);
or UO_197 (O_197,N_13967,N_14504);
or UO_198 (O_198,N_14181,N_13540);
nand UO_199 (O_199,N_14317,N_14366);
nor UO_200 (O_200,N_14963,N_14689);
nor UO_201 (O_201,N_14183,N_14596);
or UO_202 (O_202,N_13616,N_14728);
or UO_203 (O_203,N_14936,N_14002);
nor UO_204 (O_204,N_13925,N_13858);
nand UO_205 (O_205,N_13990,N_13807);
nor UO_206 (O_206,N_14072,N_14343);
or UO_207 (O_207,N_14574,N_14424);
and UO_208 (O_208,N_13798,N_14514);
nand UO_209 (O_209,N_13630,N_13869);
and UO_210 (O_210,N_14890,N_14934);
and UO_211 (O_211,N_14824,N_13830);
nand UO_212 (O_212,N_14136,N_14962);
nor UO_213 (O_213,N_13611,N_13963);
and UO_214 (O_214,N_14447,N_14715);
and UO_215 (O_215,N_14521,N_14801);
or UO_216 (O_216,N_14998,N_13939);
nand UO_217 (O_217,N_14842,N_14250);
or UO_218 (O_218,N_13585,N_14029);
and UO_219 (O_219,N_14011,N_14376);
nor UO_220 (O_220,N_14808,N_13678);
or UO_221 (O_221,N_14725,N_13980);
nand UO_222 (O_222,N_13911,N_14979);
or UO_223 (O_223,N_14057,N_14151);
nor UO_224 (O_224,N_13845,N_14120);
nand UO_225 (O_225,N_14609,N_13567);
and UO_226 (O_226,N_13774,N_14629);
nor UO_227 (O_227,N_14005,N_13753);
and UO_228 (O_228,N_13932,N_14906);
or UO_229 (O_229,N_13816,N_13520);
nand UO_230 (O_230,N_14044,N_13810);
xor UO_231 (O_231,N_14697,N_14481);
or UO_232 (O_232,N_14020,N_14069);
nor UO_233 (O_233,N_14391,N_13941);
nor UO_234 (O_234,N_14225,N_14899);
nor UO_235 (O_235,N_13836,N_14721);
or UO_236 (O_236,N_14749,N_14402);
or UO_237 (O_237,N_13620,N_14537);
or UO_238 (O_238,N_14186,N_14608);
or UO_239 (O_239,N_14502,N_14340);
or UO_240 (O_240,N_13979,N_13736);
or UO_241 (O_241,N_13561,N_14757);
nand UO_242 (O_242,N_14656,N_13929);
or UO_243 (O_243,N_13697,N_14866);
nor UO_244 (O_244,N_14293,N_14067);
and UO_245 (O_245,N_14926,N_13790);
nor UO_246 (O_246,N_14956,N_14855);
or UO_247 (O_247,N_13940,N_14755);
xor UO_248 (O_248,N_13718,N_14221);
nand UO_249 (O_249,N_14390,N_14389);
or UO_250 (O_250,N_14506,N_13687);
nor UO_251 (O_251,N_13896,N_14117);
nand UO_252 (O_252,N_14436,N_14094);
nor UO_253 (O_253,N_14948,N_14644);
nor UO_254 (O_254,N_13900,N_14303);
nand UO_255 (O_255,N_13974,N_14026);
or UO_256 (O_256,N_14301,N_13700);
and UO_257 (O_257,N_14883,N_14179);
nand UO_258 (O_258,N_14957,N_14423);
or UO_259 (O_259,N_14706,N_13966);
nand UO_260 (O_260,N_14400,N_14351);
or UO_261 (O_261,N_13832,N_14524);
and UO_262 (O_262,N_13570,N_13599);
nor UO_263 (O_263,N_14258,N_14263);
or UO_264 (O_264,N_14013,N_14233);
nor UO_265 (O_265,N_14161,N_14116);
nor UO_266 (O_266,N_13635,N_14856);
nand UO_267 (O_267,N_13936,N_14175);
or UO_268 (O_268,N_14460,N_14830);
or UO_269 (O_269,N_14794,N_14540);
nand UO_270 (O_270,N_13625,N_14261);
nor UO_271 (O_271,N_14553,N_13842);
and UO_272 (O_272,N_14239,N_14052);
and UO_273 (O_273,N_14070,N_14212);
nand UO_274 (O_274,N_14416,N_14214);
nand UO_275 (O_275,N_14255,N_13956);
and UO_276 (O_276,N_14464,N_14661);
nand UO_277 (O_277,N_14628,N_13727);
nand UO_278 (O_278,N_14396,N_14004);
or UO_279 (O_279,N_14385,N_14457);
or UO_280 (O_280,N_14681,N_14858);
nand UO_281 (O_281,N_14914,N_13614);
nand UO_282 (O_282,N_13571,N_13880);
nor UO_283 (O_283,N_14758,N_13909);
nor UO_284 (O_284,N_14021,N_14162);
and UO_285 (O_285,N_14475,N_14634);
and UO_286 (O_286,N_14220,N_14421);
nor UO_287 (O_287,N_14363,N_14211);
or UO_288 (O_288,N_14969,N_13758);
and UO_289 (O_289,N_13773,N_14298);
and UO_290 (O_290,N_13901,N_14461);
nor UO_291 (O_291,N_14565,N_13542);
nand UO_292 (O_292,N_14332,N_14454);
and UO_293 (O_293,N_13612,N_13597);
or UO_294 (O_294,N_13806,N_14315);
nor UO_295 (O_295,N_13879,N_14157);
xor UO_296 (O_296,N_14991,N_14688);
or UO_297 (O_297,N_14586,N_14707);
nor UO_298 (O_298,N_14499,N_13519);
nand UO_299 (O_299,N_14091,N_14754);
xnor UO_300 (O_300,N_14828,N_14338);
nand UO_301 (O_301,N_14719,N_14170);
or UO_302 (O_302,N_14874,N_14131);
nand UO_303 (O_303,N_13760,N_14278);
xnor UO_304 (O_304,N_14815,N_14331);
or UO_305 (O_305,N_14314,N_14260);
nand UO_306 (O_306,N_14591,N_14937);
nor UO_307 (O_307,N_14581,N_14849);
and UO_308 (O_308,N_13512,N_14203);
and UO_309 (O_309,N_13767,N_14612);
and UO_310 (O_310,N_13777,N_14913);
nor UO_311 (O_311,N_13756,N_13835);
nand UO_312 (O_312,N_13740,N_14223);
or UO_313 (O_313,N_14657,N_14163);
and UO_314 (O_314,N_14452,N_14933);
nand UO_315 (O_315,N_14901,N_14826);
or UO_316 (O_316,N_13641,N_13547);
nand UO_317 (O_317,N_14119,N_14435);
nand UO_318 (O_318,N_14900,N_13587);
nand UO_319 (O_319,N_13867,N_13942);
nand UO_320 (O_320,N_13645,N_14892);
nand UO_321 (O_321,N_14605,N_14960);
or UO_322 (O_322,N_14836,N_14046);
or UO_323 (O_323,N_14881,N_14308);
nor UO_324 (O_324,N_14894,N_14022);
xor UO_325 (O_325,N_14418,N_14101);
nor UO_326 (O_326,N_13803,N_14411);
or UO_327 (O_327,N_14827,N_14024);
and UO_328 (O_328,N_13853,N_13650);
or UO_329 (O_329,N_14542,N_13930);
nand UO_330 (O_330,N_14672,N_13800);
xnor UO_331 (O_331,N_13708,N_14413);
nand UO_332 (O_332,N_13691,N_14791);
nor UO_333 (O_333,N_13737,N_14318);
nand UO_334 (O_334,N_13623,N_14440);
nor UO_335 (O_335,N_14650,N_13831);
and UO_336 (O_336,N_13783,N_13943);
or UO_337 (O_337,N_14471,N_13511);
and UO_338 (O_338,N_13791,N_13993);
nand UO_339 (O_339,N_13795,N_14200);
or UO_340 (O_340,N_14773,N_13959);
nand UO_341 (O_341,N_13573,N_14544);
or UO_342 (O_342,N_14617,N_14085);
nand UO_343 (O_343,N_14732,N_14833);
nor UO_344 (O_344,N_14643,N_13711);
and UO_345 (O_345,N_14121,N_14804);
or UO_346 (O_346,N_14408,N_13872);
nor UO_347 (O_347,N_13589,N_14931);
and UO_348 (O_348,N_13721,N_14208);
nand UO_349 (O_349,N_14086,N_14468);
and UO_350 (O_350,N_14772,N_14924);
nand UO_351 (O_351,N_13891,N_14321);
and UO_352 (O_352,N_14994,N_14180);
nand UO_353 (O_353,N_14923,N_14156);
nand UO_354 (O_354,N_13804,N_14055);
and UO_355 (O_355,N_14124,N_14530);
or UO_356 (O_356,N_13934,N_14267);
nor UO_357 (O_357,N_14185,N_14825);
nand UO_358 (O_358,N_14473,N_13846);
or UO_359 (O_359,N_14114,N_14535);
nor UO_360 (O_360,N_13843,N_13839);
and UO_361 (O_361,N_14765,N_14252);
or UO_362 (O_362,N_13636,N_14135);
nor UO_363 (O_363,N_13778,N_14987);
and UO_364 (O_364,N_13516,N_13799);
or UO_365 (O_365,N_13588,N_13768);
nor UO_366 (O_366,N_14111,N_13595);
nand UO_367 (O_367,N_13949,N_13808);
nand UO_368 (O_368,N_14459,N_13662);
nor UO_369 (O_369,N_13648,N_14942);
or UO_370 (O_370,N_14813,N_13695);
nand UO_371 (O_371,N_14896,N_14769);
nor UO_372 (O_372,N_14105,N_13657);
and UO_373 (O_373,N_13632,N_14368);
nor UO_374 (O_374,N_14703,N_14624);
nand UO_375 (O_375,N_14271,N_14776);
nand UO_376 (O_376,N_14636,N_14799);
nor UO_377 (O_377,N_14976,N_14284);
nor UO_378 (O_378,N_13826,N_13670);
or UO_379 (O_379,N_14938,N_13962);
nand UO_380 (O_380,N_14256,N_13715);
nand UO_381 (O_381,N_14483,N_14253);
and UO_382 (O_382,N_14388,N_14740);
xnor UO_383 (O_383,N_14819,N_14510);
nor UO_384 (O_384,N_13551,N_14621);
xnor UO_385 (O_385,N_13786,N_14383);
and UO_386 (O_386,N_13841,N_13553);
and UO_387 (O_387,N_14563,N_14645);
nor UO_388 (O_388,N_14160,N_14710);
or UO_389 (O_389,N_14130,N_14789);
or UO_390 (O_390,N_13624,N_13888);
nor UO_391 (O_391,N_14860,N_13919);
nand UO_392 (O_392,N_14674,N_14275);
nor UO_393 (O_393,N_14410,N_13639);
nand UO_394 (O_394,N_13682,N_14039);
nor UO_395 (O_395,N_13859,N_13508);
nor UO_396 (O_396,N_13576,N_14653);
nand UO_397 (O_397,N_13649,N_14422);
xnor UO_398 (O_398,N_14796,N_14346);
nand UO_399 (O_399,N_14975,N_13757);
nand UO_400 (O_400,N_14311,N_13574);
and UO_401 (O_401,N_14864,N_13532);
nor UO_402 (O_402,N_13505,N_14207);
or UO_403 (O_403,N_13982,N_14793);
and UO_404 (O_404,N_14006,N_13733);
nor UO_405 (O_405,N_13535,N_14470);
and UO_406 (O_406,N_13659,N_13527);
nor UO_407 (O_407,N_14771,N_13739);
nor UO_408 (O_408,N_13698,N_14042);
and UO_409 (O_409,N_13563,N_14588);
or UO_410 (O_410,N_14154,N_13644);
or UO_411 (O_411,N_13681,N_14299);
nor UO_412 (O_412,N_14414,N_14733);
nor UO_413 (O_413,N_14184,N_13665);
nor UO_414 (O_414,N_14065,N_14083);
nand UO_415 (O_415,N_14647,N_14847);
nor UO_416 (O_416,N_14668,N_14230);
nand UO_417 (O_417,N_14361,N_14427);
and UO_418 (O_418,N_14063,N_14549);
nand UO_419 (O_419,N_13952,N_14691);
nand UO_420 (O_420,N_14916,N_14580);
nor UO_421 (O_421,N_14741,N_14748);
or UO_422 (O_422,N_14335,N_14654);
nand UO_423 (O_423,N_13559,N_14720);
or UO_424 (O_424,N_14907,N_14696);
and UO_425 (O_425,N_13784,N_13601);
and UO_426 (O_426,N_14392,N_14370);
or UO_427 (O_427,N_13781,N_13874);
nand UO_428 (O_428,N_14766,N_14622);
and UO_429 (O_429,N_14353,N_14145);
and UO_430 (O_430,N_13906,N_14992);
and UO_431 (O_431,N_13815,N_13763);
nor UO_432 (O_432,N_14444,N_14306);
or UO_433 (O_433,N_13910,N_14693);
and UO_434 (O_434,N_14218,N_13523);
nor UO_435 (O_435,N_14845,N_14242);
nand UO_436 (O_436,N_14322,N_14206);
or UO_437 (O_437,N_14615,N_13769);
or UO_438 (O_438,N_14763,N_14887);
nor UO_439 (O_439,N_14877,N_14950);
xnor UO_440 (O_440,N_14003,N_14276);
or UO_441 (O_441,N_13865,N_14294);
or UO_442 (O_442,N_14494,N_13950);
or UO_443 (O_443,N_14641,N_14977);
nand UO_444 (O_444,N_13712,N_13823);
nor UO_445 (O_445,N_14867,N_14171);
nand UO_446 (O_446,N_13833,N_14313);
nand UO_447 (O_447,N_13674,N_13738);
nor UO_448 (O_448,N_14194,N_13837);
and UO_449 (O_449,N_14861,N_13923);
nor UO_450 (O_450,N_14599,N_13522);
or UO_451 (O_451,N_14888,N_13653);
and UO_452 (O_452,N_13621,N_14164);
or UO_453 (O_453,N_14533,N_13529);
nor UO_454 (O_454,N_13500,N_14012);
or UO_455 (O_455,N_14167,N_14966);
nor UO_456 (O_456,N_14330,N_13686);
xor UO_457 (O_457,N_13732,N_13751);
nand UO_458 (O_458,N_13945,N_14488);
nor UO_459 (O_459,N_14142,N_14840);
nand UO_460 (O_460,N_14209,N_13821);
nand UO_461 (O_461,N_14625,N_13609);
nand UO_462 (O_462,N_14143,N_14669);
or UO_463 (O_463,N_14982,N_13568);
nor UO_464 (O_464,N_14680,N_13538);
and UO_465 (O_465,N_13503,N_14362);
or UO_466 (O_466,N_13507,N_14531);
nor UO_467 (O_467,N_13550,N_14060);
and UO_468 (O_468,N_14875,N_13539);
nor UO_469 (O_469,N_13717,N_14988);
nor UO_470 (O_470,N_14198,N_14337);
nand UO_471 (O_471,N_14746,N_14215);
and UO_472 (O_472,N_13579,N_14989);
nand UO_473 (O_473,N_14949,N_14897);
nor UO_474 (O_474,N_14731,N_14007);
nand UO_475 (O_475,N_13825,N_13746);
nand UO_476 (O_476,N_14677,N_14837);
nand UO_477 (O_477,N_14601,N_13775);
nand UO_478 (O_478,N_14911,N_14259);
or UO_479 (O_479,N_13881,N_14357);
nor UO_480 (O_480,N_14548,N_13569);
nand UO_481 (O_481,N_14692,N_14534);
or UO_482 (O_482,N_14507,N_14240);
or UO_483 (O_483,N_13583,N_13723);
or UO_484 (O_484,N_14280,N_14882);
or UO_485 (O_485,N_14247,N_14792);
nor UO_486 (O_486,N_14268,N_14850);
nor UO_487 (O_487,N_14584,N_14189);
nor UO_488 (O_488,N_14919,N_13702);
nor UO_489 (O_489,N_13545,N_14282);
nand UO_490 (O_490,N_14971,N_13838);
nor UO_491 (O_491,N_14980,N_13666);
nor UO_492 (O_492,N_14879,N_13747);
nand UO_493 (O_493,N_13917,N_14174);
nand UO_494 (O_494,N_13533,N_14787);
or UO_495 (O_495,N_13852,N_14148);
or UO_496 (O_496,N_14655,N_13537);
nand UO_497 (O_497,N_14216,N_13947);
or UO_498 (O_498,N_14467,N_13928);
or UO_499 (O_499,N_14399,N_14618);
and UO_500 (O_500,N_13927,N_14885);
nor UO_501 (O_501,N_13914,N_14028);
and UO_502 (O_502,N_14492,N_14545);
xor UO_503 (O_503,N_14711,N_14893);
and UO_504 (O_504,N_14382,N_13805);
nand UO_505 (O_505,N_13789,N_14285);
or UO_506 (O_506,N_14983,N_13824);
nor UO_507 (O_507,N_13638,N_14782);
nand UO_508 (O_508,N_14339,N_13530);
nand UO_509 (O_509,N_14158,N_13885);
nand UO_510 (O_510,N_14132,N_14018);
and UO_511 (O_511,N_13892,N_13578);
or UO_512 (O_512,N_14700,N_13637);
nand UO_513 (O_513,N_14649,N_14077);
or UO_514 (O_514,N_14010,N_14598);
nor UO_515 (O_515,N_14939,N_14038);
and UO_516 (O_516,N_14709,N_14035);
nor UO_517 (O_517,N_14153,N_14730);
and UO_518 (O_518,N_13864,N_13675);
or UO_519 (O_519,N_13971,N_14705);
nor UO_520 (O_520,N_13706,N_13884);
and UO_521 (O_521,N_13977,N_13703);
or UO_522 (O_522,N_14445,N_14127);
nor UO_523 (O_523,N_14973,N_14097);
nand UO_524 (O_524,N_14202,N_14310);
or UO_525 (O_525,N_14354,N_14630);
and UO_526 (O_526,N_13592,N_14802);
and UO_527 (O_527,N_14884,N_14104);
nand UO_528 (O_528,N_14326,N_14304);
or UO_529 (O_529,N_14611,N_14360);
nor UO_530 (O_530,N_13877,N_14594);
nor UO_531 (O_531,N_13844,N_14281);
or UO_532 (O_532,N_14846,N_14040);
nand UO_533 (O_533,N_13802,N_14393);
nand UO_534 (O_534,N_14638,N_13656);
nand UO_535 (O_535,N_14054,N_14463);
or UO_536 (O_536,N_14224,N_14756);
xnor UO_537 (O_537,N_13633,N_14587);
nand UO_538 (O_538,N_14290,N_13524);
nand UO_539 (O_539,N_14015,N_13922);
nor UO_540 (O_540,N_14683,N_14415);
and UO_541 (O_541,N_13772,N_14474);
xor UO_542 (O_542,N_13515,N_13948);
nor UO_543 (O_543,N_14210,N_13794);
nand UO_544 (O_544,N_14929,N_14878);
and UO_545 (O_545,N_14325,N_13647);
nor UO_546 (O_546,N_13916,N_14816);
or UO_547 (O_547,N_14166,N_14651);
nor UO_548 (O_548,N_14380,N_14642);
and UO_549 (O_549,N_14412,N_14476);
nand UO_550 (O_550,N_14562,N_14439);
or UO_551 (O_551,N_14532,N_14903);
nor UO_552 (O_552,N_14289,N_14089);
nor UO_553 (O_553,N_13964,N_13920);
nand UO_554 (O_554,N_14547,N_13602);
nand UO_555 (O_555,N_14780,N_14197);
nor UO_556 (O_556,N_14737,N_14781);
nor UO_557 (O_557,N_14662,N_14557);
and UO_558 (O_558,N_14118,N_14713);
nand UO_559 (O_559,N_13575,N_13902);
nand UO_560 (O_560,N_14873,N_14592);
and UO_561 (O_561,N_14800,N_14699);
nand UO_562 (O_562,N_14377,N_14512);
nand UO_563 (O_563,N_13728,N_14401);
nor UO_564 (O_564,N_13521,N_14751);
xnor UO_565 (O_565,N_13861,N_14550);
and UO_566 (O_566,N_14043,N_13673);
and UO_567 (O_567,N_14302,N_14403);
nor UO_568 (O_568,N_14279,N_13972);
nor UO_569 (O_569,N_14001,N_13596);
or UO_570 (O_570,N_13689,N_13679);
nand UO_571 (O_571,N_14031,N_14455);
or UO_572 (O_572,N_13953,N_14783);
nand UO_573 (O_573,N_14863,N_14438);
nor UO_574 (O_574,N_14902,N_13957);
nand UO_575 (O_575,N_14108,N_14451);
or UO_576 (O_576,N_14679,N_14324);
nor UO_577 (O_577,N_14096,N_14868);
and UO_578 (O_578,N_13544,N_13965);
nor UO_579 (O_579,N_14663,N_14222);
or UO_580 (O_580,N_14264,N_14675);
nor UO_581 (O_581,N_14272,N_14123);
nand UO_582 (O_582,N_13582,N_14964);
or UO_583 (O_583,N_14257,N_14664);
nand UO_584 (O_584,N_13898,N_14726);
nand UO_585 (O_585,N_14640,N_14918);
or UO_586 (O_586,N_14529,N_14500);
and UO_587 (O_587,N_14356,N_13696);
and UO_588 (O_588,N_14236,N_14508);
or UO_589 (O_589,N_13668,N_14169);
nand UO_590 (O_590,N_13862,N_13918);
and UO_591 (O_591,N_14659,N_14345);
nand UO_592 (O_592,N_13557,N_13594);
nor UO_593 (O_593,N_14241,N_14251);
and UO_594 (O_594,N_14694,N_13855);
and UO_595 (O_595,N_14307,N_14970);
nor UO_596 (O_596,N_14165,N_13710);
nand UO_597 (O_597,N_14371,N_14578);
nor UO_598 (O_598,N_14595,N_14248);
nand UO_599 (O_599,N_13770,N_14465);
nand UO_600 (O_600,N_14113,N_13779);
and UO_601 (O_601,N_13796,N_13685);
or UO_602 (O_602,N_14761,N_14930);
and UO_603 (O_603,N_13566,N_13933);
and UO_604 (O_604,N_14614,N_14397);
or UO_605 (O_605,N_14631,N_13693);
and UO_606 (O_606,N_14027,N_14328);
and UO_607 (O_607,N_13729,N_14928);
or UO_608 (O_608,N_14287,N_13534);
and UO_609 (O_609,N_14115,N_14821);
nor UO_610 (O_610,N_14273,N_14717);
and UO_611 (O_611,N_14552,N_14106);
nor UO_612 (O_612,N_14373,N_13759);
and UO_613 (O_613,N_14832,N_13975);
nor UO_614 (O_614,N_14788,N_13541);
nand UO_615 (O_615,N_14996,N_14478);
nand UO_616 (O_616,N_14420,N_14572);
xor UO_617 (O_617,N_14729,N_13606);
and UO_618 (O_618,N_14551,N_14103);
and UO_619 (O_619,N_14767,N_14895);
nand UO_620 (O_620,N_13986,N_13705);
and UO_621 (O_621,N_14676,N_13628);
nand UO_622 (O_622,N_14350,N_14577);
nor UO_623 (O_623,N_13549,N_14000);
nor UO_624 (O_624,N_13562,N_13985);
nor UO_625 (O_625,N_14633,N_13788);
nand UO_626 (O_626,N_13854,N_14626);
nand UO_627 (O_627,N_14334,N_14491);
and UO_628 (O_628,N_14201,N_13724);
and UO_629 (O_629,N_13660,N_13946);
or UO_630 (O_630,N_14049,N_14768);
and UO_631 (O_631,N_14144,N_14818);
nand UO_632 (O_632,N_14597,N_14419);
and UO_633 (O_633,N_13801,N_14670);
and UO_634 (O_634,N_14269,N_13793);
or UO_635 (O_635,N_13598,N_13973);
or UO_636 (O_636,N_14602,N_14646);
and UO_637 (O_637,N_14014,N_13603);
and UO_638 (O_638,N_14886,N_13552);
and UO_639 (O_639,N_13792,N_13577);
nand UO_640 (O_640,N_14172,N_13785);
nor UO_641 (O_641,N_14249,N_14482);
and UO_642 (O_642,N_13895,N_14084);
nor UO_643 (O_643,N_13978,N_13526);
and UO_644 (O_644,N_13989,N_14627);
nand UO_645 (O_645,N_13543,N_14807);
nor UO_646 (O_646,N_14869,N_14329);
or UO_647 (O_647,N_14909,N_14912);
and UO_648 (O_648,N_14442,N_14095);
nor UO_649 (O_649,N_13690,N_14109);
and UO_650 (O_650,N_14369,N_14034);
nor UO_651 (O_651,N_13780,N_14698);
nand UO_652 (O_652,N_14777,N_13870);
nor UO_653 (O_653,N_13766,N_13664);
nand UO_654 (O_654,N_13995,N_14071);
nand UO_655 (O_655,N_14093,N_14300);
and UO_656 (O_656,N_13883,N_14576);
and UO_657 (O_657,N_13868,N_14925);
or UO_658 (O_658,N_14193,N_13704);
and UO_659 (O_659,N_13661,N_13754);
and UO_660 (O_660,N_13764,N_13931);
nor UO_661 (O_661,N_13814,N_14244);
nand UO_662 (O_662,N_14945,N_14384);
nor UO_663 (O_663,N_14372,N_14870);
and UO_664 (O_664,N_14056,N_14469);
and UO_665 (O_665,N_14364,N_14616);
and UO_666 (O_666,N_14319,N_14341);
and UO_667 (O_667,N_14453,N_14759);
xor UO_668 (O_668,N_13857,N_14981);
and UO_669 (O_669,N_13983,N_14238);
nor UO_670 (O_670,N_13782,N_13907);
and UO_671 (O_671,N_14503,N_14871);
or UO_672 (O_672,N_14834,N_13935);
and UO_673 (O_673,N_14098,N_14742);
nand UO_674 (O_674,N_14462,N_14778);
nand UO_675 (O_675,N_13981,N_14336);
nor UO_676 (O_676,N_14270,N_14496);
and UO_677 (O_677,N_14947,N_13501);
and UO_678 (O_678,N_14047,N_14985);
or UO_679 (O_679,N_13716,N_13866);
and UO_680 (O_680,N_14073,N_14008);
or UO_681 (O_681,N_14889,N_14032);
nor UO_682 (O_682,N_14140,N_14603);
nand UO_683 (O_683,N_14835,N_14016);
or UO_684 (O_684,N_14134,N_14374);
nor UO_685 (O_685,N_13848,N_14226);
nand UO_686 (O_686,N_14030,N_14466);
and UO_687 (O_687,N_14619,N_14814);
and UO_688 (O_688,N_14990,N_14517);
nand UO_689 (O_689,N_13938,N_14838);
and UO_690 (O_690,N_14441,N_13688);
xor UO_691 (O_691,N_14495,N_14953);
and UO_692 (O_692,N_14519,N_14522);
nor UO_693 (O_693,N_14585,N_14037);
or UO_694 (O_694,N_14708,N_14305);
nand UO_695 (O_695,N_14854,N_14398);
nand UO_696 (O_696,N_13970,N_14671);
xnor UO_697 (O_697,N_13642,N_14922);
and UO_698 (O_698,N_14523,N_14486);
or UO_699 (O_699,N_14806,N_14489);
nor UO_700 (O_700,N_13924,N_14266);
nand UO_701 (O_701,N_13999,N_14667);
nor UO_702 (O_702,N_13960,N_14747);
nand UO_703 (O_703,N_14274,N_14348);
or UO_704 (O_704,N_14790,N_14665);
or UO_705 (O_705,N_14968,N_14583);
or UO_706 (O_706,N_14862,N_13713);
nor UO_707 (O_707,N_13976,N_14068);
nor UO_708 (O_708,N_14050,N_14283);
and UO_709 (O_709,N_14359,N_14673);
or UO_710 (O_710,N_14333,N_14606);
or UO_711 (O_711,N_14146,N_14593);
nand UO_712 (O_712,N_14917,N_14762);
nor UO_713 (O_713,N_14823,N_14569);
or UO_714 (O_714,N_14723,N_14107);
nor UO_715 (O_715,N_14568,N_14426);
nor UO_716 (O_716,N_14327,N_13926);
nor UO_717 (O_717,N_14133,N_14852);
or UO_718 (O_718,N_13684,N_14567);
and UO_719 (O_719,N_13860,N_14908);
and UO_720 (O_720,N_13742,N_14915);
nand UO_721 (O_721,N_14658,N_13863);
and UO_722 (O_722,N_13813,N_13510);
nand UO_723 (O_723,N_13894,N_14501);
nand UO_724 (O_724,N_13669,N_13692);
and UO_725 (O_725,N_13720,N_14349);
nor UO_726 (O_726,N_14961,N_13787);
nor UO_727 (O_727,N_14232,N_14429);
and UO_728 (O_728,N_14081,N_14604);
nand UO_729 (O_729,N_13873,N_13944);
and UO_730 (O_730,N_13714,N_13771);
or UO_731 (O_731,N_14652,N_13514);
or UO_732 (O_732,N_14092,N_13560);
nor UO_733 (O_733,N_14853,N_13998);
or UO_734 (O_734,N_13817,N_14059);
nand UO_735 (O_735,N_14559,N_13752);
or UO_736 (O_736,N_13994,N_14505);
or UO_737 (O_737,N_13750,N_14129);
nand UO_738 (O_738,N_14159,N_14434);
nand UO_739 (O_739,N_13997,N_14954);
nor UO_740 (O_740,N_13605,N_14965);
and UO_741 (O_741,N_13591,N_14666);
and UO_742 (O_742,N_14379,N_14023);
nand UO_743 (O_743,N_14554,N_13731);
nand UO_744 (O_744,N_13889,N_13600);
and UO_745 (O_745,N_14173,N_14610);
nor UO_746 (O_746,N_14829,N_14125);
or UO_747 (O_747,N_14295,N_14727);
xor UO_748 (O_748,N_13517,N_14493);
nand UO_749 (O_749,N_14764,N_13615);
nor UO_750 (O_750,N_14187,N_14958);
nand UO_751 (O_751,N_14894,N_13675);
nor UO_752 (O_752,N_14888,N_14162);
nand UO_753 (O_753,N_13580,N_14211);
and UO_754 (O_754,N_14159,N_14496);
nor UO_755 (O_755,N_13576,N_13532);
nand UO_756 (O_756,N_13908,N_14046);
nor UO_757 (O_757,N_14789,N_14390);
nand UO_758 (O_758,N_14072,N_14043);
or UO_759 (O_759,N_14719,N_14101);
nand UO_760 (O_760,N_14242,N_13908);
nand UO_761 (O_761,N_14893,N_14116);
or UO_762 (O_762,N_13602,N_14989);
nand UO_763 (O_763,N_14047,N_14067);
nand UO_764 (O_764,N_14647,N_14845);
or UO_765 (O_765,N_13733,N_13543);
nand UO_766 (O_766,N_13816,N_13716);
nor UO_767 (O_767,N_14844,N_13833);
xnor UO_768 (O_768,N_14261,N_13729);
or UO_769 (O_769,N_14449,N_13675);
nor UO_770 (O_770,N_13985,N_14289);
nand UO_771 (O_771,N_13701,N_13942);
nand UO_772 (O_772,N_14845,N_13711);
nand UO_773 (O_773,N_14813,N_13997);
nand UO_774 (O_774,N_14093,N_14533);
nand UO_775 (O_775,N_14268,N_14067);
nor UO_776 (O_776,N_14738,N_13933);
or UO_777 (O_777,N_14211,N_13850);
nor UO_778 (O_778,N_14801,N_14325);
nand UO_779 (O_779,N_14376,N_14018);
xnor UO_780 (O_780,N_13864,N_14165);
or UO_781 (O_781,N_14756,N_13521);
and UO_782 (O_782,N_14951,N_14875);
or UO_783 (O_783,N_14538,N_14311);
nand UO_784 (O_784,N_13542,N_13781);
nor UO_785 (O_785,N_13821,N_14447);
nor UO_786 (O_786,N_13796,N_13769);
and UO_787 (O_787,N_13647,N_14735);
nor UO_788 (O_788,N_14979,N_14801);
or UO_789 (O_789,N_13987,N_14199);
nor UO_790 (O_790,N_13795,N_14735);
or UO_791 (O_791,N_14330,N_14386);
or UO_792 (O_792,N_14269,N_13547);
nand UO_793 (O_793,N_13824,N_14852);
nand UO_794 (O_794,N_14711,N_14502);
nand UO_795 (O_795,N_14043,N_13700);
or UO_796 (O_796,N_14153,N_14021);
and UO_797 (O_797,N_14634,N_14872);
nor UO_798 (O_798,N_13864,N_14804);
nor UO_799 (O_799,N_14287,N_14201);
nand UO_800 (O_800,N_14507,N_14722);
or UO_801 (O_801,N_14650,N_14531);
and UO_802 (O_802,N_13904,N_13749);
nand UO_803 (O_803,N_14435,N_13637);
and UO_804 (O_804,N_13662,N_13980);
and UO_805 (O_805,N_14212,N_14553);
nand UO_806 (O_806,N_14667,N_14036);
nor UO_807 (O_807,N_13708,N_14562);
or UO_808 (O_808,N_14153,N_13705);
or UO_809 (O_809,N_14500,N_14703);
and UO_810 (O_810,N_13595,N_14780);
nor UO_811 (O_811,N_14483,N_13614);
or UO_812 (O_812,N_14398,N_13767);
nor UO_813 (O_813,N_13748,N_13814);
nand UO_814 (O_814,N_14848,N_14961);
nand UO_815 (O_815,N_13765,N_13614);
nor UO_816 (O_816,N_13561,N_13903);
nor UO_817 (O_817,N_14876,N_14079);
nor UO_818 (O_818,N_14628,N_13921);
and UO_819 (O_819,N_14787,N_13949);
nand UO_820 (O_820,N_14476,N_14574);
and UO_821 (O_821,N_14992,N_13884);
and UO_822 (O_822,N_14878,N_14292);
or UO_823 (O_823,N_14556,N_13526);
nor UO_824 (O_824,N_14319,N_14812);
nor UO_825 (O_825,N_14607,N_14738);
nand UO_826 (O_826,N_14443,N_14963);
nand UO_827 (O_827,N_14236,N_14759);
nor UO_828 (O_828,N_13920,N_14796);
nor UO_829 (O_829,N_14689,N_14392);
or UO_830 (O_830,N_14729,N_13751);
and UO_831 (O_831,N_14418,N_14830);
or UO_832 (O_832,N_13731,N_13804);
nand UO_833 (O_833,N_14555,N_13552);
and UO_834 (O_834,N_14161,N_14093);
and UO_835 (O_835,N_14056,N_14675);
or UO_836 (O_836,N_14452,N_14672);
nand UO_837 (O_837,N_14216,N_13607);
or UO_838 (O_838,N_13714,N_14466);
or UO_839 (O_839,N_14408,N_13805);
nor UO_840 (O_840,N_14125,N_14928);
and UO_841 (O_841,N_14767,N_14405);
nand UO_842 (O_842,N_13546,N_13971);
nand UO_843 (O_843,N_13968,N_13881);
nor UO_844 (O_844,N_14938,N_13727);
or UO_845 (O_845,N_13731,N_14899);
and UO_846 (O_846,N_14047,N_14234);
nor UO_847 (O_847,N_14987,N_14798);
and UO_848 (O_848,N_14467,N_13963);
nor UO_849 (O_849,N_13722,N_13748);
nand UO_850 (O_850,N_14917,N_13975);
nand UO_851 (O_851,N_14514,N_14865);
nor UO_852 (O_852,N_13508,N_14623);
nor UO_853 (O_853,N_14827,N_14273);
or UO_854 (O_854,N_13932,N_13832);
nand UO_855 (O_855,N_13574,N_13680);
nor UO_856 (O_856,N_14292,N_13883);
or UO_857 (O_857,N_14944,N_14308);
nand UO_858 (O_858,N_14013,N_13993);
nor UO_859 (O_859,N_13638,N_14693);
and UO_860 (O_860,N_14202,N_13733);
nand UO_861 (O_861,N_13706,N_14158);
nand UO_862 (O_862,N_14187,N_14211);
xor UO_863 (O_863,N_14664,N_14638);
and UO_864 (O_864,N_13601,N_14240);
or UO_865 (O_865,N_14523,N_14311);
or UO_866 (O_866,N_14835,N_14852);
or UO_867 (O_867,N_14984,N_13980);
nor UO_868 (O_868,N_14377,N_13652);
nand UO_869 (O_869,N_14287,N_14610);
and UO_870 (O_870,N_14709,N_14027);
nor UO_871 (O_871,N_14103,N_14559);
or UO_872 (O_872,N_14531,N_13749);
nand UO_873 (O_873,N_14631,N_14090);
or UO_874 (O_874,N_13942,N_14952);
nor UO_875 (O_875,N_14007,N_14784);
and UO_876 (O_876,N_14292,N_14278);
and UO_877 (O_877,N_13638,N_14208);
nand UO_878 (O_878,N_14675,N_13902);
and UO_879 (O_879,N_14747,N_14842);
and UO_880 (O_880,N_14915,N_14217);
or UO_881 (O_881,N_13610,N_14423);
nor UO_882 (O_882,N_14894,N_13568);
and UO_883 (O_883,N_13648,N_13722);
or UO_884 (O_884,N_13657,N_14711);
or UO_885 (O_885,N_14342,N_14157);
nor UO_886 (O_886,N_14610,N_14911);
nor UO_887 (O_887,N_13864,N_14915);
and UO_888 (O_888,N_13980,N_14760);
or UO_889 (O_889,N_14712,N_14640);
nor UO_890 (O_890,N_14708,N_14599);
or UO_891 (O_891,N_14161,N_13901);
nand UO_892 (O_892,N_13619,N_13710);
or UO_893 (O_893,N_14649,N_13517);
or UO_894 (O_894,N_14847,N_13689);
or UO_895 (O_895,N_14593,N_14452);
or UO_896 (O_896,N_14825,N_14183);
nor UO_897 (O_897,N_13709,N_14496);
and UO_898 (O_898,N_13904,N_14406);
nor UO_899 (O_899,N_14651,N_14864);
or UO_900 (O_900,N_14323,N_14191);
nand UO_901 (O_901,N_14980,N_14514);
or UO_902 (O_902,N_13769,N_14764);
and UO_903 (O_903,N_14183,N_14585);
or UO_904 (O_904,N_13563,N_14672);
nand UO_905 (O_905,N_14586,N_14138);
nand UO_906 (O_906,N_13816,N_13513);
nand UO_907 (O_907,N_14791,N_13589);
nand UO_908 (O_908,N_13596,N_13866);
and UO_909 (O_909,N_14338,N_14591);
xor UO_910 (O_910,N_13983,N_13863);
nand UO_911 (O_911,N_14057,N_13850);
or UO_912 (O_912,N_14648,N_13980);
or UO_913 (O_913,N_13662,N_14389);
nand UO_914 (O_914,N_14734,N_14648);
nand UO_915 (O_915,N_14496,N_14303);
nor UO_916 (O_916,N_14121,N_14398);
nor UO_917 (O_917,N_14533,N_13571);
or UO_918 (O_918,N_14009,N_14633);
nand UO_919 (O_919,N_13871,N_14736);
and UO_920 (O_920,N_14490,N_13695);
nand UO_921 (O_921,N_14760,N_13618);
and UO_922 (O_922,N_14233,N_14382);
nor UO_923 (O_923,N_14078,N_14886);
nand UO_924 (O_924,N_13789,N_13812);
or UO_925 (O_925,N_14710,N_14273);
and UO_926 (O_926,N_14968,N_14476);
nor UO_927 (O_927,N_13804,N_13675);
nand UO_928 (O_928,N_13986,N_14859);
xnor UO_929 (O_929,N_13975,N_13586);
nor UO_930 (O_930,N_14654,N_14430);
and UO_931 (O_931,N_14778,N_13571);
nor UO_932 (O_932,N_14818,N_13702);
nand UO_933 (O_933,N_14231,N_14544);
and UO_934 (O_934,N_14540,N_14276);
nor UO_935 (O_935,N_14753,N_13805);
nor UO_936 (O_936,N_13919,N_14732);
or UO_937 (O_937,N_14271,N_13674);
and UO_938 (O_938,N_14522,N_13708);
xnor UO_939 (O_939,N_14801,N_13508);
or UO_940 (O_940,N_13781,N_14546);
nor UO_941 (O_941,N_14098,N_13541);
nand UO_942 (O_942,N_13884,N_13716);
and UO_943 (O_943,N_14043,N_14373);
or UO_944 (O_944,N_13993,N_13707);
nand UO_945 (O_945,N_14550,N_13564);
nor UO_946 (O_946,N_13778,N_14264);
or UO_947 (O_947,N_13863,N_13754);
and UO_948 (O_948,N_13942,N_13869);
and UO_949 (O_949,N_14733,N_14651);
nor UO_950 (O_950,N_14338,N_14037);
or UO_951 (O_951,N_13702,N_13961);
xor UO_952 (O_952,N_14655,N_14578);
or UO_953 (O_953,N_14363,N_14669);
or UO_954 (O_954,N_14325,N_14465);
nand UO_955 (O_955,N_13562,N_14053);
nor UO_956 (O_956,N_13903,N_14558);
nor UO_957 (O_957,N_14752,N_13608);
and UO_958 (O_958,N_14216,N_14796);
or UO_959 (O_959,N_14235,N_13828);
nor UO_960 (O_960,N_13901,N_13998);
or UO_961 (O_961,N_13638,N_14209);
or UO_962 (O_962,N_14789,N_14886);
or UO_963 (O_963,N_13908,N_14345);
and UO_964 (O_964,N_14697,N_13859);
nor UO_965 (O_965,N_14925,N_14320);
nor UO_966 (O_966,N_13954,N_14538);
nor UO_967 (O_967,N_13632,N_14824);
or UO_968 (O_968,N_13576,N_14299);
nand UO_969 (O_969,N_13678,N_13791);
or UO_970 (O_970,N_14110,N_14758);
and UO_971 (O_971,N_13831,N_14456);
xor UO_972 (O_972,N_14202,N_14634);
or UO_973 (O_973,N_14534,N_14878);
or UO_974 (O_974,N_14539,N_14729);
nand UO_975 (O_975,N_13787,N_13893);
and UO_976 (O_976,N_13866,N_13877);
or UO_977 (O_977,N_13768,N_13932);
and UO_978 (O_978,N_14106,N_13601);
and UO_979 (O_979,N_13621,N_14882);
and UO_980 (O_980,N_14924,N_14656);
nor UO_981 (O_981,N_13519,N_14328);
or UO_982 (O_982,N_14349,N_13903);
or UO_983 (O_983,N_13619,N_13624);
and UO_984 (O_984,N_14589,N_14168);
or UO_985 (O_985,N_14491,N_14379);
or UO_986 (O_986,N_14295,N_14524);
or UO_987 (O_987,N_14271,N_14806);
nor UO_988 (O_988,N_14576,N_14558);
or UO_989 (O_989,N_14667,N_14207);
nor UO_990 (O_990,N_13862,N_13767);
nor UO_991 (O_991,N_13948,N_14598);
and UO_992 (O_992,N_14765,N_13862);
nor UO_993 (O_993,N_13775,N_14496);
and UO_994 (O_994,N_13543,N_14345);
or UO_995 (O_995,N_14970,N_14781);
nand UO_996 (O_996,N_13770,N_13736);
xnor UO_997 (O_997,N_14580,N_14138);
nor UO_998 (O_998,N_14366,N_14978);
or UO_999 (O_999,N_13974,N_13971);
or UO_1000 (O_1000,N_14740,N_14120);
nand UO_1001 (O_1001,N_14765,N_13774);
or UO_1002 (O_1002,N_13868,N_13562);
nand UO_1003 (O_1003,N_14016,N_13920);
or UO_1004 (O_1004,N_14797,N_14007);
and UO_1005 (O_1005,N_13669,N_13816);
and UO_1006 (O_1006,N_14632,N_13586);
nor UO_1007 (O_1007,N_14421,N_14533);
nand UO_1008 (O_1008,N_14845,N_13520);
and UO_1009 (O_1009,N_14310,N_14081);
nor UO_1010 (O_1010,N_14209,N_14822);
nand UO_1011 (O_1011,N_14552,N_13853);
nand UO_1012 (O_1012,N_13522,N_14891);
nand UO_1013 (O_1013,N_14269,N_14158);
and UO_1014 (O_1014,N_14345,N_14978);
xnor UO_1015 (O_1015,N_14690,N_14705);
nor UO_1016 (O_1016,N_14008,N_14595);
nand UO_1017 (O_1017,N_14658,N_14064);
and UO_1018 (O_1018,N_14456,N_13548);
and UO_1019 (O_1019,N_14121,N_14963);
nor UO_1020 (O_1020,N_13649,N_13787);
or UO_1021 (O_1021,N_13613,N_14441);
nand UO_1022 (O_1022,N_14647,N_13764);
and UO_1023 (O_1023,N_13643,N_14656);
or UO_1024 (O_1024,N_14790,N_14496);
nand UO_1025 (O_1025,N_13591,N_14344);
nand UO_1026 (O_1026,N_14374,N_13573);
nand UO_1027 (O_1027,N_14391,N_14693);
and UO_1028 (O_1028,N_13786,N_14783);
nand UO_1029 (O_1029,N_14381,N_14237);
nor UO_1030 (O_1030,N_14412,N_13791);
nor UO_1031 (O_1031,N_14237,N_14744);
or UO_1032 (O_1032,N_14150,N_13976);
nand UO_1033 (O_1033,N_14461,N_14362);
nor UO_1034 (O_1034,N_14121,N_13863);
nand UO_1035 (O_1035,N_14353,N_14839);
and UO_1036 (O_1036,N_14041,N_14813);
nor UO_1037 (O_1037,N_13530,N_14884);
or UO_1038 (O_1038,N_14950,N_14218);
or UO_1039 (O_1039,N_14897,N_14548);
nor UO_1040 (O_1040,N_14162,N_13511);
nor UO_1041 (O_1041,N_14268,N_13596);
or UO_1042 (O_1042,N_14321,N_14715);
and UO_1043 (O_1043,N_13632,N_14441);
nand UO_1044 (O_1044,N_14771,N_13519);
or UO_1045 (O_1045,N_14542,N_13639);
or UO_1046 (O_1046,N_14651,N_13846);
nand UO_1047 (O_1047,N_14008,N_14789);
nor UO_1048 (O_1048,N_13558,N_13973);
xor UO_1049 (O_1049,N_14733,N_14167);
nand UO_1050 (O_1050,N_13554,N_13800);
nor UO_1051 (O_1051,N_13944,N_14114);
and UO_1052 (O_1052,N_14492,N_14272);
nor UO_1053 (O_1053,N_13539,N_13749);
nand UO_1054 (O_1054,N_14456,N_14776);
nand UO_1055 (O_1055,N_14773,N_13597);
or UO_1056 (O_1056,N_14542,N_14270);
and UO_1057 (O_1057,N_14084,N_14993);
nand UO_1058 (O_1058,N_14456,N_14035);
nor UO_1059 (O_1059,N_14334,N_13500);
nor UO_1060 (O_1060,N_14877,N_13717);
nor UO_1061 (O_1061,N_13934,N_14367);
nor UO_1062 (O_1062,N_13500,N_14268);
and UO_1063 (O_1063,N_14198,N_14574);
or UO_1064 (O_1064,N_14554,N_13691);
or UO_1065 (O_1065,N_14377,N_13600);
nand UO_1066 (O_1066,N_14343,N_14136);
and UO_1067 (O_1067,N_14971,N_14699);
nor UO_1068 (O_1068,N_14468,N_13509);
nor UO_1069 (O_1069,N_14135,N_14007);
and UO_1070 (O_1070,N_13888,N_14258);
or UO_1071 (O_1071,N_14529,N_14870);
nand UO_1072 (O_1072,N_14874,N_14867);
nand UO_1073 (O_1073,N_13505,N_14252);
xnor UO_1074 (O_1074,N_14966,N_13728);
and UO_1075 (O_1075,N_13642,N_13619);
and UO_1076 (O_1076,N_14548,N_14641);
nand UO_1077 (O_1077,N_13944,N_14736);
and UO_1078 (O_1078,N_13739,N_14573);
nor UO_1079 (O_1079,N_14597,N_13731);
nor UO_1080 (O_1080,N_14530,N_13759);
and UO_1081 (O_1081,N_14701,N_14187);
nor UO_1082 (O_1082,N_14964,N_13519);
nor UO_1083 (O_1083,N_14453,N_14833);
xnor UO_1084 (O_1084,N_14907,N_13579);
nor UO_1085 (O_1085,N_14220,N_14012);
nor UO_1086 (O_1086,N_13596,N_13742);
xnor UO_1087 (O_1087,N_13859,N_13630);
nand UO_1088 (O_1088,N_14214,N_14013);
or UO_1089 (O_1089,N_14923,N_13504);
nand UO_1090 (O_1090,N_13902,N_14578);
and UO_1091 (O_1091,N_14940,N_14772);
or UO_1092 (O_1092,N_14451,N_14390);
and UO_1093 (O_1093,N_14299,N_14774);
and UO_1094 (O_1094,N_14246,N_14036);
and UO_1095 (O_1095,N_14247,N_14145);
and UO_1096 (O_1096,N_13948,N_14696);
nand UO_1097 (O_1097,N_14480,N_14976);
and UO_1098 (O_1098,N_13725,N_14123);
or UO_1099 (O_1099,N_13571,N_14408);
nor UO_1100 (O_1100,N_14976,N_14587);
nor UO_1101 (O_1101,N_14843,N_14144);
and UO_1102 (O_1102,N_14755,N_14330);
nor UO_1103 (O_1103,N_14856,N_13505);
or UO_1104 (O_1104,N_13926,N_14133);
nand UO_1105 (O_1105,N_13519,N_14998);
nand UO_1106 (O_1106,N_14407,N_14561);
xor UO_1107 (O_1107,N_14429,N_13672);
or UO_1108 (O_1108,N_14486,N_14146);
nor UO_1109 (O_1109,N_14394,N_14252);
nand UO_1110 (O_1110,N_13846,N_13781);
or UO_1111 (O_1111,N_14958,N_14220);
nand UO_1112 (O_1112,N_14259,N_14485);
nor UO_1113 (O_1113,N_13837,N_14408);
nor UO_1114 (O_1114,N_14208,N_14284);
nand UO_1115 (O_1115,N_14755,N_13648);
nand UO_1116 (O_1116,N_14169,N_13716);
or UO_1117 (O_1117,N_14109,N_13755);
and UO_1118 (O_1118,N_13774,N_13530);
nand UO_1119 (O_1119,N_14400,N_14457);
nand UO_1120 (O_1120,N_14758,N_14018);
and UO_1121 (O_1121,N_14694,N_13923);
and UO_1122 (O_1122,N_14247,N_14052);
nand UO_1123 (O_1123,N_13816,N_14861);
and UO_1124 (O_1124,N_14237,N_13789);
nor UO_1125 (O_1125,N_14924,N_14753);
nand UO_1126 (O_1126,N_14007,N_14816);
or UO_1127 (O_1127,N_14086,N_14446);
and UO_1128 (O_1128,N_14852,N_14152);
and UO_1129 (O_1129,N_14683,N_14576);
nand UO_1130 (O_1130,N_13856,N_13919);
or UO_1131 (O_1131,N_13903,N_14013);
xnor UO_1132 (O_1132,N_14233,N_14212);
and UO_1133 (O_1133,N_14468,N_13515);
or UO_1134 (O_1134,N_14506,N_14392);
and UO_1135 (O_1135,N_14228,N_14195);
or UO_1136 (O_1136,N_14972,N_13578);
and UO_1137 (O_1137,N_14318,N_14628);
xor UO_1138 (O_1138,N_14274,N_13792);
and UO_1139 (O_1139,N_13608,N_14075);
nor UO_1140 (O_1140,N_14854,N_14001);
nor UO_1141 (O_1141,N_14728,N_13826);
and UO_1142 (O_1142,N_14558,N_14908);
nand UO_1143 (O_1143,N_13887,N_14733);
nor UO_1144 (O_1144,N_14611,N_14890);
nand UO_1145 (O_1145,N_14450,N_14623);
and UO_1146 (O_1146,N_14568,N_13568);
nand UO_1147 (O_1147,N_14642,N_14046);
and UO_1148 (O_1148,N_14572,N_13752);
nor UO_1149 (O_1149,N_14034,N_14103);
nand UO_1150 (O_1150,N_14171,N_13761);
or UO_1151 (O_1151,N_14181,N_14624);
nand UO_1152 (O_1152,N_14654,N_13941);
nor UO_1153 (O_1153,N_14729,N_14001);
nand UO_1154 (O_1154,N_14022,N_14547);
nand UO_1155 (O_1155,N_14718,N_14333);
or UO_1156 (O_1156,N_14458,N_14829);
or UO_1157 (O_1157,N_14894,N_13983);
nor UO_1158 (O_1158,N_14642,N_14520);
and UO_1159 (O_1159,N_14295,N_14541);
nor UO_1160 (O_1160,N_14577,N_13811);
nor UO_1161 (O_1161,N_13634,N_13513);
nand UO_1162 (O_1162,N_14418,N_14045);
or UO_1163 (O_1163,N_13632,N_13538);
nand UO_1164 (O_1164,N_14230,N_14033);
or UO_1165 (O_1165,N_14902,N_14967);
or UO_1166 (O_1166,N_14459,N_13681);
nor UO_1167 (O_1167,N_13750,N_14591);
and UO_1168 (O_1168,N_13735,N_14004);
nor UO_1169 (O_1169,N_14151,N_14829);
nand UO_1170 (O_1170,N_14627,N_14273);
nor UO_1171 (O_1171,N_13742,N_13533);
nor UO_1172 (O_1172,N_13950,N_13563);
nand UO_1173 (O_1173,N_14792,N_13950);
or UO_1174 (O_1174,N_14743,N_14513);
or UO_1175 (O_1175,N_14170,N_13895);
nor UO_1176 (O_1176,N_13516,N_14695);
or UO_1177 (O_1177,N_14232,N_14070);
nand UO_1178 (O_1178,N_13790,N_14874);
nor UO_1179 (O_1179,N_14893,N_14078);
nor UO_1180 (O_1180,N_13701,N_13704);
or UO_1181 (O_1181,N_14313,N_14200);
nand UO_1182 (O_1182,N_14235,N_13681);
and UO_1183 (O_1183,N_14824,N_14816);
nand UO_1184 (O_1184,N_13815,N_14506);
and UO_1185 (O_1185,N_14179,N_14381);
and UO_1186 (O_1186,N_13668,N_14041);
nor UO_1187 (O_1187,N_14654,N_14699);
xor UO_1188 (O_1188,N_14174,N_14310);
or UO_1189 (O_1189,N_14453,N_13908);
nor UO_1190 (O_1190,N_14415,N_14339);
or UO_1191 (O_1191,N_13572,N_14001);
nor UO_1192 (O_1192,N_14516,N_14386);
nand UO_1193 (O_1193,N_14931,N_13628);
nor UO_1194 (O_1194,N_14695,N_14525);
xnor UO_1195 (O_1195,N_13808,N_14446);
xor UO_1196 (O_1196,N_13620,N_14881);
nor UO_1197 (O_1197,N_14536,N_14178);
nand UO_1198 (O_1198,N_14809,N_13523);
nor UO_1199 (O_1199,N_14852,N_14606);
and UO_1200 (O_1200,N_13775,N_14561);
or UO_1201 (O_1201,N_14684,N_14060);
nor UO_1202 (O_1202,N_13937,N_13920);
nor UO_1203 (O_1203,N_13699,N_14589);
or UO_1204 (O_1204,N_14600,N_13961);
nor UO_1205 (O_1205,N_14293,N_13514);
and UO_1206 (O_1206,N_13986,N_14098);
nor UO_1207 (O_1207,N_14423,N_14748);
nor UO_1208 (O_1208,N_14015,N_14068);
or UO_1209 (O_1209,N_13672,N_13841);
and UO_1210 (O_1210,N_14172,N_14354);
nor UO_1211 (O_1211,N_14441,N_14784);
and UO_1212 (O_1212,N_13761,N_13865);
nor UO_1213 (O_1213,N_14685,N_13942);
nand UO_1214 (O_1214,N_14216,N_13588);
or UO_1215 (O_1215,N_13879,N_14253);
nor UO_1216 (O_1216,N_14468,N_13592);
nand UO_1217 (O_1217,N_14866,N_14647);
nor UO_1218 (O_1218,N_14395,N_14216);
nand UO_1219 (O_1219,N_14599,N_14913);
nor UO_1220 (O_1220,N_14623,N_14910);
nor UO_1221 (O_1221,N_13932,N_13781);
nor UO_1222 (O_1222,N_14005,N_13994);
or UO_1223 (O_1223,N_13785,N_14260);
or UO_1224 (O_1224,N_13660,N_13829);
nor UO_1225 (O_1225,N_14227,N_14866);
nor UO_1226 (O_1226,N_13869,N_13797);
nand UO_1227 (O_1227,N_14298,N_14731);
and UO_1228 (O_1228,N_13566,N_13676);
nor UO_1229 (O_1229,N_14570,N_14668);
or UO_1230 (O_1230,N_13725,N_14088);
nor UO_1231 (O_1231,N_14571,N_14337);
or UO_1232 (O_1232,N_14527,N_14721);
nand UO_1233 (O_1233,N_14838,N_14936);
and UO_1234 (O_1234,N_14474,N_14100);
or UO_1235 (O_1235,N_13616,N_13857);
or UO_1236 (O_1236,N_14843,N_14342);
xor UO_1237 (O_1237,N_14832,N_14631);
nor UO_1238 (O_1238,N_14319,N_14971);
xor UO_1239 (O_1239,N_13613,N_14608);
or UO_1240 (O_1240,N_14980,N_14307);
nor UO_1241 (O_1241,N_13731,N_14151);
or UO_1242 (O_1242,N_14288,N_14904);
nand UO_1243 (O_1243,N_13937,N_14603);
nand UO_1244 (O_1244,N_14833,N_13758);
nand UO_1245 (O_1245,N_14282,N_13862);
nand UO_1246 (O_1246,N_14065,N_14304);
nand UO_1247 (O_1247,N_13966,N_14188);
and UO_1248 (O_1248,N_14811,N_14481);
or UO_1249 (O_1249,N_14713,N_14704);
and UO_1250 (O_1250,N_13501,N_13559);
or UO_1251 (O_1251,N_14460,N_13737);
nand UO_1252 (O_1252,N_13897,N_14274);
or UO_1253 (O_1253,N_13736,N_14094);
or UO_1254 (O_1254,N_14711,N_13777);
nand UO_1255 (O_1255,N_13888,N_14397);
and UO_1256 (O_1256,N_14775,N_13980);
or UO_1257 (O_1257,N_14969,N_13770);
and UO_1258 (O_1258,N_14353,N_13514);
and UO_1259 (O_1259,N_13758,N_14638);
nand UO_1260 (O_1260,N_14512,N_13706);
nand UO_1261 (O_1261,N_14887,N_14779);
or UO_1262 (O_1262,N_13508,N_13916);
and UO_1263 (O_1263,N_14799,N_13935);
and UO_1264 (O_1264,N_13726,N_14575);
nor UO_1265 (O_1265,N_14431,N_14271);
or UO_1266 (O_1266,N_14166,N_14540);
or UO_1267 (O_1267,N_14877,N_13909);
and UO_1268 (O_1268,N_14085,N_14697);
xor UO_1269 (O_1269,N_14959,N_13855);
or UO_1270 (O_1270,N_13552,N_14465);
nor UO_1271 (O_1271,N_13776,N_14260);
nand UO_1272 (O_1272,N_14562,N_14016);
and UO_1273 (O_1273,N_14403,N_14459);
or UO_1274 (O_1274,N_14635,N_14082);
and UO_1275 (O_1275,N_14003,N_14609);
and UO_1276 (O_1276,N_13955,N_14387);
or UO_1277 (O_1277,N_13898,N_14975);
nand UO_1278 (O_1278,N_14304,N_14393);
and UO_1279 (O_1279,N_14723,N_14637);
or UO_1280 (O_1280,N_13935,N_14906);
nor UO_1281 (O_1281,N_14367,N_13512);
nor UO_1282 (O_1282,N_13891,N_14208);
and UO_1283 (O_1283,N_14292,N_13643);
or UO_1284 (O_1284,N_13761,N_14901);
or UO_1285 (O_1285,N_13590,N_14896);
and UO_1286 (O_1286,N_14691,N_14446);
or UO_1287 (O_1287,N_13696,N_14295);
nor UO_1288 (O_1288,N_13987,N_13877);
and UO_1289 (O_1289,N_13820,N_14708);
and UO_1290 (O_1290,N_13999,N_13929);
or UO_1291 (O_1291,N_13913,N_14555);
nor UO_1292 (O_1292,N_14515,N_13823);
nand UO_1293 (O_1293,N_13751,N_14163);
or UO_1294 (O_1294,N_13843,N_13766);
nor UO_1295 (O_1295,N_14400,N_14653);
and UO_1296 (O_1296,N_14479,N_14595);
xor UO_1297 (O_1297,N_14977,N_13974);
nand UO_1298 (O_1298,N_14865,N_13977);
and UO_1299 (O_1299,N_14653,N_13985);
or UO_1300 (O_1300,N_13932,N_13589);
and UO_1301 (O_1301,N_14151,N_14056);
or UO_1302 (O_1302,N_14820,N_14834);
or UO_1303 (O_1303,N_13957,N_13721);
nand UO_1304 (O_1304,N_13577,N_14348);
or UO_1305 (O_1305,N_14380,N_14313);
nand UO_1306 (O_1306,N_13550,N_14007);
and UO_1307 (O_1307,N_14479,N_14145);
or UO_1308 (O_1308,N_13801,N_14236);
nor UO_1309 (O_1309,N_13768,N_14171);
or UO_1310 (O_1310,N_14810,N_14627);
and UO_1311 (O_1311,N_14747,N_14185);
or UO_1312 (O_1312,N_14806,N_13827);
and UO_1313 (O_1313,N_13604,N_14101);
nand UO_1314 (O_1314,N_14051,N_14923);
or UO_1315 (O_1315,N_14932,N_14416);
and UO_1316 (O_1316,N_13894,N_13790);
or UO_1317 (O_1317,N_14698,N_13569);
nor UO_1318 (O_1318,N_14012,N_14402);
xnor UO_1319 (O_1319,N_14699,N_13959);
nand UO_1320 (O_1320,N_13565,N_13723);
or UO_1321 (O_1321,N_13923,N_14126);
or UO_1322 (O_1322,N_14592,N_14827);
and UO_1323 (O_1323,N_13740,N_14924);
or UO_1324 (O_1324,N_14835,N_14073);
nor UO_1325 (O_1325,N_14999,N_14761);
nand UO_1326 (O_1326,N_13749,N_14783);
nor UO_1327 (O_1327,N_14770,N_14518);
and UO_1328 (O_1328,N_13895,N_14554);
xor UO_1329 (O_1329,N_14088,N_14241);
or UO_1330 (O_1330,N_13520,N_14644);
or UO_1331 (O_1331,N_14811,N_13828);
nor UO_1332 (O_1332,N_13616,N_14061);
nor UO_1333 (O_1333,N_14421,N_14777);
nand UO_1334 (O_1334,N_14757,N_14002);
and UO_1335 (O_1335,N_13935,N_14932);
nor UO_1336 (O_1336,N_14578,N_14992);
nor UO_1337 (O_1337,N_13795,N_14715);
nand UO_1338 (O_1338,N_14706,N_14456);
and UO_1339 (O_1339,N_14054,N_13787);
and UO_1340 (O_1340,N_14548,N_14145);
xor UO_1341 (O_1341,N_14878,N_14102);
nor UO_1342 (O_1342,N_13509,N_14880);
or UO_1343 (O_1343,N_14593,N_13500);
nand UO_1344 (O_1344,N_13811,N_14033);
and UO_1345 (O_1345,N_14748,N_14269);
nand UO_1346 (O_1346,N_14486,N_14302);
and UO_1347 (O_1347,N_14582,N_14364);
nand UO_1348 (O_1348,N_13786,N_13964);
nor UO_1349 (O_1349,N_14338,N_14085);
or UO_1350 (O_1350,N_14822,N_14668);
or UO_1351 (O_1351,N_14774,N_14868);
nor UO_1352 (O_1352,N_14788,N_14284);
nand UO_1353 (O_1353,N_14185,N_13801);
and UO_1354 (O_1354,N_14522,N_14009);
or UO_1355 (O_1355,N_14470,N_14659);
nor UO_1356 (O_1356,N_13847,N_14032);
and UO_1357 (O_1357,N_14456,N_13785);
or UO_1358 (O_1358,N_14814,N_14189);
nor UO_1359 (O_1359,N_13657,N_13663);
and UO_1360 (O_1360,N_13658,N_13735);
nand UO_1361 (O_1361,N_14280,N_14920);
nand UO_1362 (O_1362,N_13900,N_14552);
and UO_1363 (O_1363,N_14112,N_14657);
nor UO_1364 (O_1364,N_13932,N_13971);
or UO_1365 (O_1365,N_13714,N_13614);
and UO_1366 (O_1366,N_14831,N_14573);
nand UO_1367 (O_1367,N_14327,N_14725);
nand UO_1368 (O_1368,N_14367,N_14445);
or UO_1369 (O_1369,N_13612,N_14511);
and UO_1370 (O_1370,N_14271,N_14228);
and UO_1371 (O_1371,N_14163,N_13870);
nand UO_1372 (O_1372,N_14813,N_14534);
or UO_1373 (O_1373,N_14616,N_14151);
nor UO_1374 (O_1374,N_14100,N_14265);
or UO_1375 (O_1375,N_14482,N_13688);
nand UO_1376 (O_1376,N_14020,N_14398);
nand UO_1377 (O_1377,N_14173,N_14282);
or UO_1378 (O_1378,N_14485,N_14217);
nand UO_1379 (O_1379,N_13509,N_14021);
or UO_1380 (O_1380,N_14558,N_14095);
xor UO_1381 (O_1381,N_14344,N_13783);
nand UO_1382 (O_1382,N_14830,N_13775);
nand UO_1383 (O_1383,N_13669,N_14224);
or UO_1384 (O_1384,N_13560,N_14813);
and UO_1385 (O_1385,N_14560,N_14983);
and UO_1386 (O_1386,N_13734,N_13983);
nor UO_1387 (O_1387,N_14482,N_13710);
or UO_1388 (O_1388,N_14336,N_14189);
and UO_1389 (O_1389,N_13932,N_14619);
nor UO_1390 (O_1390,N_14762,N_13721);
or UO_1391 (O_1391,N_13781,N_13985);
nor UO_1392 (O_1392,N_14467,N_14105);
or UO_1393 (O_1393,N_13766,N_14604);
nor UO_1394 (O_1394,N_14086,N_14921);
xnor UO_1395 (O_1395,N_14856,N_14158);
xnor UO_1396 (O_1396,N_14333,N_14310);
xor UO_1397 (O_1397,N_14779,N_14985);
nor UO_1398 (O_1398,N_14390,N_14201);
or UO_1399 (O_1399,N_14381,N_13990);
or UO_1400 (O_1400,N_14787,N_14618);
and UO_1401 (O_1401,N_14575,N_14742);
nor UO_1402 (O_1402,N_14452,N_14285);
nor UO_1403 (O_1403,N_14895,N_14804);
nand UO_1404 (O_1404,N_14271,N_13931);
nor UO_1405 (O_1405,N_14732,N_13918);
or UO_1406 (O_1406,N_13806,N_13805);
and UO_1407 (O_1407,N_14083,N_14542);
nand UO_1408 (O_1408,N_13552,N_14476);
or UO_1409 (O_1409,N_14885,N_14368);
and UO_1410 (O_1410,N_14674,N_13876);
nand UO_1411 (O_1411,N_13696,N_14224);
or UO_1412 (O_1412,N_14434,N_14077);
or UO_1413 (O_1413,N_14314,N_14026);
and UO_1414 (O_1414,N_13862,N_13810);
or UO_1415 (O_1415,N_14301,N_14651);
nand UO_1416 (O_1416,N_13918,N_13908);
and UO_1417 (O_1417,N_14943,N_14714);
and UO_1418 (O_1418,N_14301,N_13945);
and UO_1419 (O_1419,N_14013,N_14193);
or UO_1420 (O_1420,N_14252,N_14563);
nand UO_1421 (O_1421,N_14544,N_14391);
nand UO_1422 (O_1422,N_13641,N_14437);
or UO_1423 (O_1423,N_13976,N_13521);
and UO_1424 (O_1424,N_14306,N_13737);
and UO_1425 (O_1425,N_14473,N_13916);
and UO_1426 (O_1426,N_14239,N_14002);
nor UO_1427 (O_1427,N_14677,N_13532);
nor UO_1428 (O_1428,N_14075,N_14490);
or UO_1429 (O_1429,N_13561,N_14425);
nand UO_1430 (O_1430,N_14656,N_14520);
and UO_1431 (O_1431,N_14286,N_14645);
and UO_1432 (O_1432,N_14390,N_13739);
or UO_1433 (O_1433,N_14825,N_14597);
or UO_1434 (O_1434,N_14110,N_14685);
nand UO_1435 (O_1435,N_14961,N_13734);
and UO_1436 (O_1436,N_14289,N_14408);
or UO_1437 (O_1437,N_14338,N_14379);
xnor UO_1438 (O_1438,N_13941,N_13709);
nor UO_1439 (O_1439,N_14793,N_14170);
and UO_1440 (O_1440,N_14614,N_14723);
nand UO_1441 (O_1441,N_13957,N_14747);
and UO_1442 (O_1442,N_14462,N_14148);
or UO_1443 (O_1443,N_13839,N_14556);
nand UO_1444 (O_1444,N_14441,N_14003);
or UO_1445 (O_1445,N_14180,N_14029);
nand UO_1446 (O_1446,N_14918,N_14190);
or UO_1447 (O_1447,N_14256,N_14539);
xor UO_1448 (O_1448,N_13813,N_13931);
nor UO_1449 (O_1449,N_14346,N_14001);
nand UO_1450 (O_1450,N_14391,N_14321);
and UO_1451 (O_1451,N_14610,N_13941);
xnor UO_1452 (O_1452,N_13709,N_13613);
nand UO_1453 (O_1453,N_13909,N_14082);
and UO_1454 (O_1454,N_13744,N_13877);
and UO_1455 (O_1455,N_14745,N_14841);
nor UO_1456 (O_1456,N_14259,N_14865);
or UO_1457 (O_1457,N_13726,N_13961);
or UO_1458 (O_1458,N_14773,N_14088);
xnor UO_1459 (O_1459,N_14495,N_14540);
nand UO_1460 (O_1460,N_13666,N_13985);
nand UO_1461 (O_1461,N_14827,N_14112);
nand UO_1462 (O_1462,N_14232,N_14318);
nand UO_1463 (O_1463,N_14724,N_13686);
nand UO_1464 (O_1464,N_13937,N_14120);
and UO_1465 (O_1465,N_13651,N_14859);
or UO_1466 (O_1466,N_13933,N_14682);
nor UO_1467 (O_1467,N_14521,N_14662);
nand UO_1468 (O_1468,N_13979,N_14267);
and UO_1469 (O_1469,N_13732,N_13867);
nor UO_1470 (O_1470,N_14786,N_14489);
nor UO_1471 (O_1471,N_13879,N_14769);
nor UO_1472 (O_1472,N_13562,N_14796);
and UO_1473 (O_1473,N_14771,N_14296);
nor UO_1474 (O_1474,N_14471,N_14356);
and UO_1475 (O_1475,N_13997,N_14987);
or UO_1476 (O_1476,N_14585,N_14576);
xnor UO_1477 (O_1477,N_13930,N_14653);
and UO_1478 (O_1478,N_14202,N_14105);
nor UO_1479 (O_1479,N_14923,N_13801);
or UO_1480 (O_1480,N_14278,N_14443);
nand UO_1481 (O_1481,N_13717,N_14254);
or UO_1482 (O_1482,N_14761,N_13682);
or UO_1483 (O_1483,N_14174,N_14194);
or UO_1484 (O_1484,N_14706,N_13507);
and UO_1485 (O_1485,N_14550,N_14209);
and UO_1486 (O_1486,N_13806,N_14678);
or UO_1487 (O_1487,N_14448,N_14844);
nand UO_1488 (O_1488,N_13514,N_14688);
and UO_1489 (O_1489,N_13714,N_14624);
and UO_1490 (O_1490,N_13626,N_14453);
and UO_1491 (O_1491,N_14418,N_13823);
nand UO_1492 (O_1492,N_14419,N_13815);
or UO_1493 (O_1493,N_13898,N_14992);
or UO_1494 (O_1494,N_13963,N_13733);
and UO_1495 (O_1495,N_14721,N_14731);
nand UO_1496 (O_1496,N_14934,N_14438);
nand UO_1497 (O_1497,N_14352,N_14105);
xnor UO_1498 (O_1498,N_14129,N_14549);
nand UO_1499 (O_1499,N_14223,N_14602);
nand UO_1500 (O_1500,N_14663,N_14455);
or UO_1501 (O_1501,N_14770,N_13802);
or UO_1502 (O_1502,N_14563,N_13853);
nand UO_1503 (O_1503,N_14971,N_14118);
nand UO_1504 (O_1504,N_14834,N_14285);
nor UO_1505 (O_1505,N_14295,N_13563);
nor UO_1506 (O_1506,N_14004,N_14412);
xnor UO_1507 (O_1507,N_14684,N_14280);
nand UO_1508 (O_1508,N_14376,N_14464);
nor UO_1509 (O_1509,N_14788,N_14465);
and UO_1510 (O_1510,N_14080,N_14844);
or UO_1511 (O_1511,N_14214,N_13636);
nand UO_1512 (O_1512,N_14426,N_14637);
or UO_1513 (O_1513,N_14632,N_13680);
nand UO_1514 (O_1514,N_14239,N_14659);
nand UO_1515 (O_1515,N_14582,N_14000);
nand UO_1516 (O_1516,N_13631,N_14817);
xnor UO_1517 (O_1517,N_14427,N_14718);
nor UO_1518 (O_1518,N_14541,N_14960);
and UO_1519 (O_1519,N_14335,N_14610);
or UO_1520 (O_1520,N_13679,N_13640);
and UO_1521 (O_1521,N_13768,N_13507);
or UO_1522 (O_1522,N_14861,N_14017);
and UO_1523 (O_1523,N_14559,N_14132);
and UO_1524 (O_1524,N_14895,N_14958);
nand UO_1525 (O_1525,N_13748,N_13866);
nor UO_1526 (O_1526,N_14467,N_14566);
or UO_1527 (O_1527,N_13770,N_14640);
and UO_1528 (O_1528,N_14058,N_13919);
nand UO_1529 (O_1529,N_14530,N_13542);
nor UO_1530 (O_1530,N_14345,N_13610);
or UO_1531 (O_1531,N_14925,N_14678);
nand UO_1532 (O_1532,N_14107,N_14719);
and UO_1533 (O_1533,N_14651,N_14825);
nor UO_1534 (O_1534,N_13559,N_14668);
nor UO_1535 (O_1535,N_14101,N_13812);
nor UO_1536 (O_1536,N_13922,N_14003);
nand UO_1537 (O_1537,N_14983,N_13904);
and UO_1538 (O_1538,N_13987,N_13718);
nor UO_1539 (O_1539,N_13916,N_13828);
or UO_1540 (O_1540,N_14963,N_14178);
or UO_1541 (O_1541,N_14650,N_13890);
and UO_1542 (O_1542,N_14047,N_13577);
or UO_1543 (O_1543,N_14545,N_13948);
xor UO_1544 (O_1544,N_14255,N_14801);
nor UO_1545 (O_1545,N_13967,N_14972);
nor UO_1546 (O_1546,N_13700,N_14443);
or UO_1547 (O_1547,N_13898,N_14518);
nand UO_1548 (O_1548,N_14020,N_14064);
and UO_1549 (O_1549,N_14433,N_13561);
nor UO_1550 (O_1550,N_14883,N_13969);
or UO_1551 (O_1551,N_13582,N_13591);
and UO_1552 (O_1552,N_13997,N_13659);
and UO_1553 (O_1553,N_14595,N_14405);
and UO_1554 (O_1554,N_14266,N_13838);
nor UO_1555 (O_1555,N_13965,N_14478);
and UO_1556 (O_1556,N_14296,N_14074);
and UO_1557 (O_1557,N_14934,N_14777);
and UO_1558 (O_1558,N_14121,N_14219);
or UO_1559 (O_1559,N_14580,N_14179);
and UO_1560 (O_1560,N_14772,N_13701);
nand UO_1561 (O_1561,N_14889,N_13575);
nand UO_1562 (O_1562,N_14010,N_14498);
or UO_1563 (O_1563,N_14472,N_13563);
or UO_1564 (O_1564,N_14735,N_14022);
and UO_1565 (O_1565,N_13513,N_13891);
nor UO_1566 (O_1566,N_14081,N_14184);
nor UO_1567 (O_1567,N_14317,N_14498);
and UO_1568 (O_1568,N_13972,N_14263);
and UO_1569 (O_1569,N_13897,N_14019);
or UO_1570 (O_1570,N_14867,N_14173);
nand UO_1571 (O_1571,N_14316,N_14636);
nand UO_1572 (O_1572,N_14321,N_13584);
or UO_1573 (O_1573,N_14144,N_14781);
nand UO_1574 (O_1574,N_14290,N_14573);
xor UO_1575 (O_1575,N_14645,N_14838);
nor UO_1576 (O_1576,N_14464,N_14979);
and UO_1577 (O_1577,N_13999,N_13771);
nand UO_1578 (O_1578,N_14913,N_13737);
nand UO_1579 (O_1579,N_14928,N_14802);
nand UO_1580 (O_1580,N_14616,N_14147);
or UO_1581 (O_1581,N_13525,N_13987);
or UO_1582 (O_1582,N_13990,N_14164);
nor UO_1583 (O_1583,N_14711,N_14114);
xnor UO_1584 (O_1584,N_13956,N_14915);
xor UO_1585 (O_1585,N_14865,N_13673);
nor UO_1586 (O_1586,N_13642,N_13526);
nor UO_1587 (O_1587,N_13613,N_13691);
and UO_1588 (O_1588,N_14452,N_14254);
or UO_1589 (O_1589,N_14893,N_14320);
nand UO_1590 (O_1590,N_14153,N_13536);
nand UO_1591 (O_1591,N_14434,N_13835);
and UO_1592 (O_1592,N_14073,N_13532);
nor UO_1593 (O_1593,N_14978,N_14177);
nor UO_1594 (O_1594,N_14087,N_13715);
nand UO_1595 (O_1595,N_14077,N_13865);
nor UO_1596 (O_1596,N_14892,N_14798);
or UO_1597 (O_1597,N_14140,N_13763);
or UO_1598 (O_1598,N_14906,N_13837);
and UO_1599 (O_1599,N_14362,N_14475);
and UO_1600 (O_1600,N_13701,N_14313);
nor UO_1601 (O_1601,N_14263,N_13883);
and UO_1602 (O_1602,N_14862,N_14951);
nor UO_1603 (O_1603,N_13721,N_14130);
xnor UO_1604 (O_1604,N_13900,N_14191);
nand UO_1605 (O_1605,N_14473,N_14414);
and UO_1606 (O_1606,N_14230,N_13897);
or UO_1607 (O_1607,N_13544,N_14271);
nand UO_1608 (O_1608,N_14634,N_14599);
and UO_1609 (O_1609,N_13696,N_14247);
or UO_1610 (O_1610,N_14726,N_14502);
nand UO_1611 (O_1611,N_13543,N_14862);
and UO_1612 (O_1612,N_13600,N_13680);
nor UO_1613 (O_1613,N_14916,N_13590);
xnor UO_1614 (O_1614,N_13863,N_14542);
nor UO_1615 (O_1615,N_14827,N_14602);
or UO_1616 (O_1616,N_14779,N_14003);
and UO_1617 (O_1617,N_14718,N_13812);
nand UO_1618 (O_1618,N_13651,N_13838);
and UO_1619 (O_1619,N_14771,N_14217);
nor UO_1620 (O_1620,N_14294,N_14230);
nor UO_1621 (O_1621,N_13653,N_14245);
and UO_1622 (O_1622,N_13518,N_13864);
nor UO_1623 (O_1623,N_14634,N_14052);
nor UO_1624 (O_1624,N_14257,N_14845);
and UO_1625 (O_1625,N_14165,N_14794);
or UO_1626 (O_1626,N_14916,N_13522);
nor UO_1627 (O_1627,N_14700,N_14316);
nand UO_1628 (O_1628,N_14701,N_14291);
nand UO_1629 (O_1629,N_14113,N_14498);
nand UO_1630 (O_1630,N_14403,N_14356);
nand UO_1631 (O_1631,N_13570,N_14083);
or UO_1632 (O_1632,N_13817,N_13521);
nor UO_1633 (O_1633,N_13937,N_14075);
or UO_1634 (O_1634,N_14592,N_14116);
and UO_1635 (O_1635,N_14916,N_13510);
or UO_1636 (O_1636,N_13631,N_13752);
nor UO_1637 (O_1637,N_14273,N_13868);
and UO_1638 (O_1638,N_13678,N_14488);
nand UO_1639 (O_1639,N_14187,N_13719);
nor UO_1640 (O_1640,N_14301,N_14725);
or UO_1641 (O_1641,N_13657,N_13649);
xor UO_1642 (O_1642,N_14736,N_14677);
nor UO_1643 (O_1643,N_14713,N_14832);
and UO_1644 (O_1644,N_14642,N_14928);
and UO_1645 (O_1645,N_14364,N_14192);
nor UO_1646 (O_1646,N_13518,N_13936);
nand UO_1647 (O_1647,N_14955,N_13901);
nand UO_1648 (O_1648,N_14290,N_13932);
and UO_1649 (O_1649,N_13708,N_14246);
or UO_1650 (O_1650,N_13716,N_14161);
nand UO_1651 (O_1651,N_14601,N_14135);
and UO_1652 (O_1652,N_14277,N_14509);
nand UO_1653 (O_1653,N_13815,N_14955);
nor UO_1654 (O_1654,N_14514,N_13582);
nand UO_1655 (O_1655,N_13621,N_14299);
or UO_1656 (O_1656,N_13882,N_14390);
or UO_1657 (O_1657,N_14578,N_13734);
nor UO_1658 (O_1658,N_14971,N_14964);
and UO_1659 (O_1659,N_14442,N_14353);
or UO_1660 (O_1660,N_14441,N_14865);
and UO_1661 (O_1661,N_14205,N_14040);
nand UO_1662 (O_1662,N_14974,N_14081);
nand UO_1663 (O_1663,N_13626,N_14621);
or UO_1664 (O_1664,N_14829,N_13682);
or UO_1665 (O_1665,N_14296,N_13888);
and UO_1666 (O_1666,N_14756,N_14814);
nor UO_1667 (O_1667,N_14884,N_13846);
and UO_1668 (O_1668,N_13558,N_13528);
nand UO_1669 (O_1669,N_14011,N_13790);
nand UO_1670 (O_1670,N_14597,N_14384);
or UO_1671 (O_1671,N_13542,N_14531);
nand UO_1672 (O_1672,N_13650,N_14267);
or UO_1673 (O_1673,N_14442,N_14539);
and UO_1674 (O_1674,N_14956,N_13543);
and UO_1675 (O_1675,N_13664,N_14575);
nand UO_1676 (O_1676,N_14249,N_14738);
or UO_1677 (O_1677,N_14361,N_14639);
and UO_1678 (O_1678,N_14731,N_14324);
nand UO_1679 (O_1679,N_14948,N_14233);
nand UO_1680 (O_1680,N_14739,N_14642);
and UO_1681 (O_1681,N_13635,N_14366);
or UO_1682 (O_1682,N_13511,N_14824);
nor UO_1683 (O_1683,N_14776,N_13500);
and UO_1684 (O_1684,N_14107,N_14747);
nand UO_1685 (O_1685,N_14892,N_14262);
and UO_1686 (O_1686,N_14129,N_13644);
xnor UO_1687 (O_1687,N_13953,N_14921);
nand UO_1688 (O_1688,N_14870,N_13948);
nand UO_1689 (O_1689,N_13947,N_14873);
or UO_1690 (O_1690,N_14923,N_14178);
nor UO_1691 (O_1691,N_14284,N_14394);
and UO_1692 (O_1692,N_14836,N_13906);
nand UO_1693 (O_1693,N_13547,N_14032);
or UO_1694 (O_1694,N_14951,N_14182);
nand UO_1695 (O_1695,N_13694,N_14954);
nor UO_1696 (O_1696,N_14377,N_14416);
nand UO_1697 (O_1697,N_13500,N_13552);
nand UO_1698 (O_1698,N_14771,N_13642);
nor UO_1699 (O_1699,N_14632,N_14310);
or UO_1700 (O_1700,N_14454,N_14242);
nand UO_1701 (O_1701,N_13909,N_14762);
nor UO_1702 (O_1702,N_14251,N_14552);
or UO_1703 (O_1703,N_14925,N_14266);
nand UO_1704 (O_1704,N_14805,N_14797);
nand UO_1705 (O_1705,N_13525,N_13872);
and UO_1706 (O_1706,N_14905,N_13527);
nand UO_1707 (O_1707,N_14182,N_14256);
or UO_1708 (O_1708,N_14046,N_13536);
nor UO_1709 (O_1709,N_14840,N_13716);
nor UO_1710 (O_1710,N_13501,N_14800);
nand UO_1711 (O_1711,N_14744,N_13954);
nor UO_1712 (O_1712,N_14328,N_14134);
and UO_1713 (O_1713,N_14073,N_14184);
or UO_1714 (O_1714,N_13775,N_13751);
nor UO_1715 (O_1715,N_13841,N_14999);
and UO_1716 (O_1716,N_14133,N_13614);
or UO_1717 (O_1717,N_13669,N_13584);
nor UO_1718 (O_1718,N_13607,N_14983);
or UO_1719 (O_1719,N_14399,N_14380);
nand UO_1720 (O_1720,N_14830,N_13569);
xnor UO_1721 (O_1721,N_14875,N_14976);
or UO_1722 (O_1722,N_14490,N_13752);
nand UO_1723 (O_1723,N_14100,N_14310);
nor UO_1724 (O_1724,N_14691,N_14291);
nor UO_1725 (O_1725,N_14812,N_13728);
or UO_1726 (O_1726,N_14341,N_14229);
nor UO_1727 (O_1727,N_13866,N_13894);
nand UO_1728 (O_1728,N_13994,N_13626);
or UO_1729 (O_1729,N_14349,N_14173);
or UO_1730 (O_1730,N_14552,N_13826);
or UO_1731 (O_1731,N_14675,N_14106);
nand UO_1732 (O_1732,N_14459,N_13614);
or UO_1733 (O_1733,N_14865,N_14790);
or UO_1734 (O_1734,N_13865,N_13622);
and UO_1735 (O_1735,N_14518,N_13839);
and UO_1736 (O_1736,N_13712,N_14591);
nor UO_1737 (O_1737,N_14868,N_14171);
xnor UO_1738 (O_1738,N_14347,N_13643);
and UO_1739 (O_1739,N_14260,N_14062);
nand UO_1740 (O_1740,N_14035,N_14833);
nor UO_1741 (O_1741,N_13594,N_14784);
nand UO_1742 (O_1742,N_14014,N_13695);
nor UO_1743 (O_1743,N_13894,N_13529);
nor UO_1744 (O_1744,N_14975,N_13806);
nand UO_1745 (O_1745,N_14774,N_14787);
nor UO_1746 (O_1746,N_14434,N_14026);
and UO_1747 (O_1747,N_13530,N_13829);
nor UO_1748 (O_1748,N_14866,N_14001);
nand UO_1749 (O_1749,N_14373,N_13951);
nand UO_1750 (O_1750,N_13517,N_13694);
nor UO_1751 (O_1751,N_14545,N_14805);
nand UO_1752 (O_1752,N_14039,N_14615);
nor UO_1753 (O_1753,N_13848,N_13903);
or UO_1754 (O_1754,N_14402,N_14102);
nor UO_1755 (O_1755,N_13784,N_14869);
and UO_1756 (O_1756,N_13724,N_13849);
nor UO_1757 (O_1757,N_13505,N_14681);
nor UO_1758 (O_1758,N_13673,N_13702);
nor UO_1759 (O_1759,N_13788,N_14076);
nand UO_1760 (O_1760,N_14441,N_14582);
or UO_1761 (O_1761,N_14683,N_13552);
or UO_1762 (O_1762,N_14673,N_13644);
or UO_1763 (O_1763,N_14302,N_13649);
nor UO_1764 (O_1764,N_14471,N_14814);
nor UO_1765 (O_1765,N_13753,N_14117);
and UO_1766 (O_1766,N_14116,N_13951);
or UO_1767 (O_1767,N_14365,N_14343);
and UO_1768 (O_1768,N_13533,N_13913);
or UO_1769 (O_1769,N_14846,N_14567);
and UO_1770 (O_1770,N_14490,N_14759);
nand UO_1771 (O_1771,N_13592,N_14958);
and UO_1772 (O_1772,N_14093,N_13552);
nand UO_1773 (O_1773,N_14198,N_14520);
and UO_1774 (O_1774,N_14314,N_14559);
nand UO_1775 (O_1775,N_14041,N_14451);
or UO_1776 (O_1776,N_13672,N_13868);
nor UO_1777 (O_1777,N_13515,N_13679);
and UO_1778 (O_1778,N_14709,N_13903);
xor UO_1779 (O_1779,N_14434,N_13884);
nand UO_1780 (O_1780,N_14556,N_13507);
or UO_1781 (O_1781,N_13705,N_13501);
nand UO_1782 (O_1782,N_13659,N_14434);
nand UO_1783 (O_1783,N_14027,N_14695);
nor UO_1784 (O_1784,N_14429,N_13807);
or UO_1785 (O_1785,N_14599,N_13520);
and UO_1786 (O_1786,N_14738,N_13828);
nand UO_1787 (O_1787,N_14042,N_13919);
and UO_1788 (O_1788,N_14066,N_14776);
and UO_1789 (O_1789,N_13882,N_14406);
and UO_1790 (O_1790,N_13523,N_14433);
and UO_1791 (O_1791,N_14350,N_14500);
or UO_1792 (O_1792,N_13798,N_13620);
xor UO_1793 (O_1793,N_14519,N_14323);
or UO_1794 (O_1794,N_14412,N_14486);
nand UO_1795 (O_1795,N_13962,N_14377);
and UO_1796 (O_1796,N_13784,N_13839);
and UO_1797 (O_1797,N_14430,N_13533);
or UO_1798 (O_1798,N_14450,N_14764);
or UO_1799 (O_1799,N_14078,N_14519);
and UO_1800 (O_1800,N_14794,N_14909);
nand UO_1801 (O_1801,N_13612,N_13550);
and UO_1802 (O_1802,N_14492,N_14011);
and UO_1803 (O_1803,N_14201,N_14112);
or UO_1804 (O_1804,N_14739,N_14802);
nor UO_1805 (O_1805,N_13725,N_14097);
nor UO_1806 (O_1806,N_13564,N_13765);
or UO_1807 (O_1807,N_13770,N_14251);
nand UO_1808 (O_1808,N_14508,N_13693);
or UO_1809 (O_1809,N_14710,N_14043);
nand UO_1810 (O_1810,N_14479,N_14400);
and UO_1811 (O_1811,N_14858,N_14334);
and UO_1812 (O_1812,N_14192,N_13912);
nand UO_1813 (O_1813,N_13771,N_14357);
or UO_1814 (O_1814,N_14256,N_14221);
or UO_1815 (O_1815,N_13956,N_13722);
xnor UO_1816 (O_1816,N_14292,N_13639);
or UO_1817 (O_1817,N_14763,N_13680);
nand UO_1818 (O_1818,N_14589,N_13514);
nor UO_1819 (O_1819,N_14898,N_13750);
or UO_1820 (O_1820,N_14498,N_13724);
or UO_1821 (O_1821,N_14175,N_14417);
nand UO_1822 (O_1822,N_14224,N_13839);
nor UO_1823 (O_1823,N_13707,N_13874);
or UO_1824 (O_1824,N_13752,N_14790);
nand UO_1825 (O_1825,N_14632,N_14062);
nand UO_1826 (O_1826,N_13991,N_13922);
nand UO_1827 (O_1827,N_14104,N_14117);
or UO_1828 (O_1828,N_13834,N_14924);
or UO_1829 (O_1829,N_14291,N_13580);
nand UO_1830 (O_1830,N_13801,N_13824);
nand UO_1831 (O_1831,N_14733,N_14269);
nor UO_1832 (O_1832,N_14929,N_13720);
nor UO_1833 (O_1833,N_14895,N_13693);
nand UO_1834 (O_1834,N_14712,N_14294);
nand UO_1835 (O_1835,N_14528,N_14503);
and UO_1836 (O_1836,N_14213,N_13811);
nand UO_1837 (O_1837,N_13943,N_14902);
nand UO_1838 (O_1838,N_14417,N_13800);
nor UO_1839 (O_1839,N_13952,N_13953);
or UO_1840 (O_1840,N_14467,N_13549);
nor UO_1841 (O_1841,N_13998,N_14401);
nor UO_1842 (O_1842,N_14222,N_13892);
nand UO_1843 (O_1843,N_13769,N_14679);
nand UO_1844 (O_1844,N_13877,N_14012);
or UO_1845 (O_1845,N_14041,N_13873);
and UO_1846 (O_1846,N_14013,N_14911);
or UO_1847 (O_1847,N_14492,N_14319);
nand UO_1848 (O_1848,N_14174,N_13706);
nand UO_1849 (O_1849,N_14212,N_13814);
or UO_1850 (O_1850,N_13690,N_14696);
nor UO_1851 (O_1851,N_14819,N_14228);
and UO_1852 (O_1852,N_13640,N_14229);
and UO_1853 (O_1853,N_14095,N_14658);
nand UO_1854 (O_1854,N_13683,N_14752);
or UO_1855 (O_1855,N_14871,N_14359);
nand UO_1856 (O_1856,N_13821,N_14370);
xnor UO_1857 (O_1857,N_14256,N_13905);
nand UO_1858 (O_1858,N_14131,N_13967);
xnor UO_1859 (O_1859,N_14614,N_14325);
nand UO_1860 (O_1860,N_14549,N_13517);
or UO_1861 (O_1861,N_14257,N_14067);
or UO_1862 (O_1862,N_13666,N_13900);
or UO_1863 (O_1863,N_14118,N_14174);
nand UO_1864 (O_1864,N_14798,N_14466);
and UO_1865 (O_1865,N_14373,N_14124);
nor UO_1866 (O_1866,N_13984,N_14859);
nor UO_1867 (O_1867,N_14018,N_14068);
or UO_1868 (O_1868,N_14918,N_14501);
nor UO_1869 (O_1869,N_14212,N_14374);
nand UO_1870 (O_1870,N_14043,N_14970);
nand UO_1871 (O_1871,N_13865,N_14852);
nor UO_1872 (O_1872,N_14079,N_13538);
nand UO_1873 (O_1873,N_14338,N_14822);
nand UO_1874 (O_1874,N_14438,N_14213);
or UO_1875 (O_1875,N_13938,N_14465);
nand UO_1876 (O_1876,N_14013,N_14657);
or UO_1877 (O_1877,N_13509,N_14642);
and UO_1878 (O_1878,N_14115,N_13513);
nand UO_1879 (O_1879,N_13587,N_13503);
or UO_1880 (O_1880,N_13576,N_13764);
or UO_1881 (O_1881,N_14888,N_14433);
nor UO_1882 (O_1882,N_14437,N_14708);
nor UO_1883 (O_1883,N_13573,N_13641);
or UO_1884 (O_1884,N_14633,N_13746);
nand UO_1885 (O_1885,N_13559,N_14838);
nor UO_1886 (O_1886,N_13587,N_14806);
and UO_1887 (O_1887,N_13715,N_14034);
nand UO_1888 (O_1888,N_13839,N_14884);
nand UO_1889 (O_1889,N_14054,N_14465);
and UO_1890 (O_1890,N_13765,N_14620);
and UO_1891 (O_1891,N_13828,N_14560);
or UO_1892 (O_1892,N_14339,N_13584);
and UO_1893 (O_1893,N_14223,N_14970);
and UO_1894 (O_1894,N_14903,N_14177);
nand UO_1895 (O_1895,N_14566,N_14713);
or UO_1896 (O_1896,N_13815,N_14468);
and UO_1897 (O_1897,N_13692,N_14929);
nor UO_1898 (O_1898,N_14871,N_13945);
and UO_1899 (O_1899,N_14547,N_14436);
and UO_1900 (O_1900,N_13636,N_13677);
and UO_1901 (O_1901,N_13715,N_14828);
nand UO_1902 (O_1902,N_14374,N_14295);
nand UO_1903 (O_1903,N_13798,N_14019);
nand UO_1904 (O_1904,N_14566,N_14326);
or UO_1905 (O_1905,N_13933,N_14596);
nor UO_1906 (O_1906,N_14184,N_14032);
and UO_1907 (O_1907,N_14930,N_14206);
and UO_1908 (O_1908,N_13761,N_14550);
nand UO_1909 (O_1909,N_14760,N_14168);
and UO_1910 (O_1910,N_14372,N_13989);
nand UO_1911 (O_1911,N_13912,N_14436);
or UO_1912 (O_1912,N_14982,N_13547);
or UO_1913 (O_1913,N_13673,N_13897);
nand UO_1914 (O_1914,N_14964,N_14054);
nor UO_1915 (O_1915,N_14502,N_13673);
nor UO_1916 (O_1916,N_13994,N_14795);
or UO_1917 (O_1917,N_14837,N_14275);
or UO_1918 (O_1918,N_14201,N_14378);
and UO_1919 (O_1919,N_14773,N_14361);
and UO_1920 (O_1920,N_14394,N_14658);
nor UO_1921 (O_1921,N_14782,N_14835);
or UO_1922 (O_1922,N_14214,N_14397);
and UO_1923 (O_1923,N_14118,N_14687);
nor UO_1924 (O_1924,N_14751,N_14581);
nand UO_1925 (O_1925,N_14496,N_14436);
and UO_1926 (O_1926,N_14348,N_14963);
and UO_1927 (O_1927,N_14332,N_13726);
nand UO_1928 (O_1928,N_14471,N_14264);
nor UO_1929 (O_1929,N_13949,N_14926);
and UO_1930 (O_1930,N_14697,N_13763);
and UO_1931 (O_1931,N_14353,N_13908);
nand UO_1932 (O_1932,N_14558,N_14162);
or UO_1933 (O_1933,N_14324,N_14662);
xor UO_1934 (O_1934,N_14182,N_13961);
nand UO_1935 (O_1935,N_14320,N_13637);
or UO_1936 (O_1936,N_13797,N_14762);
or UO_1937 (O_1937,N_14172,N_14280);
nor UO_1938 (O_1938,N_14047,N_13737);
and UO_1939 (O_1939,N_14211,N_14445);
nand UO_1940 (O_1940,N_14967,N_14392);
nor UO_1941 (O_1941,N_14118,N_14984);
nor UO_1942 (O_1942,N_14447,N_14054);
nor UO_1943 (O_1943,N_13831,N_13843);
nand UO_1944 (O_1944,N_14981,N_14276);
nand UO_1945 (O_1945,N_14468,N_14552);
nor UO_1946 (O_1946,N_13553,N_14088);
and UO_1947 (O_1947,N_13578,N_14663);
or UO_1948 (O_1948,N_14994,N_14582);
or UO_1949 (O_1949,N_14543,N_13981);
or UO_1950 (O_1950,N_14899,N_14608);
or UO_1951 (O_1951,N_13810,N_14578);
nor UO_1952 (O_1952,N_14881,N_14019);
nand UO_1953 (O_1953,N_14866,N_14336);
nor UO_1954 (O_1954,N_13767,N_13556);
and UO_1955 (O_1955,N_14399,N_14626);
nand UO_1956 (O_1956,N_13545,N_14400);
nand UO_1957 (O_1957,N_14662,N_14351);
or UO_1958 (O_1958,N_14749,N_14615);
nand UO_1959 (O_1959,N_13913,N_14879);
and UO_1960 (O_1960,N_13879,N_14896);
nand UO_1961 (O_1961,N_14306,N_14265);
nor UO_1962 (O_1962,N_13590,N_14510);
nor UO_1963 (O_1963,N_14040,N_14665);
nand UO_1964 (O_1964,N_14826,N_14179);
nor UO_1965 (O_1965,N_13500,N_14350);
or UO_1966 (O_1966,N_14405,N_14580);
nand UO_1967 (O_1967,N_14419,N_13709);
and UO_1968 (O_1968,N_14258,N_13807);
xnor UO_1969 (O_1969,N_14969,N_13942);
or UO_1970 (O_1970,N_14735,N_14409);
or UO_1971 (O_1971,N_14082,N_13678);
or UO_1972 (O_1972,N_13955,N_14913);
nor UO_1973 (O_1973,N_14960,N_14665);
nor UO_1974 (O_1974,N_14135,N_14259);
or UO_1975 (O_1975,N_14488,N_14434);
nand UO_1976 (O_1976,N_14462,N_14948);
nor UO_1977 (O_1977,N_14168,N_14000);
or UO_1978 (O_1978,N_14207,N_14592);
nor UO_1979 (O_1979,N_13729,N_13511);
and UO_1980 (O_1980,N_14695,N_14128);
or UO_1981 (O_1981,N_14528,N_14916);
or UO_1982 (O_1982,N_14382,N_13709);
nor UO_1983 (O_1983,N_14099,N_14010);
nor UO_1984 (O_1984,N_14647,N_14502);
nor UO_1985 (O_1985,N_14492,N_13563);
and UO_1986 (O_1986,N_14254,N_14199);
nor UO_1987 (O_1987,N_13889,N_14827);
and UO_1988 (O_1988,N_14659,N_13535);
xor UO_1989 (O_1989,N_13525,N_13896);
nor UO_1990 (O_1990,N_13836,N_14948);
nor UO_1991 (O_1991,N_13927,N_13875);
nand UO_1992 (O_1992,N_14049,N_14010);
or UO_1993 (O_1993,N_14034,N_14485);
or UO_1994 (O_1994,N_14900,N_14184);
nand UO_1995 (O_1995,N_14956,N_13944);
nor UO_1996 (O_1996,N_14567,N_14977);
nor UO_1997 (O_1997,N_14518,N_13914);
xor UO_1998 (O_1998,N_14564,N_14287);
or UO_1999 (O_1999,N_13945,N_14207);
endmodule