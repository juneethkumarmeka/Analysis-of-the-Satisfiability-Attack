module basic_3000_30000_3500_20_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1807,In_1640);
nor U1 (N_1,In_1655,In_2160);
nor U2 (N_2,In_2812,In_2501);
nand U3 (N_3,In_1231,In_2674);
and U4 (N_4,In_1465,In_2129);
nand U5 (N_5,In_584,In_1579);
nor U6 (N_6,In_2955,In_2405);
xor U7 (N_7,In_520,In_1515);
and U8 (N_8,In_2964,In_1799);
xor U9 (N_9,In_2411,In_1141);
or U10 (N_10,In_2296,In_1104);
and U11 (N_11,In_1046,In_1442);
xnor U12 (N_12,In_1957,In_458);
or U13 (N_13,In_1009,In_714);
and U14 (N_14,In_2809,In_132);
xor U15 (N_15,In_1437,In_915);
nand U16 (N_16,In_691,In_2201);
nor U17 (N_17,In_2705,In_642);
or U18 (N_18,In_1761,In_2596);
xnor U19 (N_19,In_281,In_1683);
nor U20 (N_20,In_2865,In_1066);
and U21 (N_21,In_2560,In_1914);
nor U22 (N_22,In_2617,In_1153);
nand U23 (N_23,In_262,In_1085);
nand U24 (N_24,In_983,In_1417);
xnor U25 (N_25,In_2747,In_1361);
nand U26 (N_26,In_2649,In_2268);
nand U27 (N_27,In_2307,In_2291);
nand U28 (N_28,In_122,In_2579);
nor U29 (N_29,In_2698,In_981);
or U30 (N_30,In_2357,In_2892);
xor U31 (N_31,In_1834,In_1840);
and U32 (N_32,In_1255,In_1450);
and U33 (N_33,In_652,In_2912);
or U34 (N_34,In_1200,In_1552);
or U35 (N_35,In_1239,In_1014);
xor U36 (N_36,In_865,In_615);
or U37 (N_37,In_1965,In_794);
or U38 (N_38,In_1147,In_2563);
xor U39 (N_39,In_2799,In_2039);
xnor U40 (N_40,In_2204,In_2025);
nor U41 (N_41,In_1752,In_2203);
nand U42 (N_42,In_2637,In_445);
or U43 (N_43,In_2005,In_775);
xnor U44 (N_44,In_2278,In_2722);
nor U45 (N_45,In_2101,In_918);
nor U46 (N_46,In_2800,In_2707);
or U47 (N_47,In_1942,In_561);
nand U48 (N_48,In_1839,In_411);
or U49 (N_49,In_1464,In_113);
nand U50 (N_50,In_38,In_1952);
and U51 (N_51,In_278,In_585);
nor U52 (N_52,In_1788,In_2531);
nand U53 (N_53,In_2252,In_1912);
and U54 (N_54,In_635,In_1944);
nand U55 (N_55,In_2754,In_2712);
nor U56 (N_56,In_2951,In_1340);
nand U57 (N_57,In_2830,In_2313);
nand U58 (N_58,In_607,In_677);
or U59 (N_59,In_1953,In_947);
nor U60 (N_60,In_1156,In_604);
nor U61 (N_61,In_2687,In_1859);
and U62 (N_62,In_2670,In_1630);
xor U63 (N_63,In_2123,In_2423);
nor U64 (N_64,In_1381,In_233);
or U65 (N_65,In_1501,In_1370);
nand U66 (N_66,In_455,In_2793);
xnor U67 (N_67,In_1664,In_683);
xor U68 (N_68,In_2544,In_1565);
and U69 (N_69,In_2339,In_568);
nor U70 (N_70,In_1398,In_1249);
xor U71 (N_71,In_1981,In_2012);
nor U72 (N_72,In_444,In_2390);
nor U73 (N_73,In_2285,In_24);
xor U74 (N_74,In_2728,In_2181);
xnor U75 (N_75,In_2836,In_1477);
nor U76 (N_76,In_183,In_1406);
nand U77 (N_77,In_2925,In_215);
or U78 (N_78,In_1031,In_1778);
or U79 (N_79,In_2618,In_746);
xor U80 (N_80,In_206,In_512);
or U81 (N_81,In_501,In_2169);
and U82 (N_82,In_511,In_174);
nor U83 (N_83,In_284,In_2472);
and U84 (N_84,In_196,In_2695);
and U85 (N_85,In_1117,In_2332);
and U86 (N_86,In_1876,In_1808);
nand U87 (N_87,In_1268,In_464);
nand U88 (N_88,In_1393,In_973);
xnor U89 (N_89,In_239,In_581);
and U90 (N_90,In_253,In_84);
and U91 (N_91,In_2972,In_1620);
or U92 (N_92,In_1706,In_329);
nor U93 (N_93,In_533,In_1265);
xnor U94 (N_94,In_352,In_1428);
xor U95 (N_95,In_1690,In_922);
nand U96 (N_96,In_1910,In_1182);
xor U97 (N_97,In_920,In_2262);
or U98 (N_98,In_706,In_315);
nor U99 (N_99,In_1120,In_2015);
nor U100 (N_100,In_2526,In_2042);
nand U101 (N_101,In_2509,In_1628);
nor U102 (N_102,In_2969,In_1254);
or U103 (N_103,In_1305,In_1835);
nand U104 (N_104,In_1857,In_1040);
and U105 (N_105,In_2487,In_209);
nor U106 (N_106,In_1487,In_83);
xnor U107 (N_107,In_2853,In_382);
and U108 (N_108,In_1391,In_1734);
nor U109 (N_109,In_1336,In_2067);
nand U110 (N_110,In_1415,In_2959);
and U111 (N_111,In_2701,In_251);
nor U112 (N_112,In_489,In_576);
and U113 (N_113,In_569,In_2026);
or U114 (N_114,In_1682,In_440);
xnor U115 (N_115,In_356,In_2246);
or U116 (N_116,In_1668,In_921);
xnor U117 (N_117,In_15,In_468);
xnor U118 (N_118,In_147,In_2207);
and U119 (N_119,In_1351,In_620);
xnor U120 (N_120,In_2831,In_1161);
xnor U121 (N_121,In_1257,In_2446);
nor U122 (N_122,In_1926,In_96);
nand U123 (N_123,In_2982,In_1824);
and U124 (N_124,In_8,In_1800);
or U125 (N_125,In_2003,In_2240);
and U126 (N_126,In_3,In_142);
nand U127 (N_127,In_1679,In_2182);
nor U128 (N_128,In_1403,In_854);
and U129 (N_129,In_1791,In_2073);
nor U130 (N_130,In_828,In_1897);
or U131 (N_131,In_2915,In_1606);
and U132 (N_132,In_2779,In_2211);
nand U133 (N_133,In_2088,In_228);
xnor U134 (N_134,In_1865,In_2055);
xor U135 (N_135,In_293,In_1158);
nor U136 (N_136,In_1976,In_2612);
and U137 (N_137,In_1137,In_1502);
nand U138 (N_138,In_807,In_28);
nand U139 (N_139,In_1353,In_2166);
xnor U140 (N_140,In_1478,In_645);
and U141 (N_141,In_1138,In_1537);
and U142 (N_142,In_686,In_1469);
or U143 (N_143,In_2994,In_1637);
nor U144 (N_144,In_2842,In_1073);
nor U145 (N_145,In_617,In_2510);
nor U146 (N_146,In_2774,In_1726);
nand U147 (N_147,In_968,In_1877);
xor U148 (N_148,In_388,In_109);
and U149 (N_149,In_2691,In_119);
xnor U150 (N_150,In_2205,In_1033);
or U151 (N_151,In_1258,In_1235);
and U152 (N_152,In_780,In_210);
or U153 (N_153,In_1320,In_274);
nand U154 (N_154,In_705,In_2826);
xor U155 (N_155,In_2217,In_2881);
or U156 (N_156,In_149,In_949);
or U157 (N_157,In_1619,In_2931);
nor U158 (N_158,In_2180,In_1260);
xnor U159 (N_159,In_1773,In_773);
nand U160 (N_160,In_847,In_2730);
nor U161 (N_161,In_2578,In_924);
nand U162 (N_162,In_186,In_2079);
nand U163 (N_163,In_791,In_2932);
nor U164 (N_164,In_1636,In_78);
or U165 (N_165,In_936,In_1961);
nand U166 (N_166,In_2330,In_2938);
nor U167 (N_167,In_1938,In_806);
and U168 (N_168,In_504,In_1987);
nor U169 (N_169,In_1722,In_127);
nand U170 (N_170,In_2421,In_135);
nand U171 (N_171,In_1899,In_2046);
xor U172 (N_172,In_1850,In_1584);
xor U173 (N_173,In_1764,In_2970);
or U174 (N_174,In_379,In_788);
nor U175 (N_175,In_2795,In_1823);
and U176 (N_176,In_942,In_1357);
nand U177 (N_177,In_2383,In_463);
nand U178 (N_178,In_1038,In_2045);
xnor U179 (N_179,In_2667,In_808);
nand U180 (N_180,In_1844,In_1184);
and U181 (N_181,In_157,In_19);
and U182 (N_182,In_2576,In_1276);
xor U183 (N_183,In_2097,In_1385);
or U184 (N_184,In_600,In_245);
or U185 (N_185,In_2369,In_2197);
nand U186 (N_186,In_1646,In_2402);
xnor U187 (N_187,In_731,In_744);
and U188 (N_188,In_249,In_1697);
nand U189 (N_189,In_2610,In_2115);
nand U190 (N_190,In_970,In_179);
and U191 (N_191,In_1941,In_650);
and U192 (N_192,In_2273,In_2384);
and U193 (N_193,In_1724,In_128);
xor U194 (N_194,In_451,In_2414);
and U195 (N_195,In_760,In_2876);
xnor U196 (N_196,In_2124,In_2480);
xor U197 (N_197,In_2671,In_2403);
or U198 (N_198,In_335,In_2630);
xor U199 (N_199,In_449,In_2469);
nor U200 (N_200,In_1321,In_161);
or U201 (N_201,In_1448,In_955);
or U202 (N_202,In_1443,In_137);
nor U203 (N_203,In_442,In_2893);
or U204 (N_204,In_1185,In_1191);
nand U205 (N_205,In_2785,In_400);
or U206 (N_206,In_2080,In_2622);
and U207 (N_207,In_1407,In_2658);
nand U208 (N_208,In_567,In_1974);
xnor U209 (N_209,In_82,In_1744);
nand U210 (N_210,In_1253,In_2839);
or U211 (N_211,In_1713,In_1476);
xnor U212 (N_212,In_897,In_1095);
nor U213 (N_213,In_1146,In_402);
nand U214 (N_214,In_2214,In_2266);
or U215 (N_215,In_2766,In_2334);
xnor U216 (N_216,In_2483,In_2723);
nor U217 (N_217,In_2492,In_181);
or U218 (N_218,In_2855,In_1400);
nand U219 (N_219,In_2318,In_553);
and U220 (N_220,In_2133,In_1310);
and U221 (N_221,In_2693,In_996);
and U222 (N_222,In_2535,In_2961);
or U223 (N_223,In_2121,In_1090);
and U224 (N_224,In_1853,In_2755);
nand U225 (N_225,In_597,In_658);
nor U226 (N_226,In_241,In_551);
and U227 (N_227,In_832,In_2586);
nand U228 (N_228,In_1661,In_301);
xor U229 (N_229,In_2780,In_474);
nor U230 (N_230,In_713,In_2742);
xor U231 (N_231,In_1447,In_1498);
xnor U232 (N_232,In_1580,In_1226);
and U233 (N_233,In_1607,In_289);
nor U234 (N_234,In_528,In_1463);
nand U235 (N_235,In_1078,In_2632);
xor U236 (N_236,In_815,In_362);
or U237 (N_237,In_1955,In_2430);
nand U238 (N_238,In_261,In_2297);
and U239 (N_239,In_1044,In_1013);
nor U240 (N_240,In_1885,In_2222);
or U241 (N_241,In_1317,In_1525);
xor U242 (N_242,In_2344,In_934);
or U243 (N_243,In_27,In_1071);
or U244 (N_244,In_2634,In_2271);
or U245 (N_245,In_2615,In_2434);
xor U246 (N_246,In_177,In_795);
xor U247 (N_247,In_1803,In_2335);
nand U248 (N_248,In_861,In_2275);
nand U249 (N_249,In_2752,In_1238);
xnor U250 (N_250,In_1227,In_1083);
nor U251 (N_251,In_2984,In_348);
nand U252 (N_252,In_1805,In_152);
or U253 (N_253,In_2293,In_2870);
or U254 (N_254,In_1759,In_91);
nor U255 (N_255,In_66,In_2758);
nor U256 (N_256,In_1248,In_491);
nor U257 (N_257,In_2543,In_280);
xor U258 (N_258,In_1990,In_2888);
or U259 (N_259,In_2212,In_679);
and U260 (N_260,In_220,In_2466);
and U261 (N_261,In_1197,In_1010);
xor U262 (N_262,In_1963,In_769);
nand U263 (N_263,In_232,In_1927);
nor U264 (N_264,In_2896,In_1451);
xnor U265 (N_265,In_763,In_782);
xnor U266 (N_266,In_116,In_2161);
xnor U267 (N_267,In_264,In_1563);
nand U268 (N_268,In_1416,In_2355);
or U269 (N_269,In_1294,In_1700);
nand U270 (N_270,In_2873,In_2602);
or U271 (N_271,In_1982,In_820);
xnor U272 (N_272,In_2993,In_1766);
and U273 (N_273,In_979,In_1680);
nor U274 (N_274,In_1745,In_2497);
xnor U275 (N_275,In_523,In_2781);
nor U276 (N_276,In_2852,In_2810);
nand U277 (N_277,In_2152,In_418);
xnor U278 (N_278,In_68,In_2192);
nand U279 (N_279,In_2044,In_1298);
xnor U280 (N_280,In_1500,In_1711);
nand U281 (N_281,In_219,In_1190);
nor U282 (N_282,In_1002,In_764);
and U283 (N_283,In_2484,In_1937);
xnor U284 (N_284,In_2768,In_2775);
or U285 (N_285,In_2032,In_2762);
or U286 (N_286,In_130,In_2269);
xnor U287 (N_287,In_1519,In_2744);
or U288 (N_288,In_818,In_257);
or U289 (N_289,In_333,In_1650);
or U290 (N_290,In_419,In_1827);
nor U291 (N_291,In_1207,In_208);
and U292 (N_292,In_287,In_1131);
xor U293 (N_293,In_2452,In_1828);
or U294 (N_294,In_1060,In_1180);
nor U295 (N_295,In_2627,In_882);
xor U296 (N_296,In_2651,In_1316);
nand U297 (N_297,In_1420,In_336);
xnor U298 (N_298,In_154,In_2159);
nand U299 (N_299,In_2022,In_1424);
xnor U300 (N_300,In_1780,In_1929);
nor U301 (N_301,In_1318,In_2569);
and U302 (N_302,In_1301,In_2745);
nand U303 (N_303,In_1196,In_2949);
and U304 (N_304,In_354,In_361);
or U305 (N_305,In_1728,In_2004);
and U306 (N_306,In_235,In_2131);
xnor U307 (N_307,In_1849,In_656);
or U308 (N_308,In_212,In_950);
xor U309 (N_309,In_2567,In_2624);
nor U310 (N_310,In_2224,In_1194);
nand U311 (N_311,In_1003,In_260);
nand U312 (N_312,In_187,In_2682);
xnor U313 (N_313,In_1577,In_1287);
or U314 (N_314,In_2903,In_509);
or U315 (N_315,In_2021,In_709);
nor U316 (N_316,In_1529,In_325);
and U317 (N_317,In_614,In_880);
and U318 (N_318,In_95,In_640);
and U319 (N_319,In_631,In_459);
nand U320 (N_320,In_1064,In_2422);
nor U321 (N_321,In_870,In_2155);
nand U322 (N_322,In_1118,In_2690);
and U323 (N_323,In_1608,In_1947);
nor U324 (N_324,In_1466,In_1719);
or U325 (N_325,In_2248,In_125);
nand U326 (N_326,In_2909,In_1684);
nand U327 (N_327,In_2570,In_2054);
xnor U328 (N_328,In_805,In_609);
or U329 (N_329,In_1241,In_410);
nor U330 (N_330,In_2595,In_1402);
or U331 (N_331,In_1335,In_1916);
or U332 (N_332,In_2660,In_2528);
or U333 (N_333,In_2188,In_1647);
nand U334 (N_334,In_708,In_1059);
nor U335 (N_335,In_193,In_790);
nor U336 (N_336,In_1022,In_376);
nand U337 (N_337,In_560,In_1485);
nor U338 (N_338,In_2902,In_1562);
or U339 (N_339,In_2106,In_156);
or U340 (N_340,In_2257,In_1667);
nand U341 (N_341,In_23,In_1432);
nor U342 (N_342,In_1838,In_2144);
nand U343 (N_343,In_1509,In_31);
nor U344 (N_344,In_563,In_1052);
or U345 (N_345,In_589,In_108);
nor U346 (N_346,In_342,In_1069);
or U347 (N_347,In_2213,In_1244);
nor U348 (N_348,In_2232,In_2153);
nand U349 (N_349,In_55,In_2037);
xnor U350 (N_350,In_0,In_1781);
nand U351 (N_351,In_2559,In_2347);
xnor U352 (N_352,In_2817,In_63);
and U353 (N_353,In_732,In_2065);
xor U354 (N_354,In_1496,In_1288);
and U355 (N_355,In_188,In_1396);
nand U356 (N_356,In_761,In_197);
and U357 (N_357,In_518,In_2735);
or U358 (N_358,In_2898,In_1341);
xor U359 (N_359,In_1209,In_2546);
and U360 (N_360,In_727,In_200);
nand U361 (N_361,In_701,In_2713);
nor U362 (N_362,In_1600,In_1218);
and U363 (N_363,In_2479,In_437);
xnor U364 (N_364,In_1538,In_1864);
or U365 (N_365,In_1387,In_283);
xnor U366 (N_366,In_2024,In_1930);
nand U367 (N_367,In_2465,In_2132);
nor U368 (N_368,In_999,In_496);
xnor U369 (N_369,In_676,In_2103);
nand U370 (N_370,In_2074,In_1481);
or U371 (N_371,In_1792,In_2765);
nand U372 (N_372,In_2680,In_982);
nor U373 (N_373,In_2791,In_2401);
or U374 (N_374,In_2813,In_2070);
nor U375 (N_375,In_1887,In_505);
nand U376 (N_376,In_1793,In_1959);
nor U377 (N_377,In_1629,In_670);
nand U378 (N_378,In_374,In_1913);
and U379 (N_379,In_2895,In_2573);
xnor U380 (N_380,In_2478,In_1280);
and U381 (N_381,In_2322,In_2066);
nand U382 (N_382,In_1625,In_2580);
nor U383 (N_383,In_2756,In_371);
nor U384 (N_384,In_867,In_2867);
nor U385 (N_385,In_644,In_1568);
xnor U386 (N_386,In_1873,In_2125);
nand U387 (N_387,In_2767,In_2191);
nand U388 (N_388,In_1704,In_857);
or U389 (N_389,In_1948,In_1893);
xor U390 (N_390,In_1454,In_9);
and U391 (N_391,In_2393,In_180);
or U392 (N_392,In_414,In_2738);
nor U393 (N_393,In_2283,In_1545);
or U394 (N_394,In_236,In_1199);
or U395 (N_395,In_2841,In_2261);
or U396 (N_396,In_346,In_1030);
nor U397 (N_397,In_2824,In_508);
nor U398 (N_398,In_2729,In_1074);
nand U399 (N_399,In_1776,In_923);
or U400 (N_400,In_1931,In_347);
xor U401 (N_401,In_2477,In_433);
nor U402 (N_402,In_1845,In_2163);
nor U403 (N_403,In_1323,In_655);
nor U404 (N_404,In_139,In_2921);
or U405 (N_405,In_311,In_695);
nor U406 (N_406,In_291,In_1405);
nor U407 (N_407,In_1097,In_961);
and U408 (N_408,In_2195,In_1050);
and U409 (N_409,In_2018,In_1693);
and U410 (N_410,In_1047,In_2808);
nand U411 (N_411,In_1289,In_1998);
nor U412 (N_412,In_2315,In_303);
nand U413 (N_413,In_1343,In_25);
nand U414 (N_414,In_1539,In_793);
xor U415 (N_415,In_2600,In_2241);
and U416 (N_416,In_380,In_2397);
nand U417 (N_417,In_477,In_1004);
xnor U418 (N_418,In_951,In_851);
nand U419 (N_419,In_2284,In_1034);
nor U420 (N_420,In_1907,In_357);
and U421 (N_421,In_1846,In_1115);
xor U422 (N_422,In_1750,In_2720);
or U423 (N_423,In_1904,In_2875);
xnor U424 (N_424,In_2663,In_2706);
or U425 (N_425,In_1512,In_1497);
or U426 (N_426,In_2760,In_2179);
or U427 (N_427,In_2256,In_1205);
xnor U428 (N_428,In_1270,In_1215);
nor U429 (N_429,In_487,In_2416);
xor U430 (N_430,In_910,In_1526);
and U431 (N_431,In_1855,In_2331);
nor U432 (N_432,In_877,In_1087);
or U433 (N_433,In_165,In_513);
and U434 (N_434,In_2684,In_138);
or U435 (N_435,In_1359,In_2008);
and U436 (N_436,In_800,In_2525);
xor U437 (N_437,In_2116,In_1493);
nand U438 (N_438,In_429,In_515);
and U439 (N_439,In_723,In_2611);
xnor U440 (N_440,In_184,In_637);
or U441 (N_441,In_2126,In_2597);
xor U442 (N_442,In_292,In_2514);
nand U443 (N_443,In_612,In_2451);
and U444 (N_444,In_730,In_1483);
or U445 (N_445,In_948,In_2776);
nand U446 (N_446,In_571,In_1614);
nand U447 (N_447,In_634,In_954);
and U448 (N_448,In_579,In_1434);
or U449 (N_449,In_667,In_1126);
nand U450 (N_450,In_1832,In_1154);
nand U451 (N_451,In_1354,In_517);
or U452 (N_452,In_2249,In_1753);
nor U453 (N_453,In_830,In_499);
xnor U454 (N_454,In_2154,In_757);
nand U455 (N_455,In_2619,In_1548);
nand U456 (N_456,In_1589,In_2081);
and U457 (N_457,In_2272,In_1594);
xor U458 (N_458,In_839,In_1993);
or U459 (N_459,In_1966,In_875);
nand U460 (N_460,In_488,In_558);
or U461 (N_461,In_2977,In_2060);
xor U462 (N_462,In_755,In_1747);
xor U463 (N_463,In_1124,In_243);
and U464 (N_464,In_1346,In_456);
or U465 (N_465,In_2894,In_136);
nand U466 (N_466,In_1277,In_1676);
and U467 (N_467,In_1080,In_1702);
and U468 (N_468,In_548,In_2862);
or U469 (N_469,In_2613,In_2105);
and U470 (N_470,In_2467,In_919);
nor U471 (N_471,In_1394,In_492);
or U472 (N_472,In_461,In_1135);
nor U473 (N_473,In_2242,In_1103);
and U474 (N_474,In_205,In_2226);
nor U475 (N_475,In_1348,In_168);
nand U476 (N_476,In_1475,In_1574);
and U477 (N_477,In_1678,In_539);
xor U478 (N_478,In_1240,In_2035);
and U479 (N_479,In_1583,In_1486);
xor U480 (N_480,In_1414,In_1171);
or U481 (N_481,In_2410,In_965);
nor U482 (N_482,In_1572,In_2996);
xnor U483 (N_483,In_2082,In_2555);
nor U484 (N_484,In_1866,In_1430);
and U485 (N_485,In_945,In_2904);
or U486 (N_486,In_72,In_669);
and U487 (N_487,In_2235,In_2554);
and U488 (N_488,In_1232,In_65);
nand U489 (N_489,In_1889,In_689);
or U490 (N_490,In_747,In_1128);
nor U491 (N_491,In_534,In_1063);
or U492 (N_492,In_17,In_884);
xnor U493 (N_493,In_1968,In_1804);
or U494 (N_494,In_783,In_373);
nand U495 (N_495,In_1677,In_1397);
xor U496 (N_496,In_1737,In_833);
and U497 (N_497,In_2556,In_1311);
xnor U498 (N_498,In_736,In_1670);
xor U499 (N_499,In_1108,In_2537);
or U500 (N_500,In_2225,In_1020);
or U501 (N_501,In_2547,In_39);
xnor U502 (N_502,In_49,In_1878);
nor U503 (N_503,In_792,In_201);
nor U504 (N_504,In_2916,In_1796);
xnor U505 (N_505,In_2944,In_2620);
xnor U506 (N_506,In_2845,In_1132);
or U507 (N_507,In_1275,In_1170);
nand U508 (N_508,In_2957,In_2529);
xor U509 (N_509,In_2084,In_2930);
nand U510 (N_510,In_2749,In_1174);
nor U511 (N_511,In_1723,In_564);
nor U512 (N_512,In_331,In_1109);
xor U513 (N_513,In_1474,In_1383);
nor U514 (N_514,In_1658,In_1935);
xnor U515 (N_515,In_858,In_428);
nand U516 (N_516,In_2142,In_993);
xor U517 (N_517,In_1429,In_1179);
or U518 (N_518,In_2697,In_1656);
and U519 (N_519,In_1898,In_1851);
nor U520 (N_520,In_1918,In_1695);
nor U521 (N_521,In_227,In_1817);
nor U522 (N_522,In_2743,In_408);
xor U523 (N_523,In_1144,In_1672);
or U524 (N_524,In_29,In_481);
xor U525 (N_525,In_577,In_1217);
nor U526 (N_526,In_404,In_2608);
and U527 (N_527,In_653,In_151);
xnor U528 (N_528,In_2127,In_1616);
xor U529 (N_529,In_1624,In_860);
xnor U530 (N_530,In_288,In_2750);
nand U531 (N_531,In_204,In_1426);
xnor U532 (N_532,In_738,In_2678);
nor U533 (N_533,In_559,In_2486);
or U534 (N_534,In_2040,In_1911);
and U535 (N_535,In_1740,In_827);
nand U536 (N_536,In_1622,In_1112);
nand U537 (N_537,In_1758,In_562);
nor U538 (N_538,In_1376,In_2251);
xnor U539 (N_539,In_2981,In_2375);
nand U540 (N_540,In_1511,In_1334);
xnor U541 (N_541,In_1304,In_2072);
nor U542 (N_542,In_285,In_2491);
and U543 (N_543,In_310,In_2797);
nor U544 (N_544,In_1041,In_2215);
or U545 (N_545,In_146,In_1905);
or U546 (N_546,In_1084,In_494);
and U547 (N_547,In_740,In_2281);
and U548 (N_548,In_471,In_1023);
xor U549 (N_549,In_248,In_409);
xnor U550 (N_550,In_985,In_150);
or U551 (N_551,In_962,In_2023);
nand U552 (N_552,In_2987,In_1322);
and U553 (N_553,In_2886,In_163);
and U554 (N_554,In_2816,In_1774);
and U555 (N_555,In_1026,In_2638);
and U556 (N_556,In_543,In_524);
or U557 (N_557,In_1012,In_1735);
xnor U558 (N_558,In_2498,In_1547);
or U559 (N_559,In_1150,In_231);
and U560 (N_560,In_2095,In_1715);
and U561 (N_561,In_2098,In_592);
xor U562 (N_562,In_698,In_852);
nand U563 (N_563,In_267,In_2711);
or U564 (N_564,In_2923,In_1130);
xor U565 (N_565,In_211,In_1193);
nor U566 (N_566,In_1830,In_1362);
and U567 (N_567,In_1139,In_2801);
nand U568 (N_568,In_1561,In_1230);
nor U569 (N_569,In_904,In_2990);
and U570 (N_570,In_2884,In_1975);
nor U571 (N_571,In_102,In_2041);
nand U572 (N_572,In_977,In_1833);
or U573 (N_573,In_1582,In_664);
or U574 (N_574,In_117,In_1569);
nand U575 (N_575,In_711,In_61);
and U576 (N_576,In_1291,In_2255);
and U577 (N_577,In_1571,In_1843);
and U578 (N_578,In_1992,In_1223);
nand U579 (N_579,In_2519,In_619);
or U580 (N_580,In_1102,In_2939);
xnor U581 (N_581,In_502,In_1809);
nor U582 (N_582,In_2463,In_2878);
or U583 (N_583,In_2454,In_1599);
xor U584 (N_584,In_1769,In_2843);
or U585 (N_585,In_802,In_2764);
nor U586 (N_586,In_2216,In_2833);
and U587 (N_587,In_372,In_2995);
nor U588 (N_588,In_2059,In_1555);
or U589 (N_589,In_2891,In_1757);
nand U590 (N_590,In_855,In_42);
nand U591 (N_591,In_2521,In_1039);
xor U592 (N_592,In_943,In_889);
xor U593 (N_593,In_2424,In_2926);
or U594 (N_594,In_2811,In_2819);
nand U595 (N_595,In_2184,In_308);
xnor U596 (N_596,In_1558,In_282);
nand U597 (N_597,In_2540,In_912);
nand U598 (N_598,In_2748,In_294);
and U599 (N_599,In_1732,In_396);
nand U600 (N_600,In_2636,In_1105);
or U601 (N_601,In_2605,In_2709);
nand U602 (N_602,In_2052,In_2259);
xor U603 (N_603,In_1559,In_1906);
and U604 (N_604,In_2360,In_2539);
or U605 (N_605,In_1399,In_570);
nor U606 (N_606,In_1527,In_1167);
or U607 (N_607,In_734,In_2309);
xor U608 (N_608,In_2979,In_2953);
nand U609 (N_609,In_1575,In_222);
and U610 (N_610,In_2488,In_2899);
nor U611 (N_611,In_2802,In_2379);
and U612 (N_612,In_324,In_2848);
nand U613 (N_613,In_881,In_1263);
nand U614 (N_614,In_587,In_630);
xnor U615 (N_615,In_1532,In_2724);
and U616 (N_616,In_1164,In_2726);
nor U617 (N_617,In_1903,In_521);
or U618 (N_618,In_266,In_32);
and U619 (N_619,In_2635,In_365);
nand U620 (N_620,In_172,In_62);
nor U621 (N_621,In_2464,In_1507);
xnor U622 (N_622,In_772,In_2361);
nor U623 (N_623,In_424,In_687);
nor U624 (N_624,In_2731,In_1412);
nand U625 (N_625,In_263,In_467);
nor U626 (N_626,In_1011,In_2274);
xnor U627 (N_627,In_510,In_2370);
xor U628 (N_628,In_2849,In_1615);
or U629 (N_629,In_2316,In_1533);
nor U630 (N_630,In_1324,In_195);
nand U631 (N_631,In_850,In_2599);
and U632 (N_632,In_547,In_1553);
and U633 (N_633,In_1924,In_2960);
nand U634 (N_634,In_1473,In_911);
nor U635 (N_635,In_1365,In_1770);
nand U636 (N_636,In_2069,In_2178);
nor U637 (N_637,In_649,In_298);
xor U638 (N_638,In_1222,In_964);
and U639 (N_639,In_1256,In_353);
nand U640 (N_640,In_821,In_871);
and U641 (N_641,In_2439,In_971);
nand U642 (N_642,In_2270,In_2700);
xor U643 (N_643,In_2631,In_1570);
or U644 (N_644,In_18,In_2461);
or U645 (N_645,In_2263,In_2146);
xor U646 (N_646,In_931,In_835);
or U647 (N_647,In_2897,In_2918);
or U648 (N_648,In_99,In_1890);
nor U649 (N_649,In_2299,In_1659);
and U650 (N_650,In_1564,In_2662);
or U651 (N_651,In_672,In_2582);
or U652 (N_652,In_2208,In_532);
xor U653 (N_653,In_1880,In_2087);
and U654 (N_654,In_2545,In_22);
xnor U655 (N_655,In_2376,In_495);
nor U656 (N_656,In_2173,In_1264);
or U657 (N_657,In_2666,In_2011);
and U658 (N_658,In_2171,In_493);
or U659 (N_659,In_485,In_842);
xnor U660 (N_660,In_1247,In_1303);
xor U661 (N_661,In_1211,In_1366);
nor U662 (N_662,In_879,In_1456);
nand U663 (N_663,In_2900,In_140);
or U664 (N_664,In_778,In_966);
or U665 (N_665,In_2495,In_2639);
or U666 (N_666,In_4,In_1524);
or U667 (N_667,In_2077,In_2685);
and U668 (N_668,In_2085,In_384);
and U669 (N_669,In_2502,In_2524);
nor U670 (N_670,In_682,In_2258);
xnor U671 (N_671,In_2389,In_2992);
xnor U672 (N_672,In_2139,In_2356);
xnor U673 (N_673,In_838,In_1915);
xor U674 (N_674,In_2288,In_2948);
nor U675 (N_675,In_141,In_900);
xnor U676 (N_676,In_1035,In_1368);
nand U677 (N_677,In_321,In_213);
and U678 (N_678,In_1902,In_742);
or U679 (N_679,In_665,In_990);
nand U680 (N_680,In_1861,In_728);
nand U681 (N_681,In_394,In_415);
or U682 (N_682,In_2305,In_2387);
nand U683 (N_683,In_100,In_2920);
and U684 (N_684,In_837,In_566);
xor U685 (N_685,In_927,In_2736);
xor U686 (N_686,In_1446,In_639);
xnor U687 (N_687,In_1560,In_2857);
and U688 (N_688,In_2966,In_1418);
xor U689 (N_689,In_2815,In_1272);
xor U690 (N_690,In_1113,In_1841);
nand U691 (N_691,In_71,In_2174);
or U692 (N_692,In_1203,In_2435);
xnor U693 (N_693,In_2719,In_1516);
and U694 (N_694,In_2388,In_2277);
and U695 (N_695,In_1077,In_1663);
nand U696 (N_696,In_1557,In_2450);
nand U697 (N_697,In_674,In_2936);
or U698 (N_698,In_1954,In_1198);
nand U699 (N_699,In_2985,In_2943);
nor U700 (N_700,In_2051,In_503);
xnor U701 (N_701,In_2607,In_2565);
and U702 (N_702,In_318,In_462);
xor U703 (N_703,In_2189,In_2165);
nand U704 (N_704,In_2020,In_317);
xnor U705 (N_705,In_1848,In_1922);
nand U706 (N_706,In_1513,In_430);
or U707 (N_707,In_1160,In_878);
or U708 (N_708,In_1494,In_1751);
nor U709 (N_709,In_2820,In_334);
xor U710 (N_710,In_2686,In_339);
nand U711 (N_711,In_608,In_1243);
and U712 (N_712,In_601,In_729);
xnor U713 (N_713,In_1435,In_2407);
and U714 (N_714,In_1739,In_2788);
nand U715 (N_715,In_2557,In_1891);
or U716 (N_716,In_1760,In_516);
xor U717 (N_717,In_115,In_1999);
and U718 (N_718,In_606,In_1266);
nand U719 (N_719,In_2286,In_685);
nand U720 (N_720,In_2928,In_1587);
or U721 (N_721,In_2646,In_840);
nand U722 (N_722,In_2534,In_2522);
nor U723 (N_723,In_216,In_1674);
nor U724 (N_724,In_1567,In_2583);
nand U725 (N_725,In_2075,In_550);
or U726 (N_726,In_2947,In_2243);
or U727 (N_727,In_93,In_2606);
xor U728 (N_728,In_443,In_2584);
and U729 (N_729,In_1802,In_2230);
and U730 (N_730,In_2428,In_2119);
nor U731 (N_731,In_960,In_873);
or U732 (N_732,In_134,In_1236);
xor U733 (N_733,In_932,In_1813);
xnor U734 (N_734,In_1595,In_1505);
nand U735 (N_735,In_2295,In_2199);
or U736 (N_736,In_2805,In_182);
nand U737 (N_737,In_2043,In_1721);
nand U738 (N_738,In_2517,In_240);
xor U739 (N_739,In_57,In_319);
or U740 (N_740,In_2100,In_1213);
nand U741 (N_741,In_2250,In_2757);
and U742 (N_742,In_2238,In_1462);
or U743 (N_743,In_2512,In_1342);
or U744 (N_744,In_1610,In_190);
nand U745 (N_745,In_2507,In_2721);
xor U746 (N_746,In_2542,In_2352);
xnor U747 (N_747,In_1578,In_2562);
nand U748 (N_748,In_2209,In_814);
and U749 (N_749,In_2033,In_2905);
nand U750 (N_750,In_279,In_81);
nand U751 (N_751,In_2838,In_2394);
xor U752 (N_752,In_725,In_1186);
and U753 (N_753,In_2028,In_2504);
nor U754 (N_754,In_2550,In_845);
nand U755 (N_755,In_2798,In_1716);
nor U756 (N_756,In_739,In_1358);
nor U757 (N_757,In_104,In_1053);
or U758 (N_758,In_1106,In_819);
and U759 (N_759,In_765,In_431);
nand U760 (N_760,In_1482,In_1638);
and U761 (N_761,In_831,In_398);
nand U762 (N_762,In_1140,In_230);
and U763 (N_763,In_716,In_1088);
nand U764 (N_764,In_2437,In_1612);
xor U765 (N_765,In_386,In_1472);
nor U766 (N_766,In_2858,In_2496);
xor U767 (N_767,In_869,In_123);
or U768 (N_768,In_2642,In_2641);
and U769 (N_769,In_453,In_1008);
nor U770 (N_770,In_2458,In_896);
nand U771 (N_771,In_972,In_2922);
xnor U772 (N_772,In_1756,In_2956);
and U773 (N_773,In_627,In_1632);
or U774 (N_774,In_1945,In_2320);
and U775 (N_775,In_121,In_2846);
nand U776 (N_776,In_2732,In_1777);
xnor U777 (N_777,In_1986,In_97);
xor U778 (N_778,In_1148,In_2715);
or U779 (N_779,In_1811,In_479);
nand U780 (N_780,In_994,In_544);
nand U781 (N_781,In_306,In_1605);
xor U782 (N_782,In_2298,In_420);
or U783 (N_783,In_1504,In_1292);
nor U784 (N_784,In_2112,In_1510);
xor U785 (N_785,In_768,In_610);
nor U786 (N_786,In_1554,In_2362);
or U787 (N_787,In_785,In_207);
and U788 (N_788,In_1593,In_191);
nor U789 (N_789,In_1908,In_1731);
nor U790 (N_790,In_1815,In_2564);
or U791 (N_791,In_632,In_2367);
and U792 (N_792,In_2363,In_1590);
nand U793 (N_793,In_2239,In_2076);
nand U794 (N_794,In_1847,In_2418);
nor U795 (N_795,In_272,In_1712);
xor U796 (N_796,In_1862,In_144);
nor U797 (N_797,In_753,In_641);
nand U798 (N_798,In_12,In_1413);
nand U799 (N_799,In_1951,In_159);
xnor U800 (N_800,In_2777,In_1576);
nor U801 (N_801,In_2854,In_626);
or U802 (N_802,In_166,In_2433);
nor U803 (N_803,In_2002,In_1444);
nor U804 (N_804,In_699,In_1237);
nand U805 (N_805,In_913,In_358);
or U806 (N_806,In_939,In_2476);
or U807 (N_807,In_2941,In_7);
nor U808 (N_808,In_1079,In_2092);
xnor U809 (N_809,In_1892,In_995);
and U810 (N_810,In_1259,In_1173);
and U811 (N_811,In_1302,In_1488);
and U812 (N_812,In_2759,In_369);
or U813 (N_813,In_2459,In_2104);
xor U814 (N_814,In_403,In_1685);
or U815 (N_815,In_2739,In_565);
and U816 (N_816,In_1329,In_2460);
xnor U817 (N_817,In_1119,In_1379);
or U818 (N_818,In_1871,In_1950);
xor U819 (N_819,In_1086,In_2772);
and U820 (N_820,In_1364,In_2061);
and U821 (N_821,In_998,In_2210);
xor U822 (N_822,In_2017,In_160);
and U823 (N_823,In_1214,In_1729);
nor U824 (N_824,In_762,In_169);
and U825 (N_825,In_76,In_2447);
nand U826 (N_826,In_2792,In_452);
xnor U827 (N_827,In_822,In_552);
or U828 (N_828,In_2863,In_1643);
nor U829 (N_829,In_2371,In_2378);
xnor U830 (N_830,In_2789,In_2382);
and U831 (N_831,In_2594,In_69);
or U832 (N_832,In_1204,In_1517);
xor U833 (N_833,In_1461,In_254);
or U834 (N_834,In_2485,In_2019);
nor U835 (N_835,In_754,In_527);
nor U836 (N_836,In_1228,In_2561);
nor U837 (N_837,In_170,In_2999);
nor U838 (N_838,In_1151,In_1995);
or U839 (N_839,In_1956,In_1772);
xor U840 (N_840,In_185,In_2654);
and U841 (N_841,In_2392,In_2187);
nor U842 (N_842,In_1453,In_2001);
and U843 (N_843,In_1814,In_2645);
or U844 (N_844,In_2050,In_1727);
nand U845 (N_845,In_1172,In_2558);
or U846 (N_846,In_2592,In_265);
nand U847 (N_847,In_327,In_663);
nand U848 (N_848,In_2218,In_2530);
and U849 (N_849,In_2183,In_824);
or U850 (N_850,In_605,In_2157);
or U851 (N_851,In_2727,In_675);
xor U852 (N_852,In_1642,In_1297);
or U853 (N_853,In_74,In_717);
nand U854 (N_854,In_623,In_2300);
or U855 (N_855,In_2058,In_863);
xor U856 (N_856,In_1495,In_454);
nand U857 (N_857,In_2343,In_1681);
nand U858 (N_858,In_2952,In_2448);
and U859 (N_859,In_2358,In_2503);
xnor U860 (N_860,In_1920,In_1645);
nor U861 (N_861,In_1345,In_229);
or U862 (N_862,In_1175,In_2566);
and U863 (N_863,In_2228,In_1627);
xnor U864 (N_864,In_789,In_85);
nor U865 (N_865,In_959,In_1534);
nor U866 (N_866,In_2099,In_385);
or U867 (N_867,In_412,In_90);
and U868 (N_868,In_2267,In_2834);
nor U869 (N_869,In_2482,In_1870);
and U870 (N_870,In_2337,In_1360);
xor U871 (N_871,In_648,In_519);
and U872 (N_872,In_2761,In_531);
or U873 (N_873,In_89,In_1344);
nand U874 (N_874,In_2141,In_2014);
xor U875 (N_875,In_953,In_2629);
or U876 (N_876,In_1609,In_1480);
nand U877 (N_877,In_2289,In_2538);
and U878 (N_878,In_390,In_1282);
xor U879 (N_879,In_107,In_1404);
and U880 (N_880,In_834,In_1273);
xor U881 (N_881,In_46,In_290);
xor U882 (N_882,In_1449,In_628);
xor U883 (N_883,In_1708,In_1054);
or U884 (N_884,In_2167,In_1644);
nand U885 (N_885,In_2441,In_2333);
or U886 (N_886,In_1278,In_1717);
or U887 (N_887,In_2086,In_929);
and U888 (N_888,In_1015,In_158);
nor U889 (N_889,In_35,In_178);
nor U890 (N_890,In_164,In_1588);
or U891 (N_891,In_2233,In_1738);
nand U892 (N_892,In_2782,In_2443);
or U893 (N_893,In_1556,In_1017);
nand U894 (N_894,In_1221,In_417);
xnor U895 (N_895,In_1518,In_2954);
and U896 (N_896,In_530,In_1967);
nand U897 (N_897,In_475,In_872);
or U898 (N_898,In_2176,In_901);
or U899 (N_899,In_1900,In_1049);
xor U900 (N_900,In_1573,In_590);
or U901 (N_901,In_595,In_1374);
nor U902 (N_902,In_1623,In_483);
nand U903 (N_903,In_2536,In_2552);
and U904 (N_904,In_37,In_51);
nand U905 (N_905,In_2493,In_2659);
nand U906 (N_906,In_555,In_1422);
or U907 (N_907,In_980,In_2168);
and U908 (N_908,In_1092,In_2971);
or U909 (N_909,In_522,In_349);
xor U910 (N_910,In_598,In_1081);
nor U911 (N_911,In_1536,In_2147);
xnor U912 (N_912,In_1881,In_322);
and U913 (N_913,In_6,In_448);
and U914 (N_914,In_1943,In_399);
nand U915 (N_915,In_2710,In_276);
nand U916 (N_916,In_2609,In_155);
nor U917 (N_917,In_2997,In_34);
nand U918 (N_918,In_2672,In_2962);
or U919 (N_919,In_2541,In_225);
and U920 (N_920,In_59,In_101);
nor U921 (N_921,In_1072,In_2062);
nor U922 (N_922,In_2364,In_1831);
nor U923 (N_923,In_1202,In_1427);
xnor U924 (N_924,In_1821,In_124);
nor U925 (N_925,In_1991,In_1604);
or U926 (N_926,In_743,In_1208);
xnor U927 (N_927,In_2864,In_2940);
and U928 (N_928,In_1025,In_1458);
nor U929 (N_929,In_2590,In_2089);
nand U930 (N_930,In_176,In_2010);
nor U931 (N_931,In_1401,In_88);
nand U932 (N_932,In_2237,In_391);
and U933 (N_933,In_2359,In_221);
nor U934 (N_934,In_1,In_2500);
xnor U935 (N_935,In_2432,In_2818);
xor U936 (N_936,In_694,In_903);
nor U937 (N_937,In_1836,In_2151);
nand U938 (N_938,In_2633,In_1471);
xor U939 (N_939,In_2889,In_238);
and U940 (N_940,In_797,In_167);
or U941 (N_941,In_1932,In_226);
xnor U942 (N_942,In_94,In_2314);
nor U943 (N_943,In_666,In_1633);
nor U944 (N_944,In_1988,In_907);
nor U945 (N_945,In_2490,In_1585);
or U946 (N_946,In_2130,In_1188);
xor U947 (N_947,In_2883,In_2655);
xor U948 (N_948,In_2880,In_302);
nand U949 (N_949,In_2551,In_1566);
xnor U950 (N_950,In_312,In_849);
nand U951 (N_951,In_1029,In_490);
xor U952 (N_952,In_591,In_2380);
or U953 (N_953,In_2134,In_1242);
xor U954 (N_954,In_659,In_2122);
xor U955 (N_955,In_853,In_2440);
xnor U956 (N_956,In_2471,In_64);
nor U957 (N_957,In_77,In_217);
nand U958 (N_958,In_1790,In_1395);
nand U959 (N_959,In_244,In_1856);
nand U960 (N_960,In_988,In_890);
and U961 (N_961,In_940,In_767);
and U962 (N_962,In_2621,In_2282);
nand U963 (N_963,In_255,In_2664);
xor U964 (N_964,In_2455,In_749);
nand U965 (N_965,In_1919,In_787);
nor U966 (N_966,In_2264,In_1598);
xnor U967 (N_967,In_2740,In_1549);
or U968 (N_968,In_1613,In_796);
and U969 (N_969,In_1467,In_2647);
xor U970 (N_970,In_1535,In_2229);
nand U971 (N_971,In_572,In_1768);
or U972 (N_972,In_2198,In_1129);
and U973 (N_973,In_2657,In_1523);
nand U974 (N_974,In_2821,In_1826);
xnor U975 (N_975,In_473,In_2354);
and U976 (N_976,In_1382,In_2007);
and U977 (N_977,In_1315,In_1979);
nor U978 (N_978,In_898,In_1367);
xor U979 (N_979,In_1994,In_1155);
nor U980 (N_980,In_1933,In_1094);
or U981 (N_981,In_1296,In_378);
nand U982 (N_982,In_784,In_1392);
and U983 (N_983,In_1962,In_1894);
nor U984 (N_984,In_874,In_54);
and U985 (N_985,In_2325,In_616);
nor U986 (N_986,In_735,In_1816);
or U987 (N_987,In_199,In_110);
nor U988 (N_988,In_1958,In_975);
xnor U989 (N_989,In_696,In_2489);
nand U990 (N_990,In_1784,In_1423);
nand U991 (N_991,In_129,In_1441);
or U992 (N_992,In_2998,In_246);
and U993 (N_993,In_1818,In_1246);
and U994 (N_994,In_1300,In_1262);
nor U995 (N_995,In_202,In_1746);
nand U996 (N_996,In_1971,In_2689);
or U997 (N_997,In_1372,In_469);
and U998 (N_998,In_1872,In_2350);
nand U999 (N_999,In_1460,In_647);
nand U1000 (N_1000,In_541,In_476);
nor U1001 (N_1001,In_377,In_1867);
nor U1002 (N_1002,In_1436,In_1168);
and U1003 (N_1003,In_991,In_2470);
xnor U1004 (N_1004,In_2038,In_1854);
nor U1005 (N_1005,In_53,In_941);
nand U1006 (N_1006,In_2196,In_602);
nor U1007 (N_1007,In_2400,In_2223);
xor U1008 (N_1008,In_2345,In_596);
nand U1009 (N_1009,In_1662,In_1284);
nor U1010 (N_1010,In_697,In_2351);
nor U1011 (N_1011,In_2532,In_105);
nor U1012 (N_1012,In_1005,In_2053);
or U1013 (N_1013,In_2431,In_1032);
and U1014 (N_1014,In_657,In_816);
nor U1015 (N_1015,In_148,In_401);
nand U1016 (N_1016,In_2717,In_2253);
and U1017 (N_1017,In_935,In_526);
nor U1018 (N_1018,In_2786,In_712);
nand U1019 (N_1019,In_2585,In_92);
and U1020 (N_1020,In_2111,In_2699);
or U1021 (N_1021,In_26,In_2924);
xor U1022 (N_1022,In_234,In_1133);
xnor U1023 (N_1023,In_967,In_693);
and U1024 (N_1024,In_44,In_337);
xor U1025 (N_1025,In_79,In_1229);
and U1026 (N_1026,In_1795,In_1765);
xnor U1027 (N_1027,In_427,In_1985);
xnor U1028 (N_1028,In_2399,In_426);
or U1029 (N_1029,In_383,In_986);
xor U1030 (N_1030,In_1983,In_1057);
nor U1031 (N_1031,In_894,In_2148);
and U1032 (N_1032,In_2327,In_1783);
xnor U1033 (N_1033,In_2860,In_1626);
or U1034 (N_1034,In_1274,In_1806);
and U1035 (N_1035,In_198,In_1489);
or U1036 (N_1036,In_557,In_1692);
nor U1037 (N_1037,In_1470,In_343);
and U1038 (N_1038,In_588,In_1299);
nand U1039 (N_1039,In_2917,In_1388);
xnor U1040 (N_1040,In_2329,In_2869);
or U1041 (N_1041,In_1352,In_1787);
nand U1042 (N_1042,In_1934,In_2934);
and U1043 (N_1043,In_242,In_2279);
or U1044 (N_1044,In_2725,In_750);
xnor U1045 (N_1045,In_2219,In_1220);
or U1046 (N_1046,In_963,In_2234);
nor U1047 (N_1047,In_48,In_2877);
xor U1048 (N_1048,In_618,In_439);
xor U1049 (N_1049,In_908,In_2457);
nand U1050 (N_1050,In_1347,In_599);
or U1051 (N_1051,In_1720,In_1093);
and U1052 (N_1052,In_680,In_2828);
nand U1053 (N_1053,In_1225,In_340);
nor U1054 (N_1054,In_1603,In_506);
xor U1055 (N_1055,In_2598,In_2518);
and U1056 (N_1056,In_425,In_1540);
nor U1057 (N_1057,In_2694,In_1024);
or U1058 (N_1058,In_466,In_2704);
nand U1059 (N_1059,In_1528,In_2374);
or U1060 (N_1060,In_2653,In_1586);
xor U1061 (N_1061,In_583,In_1159);
or U1062 (N_1062,In_120,In_2000);
nor U1063 (N_1063,In_1675,In_1439);
and U1064 (N_1064,In_1852,In_307);
or U1065 (N_1065,In_892,In_1786);
nor U1066 (N_1066,In_2419,In_525);
xnor U1067 (N_1067,In_2911,In_275);
nor U1068 (N_1068,In_1858,In_2481);
nand U1069 (N_1069,In_360,In_2986);
nand U1070 (N_1070,In_748,In_189);
nand U1071 (N_1071,In_434,In_1062);
nor U1072 (N_1072,In_2588,In_2113);
nand U1073 (N_1073,In_256,In_1378);
nand U1074 (N_1074,In_2803,In_681);
xnor U1075 (N_1075,In_876,In_351);
xor U1076 (N_1076,In_2308,In_540);
xnor U1077 (N_1077,In_2406,In_2135);
and U1078 (N_1078,In_1409,In_1195);
and U1079 (N_1079,In_1883,In_2221);
nor U1080 (N_1080,In_1166,In_10);
and U1081 (N_1081,In_11,In_2974);
nor U1082 (N_1082,In_316,In_722);
xor U1083 (N_1083,In_1251,In_2593);
or U1084 (N_1084,In_1056,In_1269);
nor U1085 (N_1085,In_2603,In_2429);
xor U1086 (N_1086,In_2338,In_2840);
or U1087 (N_1087,In_1936,In_332);
and U1088 (N_1088,In_2254,In_2164);
nor U1089 (N_1089,In_2475,In_436);
or U1090 (N_1090,In_2702,In_395);
and U1091 (N_1091,In_1319,In_2859);
nand U1092 (N_1092,In_286,In_314);
nand U1093 (N_1093,In_2988,In_2445);
nor U1094 (N_1094,In_593,In_330);
nor U1095 (N_1095,In_2326,In_2668);
xor U1096 (N_1096,In_2391,In_974);
nand U1097 (N_1097,In_1688,In_536);
nand U1098 (N_1098,In_1810,In_883);
xor U1099 (N_1099,In_1111,In_2136);
nand U1100 (N_1100,In_1333,In_804);
and U1101 (N_1101,In_2652,In_1307);
nand U1102 (N_1102,In_2373,In_2901);
or U1103 (N_1103,In_629,In_2310);
xor U1104 (N_1104,In_145,In_497);
and U1105 (N_1105,In_1641,In_1468);
nor U1106 (N_1106,In_984,In_224);
and U1107 (N_1107,In_1718,In_2581);
and U1108 (N_1108,In_2290,In_578);
nor U1109 (N_1109,In_1165,In_702);
or U1110 (N_1110,In_2887,In_2027);
and U1111 (N_1111,In_2034,In_1698);
or U1112 (N_1112,In_1355,In_1875);
or U1113 (N_1113,In_1541,In_549);
and U1114 (N_1114,In_359,In_2120);
and U1115 (N_1115,In_636,In_1313);
or U1116 (N_1116,In_726,In_268);
nor U1117 (N_1117,In_2778,In_2827);
nand U1118 (N_1118,In_397,In_2381);
or U1119 (N_1119,In_1581,In_1782);
and U1120 (N_1120,In_2395,In_556);
nor U1121 (N_1121,In_2679,In_1001);
nand U1122 (N_1122,In_1061,In_1520);
xnor U1123 (N_1123,In_2933,In_1252);
nor U1124 (N_1124,In_367,In_976);
and U1125 (N_1125,In_214,In_586);
xor U1126 (N_1126,In_1390,In_1070);
nor U1127 (N_1127,In_2427,In_2499);
and U1128 (N_1128,In_646,In_1884);
or U1129 (N_1129,In_87,In_1789);
nand U1130 (N_1130,In_700,In_1492);
or U1131 (N_1131,In_1921,In_2734);
or U1132 (N_1132,In_1696,In_917);
or U1133 (N_1133,In_2444,In_2676);
and U1134 (N_1134,In_1162,In_2906);
nor U1135 (N_1135,In_535,In_2677);
and U1136 (N_1136,In_2342,In_1363);
or U1137 (N_1137,In_2319,In_368);
nand U1138 (N_1138,In_2688,In_2083);
xor U1139 (N_1139,In_2473,In_1419);
and U1140 (N_1140,In_1068,In_2737);
and U1141 (N_1141,In_1710,In_2078);
nor U1142 (N_1142,In_2006,In_393);
or U1143 (N_1143,In_2276,In_126);
nand U1144 (N_1144,In_2438,In_1521);
xor U1145 (N_1145,In_2980,In_1386);
nor U1146 (N_1146,In_1514,In_826);
nand U1147 (N_1147,In_2929,In_2616);
nor U1148 (N_1148,In_2220,In_2102);
nor U1149 (N_1149,In_703,In_1686);
and U1150 (N_1150,In_2149,In_2822);
xor U1151 (N_1151,In_1551,In_1410);
and U1152 (N_1152,In_2,In_1027);
nand U1153 (N_1153,In_733,In_1350);
nand U1154 (N_1154,In_50,In_1785);
and U1155 (N_1155,In_2064,In_1960);
nor U1156 (N_1156,In_1709,In_766);
nand U1157 (N_1157,In_957,In_2829);
and U1158 (N_1158,In_250,In_1192);
or U1159 (N_1159,In_2426,In_2306);
nor U1160 (N_1160,In_2625,In_2090);
xor U1161 (N_1161,In_2409,In_2404);
and U1162 (N_1162,In_2280,In_684);
nor U1163 (N_1163,In_2968,In_2436);
xor U1164 (N_1164,In_933,In_1544);
or U1165 (N_1165,In_2574,In_2303);
xor U1166 (N_1166,In_323,In_1771);
xnor U1167 (N_1167,In_2589,In_2096);
nand U1168 (N_1168,In_2348,In_2991);
nand U1169 (N_1169,In_856,In_2825);
nand U1170 (N_1170,In_1691,In_1018);
nand U1171 (N_1171,In_914,In_2398);
nand U1172 (N_1172,In_1048,In_1705);
nor U1173 (N_1173,In_465,In_2453);
xor U1174 (N_1174,In_441,In_613);
xor U1175 (N_1175,In_868,In_1797);
or U1176 (N_1176,In_573,In_2835);
xnor U1177 (N_1177,In_1882,In_2244);
and U1178 (N_1178,In_710,In_1874);
xor U1179 (N_1179,In_2511,In_721);
and U1180 (N_1180,In_2946,In_73);
or U1181 (N_1181,In_643,In_2733);
nand U1182 (N_1182,In_143,In_277);
nand U1183 (N_1183,In_2769,In_2548);
nor U1184 (N_1184,In_2945,In_70);
xnor U1185 (N_1185,In_295,In_1187);
nor U1186 (N_1186,In_2047,In_774);
nand U1187 (N_1187,In_1660,In_1408);
or U1188 (N_1188,In_2796,In_1479);
nand U1189 (N_1189,In_1666,In_1621);
nor U1190 (N_1190,In_661,In_1651);
nor U1191 (N_1191,In_2094,In_326);
or U1192 (N_1192,In_654,In_624);
nand U1193 (N_1193,In_422,In_106);
nor U1194 (N_1194,In_1101,In_375);
or U1195 (N_1195,In_758,In_2919);
nand U1196 (N_1196,In_2696,In_1689);
nor U1197 (N_1197,In_2804,In_2771);
or U1198 (N_1198,In_1901,In_690);
xnor U1199 (N_1199,In_2644,In_1245);
and U1200 (N_1200,In_1989,In_1051);
nor U1201 (N_1201,In_770,In_1964);
nand U1202 (N_1202,In_2967,In_2673);
or U1203 (N_1203,In_622,In_2158);
nor U1204 (N_1204,In_2753,In_2914);
nand U1205 (N_1205,In_381,In_2879);
or U1206 (N_1206,In_958,In_370);
and U1207 (N_1207,In_2770,In_1445);
nor U1208 (N_1208,In_2412,In_14);
or U1209 (N_1209,In_2844,In_1596);
and U1210 (N_1210,In_472,In_1531);
nor U1211 (N_1211,In_1114,In_1794);
nor U1212 (N_1212,In_269,In_2117);
xnor U1213 (N_1213,In_724,In_2950);
nand U1214 (N_1214,In_2145,In_2708);
and U1215 (N_1215,In_2036,In_446);
or U1216 (N_1216,In_2872,In_720);
nor U1217 (N_1217,In_2882,In_363);
nand U1218 (N_1218,In_2172,In_554);
nor U1219 (N_1219,In_1970,In_480);
and U1220 (N_1220,In_111,In_309);
and U1221 (N_1221,In_2508,In_2983);
and U1222 (N_1222,In_937,In_2975);
xnor U1223 (N_1223,In_1984,In_1371);
nand U1224 (N_1224,In_2669,In_2505);
nand U1225 (N_1225,In_671,In_2260);
nand U1226 (N_1226,In_786,In_719);
and U1227 (N_1227,In_1349,In_457);
xnor U1228 (N_1228,In_2965,In_987);
nor U1229 (N_1229,In_1923,In_752);
xor U1230 (N_1230,In_1736,In_2301);
nor U1231 (N_1231,In_328,In_297);
or U1232 (N_1232,In_1007,In_2137);
xor U1233 (N_1233,In_2311,In_1021);
xnor U1234 (N_1234,In_114,In_829);
or U1235 (N_1235,In_1281,In_1503);
nand U1236 (N_1236,In_1145,In_438);
or U1237 (N_1237,In_1216,In_41);
nand U1238 (N_1238,In_1699,In_1431);
nor U1239 (N_1239,In_2866,In_859);
xnor U1240 (N_1240,In_16,In_52);
nor U1241 (N_1241,In_173,In_1037);
nor U1242 (N_1242,In_823,In_1648);
or U1243 (N_1243,In_500,In_1542);
nand U1244 (N_1244,In_1306,In_1863);
xnor U1245 (N_1245,In_1261,In_1639);
and U1246 (N_1246,In_801,In_2175);
or U1247 (N_1247,In_1822,In_611);
nor U1248 (N_1248,In_2177,In_2571);
and U1249 (N_1249,In_486,In_67);
and U1250 (N_1250,In_866,In_271);
xor U1251 (N_1251,In_1176,In_338);
and U1252 (N_1252,In_1879,In_1377);
nor U1253 (N_1253,In_1271,In_1925);
nand U1254 (N_1254,In_1136,In_447);
nand U1255 (N_1255,In_2958,In_1707);
nand U1256 (N_1256,In_1212,In_1286);
nand U1257 (N_1257,In_484,In_745);
nand U1258 (N_1258,In_2963,In_2577);
nand U1259 (N_1259,In_844,In_432);
or U1260 (N_1260,In_1842,In_2442);
and U1261 (N_1261,In_1036,In_2372);
nand U1262 (N_1262,In_1714,In_1201);
nand U1263 (N_1263,In_2591,In_389);
nor U1264 (N_1264,In_2716,In_2935);
nor U1265 (N_1265,In_1091,In_633);
xnor U1266 (N_1266,In_1652,In_2506);
and U1267 (N_1267,In_259,In_2206);
nor U1268 (N_1268,In_2186,In_1973);
xnor U1269 (N_1269,In_1909,In_2533);
nor U1270 (N_1270,In_247,In_2304);
and U1271 (N_1271,In_2193,In_1499);
nand U1272 (N_1272,In_2287,In_1055);
or U1273 (N_1273,In_862,In_660);
or U1274 (N_1274,In_1177,In_1597);
nand U1275 (N_1275,In_1631,In_1801);
or U1276 (N_1276,In_2913,In_2170);
and U1277 (N_1277,In_1869,In_20);
nor U1278 (N_1278,In_507,In_2114);
nand U1279 (N_1279,In_1142,In_21);
nor U1280 (N_1280,In_2643,In_2323);
or U1281 (N_1281,In_2806,In_2194);
or U1282 (N_1282,In_946,In_1384);
and U1283 (N_1283,In_2927,In_1224);
nor U1284 (N_1284,In_2474,In_1308);
xnor U1285 (N_1285,In_1978,In_2425);
and U1286 (N_1286,In_2516,In_2048);
nand U1287 (N_1287,In_36,In_2368);
nand U1288 (N_1288,In_956,In_1665);
xnor U1289 (N_1289,In_1617,In_542);
nor U1290 (N_1290,In_1178,In_2890);
and U1291 (N_1291,In_2850,In_1657);
or U1292 (N_1292,In_799,In_1940);
nor U1293 (N_1293,In_2200,In_1618);
or U1294 (N_1294,In_916,In_1127);
and U1295 (N_1295,In_1694,In_2523);
nand U1296 (N_1296,In_1338,In_514);
nand U1297 (N_1297,In_2140,In_1089);
or U1298 (N_1298,In_407,In_812);
xnor U1299 (N_1299,In_2057,In_928);
xnor U1300 (N_1300,In_2910,In_678);
nand U1301 (N_1301,In_2162,In_1267);
nand U1302 (N_1302,In_574,In_580);
or U1303 (N_1303,In_1762,In_2413);
nand U1304 (N_1304,In_273,In_2549);
or U1305 (N_1305,In_5,In_45);
and U1306 (N_1306,In_1210,In_1969);
and U1307 (N_1307,In_1043,In_482);
nand U1308 (N_1308,In_56,In_841);
nor U1309 (N_1309,In_1860,In_1328);
and U1310 (N_1310,In_1380,In_2292);
and U1311 (N_1311,In_885,In_1741);
or U1312 (N_1312,In_1754,In_1457);
or U1313 (N_1313,In_1530,In_2294);
or U1314 (N_1314,In_305,In_2640);
nand U1315 (N_1315,In_1152,In_2202);
xnor U1316 (N_1316,In_86,In_2973);
nor U1317 (N_1317,In_944,In_1455);
xnor U1318 (N_1318,In_1980,In_2328);
xor U1319 (N_1319,In_737,In_421);
xor U1320 (N_1320,In_759,In_2628);
or U1321 (N_1321,In_2396,In_1065);
and U1322 (N_1322,In_1183,In_2016);
or U1323 (N_1323,In_2520,In_2794);
and U1324 (N_1324,In_1669,In_112);
nor U1325 (N_1325,In_621,In_1602);
or U1326 (N_1326,In_1314,In_1309);
nand U1327 (N_1327,In_2420,In_1331);
or U1328 (N_1328,In_2190,In_2185);
and U1329 (N_1329,In_2568,In_2656);
nand U1330 (N_1330,In_350,In_2692);
or U1331 (N_1331,In_416,In_751);
nand U1332 (N_1332,In_930,In_1506);
nand U1333 (N_1333,In_218,In_938);
and U1334 (N_1334,In_756,In_625);
xnor U1335 (N_1335,In_2385,In_1601);
nor U1336 (N_1336,In_776,In_1045);
nand U1337 (N_1337,In_1433,In_1725);
and U1338 (N_1338,In_2336,In_194);
nor U1339 (N_1339,In_906,In_252);
nor U1340 (N_1340,In_848,In_1748);
xnor U1341 (N_1341,In_1917,In_1356);
and U1342 (N_1342,In_2907,In_2553);
nor U1343 (N_1343,In_1755,In_1019);
and U1344 (N_1344,In_450,In_825);
xor U1345 (N_1345,In_13,In_1411);
and U1346 (N_1346,In_909,In_741);
nand U1347 (N_1347,In_2366,In_2417);
and U1348 (N_1348,In_2377,In_2513);
xor U1349 (N_1349,In_2868,In_1076);
nor U1350 (N_1350,In_575,In_364);
nand U1351 (N_1351,In_47,In_2787);
nor U1352 (N_1352,In_118,In_2703);
and U1353 (N_1353,In_704,In_2575);
or U1354 (N_1354,In_2650,In_1798);
nor U1355 (N_1355,In_2009,In_1673);
xor U1356 (N_1356,In_1763,In_1285);
xnor U1357 (N_1357,In_969,In_688);
or U1358 (N_1358,In_2908,In_2093);
or U1359 (N_1359,In_98,In_1075);
nor U1360 (N_1360,In_2365,In_2604);
xor U1361 (N_1361,In_1868,In_2661);
nor U1362 (N_1362,In_715,In_895);
nand U1363 (N_1363,In_2247,In_320);
nand U1364 (N_1364,In_1116,In_1000);
nand U1365 (N_1365,In_2790,In_1325);
nand U1366 (N_1366,In_2068,In_2614);
nand U1367 (N_1367,In_2340,In_2773);
or U1368 (N_1368,In_366,In_392);
and U1369 (N_1369,In_2029,In_1181);
or U1370 (N_1370,In_2386,In_978);
nor U1371 (N_1371,In_1825,In_1327);
nor U1372 (N_1372,In_1143,In_1125);
and U1373 (N_1373,In_1820,In_1671);
nand U1374 (N_1374,In_1649,In_2683);
or U1375 (N_1375,In_2265,In_80);
xor U1376 (N_1376,In_651,In_2832);
xnor U1377 (N_1377,In_2942,In_258);
and U1378 (N_1378,In_133,In_545);
xnor U1379 (N_1379,In_341,In_171);
and U1380 (N_1380,In_2572,In_1508);
or U1381 (N_1381,In_2346,In_1369);
and U1382 (N_1382,In_582,In_103);
or U1383 (N_1383,In_1997,In_2091);
or U1384 (N_1384,In_2527,In_2456);
or U1385 (N_1385,In_1337,In_153);
nand U1386 (N_1386,In_2415,In_313);
xor U1387 (N_1387,In_817,In_2851);
and U1388 (N_1388,In_779,In_594);
nor U1389 (N_1389,In_460,In_1635);
nor U1390 (N_1390,In_662,In_2871);
xnor U1391 (N_1391,In_2071,In_2231);
xnor U1392 (N_1392,In_2049,In_2494);
or U1393 (N_1393,In_355,In_2665);
nand U1394 (N_1394,In_1459,In_989);
nor U1395 (N_1395,In_1233,In_2784);
xor U1396 (N_1396,In_1425,In_1326);
nand U1397 (N_1397,In_296,In_811);
nor U1398 (N_1398,In_33,In_2741);
or U1399 (N_1399,In_846,In_1779);
nand U1400 (N_1400,In_2324,In_1733);
or U1401 (N_1401,In_2937,In_1100);
nor U1402 (N_1402,In_2675,In_2856);
nand U1403 (N_1403,In_1332,In_992);
nand U1404 (N_1404,In_1742,In_537);
xor U1405 (N_1405,In_1389,In_1110);
nor U1406 (N_1406,In_809,In_1701);
nor U1407 (N_1407,In_304,In_2718);
xor U1408 (N_1408,In_893,In_707);
or U1409 (N_1409,In_435,In_1121);
nor U1410 (N_1410,In_1490,In_843);
nand U1411 (N_1411,In_777,In_1157);
or U1412 (N_1412,In_1312,In_1837);
xnor U1413 (N_1413,In_1149,In_1421);
nor U1414 (N_1414,In_1812,In_1611);
and U1415 (N_1415,In_2837,In_2587);
or U1416 (N_1416,In_1169,In_1928);
nor U1417 (N_1417,In_2107,In_1099);
nor U1418 (N_1418,In_1743,In_423);
nor U1419 (N_1419,In_300,In_1491);
xor U1420 (N_1420,In_405,In_1977);
xnor U1421 (N_1421,In_1042,In_2353);
nor U1422 (N_1422,In_478,In_1107);
nand U1423 (N_1423,In_1946,In_952);
nor U1424 (N_1424,In_1896,In_2143);
nand U1425 (N_1425,In_1634,In_2989);
or U1426 (N_1426,In_1189,In_2227);
nand U1427 (N_1427,In_270,In_2515);
nor U1428 (N_1428,In_1234,In_2063);
nand U1429 (N_1429,In_1895,In_2814);
or U1430 (N_1430,In_1592,In_2601);
xnor U1431 (N_1431,In_1028,In_1543);
nor U1432 (N_1432,In_864,In_30);
or U1433 (N_1433,In_810,In_2751);
and U1434 (N_1434,In_2976,In_75);
and U1435 (N_1435,In_344,In_1653);
nand U1436 (N_1436,In_1703,In_2462);
and U1437 (N_1437,In_413,In_925);
xnor U1438 (N_1438,In_60,In_603);
xor U1439 (N_1439,In_1996,In_1250);
nor U1440 (N_1440,In_836,In_1546);
nor U1441 (N_1441,In_1886,In_781);
nor U1442 (N_1442,In_387,In_1134);
nor U1443 (N_1443,In_1123,In_345);
and U1444 (N_1444,In_1687,In_2746);
or U1445 (N_1445,In_1767,In_1219);
xnor U1446 (N_1446,In_902,In_997);
and U1447 (N_1447,In_2156,In_887);
nand U1448 (N_1448,In_1939,In_223);
and U1449 (N_1449,In_2150,In_2763);
nor U1450 (N_1450,In_2031,In_1749);
nor U1451 (N_1451,In_1375,In_2030);
and U1452 (N_1452,In_1098,In_2349);
and U1453 (N_1453,In_1082,In_2312);
and U1454 (N_1454,In_1122,In_2408);
nor U1455 (N_1455,In_1522,In_2128);
and U1456 (N_1456,In_2714,In_131);
or U1457 (N_1457,In_2626,In_1484);
nor U1458 (N_1458,In_1775,In_1888);
xnor U1459 (N_1459,In_1096,In_192);
or U1460 (N_1460,In_2245,In_1972);
nor U1461 (N_1461,In_2138,In_299);
xor U1462 (N_1462,In_2302,In_1373);
xor U1463 (N_1463,In_162,In_899);
xor U1464 (N_1464,In_718,In_406);
nand U1465 (N_1465,In_2623,In_2110);
xnor U1466 (N_1466,In_2861,In_813);
and U1467 (N_1467,In_2317,In_2874);
or U1468 (N_1468,In_771,In_1006);
nor U1469 (N_1469,In_798,In_237);
and U1470 (N_1470,In_2468,In_2807);
or U1471 (N_1471,In_2681,In_1295);
nor U1472 (N_1472,In_470,In_2013);
and U1473 (N_1473,In_2885,In_58);
and U1474 (N_1474,In_1283,In_1591);
nand U1475 (N_1475,In_1058,In_2449);
nand U1476 (N_1476,In_692,In_2341);
nor U1477 (N_1477,In_891,In_2978);
nor U1478 (N_1478,In_668,In_40);
and U1479 (N_1479,In_1290,In_638);
and U1480 (N_1480,In_1279,In_1293);
nand U1481 (N_1481,In_498,In_2109);
or U1482 (N_1482,In_2118,In_2847);
nor U1483 (N_1483,In_1550,In_1206);
xor U1484 (N_1484,In_926,In_175);
xor U1485 (N_1485,In_1452,In_1819);
nand U1486 (N_1486,In_203,In_2108);
or U1487 (N_1487,In_1016,In_43);
and U1488 (N_1488,In_1438,In_2236);
xnor U1489 (N_1489,In_1339,In_2648);
xnor U1490 (N_1490,In_546,In_538);
nor U1491 (N_1491,In_905,In_2783);
or U1492 (N_1492,In_1730,In_803);
nor U1493 (N_1493,In_2056,In_1067);
and U1494 (N_1494,In_1829,In_1440);
xnor U1495 (N_1495,In_2321,In_1330);
nand U1496 (N_1496,In_886,In_2823);
or U1497 (N_1497,In_888,In_1949);
xor U1498 (N_1498,In_1163,In_529);
or U1499 (N_1499,In_1654,In_673);
xnor U1500 (N_1500,N_1399,N_1414);
and U1501 (N_1501,N_990,N_395);
or U1502 (N_1502,N_1073,N_854);
nor U1503 (N_1503,N_1053,N_191);
nor U1504 (N_1504,N_210,N_241);
nand U1505 (N_1505,N_1068,N_575);
xnor U1506 (N_1506,N_1452,N_209);
nor U1507 (N_1507,N_1358,N_1361);
xor U1508 (N_1508,N_810,N_110);
nand U1509 (N_1509,N_778,N_1075);
and U1510 (N_1510,N_378,N_552);
and U1511 (N_1511,N_1220,N_1302);
nand U1512 (N_1512,N_512,N_219);
and U1513 (N_1513,N_1014,N_187);
nand U1514 (N_1514,N_1336,N_1359);
nand U1515 (N_1515,N_6,N_518);
nor U1516 (N_1516,N_253,N_1439);
or U1517 (N_1517,N_1006,N_477);
or U1518 (N_1518,N_272,N_742);
or U1519 (N_1519,N_350,N_177);
xnor U1520 (N_1520,N_1033,N_855);
nor U1521 (N_1521,N_1298,N_417);
nor U1522 (N_1522,N_408,N_1477);
or U1523 (N_1523,N_326,N_1032);
nand U1524 (N_1524,N_324,N_967);
xnor U1525 (N_1525,N_1065,N_1363);
and U1526 (N_1526,N_172,N_308);
or U1527 (N_1527,N_182,N_681);
nor U1528 (N_1528,N_971,N_933);
nor U1529 (N_1529,N_74,N_767);
nor U1530 (N_1530,N_962,N_638);
xor U1531 (N_1531,N_1378,N_1262);
and U1532 (N_1532,N_36,N_1013);
xnor U1533 (N_1533,N_802,N_838);
xor U1534 (N_1534,N_906,N_874);
or U1535 (N_1535,N_1029,N_514);
or U1536 (N_1536,N_574,N_687);
xor U1537 (N_1537,N_865,N_118);
or U1538 (N_1538,N_522,N_1016);
and U1539 (N_1539,N_487,N_712);
and U1540 (N_1540,N_673,N_317);
or U1541 (N_1541,N_839,N_136);
or U1542 (N_1542,N_69,N_1097);
nand U1543 (N_1543,N_938,N_318);
nor U1544 (N_1544,N_884,N_746);
nand U1545 (N_1545,N_1417,N_616);
and U1546 (N_1546,N_877,N_1171);
or U1547 (N_1547,N_328,N_1481);
or U1548 (N_1548,N_1374,N_1400);
or U1549 (N_1549,N_785,N_516);
nand U1550 (N_1550,N_627,N_790);
xnor U1551 (N_1551,N_1407,N_557);
nor U1552 (N_1552,N_1401,N_1288);
or U1553 (N_1553,N_66,N_342);
and U1554 (N_1554,N_832,N_335);
nor U1555 (N_1555,N_1486,N_1);
nor U1556 (N_1556,N_1311,N_1163);
nor U1557 (N_1557,N_1069,N_213);
xor U1558 (N_1558,N_615,N_911);
xor U1559 (N_1559,N_1460,N_336);
or U1560 (N_1560,N_331,N_347);
or U1561 (N_1561,N_1416,N_57);
xnor U1562 (N_1562,N_282,N_1464);
and U1563 (N_1563,N_1057,N_142);
nand U1564 (N_1564,N_887,N_101);
nand U1565 (N_1565,N_84,N_885);
and U1566 (N_1566,N_761,N_745);
or U1567 (N_1567,N_256,N_920);
or U1568 (N_1568,N_502,N_783);
xor U1569 (N_1569,N_406,N_1027);
nor U1570 (N_1570,N_1076,N_530);
xnor U1571 (N_1571,N_642,N_83);
nand U1572 (N_1572,N_1349,N_1397);
nand U1573 (N_1573,N_416,N_115);
and U1574 (N_1574,N_992,N_1461);
or U1575 (N_1575,N_538,N_734);
nor U1576 (N_1576,N_592,N_246);
nand U1577 (N_1577,N_1131,N_462);
and U1578 (N_1578,N_1447,N_438);
and U1579 (N_1579,N_702,N_31);
nor U1580 (N_1580,N_201,N_1042);
or U1581 (N_1581,N_1296,N_650);
and U1582 (N_1582,N_1007,N_49);
nor U1583 (N_1583,N_504,N_1487);
nand U1584 (N_1584,N_124,N_1320);
nand U1585 (N_1585,N_1081,N_679);
and U1586 (N_1586,N_402,N_1498);
nor U1587 (N_1587,N_1205,N_671);
xnor U1588 (N_1588,N_1157,N_1213);
or U1589 (N_1589,N_1022,N_1269);
or U1590 (N_1590,N_410,N_85);
nand U1591 (N_1591,N_194,N_781);
nand U1592 (N_1592,N_44,N_38);
xor U1593 (N_1593,N_307,N_978);
nor U1594 (N_1594,N_735,N_506);
nand U1595 (N_1595,N_1389,N_52);
or U1596 (N_1596,N_398,N_848);
nor U1597 (N_1597,N_455,N_10);
xor U1598 (N_1598,N_1338,N_291);
nand U1599 (N_1599,N_461,N_711);
nand U1600 (N_1600,N_842,N_714);
or U1601 (N_1601,N_663,N_1412);
nor U1602 (N_1602,N_1138,N_491);
xnor U1603 (N_1603,N_1404,N_351);
nand U1604 (N_1604,N_1125,N_1118);
and U1605 (N_1605,N_19,N_1335);
xor U1606 (N_1606,N_7,N_1038);
xor U1607 (N_1607,N_773,N_76);
or U1608 (N_1608,N_1054,N_665);
nor U1609 (N_1609,N_1214,N_1370);
and U1610 (N_1610,N_28,N_130);
nand U1611 (N_1611,N_190,N_1207);
nor U1612 (N_1612,N_257,N_91);
xor U1613 (N_1613,N_928,N_176);
xor U1614 (N_1614,N_27,N_131);
xor U1615 (N_1615,N_1462,N_1367);
xor U1616 (N_1616,N_814,N_1492);
nor U1617 (N_1617,N_1329,N_520);
or U1618 (N_1618,N_1406,N_591);
and U1619 (N_1619,N_385,N_141);
or U1620 (N_1620,N_708,N_313);
xor U1621 (N_1621,N_644,N_242);
and U1622 (N_1622,N_703,N_180);
nor U1623 (N_1623,N_1419,N_886);
and U1624 (N_1624,N_479,N_46);
and U1625 (N_1625,N_1059,N_102);
nor U1626 (N_1626,N_433,N_929);
or U1627 (N_1627,N_547,N_1255);
or U1628 (N_1628,N_295,N_1484);
and U1629 (N_1629,N_1395,N_910);
xnor U1630 (N_1630,N_404,N_1490);
xnor U1631 (N_1631,N_473,N_364);
and U1632 (N_1632,N_713,N_1450);
or U1633 (N_1633,N_409,N_375);
nor U1634 (N_1634,N_1170,N_890);
nor U1635 (N_1635,N_576,N_608);
and U1636 (N_1636,N_1119,N_654);
and U1637 (N_1637,N_259,N_1150);
xor U1638 (N_1638,N_1441,N_541);
and U1639 (N_1639,N_693,N_1135);
nand U1640 (N_1640,N_1434,N_279);
or U1641 (N_1641,N_863,N_826);
and U1642 (N_1642,N_828,N_106);
nor U1643 (N_1643,N_78,N_896);
or U1644 (N_1644,N_2,N_927);
nor U1645 (N_1645,N_1117,N_258);
nor U1646 (N_1646,N_862,N_769);
or U1647 (N_1647,N_450,N_1390);
and U1648 (N_1648,N_723,N_63);
xnor U1649 (N_1649,N_144,N_70);
nor U1650 (N_1650,N_595,N_777);
xnor U1651 (N_1651,N_1074,N_1306);
and U1652 (N_1652,N_1377,N_1200);
xor U1653 (N_1653,N_87,N_1274);
and U1654 (N_1654,N_904,N_1301);
nand U1655 (N_1655,N_271,N_186);
nand U1656 (N_1656,N_218,N_747);
nand U1657 (N_1657,N_951,N_900);
or U1658 (N_1658,N_1112,N_212);
and U1659 (N_1659,N_156,N_200);
or U1660 (N_1660,N_1266,N_273);
nor U1661 (N_1661,N_1479,N_1483);
and U1662 (N_1662,N_803,N_602);
or U1663 (N_1663,N_695,N_355);
xor U1664 (N_1664,N_1287,N_389);
xor U1665 (N_1665,N_830,N_550);
nor U1666 (N_1666,N_1313,N_1391);
nor U1667 (N_1667,N_543,N_1062);
or U1668 (N_1668,N_1149,N_198);
nand U1669 (N_1669,N_228,N_744);
nand U1670 (N_1670,N_1355,N_1257);
nor U1671 (N_1671,N_590,N_961);
xnor U1672 (N_1672,N_423,N_26);
and U1673 (N_1673,N_1373,N_353);
nand U1674 (N_1674,N_1428,N_721);
xor U1675 (N_1675,N_1384,N_709);
nor U1676 (N_1676,N_605,N_1037);
or U1677 (N_1677,N_738,N_1433);
and U1678 (N_1678,N_816,N_157);
xor U1679 (N_1679,N_812,N_283);
nand U1680 (N_1680,N_625,N_275);
nor U1681 (N_1681,N_749,N_357);
nor U1682 (N_1682,N_316,N_1051);
xnor U1683 (N_1683,N_684,N_883);
or U1684 (N_1684,N_1045,N_1246);
nor U1685 (N_1685,N_622,N_857);
xnor U1686 (N_1686,N_934,N_924);
xnor U1687 (N_1687,N_1225,N_722);
and U1688 (N_1688,N_980,N_1195);
nand U1689 (N_1689,N_319,N_1031);
nand U1690 (N_1690,N_252,N_1156);
or U1691 (N_1691,N_1431,N_123);
nand U1692 (N_1692,N_158,N_486);
or U1693 (N_1693,N_798,N_728);
xnor U1694 (N_1694,N_9,N_901);
nor U1695 (N_1695,N_233,N_941);
and U1696 (N_1696,N_856,N_12);
nor U1697 (N_1697,N_215,N_22);
nand U1698 (N_1698,N_1242,N_226);
xnor U1699 (N_1699,N_999,N_1368);
xnor U1700 (N_1700,N_1472,N_236);
or U1701 (N_1701,N_1020,N_809);
and U1702 (N_1702,N_1418,N_1388);
and U1703 (N_1703,N_249,N_1325);
nand U1704 (N_1704,N_556,N_606);
xor U1705 (N_1705,N_1303,N_67);
or U1706 (N_1706,N_1383,N_689);
or U1707 (N_1707,N_1328,N_459);
and U1708 (N_1708,N_1025,N_1048);
or U1709 (N_1709,N_680,N_1233);
or U1710 (N_1710,N_1174,N_572);
or U1711 (N_1711,N_942,N_548);
nor U1712 (N_1712,N_1426,N_1348);
xor U1713 (N_1713,N_947,N_1279);
or U1714 (N_1714,N_222,N_15);
xnor U1715 (N_1715,N_573,N_765);
xnor U1716 (N_1716,N_771,N_536);
xnor U1717 (N_1717,N_607,N_1470);
and U1718 (N_1718,N_500,N_1111);
nand U1719 (N_1719,N_813,N_359);
nor U1720 (N_1720,N_1432,N_11);
xnor U1721 (N_1721,N_628,N_1113);
or U1722 (N_1722,N_549,N_1276);
xnor U1723 (N_1723,N_694,N_276);
nor U1724 (N_1724,N_18,N_1114);
nand U1725 (N_1725,N_535,N_766);
nor U1726 (N_1726,N_61,N_1012);
xnor U1727 (N_1727,N_1275,N_898);
or U1728 (N_1728,N_337,N_105);
nor U1729 (N_1729,N_1376,N_488);
nor U1730 (N_1730,N_1206,N_1124);
or U1731 (N_1731,N_989,N_1001);
or U1732 (N_1732,N_160,N_675);
or U1733 (N_1733,N_358,N_955);
nand U1734 (N_1734,N_1425,N_1226);
nand U1735 (N_1735,N_56,N_1413);
nand U1736 (N_1736,N_779,N_823);
and U1737 (N_1737,N_82,N_1091);
nand U1738 (N_1738,N_1175,N_780);
or U1739 (N_1739,N_1291,N_293);
or U1740 (N_1740,N_20,N_988);
nand U1741 (N_1741,N_401,N_819);
xor U1742 (N_1742,N_844,N_822);
xor U1743 (N_1743,N_21,N_274);
xor U1744 (N_1744,N_649,N_991);
nand U1745 (N_1745,N_62,N_1443);
nor U1746 (N_1746,N_1292,N_1201);
xnor U1747 (N_1747,N_254,N_1493);
nor U1748 (N_1748,N_1203,N_604);
and U1749 (N_1749,N_774,N_935);
nor U1750 (N_1750,N_891,N_1099);
or U1751 (N_1751,N_662,N_850);
and U1752 (N_1752,N_418,N_1382);
nand U1753 (N_1753,N_205,N_882);
and U1754 (N_1754,N_250,N_1438);
or U1755 (N_1755,N_1356,N_1093);
or U1756 (N_1756,N_381,N_1371);
or U1757 (N_1757,N_1415,N_237);
or U1758 (N_1758,N_1307,N_352);
or U1759 (N_1759,N_425,N_1046);
nor U1760 (N_1760,N_845,N_97);
and U1761 (N_1761,N_388,N_1066);
xnor U1762 (N_1762,N_464,N_852);
or U1763 (N_1763,N_588,N_1247);
nor U1764 (N_1764,N_878,N_469);
or U1765 (N_1765,N_1326,N_474);
nor U1766 (N_1766,N_719,N_45);
nand U1767 (N_1767,N_1224,N_655);
or U1768 (N_1768,N_944,N_303);
xnor U1769 (N_1769,N_902,N_659);
xnor U1770 (N_1770,N_508,N_1421);
nor U1771 (N_1771,N_346,N_1345);
nand U1772 (N_1772,N_413,N_305);
or U1773 (N_1773,N_544,N_1386);
or U1774 (N_1774,N_578,N_584);
nand U1775 (N_1775,N_1259,N_676);
nand U1776 (N_1776,N_637,N_599);
and U1777 (N_1777,N_922,N_245);
and U1778 (N_1778,N_1314,N_292);
and U1779 (N_1779,N_1495,N_881);
nand U1780 (N_1780,N_970,N_784);
nand U1781 (N_1781,N_419,N_1465);
or U1782 (N_1782,N_1197,N_179);
xnor U1783 (N_1783,N_384,N_312);
nand U1784 (N_1784,N_1047,N_390);
nand U1785 (N_1785,N_1109,N_894);
nor U1786 (N_1786,N_93,N_529);
nand U1787 (N_1787,N_53,N_634);
and U1788 (N_1788,N_1256,N_788);
and U1789 (N_1789,N_1366,N_231);
xor U1790 (N_1790,N_152,N_1482);
nand U1791 (N_1791,N_1004,N_1172);
or U1792 (N_1792,N_973,N_993);
xor U1793 (N_1793,N_1337,N_453);
xnor U1794 (N_1794,N_1267,N_1188);
and U1795 (N_1795,N_1300,N_482);
nor U1796 (N_1796,N_859,N_1082);
and U1797 (N_1797,N_248,N_800);
xor U1798 (N_1798,N_580,N_1077);
xor U1799 (N_1799,N_869,N_161);
nor U1800 (N_1800,N_782,N_736);
and U1801 (N_1801,N_162,N_165);
nor U1802 (N_1802,N_341,N_64);
nand U1803 (N_1803,N_908,N_1078);
and U1804 (N_1804,N_847,N_875);
nor U1805 (N_1805,N_1160,N_1339);
or U1806 (N_1806,N_1238,N_452);
nand U1807 (N_1807,N_619,N_299);
or U1808 (N_1808,N_964,N_1126);
or U1809 (N_1809,N_1222,N_72);
or U1810 (N_1810,N_369,N_1227);
xnor U1811 (N_1811,N_463,N_1129);
and U1812 (N_1812,N_1088,N_808);
and U1813 (N_1813,N_873,N_1079);
nand U1814 (N_1814,N_125,N_1295);
xor U1815 (N_1815,N_447,N_925);
xor U1816 (N_1816,N_569,N_23);
or U1817 (N_1817,N_60,N_278);
nor U1818 (N_1818,N_428,N_240);
nand U1819 (N_1819,N_265,N_0);
nor U1820 (N_1820,N_772,N_757);
xor U1821 (N_1821,N_135,N_14);
xor U1822 (N_1822,N_1489,N_111);
nor U1823 (N_1823,N_497,N_1310);
or U1824 (N_1824,N_239,N_716);
or U1825 (N_1825,N_349,N_1084);
nand U1826 (N_1826,N_492,N_1488);
xnor U1827 (N_1827,N_95,N_432);
nor U1828 (N_1828,N_979,N_1278);
xor U1829 (N_1829,N_566,N_907);
xnor U1830 (N_1830,N_1009,N_840);
and U1831 (N_1831,N_140,N_16);
nor U1832 (N_1832,N_167,N_1183);
nor U1833 (N_1833,N_214,N_325);
or U1834 (N_1834,N_1058,N_414);
and U1835 (N_1835,N_755,N_1245);
nand U1836 (N_1836,N_168,N_1420);
and U1837 (N_1837,N_1333,N_515);
and U1838 (N_1838,N_129,N_1185);
xor U1839 (N_1839,N_1189,N_34);
nand U1840 (N_1840,N_481,N_794);
xnor U1841 (N_1841,N_143,N_546);
nor U1842 (N_1842,N_1261,N_465);
xnor U1843 (N_1843,N_367,N_611);
or U1844 (N_1844,N_563,N_224);
nand U1845 (N_1845,N_173,N_1318);
xor U1846 (N_1846,N_297,N_499);
and U1847 (N_1847,N_682,N_183);
nor U1848 (N_1848,N_903,N_1162);
and U1849 (N_1849,N_952,N_1392);
xor U1850 (N_1850,N_623,N_1403);
xnor U1851 (N_1851,N_334,N_1215);
nand U1852 (N_1852,N_498,N_889);
or U1853 (N_1853,N_507,N_1110);
and U1854 (N_1854,N_1398,N_705);
nand U1855 (N_1855,N_931,N_1272);
nand U1856 (N_1856,N_1080,N_641);
or U1857 (N_1857,N_54,N_327);
xor U1858 (N_1858,N_581,N_1396);
and U1859 (N_1859,N_8,N_260);
nand U1860 (N_1860,N_976,N_128);
or U1861 (N_1861,N_227,N_1381);
nor U1862 (N_1862,N_470,N_108);
nand U1863 (N_1863,N_1448,N_119);
nor U1864 (N_1864,N_446,N_332);
nand U1865 (N_1865,N_298,N_539);
nand U1866 (N_1866,N_617,N_585);
nor U1867 (N_1867,N_791,N_633);
or U1868 (N_1868,N_1064,N_759);
or U1869 (N_1869,N_731,N_821);
or U1870 (N_1870,N_526,N_396);
xor U1871 (N_1871,N_1260,N_354);
nand U1872 (N_1872,N_914,N_1043);
xnor U1873 (N_1873,N_1457,N_1322);
xnor U1874 (N_1874,N_1144,N_743);
nor U1875 (N_1875,N_1121,N_612);
nor U1876 (N_1876,N_1332,N_571);
xnor U1877 (N_1877,N_262,N_41);
nor U1878 (N_1878,N_287,N_1430);
and U1879 (N_1879,N_1408,N_277);
nor U1880 (N_1880,N_741,N_510);
and U1881 (N_1881,N_589,N_344);
xor U1882 (N_1882,N_368,N_1060);
nor U1883 (N_1883,N_525,N_1342);
xnor U1884 (N_1884,N_727,N_730);
xor U1885 (N_1885,N_361,N_1083);
and U1886 (N_1886,N_912,N_1094);
nand U1887 (N_1887,N_706,N_387);
nor U1888 (N_1888,N_923,N_1141);
xnor U1889 (N_1889,N_1351,N_554);
or U1890 (N_1890,N_468,N_251);
nor U1891 (N_1891,N_1052,N_517);
xor U1892 (N_1892,N_752,N_764);
nor U1893 (N_1893,N_496,N_846);
nor U1894 (N_1894,N_820,N_397);
or U1895 (N_1895,N_1235,N_943);
nor U1896 (N_1896,N_1100,N_753);
and U1897 (N_1897,N_1293,N_1169);
nand U1898 (N_1898,N_1273,N_690);
and U1899 (N_1899,N_946,N_1089);
or U1900 (N_1900,N_304,N_429);
nand U1901 (N_1901,N_372,N_661);
nand U1902 (N_1902,N_284,N_109);
nand U1903 (N_1903,N_365,N_1123);
nor U1904 (N_1904,N_1194,N_523);
or U1905 (N_1905,N_677,N_567);
nor U1906 (N_1906,N_280,N_1281);
or U1907 (N_1907,N_1466,N_645);
xnor U1908 (N_1908,N_1280,N_932);
nor U1909 (N_1909,N_285,N_1164);
nand U1910 (N_1910,N_185,N_1440);
nor U1911 (N_1911,N_1070,N_127);
nand U1912 (N_1912,N_1107,N_51);
and U1913 (N_1913,N_1103,N_763);
nor U1914 (N_1914,N_1308,N_1133);
and U1915 (N_1915,N_740,N_25);
and U1916 (N_1916,N_1485,N_658);
nor U1917 (N_1917,N_1198,N_751);
or U1918 (N_1918,N_1211,N_163);
xor U1919 (N_1919,N_949,N_521);
nor U1920 (N_1920,N_126,N_919);
nand U1921 (N_1921,N_597,N_963);
xor U1922 (N_1922,N_825,N_833);
and U1923 (N_1923,N_1268,N_513);
and U1924 (N_1924,N_996,N_422);
or U1925 (N_1925,N_220,N_1202);
nor U1926 (N_1926,N_1158,N_90);
or U1927 (N_1927,N_1067,N_691);
nor U1928 (N_1928,N_542,N_100);
and U1929 (N_1929,N_948,N_164);
and U1930 (N_1930,N_1044,N_870);
nor U1931 (N_1931,N_475,N_399);
nor U1932 (N_1932,N_1271,N_787);
nand U1933 (N_1933,N_151,N_899);
xnor U1934 (N_1934,N_797,N_620);
nand U1935 (N_1935,N_799,N_79);
nand U1936 (N_1936,N_564,N_975);
nand U1937 (N_1937,N_314,N_1405);
and U1938 (N_1938,N_1146,N_1341);
nor U1939 (N_1939,N_269,N_1139);
or U1940 (N_1940,N_577,N_598);
nand U1941 (N_1941,N_770,N_1353);
and U1942 (N_1942,N_138,N_897);
and U1943 (N_1943,N_1340,N_412);
nand U1944 (N_1944,N_1243,N_137);
or U1945 (N_1945,N_420,N_1343);
xnor U1946 (N_1946,N_235,N_1499);
nor U1947 (N_1947,N_225,N_55);
or U1948 (N_1948,N_68,N_699);
and U1949 (N_1949,N_3,N_648);
nor U1950 (N_1950,N_715,N_1444);
nor U1951 (N_1951,N_653,N_704);
nand U1952 (N_1952,N_217,N_905);
and U1953 (N_1953,N_148,N_534);
and U1954 (N_1954,N_1241,N_593);
xor U1955 (N_1955,N_1134,N_1334);
and U1956 (N_1956,N_1354,N_1496);
and U1957 (N_1957,N_1264,N_930);
or U1958 (N_1958,N_221,N_1072);
xor U1959 (N_1959,N_868,N_707);
nor U1960 (N_1960,N_435,N_1309);
and U1961 (N_1961,N_939,N_441);
nor U1962 (N_1962,N_1315,N_306);
or U1963 (N_1963,N_267,N_1265);
nor U1964 (N_1964,N_1263,N_1250);
or U1965 (N_1965,N_801,N_1372);
or U1966 (N_1966,N_207,N_1459);
nand U1967 (N_1967,N_437,N_1176);
xnor U1968 (N_1968,N_737,N_892);
xor U1969 (N_1969,N_594,N_916);
and U1970 (N_1970,N_466,N_668);
and U1971 (N_1971,N_1491,N_405);
or U1972 (N_1972,N_540,N_178);
nor U1973 (N_1973,N_471,N_1148);
and U1974 (N_1974,N_796,N_1063);
nand U1975 (N_1975,N_1327,N_343);
nand U1976 (N_1976,N_1330,N_113);
and U1977 (N_1977,N_1347,N_621);
xor U1978 (N_1978,N_528,N_1153);
and U1979 (N_1979,N_1357,N_1365);
or U1980 (N_1980,N_1231,N_1240);
nor U1981 (N_1981,N_407,N_467);
nand U1982 (N_1982,N_92,N_133);
or U1983 (N_1983,N_1092,N_997);
xor U1984 (N_1984,N_974,N_289);
nand U1985 (N_1985,N_4,N_876);
nand U1986 (N_1986,N_270,N_88);
xor U1987 (N_1987,N_59,N_841);
or U1988 (N_1988,N_789,N_65);
and U1989 (N_1989,N_1344,N_732);
nor U1990 (N_1990,N_202,N_685);
nand U1991 (N_1991,N_1364,N_553);
nand U1992 (N_1992,N_630,N_445);
or U1993 (N_1993,N_189,N_871);
nor U1994 (N_1994,N_1402,N_363);
xnor U1995 (N_1995,N_374,N_1244);
xor U1996 (N_1996,N_243,N_103);
and U1997 (N_1997,N_340,N_639);
nor U1998 (N_1998,N_555,N_94);
nor U1999 (N_1999,N_73,N_956);
nor U2000 (N_2000,N_1437,N_836);
and U2001 (N_2001,N_701,N_579);
nor U2002 (N_2002,N_674,N_1218);
or U2003 (N_2003,N_146,N_37);
or U2004 (N_2004,N_1192,N_503);
nand U2005 (N_2005,N_968,N_48);
or U2006 (N_2006,N_1283,N_696);
nor U2007 (N_2007,N_643,N_1290);
xor U2008 (N_2008,N_626,N_174);
nor U2009 (N_2009,N_13,N_383);
nand U2010 (N_2010,N_1017,N_483);
nand U2011 (N_2011,N_853,N_345);
nand U2012 (N_2012,N_1497,N_1108);
xnor U2013 (N_2013,N_371,N_1005);
or U2014 (N_2014,N_263,N_1061);
or U2015 (N_2015,N_47,N_632);
nor U2016 (N_2016,N_460,N_1229);
xnor U2017 (N_2017,N_533,N_1116);
and U2018 (N_2018,N_718,N_1427);
nor U2019 (N_2019,N_618,N_117);
nand U2020 (N_2020,N_983,N_1180);
nand U2021 (N_2021,N_159,N_139);
or U2022 (N_2022,N_614,N_1297);
xnor U2023 (N_2023,N_232,N_953);
or U2024 (N_2024,N_866,N_112);
xor U2025 (N_2025,N_1098,N_1028);
nand U2026 (N_2026,N_1234,N_1182);
xor U2027 (N_2027,N_726,N_1317);
xnor U2028 (N_2028,N_264,N_1305);
nand U2029 (N_2029,N_321,N_1480);
or U2030 (N_2030,N_149,N_81);
nor U2031 (N_2031,N_1467,N_1324);
and U2032 (N_2032,N_926,N_669);
nor U2033 (N_2033,N_1105,N_444);
and U2034 (N_2034,N_1237,N_1212);
and U2035 (N_2035,N_945,N_315);
nand U2036 (N_2036,N_562,N_559);
or U2037 (N_2037,N_443,N_472);
nand U2038 (N_2038,N_391,N_153);
xor U2039 (N_2039,N_1178,N_1204);
nand U2040 (N_2040,N_451,N_1216);
xnor U2041 (N_2041,N_670,N_985);
nor U2042 (N_2042,N_1446,N_1087);
or U2043 (N_2043,N_1375,N_966);
xnor U2044 (N_2044,N_1471,N_1451);
and U2045 (N_2045,N_750,N_107);
and U2046 (N_2046,N_805,N_1010);
xor U2047 (N_2047,N_457,N_601);
nand U2048 (N_2048,N_1019,N_188);
xor U2049 (N_2049,N_29,N_449);
or U2050 (N_2050,N_1115,N_986);
and U2051 (N_2051,N_994,N_1254);
nand U2052 (N_2052,N_288,N_403);
nand U2053 (N_2053,N_1186,N_829);
and U2054 (N_2054,N_223,N_1130);
nor U2055 (N_2055,N_1041,N_478);
nor U2056 (N_2056,N_430,N_454);
nor U2057 (N_2057,N_489,N_688);
xor U2058 (N_2058,N_458,N_1039);
nand U2059 (N_2059,N_394,N_867);
nor U2060 (N_2060,N_807,N_1219);
nand U2061 (N_2061,N_204,N_982);
nand U2062 (N_2062,N_1040,N_400);
or U2063 (N_2063,N_1230,N_1024);
xor U2064 (N_2064,N_568,N_1136);
or U2065 (N_2065,N_1168,N_739);
and U2066 (N_2066,N_1282,N_366);
or U2067 (N_2067,N_1350,N_150);
nor U2068 (N_2068,N_918,N_1217);
or U2069 (N_2069,N_717,N_603);
xnor U2070 (N_2070,N_476,N_247);
nand U2071 (N_2071,N_1002,N_1454);
xor U2072 (N_2072,N_957,N_1277);
xor U2073 (N_2073,N_879,N_77);
and U2074 (N_2074,N_1449,N_1196);
nand U2075 (N_2075,N_843,N_629);
nor U2076 (N_2076,N_1323,N_995);
and U2077 (N_2077,N_43,N_1422);
or U2078 (N_2078,N_255,N_1071);
and U2079 (N_2079,N_42,N_1253);
or U2080 (N_2080,N_1122,N_442);
nor U2081 (N_2081,N_104,N_537);
or U2082 (N_2082,N_1362,N_322);
nor U2083 (N_2083,N_193,N_490);
and U2084 (N_2084,N_1161,N_667);
nand U2085 (N_2085,N_448,N_917);
and U2086 (N_2086,N_1463,N_1023);
xnor U2087 (N_2087,N_348,N_1147);
or U2088 (N_2088,N_551,N_1409);
nand U2089 (N_2089,N_806,N_379);
and U2090 (N_2090,N_837,N_646);
nand U2091 (N_2091,N_1209,N_698);
nor U2092 (N_2092,N_1035,N_972);
nand U2093 (N_2093,N_1442,N_1424);
and U2094 (N_2094,N_710,N_309);
nor U2095 (N_2095,N_1165,N_1455);
xor U2096 (N_2096,N_196,N_1475);
nor U2097 (N_2097,N_32,N_880);
xnor U2098 (N_2098,N_565,N_959);
and U2099 (N_2099,N_380,N_1352);
and U2100 (N_2100,N_281,N_339);
or U2101 (N_2101,N_570,N_300);
or U2102 (N_2102,N_921,N_373);
nor U2103 (N_2103,N_827,N_1369);
nor U2104 (N_2104,N_166,N_1410);
or U2105 (N_2105,N_1036,N_1187);
nor U2106 (N_2106,N_1179,N_195);
or U2107 (N_2107,N_960,N_1140);
nand U2108 (N_2108,N_485,N_977);
xor U2109 (N_2109,N_672,N_360);
nand U2110 (N_2110,N_748,N_1312);
nor U2111 (N_2111,N_216,N_724);
xnor U2112 (N_2112,N_456,N_484);
xnor U2113 (N_2113,N_1142,N_96);
xor U2114 (N_2114,N_1166,N_1191);
nand U2115 (N_2115,N_758,N_1304);
xnor U2116 (N_2116,N_376,N_171);
xnor U2117 (N_2117,N_1193,N_392);
nand U2118 (N_2118,N_301,N_1385);
and U2119 (N_2119,N_969,N_1294);
and U2120 (N_2120,N_1049,N_1270);
or U2121 (N_2121,N_1102,N_651);
nor U2122 (N_2122,N_80,N_1152);
nand U2123 (N_2123,N_817,N_1346);
xnor U2124 (N_2124,N_206,N_208);
or U2125 (N_2125,N_424,N_330);
nand U2126 (N_2126,N_1155,N_1251);
or U2127 (N_2127,N_132,N_656);
and U2128 (N_2128,N_71,N_24);
and U2129 (N_2129,N_954,N_333);
xor U2130 (N_2130,N_610,N_505);
nand U2131 (N_2131,N_1018,N_431);
or U2132 (N_2132,N_120,N_244);
or U2133 (N_2133,N_582,N_635);
and U2134 (N_2134,N_600,N_647);
or U2135 (N_2135,N_362,N_480);
and U2136 (N_2136,N_524,N_652);
nor U2137 (N_2137,N_75,N_1299);
nand U2138 (N_2138,N_169,N_1223);
or U2139 (N_2139,N_561,N_636);
nor U2140 (N_2140,N_311,N_145);
nand U2141 (N_2141,N_729,N_211);
xnor U2142 (N_2142,N_1137,N_286);
nor U2143 (N_2143,N_1232,N_895);
or U2144 (N_2144,N_1387,N_1101);
nand U2145 (N_2145,N_1319,N_1456);
nor U2146 (N_2146,N_965,N_786);
or U2147 (N_2147,N_1145,N_30);
nor U2148 (N_2148,N_532,N_760);
or U2149 (N_2149,N_1177,N_697);
and U2150 (N_2150,N_720,N_495);
or U2151 (N_2151,N_1468,N_1000);
xnor U2152 (N_2152,N_1393,N_439);
and U2153 (N_2153,N_586,N_261);
nand U2154 (N_2154,N_657,N_1096);
xnor U2155 (N_2155,N_835,N_913);
nor U2156 (N_2156,N_33,N_678);
nand U2157 (N_2157,N_768,N_1210);
nand U2158 (N_2158,N_229,N_427);
and U2159 (N_2159,N_519,N_147);
nor U2160 (N_2160,N_329,N_596);
nand U2161 (N_2161,N_1208,N_199);
and U2162 (N_2162,N_415,N_421);
nand U2163 (N_2163,N_858,N_1015);
nand U2164 (N_2164,N_1154,N_664);
or U2165 (N_2165,N_583,N_1436);
xnor U2166 (N_2166,N_122,N_1167);
nor U2167 (N_2167,N_509,N_1411);
xor U2168 (N_2168,N_1453,N_1249);
or U2169 (N_2169,N_1445,N_386);
xor U2170 (N_2170,N_849,N_1085);
or U2171 (N_2171,N_940,N_631);
nand U2172 (N_2172,N_776,N_613);
xor U2173 (N_2173,N_1159,N_203);
and U2174 (N_2174,N_501,N_266);
and U2175 (N_2175,N_560,N_950);
nand U2176 (N_2176,N_692,N_234);
nor U2177 (N_2177,N_1132,N_50);
and U2178 (N_2178,N_733,N_175);
nand U2179 (N_2179,N_804,N_1128);
nor U2180 (N_2180,N_609,N_1173);
or U2181 (N_2181,N_1478,N_1429);
nor U2182 (N_2182,N_1011,N_494);
xnor U2183 (N_2183,N_1248,N_1331);
nand U2184 (N_2184,N_377,N_356);
xor U2185 (N_2185,N_861,N_99);
and U2186 (N_2186,N_238,N_1055);
xnor U2187 (N_2187,N_893,N_1184);
or U2188 (N_2188,N_121,N_660);
xnor U2189 (N_2189,N_754,N_1360);
nand U2190 (N_2190,N_5,N_17);
or U2191 (N_2191,N_338,N_1190);
nor U2192 (N_2192,N_1423,N_1086);
nand U2193 (N_2193,N_1494,N_527);
and U2194 (N_2194,N_1056,N_1379);
and U2195 (N_2195,N_864,N_1050);
nand U2196 (N_2196,N_811,N_795);
nand U2197 (N_2197,N_624,N_1003);
or U2198 (N_2198,N_815,N_268);
nand U2199 (N_2199,N_434,N_511);
or U2200 (N_2200,N_310,N_1026);
nor U2201 (N_2201,N_1435,N_40);
and U2202 (N_2202,N_493,N_411);
or U2203 (N_2203,N_323,N_1239);
and U2204 (N_2204,N_1034,N_756);
nand U2205 (N_2205,N_1008,N_192);
nor U2206 (N_2206,N_1469,N_1394);
nor U2207 (N_2207,N_888,N_1021);
xor U2208 (N_2208,N_793,N_89);
and U2209 (N_2209,N_1473,N_1127);
nand U2210 (N_2210,N_958,N_1120);
nor U2211 (N_2211,N_1104,N_987);
nand U2212 (N_2212,N_558,N_39);
or U2213 (N_2213,N_370,N_683);
and U2214 (N_2214,N_762,N_393);
nor U2215 (N_2215,N_818,N_98);
nand U2216 (N_2216,N_792,N_436);
and U2217 (N_2217,N_531,N_184);
nor U2218 (N_2218,N_1151,N_1289);
nor U2219 (N_2219,N_1236,N_872);
nand U2220 (N_2220,N_114,N_1458);
xor U2221 (N_2221,N_382,N_302);
xor U2222 (N_2222,N_1199,N_915);
and U2223 (N_2223,N_1316,N_1221);
xnor U2224 (N_2224,N_426,N_984);
and U2225 (N_2225,N_640,N_86);
and U2226 (N_2226,N_936,N_134);
nor U2227 (N_2227,N_909,N_860);
nand U2228 (N_2228,N_1380,N_230);
nor U2229 (N_2229,N_116,N_1285);
nor U2230 (N_2230,N_1252,N_981);
nand U2231 (N_2231,N_154,N_197);
nor U2232 (N_2232,N_998,N_700);
and U2233 (N_2233,N_1321,N_1181);
xnor U2234 (N_2234,N_1090,N_1106);
xor U2235 (N_2235,N_155,N_294);
and U2236 (N_2236,N_170,N_1228);
or U2237 (N_2237,N_1284,N_320);
xnor U2238 (N_2238,N_440,N_1258);
xnor U2239 (N_2239,N_725,N_1095);
nor U2240 (N_2240,N_851,N_545);
and U2241 (N_2241,N_775,N_824);
xor U2242 (N_2242,N_834,N_1476);
nand U2243 (N_2243,N_1286,N_1474);
or U2244 (N_2244,N_666,N_1030);
nor U2245 (N_2245,N_587,N_181);
nor U2246 (N_2246,N_58,N_937);
or U2247 (N_2247,N_35,N_1143);
or U2248 (N_2248,N_686,N_831);
nor U2249 (N_2249,N_290,N_296);
and U2250 (N_2250,N_1199,N_199);
nand U2251 (N_2251,N_173,N_590);
nand U2252 (N_2252,N_937,N_443);
xor U2253 (N_2253,N_1143,N_763);
nor U2254 (N_2254,N_1017,N_227);
nor U2255 (N_2255,N_896,N_1206);
nand U2256 (N_2256,N_1007,N_1225);
nor U2257 (N_2257,N_202,N_868);
xnor U2258 (N_2258,N_378,N_1466);
xnor U2259 (N_2259,N_902,N_1334);
and U2260 (N_2260,N_124,N_858);
nand U2261 (N_2261,N_1114,N_188);
or U2262 (N_2262,N_1477,N_700);
xor U2263 (N_2263,N_1368,N_913);
and U2264 (N_2264,N_1419,N_302);
or U2265 (N_2265,N_309,N_505);
and U2266 (N_2266,N_150,N_927);
or U2267 (N_2267,N_683,N_448);
or U2268 (N_2268,N_542,N_303);
and U2269 (N_2269,N_178,N_267);
or U2270 (N_2270,N_1043,N_575);
and U2271 (N_2271,N_171,N_671);
nor U2272 (N_2272,N_951,N_442);
nand U2273 (N_2273,N_490,N_979);
nand U2274 (N_2274,N_279,N_918);
and U2275 (N_2275,N_379,N_988);
xor U2276 (N_2276,N_1135,N_838);
nor U2277 (N_2277,N_1382,N_1393);
xnor U2278 (N_2278,N_1135,N_821);
xnor U2279 (N_2279,N_68,N_1392);
nand U2280 (N_2280,N_1031,N_639);
nor U2281 (N_2281,N_1171,N_1145);
and U2282 (N_2282,N_24,N_1281);
xnor U2283 (N_2283,N_1442,N_1326);
and U2284 (N_2284,N_374,N_22);
nand U2285 (N_2285,N_1206,N_242);
nor U2286 (N_2286,N_1350,N_691);
or U2287 (N_2287,N_92,N_1398);
nor U2288 (N_2288,N_572,N_1336);
or U2289 (N_2289,N_1024,N_225);
nor U2290 (N_2290,N_880,N_753);
nor U2291 (N_2291,N_1291,N_966);
or U2292 (N_2292,N_662,N_549);
nor U2293 (N_2293,N_862,N_497);
and U2294 (N_2294,N_942,N_1307);
or U2295 (N_2295,N_878,N_501);
nand U2296 (N_2296,N_1485,N_668);
xnor U2297 (N_2297,N_955,N_238);
and U2298 (N_2298,N_60,N_51);
nand U2299 (N_2299,N_1206,N_824);
nor U2300 (N_2300,N_732,N_176);
nand U2301 (N_2301,N_903,N_834);
xnor U2302 (N_2302,N_511,N_683);
nand U2303 (N_2303,N_320,N_938);
nand U2304 (N_2304,N_629,N_305);
nand U2305 (N_2305,N_358,N_1333);
and U2306 (N_2306,N_653,N_1323);
nand U2307 (N_2307,N_1178,N_89);
or U2308 (N_2308,N_984,N_190);
or U2309 (N_2309,N_1029,N_737);
xnor U2310 (N_2310,N_1105,N_1077);
or U2311 (N_2311,N_206,N_47);
nor U2312 (N_2312,N_643,N_1498);
nor U2313 (N_2313,N_327,N_367);
xnor U2314 (N_2314,N_577,N_177);
and U2315 (N_2315,N_1173,N_295);
and U2316 (N_2316,N_693,N_742);
nand U2317 (N_2317,N_738,N_1010);
xnor U2318 (N_2318,N_1323,N_1053);
and U2319 (N_2319,N_369,N_664);
nor U2320 (N_2320,N_1006,N_529);
nand U2321 (N_2321,N_469,N_318);
and U2322 (N_2322,N_168,N_568);
or U2323 (N_2323,N_707,N_637);
xnor U2324 (N_2324,N_527,N_270);
xnor U2325 (N_2325,N_64,N_1473);
xnor U2326 (N_2326,N_664,N_1477);
xor U2327 (N_2327,N_650,N_981);
or U2328 (N_2328,N_1005,N_188);
xor U2329 (N_2329,N_506,N_761);
nand U2330 (N_2330,N_1383,N_1401);
nor U2331 (N_2331,N_541,N_1307);
nor U2332 (N_2332,N_490,N_187);
xnor U2333 (N_2333,N_341,N_967);
and U2334 (N_2334,N_722,N_658);
or U2335 (N_2335,N_1090,N_1427);
nand U2336 (N_2336,N_31,N_1426);
and U2337 (N_2337,N_931,N_602);
and U2338 (N_2338,N_20,N_1118);
nand U2339 (N_2339,N_457,N_927);
and U2340 (N_2340,N_1179,N_112);
or U2341 (N_2341,N_1166,N_532);
nor U2342 (N_2342,N_1303,N_1025);
and U2343 (N_2343,N_538,N_1117);
nor U2344 (N_2344,N_209,N_1393);
nand U2345 (N_2345,N_1163,N_572);
or U2346 (N_2346,N_1154,N_1057);
nand U2347 (N_2347,N_1349,N_1118);
xor U2348 (N_2348,N_1495,N_1342);
nor U2349 (N_2349,N_13,N_58);
nand U2350 (N_2350,N_1430,N_923);
or U2351 (N_2351,N_432,N_904);
xor U2352 (N_2352,N_616,N_473);
or U2353 (N_2353,N_708,N_283);
xor U2354 (N_2354,N_279,N_61);
xnor U2355 (N_2355,N_1198,N_359);
or U2356 (N_2356,N_1497,N_394);
and U2357 (N_2357,N_943,N_1209);
nand U2358 (N_2358,N_1329,N_211);
nor U2359 (N_2359,N_467,N_351);
and U2360 (N_2360,N_1375,N_310);
xnor U2361 (N_2361,N_677,N_482);
nor U2362 (N_2362,N_1049,N_222);
and U2363 (N_2363,N_642,N_959);
nor U2364 (N_2364,N_241,N_1095);
xor U2365 (N_2365,N_921,N_1335);
xnor U2366 (N_2366,N_685,N_738);
or U2367 (N_2367,N_715,N_980);
and U2368 (N_2368,N_262,N_784);
xnor U2369 (N_2369,N_609,N_865);
xnor U2370 (N_2370,N_788,N_949);
and U2371 (N_2371,N_1315,N_1);
and U2372 (N_2372,N_1381,N_981);
or U2373 (N_2373,N_204,N_1061);
or U2374 (N_2374,N_967,N_608);
xor U2375 (N_2375,N_401,N_557);
nand U2376 (N_2376,N_165,N_655);
xor U2377 (N_2377,N_182,N_276);
nor U2378 (N_2378,N_258,N_313);
or U2379 (N_2379,N_428,N_742);
nand U2380 (N_2380,N_613,N_248);
nand U2381 (N_2381,N_1238,N_876);
or U2382 (N_2382,N_923,N_809);
and U2383 (N_2383,N_1159,N_389);
nor U2384 (N_2384,N_943,N_892);
nor U2385 (N_2385,N_1058,N_638);
nand U2386 (N_2386,N_510,N_116);
and U2387 (N_2387,N_1104,N_58);
or U2388 (N_2388,N_571,N_863);
nor U2389 (N_2389,N_1083,N_1399);
nor U2390 (N_2390,N_1140,N_264);
or U2391 (N_2391,N_235,N_703);
xor U2392 (N_2392,N_616,N_373);
or U2393 (N_2393,N_133,N_37);
nand U2394 (N_2394,N_1331,N_970);
and U2395 (N_2395,N_560,N_325);
and U2396 (N_2396,N_144,N_1327);
nor U2397 (N_2397,N_1147,N_98);
nor U2398 (N_2398,N_726,N_1067);
and U2399 (N_2399,N_188,N_959);
nor U2400 (N_2400,N_238,N_1433);
and U2401 (N_2401,N_977,N_824);
and U2402 (N_2402,N_1483,N_1344);
and U2403 (N_2403,N_1277,N_1063);
or U2404 (N_2404,N_1254,N_110);
or U2405 (N_2405,N_629,N_620);
nor U2406 (N_2406,N_164,N_1166);
nor U2407 (N_2407,N_375,N_5);
nand U2408 (N_2408,N_686,N_395);
and U2409 (N_2409,N_1000,N_1137);
nand U2410 (N_2410,N_1430,N_1080);
xor U2411 (N_2411,N_433,N_1019);
xnor U2412 (N_2412,N_29,N_324);
xor U2413 (N_2413,N_107,N_1371);
xor U2414 (N_2414,N_977,N_60);
nor U2415 (N_2415,N_650,N_1031);
and U2416 (N_2416,N_1172,N_1456);
or U2417 (N_2417,N_851,N_427);
or U2418 (N_2418,N_658,N_324);
xor U2419 (N_2419,N_1053,N_855);
and U2420 (N_2420,N_85,N_1354);
xor U2421 (N_2421,N_963,N_1188);
xnor U2422 (N_2422,N_82,N_37);
xor U2423 (N_2423,N_1106,N_255);
or U2424 (N_2424,N_1042,N_1314);
or U2425 (N_2425,N_748,N_1251);
nand U2426 (N_2426,N_959,N_1108);
xor U2427 (N_2427,N_1380,N_153);
and U2428 (N_2428,N_93,N_457);
or U2429 (N_2429,N_956,N_275);
nor U2430 (N_2430,N_756,N_559);
nor U2431 (N_2431,N_117,N_878);
nor U2432 (N_2432,N_44,N_1406);
or U2433 (N_2433,N_1355,N_346);
or U2434 (N_2434,N_558,N_729);
or U2435 (N_2435,N_979,N_917);
nor U2436 (N_2436,N_399,N_1322);
or U2437 (N_2437,N_872,N_854);
or U2438 (N_2438,N_75,N_471);
nor U2439 (N_2439,N_56,N_335);
nor U2440 (N_2440,N_1027,N_28);
xor U2441 (N_2441,N_1071,N_51);
nor U2442 (N_2442,N_1046,N_457);
nor U2443 (N_2443,N_877,N_331);
or U2444 (N_2444,N_1249,N_737);
xor U2445 (N_2445,N_752,N_379);
or U2446 (N_2446,N_1280,N_1433);
xnor U2447 (N_2447,N_150,N_569);
xnor U2448 (N_2448,N_1251,N_527);
xnor U2449 (N_2449,N_1263,N_75);
nor U2450 (N_2450,N_144,N_510);
and U2451 (N_2451,N_692,N_998);
nor U2452 (N_2452,N_1116,N_506);
nand U2453 (N_2453,N_441,N_1370);
or U2454 (N_2454,N_608,N_403);
nor U2455 (N_2455,N_1493,N_857);
or U2456 (N_2456,N_1155,N_889);
nor U2457 (N_2457,N_921,N_1258);
nand U2458 (N_2458,N_736,N_272);
xnor U2459 (N_2459,N_1167,N_601);
nor U2460 (N_2460,N_1248,N_949);
xor U2461 (N_2461,N_866,N_893);
nand U2462 (N_2462,N_958,N_1276);
nor U2463 (N_2463,N_532,N_154);
nor U2464 (N_2464,N_391,N_586);
xnor U2465 (N_2465,N_451,N_250);
and U2466 (N_2466,N_1197,N_191);
or U2467 (N_2467,N_2,N_336);
and U2468 (N_2468,N_310,N_198);
or U2469 (N_2469,N_1221,N_1324);
nor U2470 (N_2470,N_962,N_827);
or U2471 (N_2471,N_308,N_349);
xnor U2472 (N_2472,N_537,N_189);
nand U2473 (N_2473,N_86,N_214);
or U2474 (N_2474,N_194,N_1219);
nor U2475 (N_2475,N_1346,N_1032);
and U2476 (N_2476,N_168,N_470);
nor U2477 (N_2477,N_494,N_1353);
nor U2478 (N_2478,N_329,N_1085);
nor U2479 (N_2479,N_1237,N_540);
or U2480 (N_2480,N_1152,N_1270);
or U2481 (N_2481,N_434,N_126);
nor U2482 (N_2482,N_8,N_244);
nor U2483 (N_2483,N_1488,N_244);
or U2484 (N_2484,N_537,N_1203);
xnor U2485 (N_2485,N_1327,N_1365);
nand U2486 (N_2486,N_796,N_169);
or U2487 (N_2487,N_229,N_139);
nand U2488 (N_2488,N_1037,N_431);
nand U2489 (N_2489,N_263,N_471);
nor U2490 (N_2490,N_1040,N_408);
and U2491 (N_2491,N_82,N_1426);
and U2492 (N_2492,N_656,N_378);
or U2493 (N_2493,N_312,N_202);
and U2494 (N_2494,N_602,N_1023);
xor U2495 (N_2495,N_134,N_756);
nor U2496 (N_2496,N_995,N_1238);
nor U2497 (N_2497,N_744,N_483);
xor U2498 (N_2498,N_423,N_1411);
and U2499 (N_2499,N_918,N_1297);
nor U2500 (N_2500,N_667,N_34);
nand U2501 (N_2501,N_1474,N_997);
nor U2502 (N_2502,N_206,N_1);
nor U2503 (N_2503,N_1429,N_461);
or U2504 (N_2504,N_402,N_1472);
and U2505 (N_2505,N_1489,N_1094);
xor U2506 (N_2506,N_446,N_995);
xnor U2507 (N_2507,N_1276,N_736);
nor U2508 (N_2508,N_1473,N_989);
and U2509 (N_2509,N_1003,N_280);
xor U2510 (N_2510,N_751,N_110);
xor U2511 (N_2511,N_498,N_586);
nor U2512 (N_2512,N_667,N_1043);
nand U2513 (N_2513,N_1062,N_1268);
or U2514 (N_2514,N_14,N_54);
or U2515 (N_2515,N_891,N_90);
nand U2516 (N_2516,N_539,N_1038);
or U2517 (N_2517,N_625,N_839);
or U2518 (N_2518,N_961,N_447);
nand U2519 (N_2519,N_326,N_641);
and U2520 (N_2520,N_141,N_150);
nand U2521 (N_2521,N_580,N_152);
nor U2522 (N_2522,N_679,N_878);
and U2523 (N_2523,N_1000,N_1172);
nor U2524 (N_2524,N_113,N_1083);
and U2525 (N_2525,N_583,N_37);
or U2526 (N_2526,N_520,N_1051);
or U2527 (N_2527,N_552,N_214);
nor U2528 (N_2528,N_177,N_108);
and U2529 (N_2529,N_757,N_784);
nor U2530 (N_2530,N_38,N_1082);
nand U2531 (N_2531,N_82,N_187);
and U2532 (N_2532,N_1407,N_1474);
nor U2533 (N_2533,N_131,N_320);
nand U2534 (N_2534,N_1149,N_450);
and U2535 (N_2535,N_658,N_1133);
nand U2536 (N_2536,N_791,N_178);
xor U2537 (N_2537,N_1286,N_1252);
nor U2538 (N_2538,N_54,N_1391);
or U2539 (N_2539,N_638,N_278);
or U2540 (N_2540,N_148,N_604);
and U2541 (N_2541,N_1258,N_1292);
or U2542 (N_2542,N_1264,N_1098);
and U2543 (N_2543,N_1038,N_109);
or U2544 (N_2544,N_1334,N_609);
nand U2545 (N_2545,N_1118,N_184);
xnor U2546 (N_2546,N_1056,N_682);
nand U2547 (N_2547,N_421,N_900);
xnor U2548 (N_2548,N_665,N_834);
nand U2549 (N_2549,N_1073,N_42);
nand U2550 (N_2550,N_41,N_63);
or U2551 (N_2551,N_404,N_866);
and U2552 (N_2552,N_164,N_475);
nor U2553 (N_2553,N_1162,N_479);
or U2554 (N_2554,N_775,N_1196);
nor U2555 (N_2555,N_228,N_232);
or U2556 (N_2556,N_491,N_1066);
xor U2557 (N_2557,N_421,N_1005);
nor U2558 (N_2558,N_907,N_991);
and U2559 (N_2559,N_1134,N_32);
nand U2560 (N_2560,N_1241,N_882);
xnor U2561 (N_2561,N_774,N_1364);
nand U2562 (N_2562,N_1066,N_179);
xnor U2563 (N_2563,N_294,N_657);
and U2564 (N_2564,N_1033,N_142);
nor U2565 (N_2565,N_1371,N_962);
and U2566 (N_2566,N_250,N_717);
nor U2567 (N_2567,N_1291,N_715);
nor U2568 (N_2568,N_365,N_1307);
and U2569 (N_2569,N_1459,N_524);
nand U2570 (N_2570,N_575,N_1259);
nor U2571 (N_2571,N_1445,N_1314);
nand U2572 (N_2572,N_802,N_800);
nor U2573 (N_2573,N_63,N_430);
nand U2574 (N_2574,N_303,N_1353);
and U2575 (N_2575,N_80,N_726);
nor U2576 (N_2576,N_459,N_62);
xor U2577 (N_2577,N_734,N_1109);
nand U2578 (N_2578,N_1383,N_576);
and U2579 (N_2579,N_711,N_323);
or U2580 (N_2580,N_376,N_747);
and U2581 (N_2581,N_184,N_725);
xnor U2582 (N_2582,N_663,N_159);
xor U2583 (N_2583,N_712,N_1144);
or U2584 (N_2584,N_627,N_1030);
nor U2585 (N_2585,N_276,N_222);
or U2586 (N_2586,N_1121,N_781);
or U2587 (N_2587,N_254,N_591);
and U2588 (N_2588,N_564,N_1093);
nor U2589 (N_2589,N_1201,N_155);
nand U2590 (N_2590,N_98,N_830);
nor U2591 (N_2591,N_851,N_1365);
nor U2592 (N_2592,N_1049,N_932);
and U2593 (N_2593,N_1468,N_609);
or U2594 (N_2594,N_1320,N_605);
xor U2595 (N_2595,N_395,N_326);
nor U2596 (N_2596,N_602,N_1280);
or U2597 (N_2597,N_423,N_658);
or U2598 (N_2598,N_821,N_1306);
xor U2599 (N_2599,N_1371,N_1111);
or U2600 (N_2600,N_394,N_746);
nor U2601 (N_2601,N_969,N_1496);
xnor U2602 (N_2602,N_235,N_10);
nor U2603 (N_2603,N_225,N_889);
nor U2604 (N_2604,N_637,N_453);
and U2605 (N_2605,N_229,N_880);
xor U2606 (N_2606,N_189,N_841);
or U2607 (N_2607,N_1216,N_526);
nand U2608 (N_2608,N_658,N_1227);
nor U2609 (N_2609,N_1157,N_576);
nor U2610 (N_2610,N_220,N_23);
and U2611 (N_2611,N_355,N_536);
xnor U2612 (N_2612,N_1241,N_1327);
nand U2613 (N_2613,N_227,N_1343);
or U2614 (N_2614,N_934,N_461);
nor U2615 (N_2615,N_460,N_103);
nand U2616 (N_2616,N_992,N_993);
nand U2617 (N_2617,N_1456,N_559);
nor U2618 (N_2618,N_842,N_357);
and U2619 (N_2619,N_982,N_207);
and U2620 (N_2620,N_322,N_1427);
nand U2621 (N_2621,N_135,N_428);
nor U2622 (N_2622,N_952,N_923);
xnor U2623 (N_2623,N_449,N_1048);
or U2624 (N_2624,N_584,N_899);
or U2625 (N_2625,N_223,N_103);
or U2626 (N_2626,N_806,N_1296);
and U2627 (N_2627,N_1185,N_1078);
nand U2628 (N_2628,N_487,N_1354);
and U2629 (N_2629,N_261,N_439);
nor U2630 (N_2630,N_555,N_259);
xor U2631 (N_2631,N_773,N_1082);
and U2632 (N_2632,N_840,N_187);
or U2633 (N_2633,N_191,N_1060);
xor U2634 (N_2634,N_1148,N_1073);
or U2635 (N_2635,N_282,N_1160);
or U2636 (N_2636,N_1342,N_181);
nand U2637 (N_2637,N_1056,N_1161);
nand U2638 (N_2638,N_59,N_698);
or U2639 (N_2639,N_1275,N_141);
nor U2640 (N_2640,N_1279,N_189);
nor U2641 (N_2641,N_924,N_1428);
and U2642 (N_2642,N_501,N_617);
and U2643 (N_2643,N_602,N_1338);
nor U2644 (N_2644,N_1356,N_994);
or U2645 (N_2645,N_227,N_1292);
xnor U2646 (N_2646,N_136,N_1224);
xor U2647 (N_2647,N_150,N_56);
nor U2648 (N_2648,N_1388,N_151);
nand U2649 (N_2649,N_803,N_194);
xnor U2650 (N_2650,N_1458,N_1092);
and U2651 (N_2651,N_484,N_150);
xor U2652 (N_2652,N_1200,N_362);
or U2653 (N_2653,N_921,N_685);
nor U2654 (N_2654,N_1345,N_985);
and U2655 (N_2655,N_956,N_1207);
and U2656 (N_2656,N_835,N_563);
and U2657 (N_2657,N_35,N_1429);
nor U2658 (N_2658,N_783,N_1081);
or U2659 (N_2659,N_761,N_113);
nor U2660 (N_2660,N_1008,N_265);
and U2661 (N_2661,N_1290,N_501);
nor U2662 (N_2662,N_1440,N_1043);
nand U2663 (N_2663,N_264,N_589);
and U2664 (N_2664,N_1158,N_403);
nand U2665 (N_2665,N_928,N_85);
and U2666 (N_2666,N_170,N_1253);
or U2667 (N_2667,N_1451,N_1310);
and U2668 (N_2668,N_511,N_1205);
xnor U2669 (N_2669,N_1034,N_1299);
xnor U2670 (N_2670,N_1249,N_584);
nor U2671 (N_2671,N_1288,N_1105);
xnor U2672 (N_2672,N_1240,N_767);
nand U2673 (N_2673,N_43,N_691);
xnor U2674 (N_2674,N_180,N_1242);
nand U2675 (N_2675,N_205,N_209);
xor U2676 (N_2676,N_110,N_12);
and U2677 (N_2677,N_553,N_208);
and U2678 (N_2678,N_392,N_1012);
nor U2679 (N_2679,N_598,N_341);
nand U2680 (N_2680,N_274,N_339);
and U2681 (N_2681,N_137,N_1040);
xnor U2682 (N_2682,N_1330,N_1181);
and U2683 (N_2683,N_81,N_490);
xnor U2684 (N_2684,N_781,N_432);
nand U2685 (N_2685,N_1141,N_1059);
nand U2686 (N_2686,N_104,N_324);
and U2687 (N_2687,N_684,N_1100);
nor U2688 (N_2688,N_1023,N_449);
nor U2689 (N_2689,N_985,N_39);
nand U2690 (N_2690,N_49,N_1016);
nand U2691 (N_2691,N_736,N_1428);
or U2692 (N_2692,N_346,N_823);
or U2693 (N_2693,N_668,N_429);
and U2694 (N_2694,N_413,N_1442);
and U2695 (N_2695,N_629,N_1301);
nand U2696 (N_2696,N_598,N_18);
nand U2697 (N_2697,N_209,N_1223);
or U2698 (N_2698,N_233,N_1204);
and U2699 (N_2699,N_106,N_976);
nand U2700 (N_2700,N_419,N_1308);
and U2701 (N_2701,N_15,N_1246);
xnor U2702 (N_2702,N_339,N_334);
xor U2703 (N_2703,N_2,N_640);
xor U2704 (N_2704,N_707,N_775);
and U2705 (N_2705,N_239,N_1445);
nand U2706 (N_2706,N_1487,N_994);
nor U2707 (N_2707,N_1027,N_1074);
nand U2708 (N_2708,N_604,N_1479);
and U2709 (N_2709,N_718,N_558);
nand U2710 (N_2710,N_545,N_1406);
or U2711 (N_2711,N_992,N_298);
or U2712 (N_2712,N_385,N_713);
nor U2713 (N_2713,N_569,N_1065);
xor U2714 (N_2714,N_1160,N_1326);
nand U2715 (N_2715,N_112,N_220);
xor U2716 (N_2716,N_539,N_70);
or U2717 (N_2717,N_292,N_253);
xnor U2718 (N_2718,N_1235,N_1180);
or U2719 (N_2719,N_570,N_815);
nor U2720 (N_2720,N_191,N_1207);
xor U2721 (N_2721,N_1395,N_844);
xnor U2722 (N_2722,N_846,N_93);
xnor U2723 (N_2723,N_1312,N_65);
xor U2724 (N_2724,N_503,N_1175);
nand U2725 (N_2725,N_406,N_237);
and U2726 (N_2726,N_912,N_1447);
nor U2727 (N_2727,N_875,N_1174);
nor U2728 (N_2728,N_363,N_1064);
nor U2729 (N_2729,N_1293,N_1219);
nand U2730 (N_2730,N_33,N_431);
xnor U2731 (N_2731,N_701,N_995);
nand U2732 (N_2732,N_550,N_381);
xor U2733 (N_2733,N_801,N_268);
xor U2734 (N_2734,N_36,N_1453);
or U2735 (N_2735,N_890,N_875);
nand U2736 (N_2736,N_867,N_503);
nand U2737 (N_2737,N_231,N_65);
and U2738 (N_2738,N_1192,N_1397);
nand U2739 (N_2739,N_585,N_923);
or U2740 (N_2740,N_1148,N_214);
or U2741 (N_2741,N_935,N_728);
nand U2742 (N_2742,N_732,N_888);
xnor U2743 (N_2743,N_1091,N_178);
and U2744 (N_2744,N_626,N_1367);
xnor U2745 (N_2745,N_154,N_1127);
nor U2746 (N_2746,N_807,N_698);
and U2747 (N_2747,N_1462,N_989);
xor U2748 (N_2748,N_921,N_736);
xnor U2749 (N_2749,N_263,N_97);
and U2750 (N_2750,N_561,N_276);
or U2751 (N_2751,N_706,N_197);
nor U2752 (N_2752,N_971,N_1247);
xor U2753 (N_2753,N_180,N_931);
nand U2754 (N_2754,N_462,N_289);
xnor U2755 (N_2755,N_285,N_1154);
nand U2756 (N_2756,N_285,N_521);
nor U2757 (N_2757,N_808,N_777);
or U2758 (N_2758,N_709,N_1320);
nor U2759 (N_2759,N_386,N_757);
nand U2760 (N_2760,N_925,N_97);
and U2761 (N_2761,N_1399,N_908);
xnor U2762 (N_2762,N_756,N_1207);
nor U2763 (N_2763,N_742,N_662);
nand U2764 (N_2764,N_554,N_861);
xnor U2765 (N_2765,N_753,N_679);
nor U2766 (N_2766,N_654,N_368);
or U2767 (N_2767,N_549,N_342);
and U2768 (N_2768,N_1090,N_906);
nor U2769 (N_2769,N_1275,N_1087);
and U2770 (N_2770,N_276,N_979);
or U2771 (N_2771,N_1174,N_659);
nand U2772 (N_2772,N_1373,N_629);
and U2773 (N_2773,N_412,N_1401);
xnor U2774 (N_2774,N_1229,N_779);
nand U2775 (N_2775,N_1023,N_1367);
nand U2776 (N_2776,N_463,N_1298);
or U2777 (N_2777,N_775,N_508);
xnor U2778 (N_2778,N_762,N_453);
and U2779 (N_2779,N_63,N_815);
or U2780 (N_2780,N_1319,N_252);
and U2781 (N_2781,N_49,N_442);
xnor U2782 (N_2782,N_900,N_384);
and U2783 (N_2783,N_881,N_271);
nand U2784 (N_2784,N_291,N_463);
nand U2785 (N_2785,N_359,N_1435);
and U2786 (N_2786,N_1019,N_588);
nand U2787 (N_2787,N_139,N_792);
xnor U2788 (N_2788,N_1322,N_798);
xnor U2789 (N_2789,N_1075,N_794);
xor U2790 (N_2790,N_851,N_1119);
xor U2791 (N_2791,N_608,N_1452);
or U2792 (N_2792,N_498,N_299);
and U2793 (N_2793,N_844,N_694);
xnor U2794 (N_2794,N_125,N_808);
nand U2795 (N_2795,N_812,N_528);
nor U2796 (N_2796,N_890,N_282);
xnor U2797 (N_2797,N_936,N_1277);
xnor U2798 (N_2798,N_1499,N_81);
or U2799 (N_2799,N_1466,N_1038);
nand U2800 (N_2800,N_1479,N_174);
nand U2801 (N_2801,N_86,N_480);
nor U2802 (N_2802,N_946,N_97);
xnor U2803 (N_2803,N_57,N_1487);
nor U2804 (N_2804,N_527,N_767);
xnor U2805 (N_2805,N_241,N_303);
nor U2806 (N_2806,N_427,N_551);
nand U2807 (N_2807,N_1233,N_1087);
xnor U2808 (N_2808,N_1131,N_1415);
nand U2809 (N_2809,N_1077,N_44);
and U2810 (N_2810,N_1317,N_107);
or U2811 (N_2811,N_1064,N_1427);
nor U2812 (N_2812,N_25,N_1489);
nor U2813 (N_2813,N_937,N_1273);
nor U2814 (N_2814,N_1378,N_709);
nor U2815 (N_2815,N_1277,N_1280);
or U2816 (N_2816,N_348,N_524);
or U2817 (N_2817,N_1310,N_247);
nor U2818 (N_2818,N_1319,N_1499);
xor U2819 (N_2819,N_1187,N_1033);
or U2820 (N_2820,N_317,N_1008);
xor U2821 (N_2821,N_736,N_841);
xor U2822 (N_2822,N_792,N_848);
nand U2823 (N_2823,N_181,N_208);
or U2824 (N_2824,N_885,N_159);
nand U2825 (N_2825,N_1456,N_232);
xor U2826 (N_2826,N_1280,N_187);
and U2827 (N_2827,N_1262,N_115);
or U2828 (N_2828,N_937,N_500);
or U2829 (N_2829,N_1232,N_90);
nand U2830 (N_2830,N_1028,N_688);
or U2831 (N_2831,N_619,N_116);
and U2832 (N_2832,N_720,N_733);
and U2833 (N_2833,N_385,N_214);
nand U2834 (N_2834,N_884,N_750);
xnor U2835 (N_2835,N_699,N_1369);
xor U2836 (N_2836,N_334,N_206);
nand U2837 (N_2837,N_1240,N_1192);
and U2838 (N_2838,N_1365,N_795);
nand U2839 (N_2839,N_1457,N_1200);
and U2840 (N_2840,N_1252,N_654);
xor U2841 (N_2841,N_1213,N_120);
nand U2842 (N_2842,N_1474,N_480);
nor U2843 (N_2843,N_1281,N_1351);
or U2844 (N_2844,N_363,N_648);
xor U2845 (N_2845,N_1406,N_340);
or U2846 (N_2846,N_416,N_174);
xnor U2847 (N_2847,N_23,N_624);
or U2848 (N_2848,N_111,N_1094);
nand U2849 (N_2849,N_493,N_519);
and U2850 (N_2850,N_839,N_570);
nand U2851 (N_2851,N_544,N_1250);
or U2852 (N_2852,N_1331,N_554);
or U2853 (N_2853,N_876,N_784);
and U2854 (N_2854,N_1231,N_741);
xor U2855 (N_2855,N_401,N_835);
or U2856 (N_2856,N_1309,N_913);
xnor U2857 (N_2857,N_399,N_926);
xor U2858 (N_2858,N_334,N_827);
nand U2859 (N_2859,N_997,N_1436);
nor U2860 (N_2860,N_714,N_1333);
nand U2861 (N_2861,N_271,N_813);
nand U2862 (N_2862,N_768,N_965);
xor U2863 (N_2863,N_340,N_409);
and U2864 (N_2864,N_1041,N_991);
nand U2865 (N_2865,N_1209,N_679);
and U2866 (N_2866,N_178,N_455);
xor U2867 (N_2867,N_1491,N_1248);
or U2868 (N_2868,N_1277,N_1372);
nor U2869 (N_2869,N_833,N_1183);
nand U2870 (N_2870,N_640,N_140);
and U2871 (N_2871,N_1480,N_1358);
nor U2872 (N_2872,N_84,N_505);
xor U2873 (N_2873,N_1167,N_442);
nor U2874 (N_2874,N_919,N_1244);
nand U2875 (N_2875,N_351,N_204);
and U2876 (N_2876,N_961,N_725);
xor U2877 (N_2877,N_114,N_899);
nand U2878 (N_2878,N_831,N_1327);
xor U2879 (N_2879,N_766,N_1370);
xnor U2880 (N_2880,N_401,N_851);
nand U2881 (N_2881,N_324,N_318);
nand U2882 (N_2882,N_1018,N_1385);
and U2883 (N_2883,N_1291,N_1415);
xnor U2884 (N_2884,N_1112,N_618);
nor U2885 (N_2885,N_1125,N_43);
xor U2886 (N_2886,N_714,N_1416);
xor U2887 (N_2887,N_407,N_1406);
xor U2888 (N_2888,N_1217,N_832);
xor U2889 (N_2889,N_869,N_1137);
nor U2890 (N_2890,N_1125,N_943);
nand U2891 (N_2891,N_1117,N_162);
nor U2892 (N_2892,N_144,N_362);
xnor U2893 (N_2893,N_224,N_1408);
or U2894 (N_2894,N_1141,N_742);
and U2895 (N_2895,N_443,N_984);
or U2896 (N_2896,N_826,N_1006);
nor U2897 (N_2897,N_74,N_25);
nor U2898 (N_2898,N_339,N_765);
nand U2899 (N_2899,N_857,N_1294);
xor U2900 (N_2900,N_962,N_495);
nor U2901 (N_2901,N_1430,N_743);
nor U2902 (N_2902,N_1041,N_1100);
nand U2903 (N_2903,N_461,N_387);
nor U2904 (N_2904,N_1201,N_610);
nor U2905 (N_2905,N_101,N_1166);
nor U2906 (N_2906,N_1155,N_561);
nor U2907 (N_2907,N_342,N_1490);
and U2908 (N_2908,N_265,N_389);
nor U2909 (N_2909,N_1129,N_1110);
and U2910 (N_2910,N_606,N_1026);
nor U2911 (N_2911,N_1240,N_856);
xor U2912 (N_2912,N_1210,N_1198);
nand U2913 (N_2913,N_1443,N_1200);
nor U2914 (N_2914,N_288,N_113);
and U2915 (N_2915,N_380,N_156);
or U2916 (N_2916,N_952,N_1169);
nor U2917 (N_2917,N_347,N_758);
and U2918 (N_2918,N_684,N_753);
xnor U2919 (N_2919,N_1465,N_1058);
nor U2920 (N_2920,N_3,N_904);
or U2921 (N_2921,N_1173,N_943);
nor U2922 (N_2922,N_437,N_1401);
nor U2923 (N_2923,N_145,N_1041);
xor U2924 (N_2924,N_253,N_1375);
nor U2925 (N_2925,N_570,N_855);
or U2926 (N_2926,N_1228,N_1285);
nor U2927 (N_2927,N_818,N_975);
nand U2928 (N_2928,N_586,N_537);
xnor U2929 (N_2929,N_997,N_474);
nor U2930 (N_2930,N_1193,N_794);
or U2931 (N_2931,N_1160,N_1427);
and U2932 (N_2932,N_812,N_1434);
nand U2933 (N_2933,N_174,N_171);
xor U2934 (N_2934,N_216,N_1497);
nor U2935 (N_2935,N_936,N_707);
nand U2936 (N_2936,N_173,N_1208);
or U2937 (N_2937,N_370,N_1417);
nor U2938 (N_2938,N_123,N_905);
or U2939 (N_2939,N_79,N_642);
or U2940 (N_2940,N_587,N_203);
and U2941 (N_2941,N_39,N_1021);
and U2942 (N_2942,N_1065,N_243);
nand U2943 (N_2943,N_642,N_819);
or U2944 (N_2944,N_1197,N_13);
or U2945 (N_2945,N_1143,N_1237);
and U2946 (N_2946,N_1469,N_766);
xnor U2947 (N_2947,N_360,N_1381);
nor U2948 (N_2948,N_1063,N_1439);
and U2949 (N_2949,N_1376,N_1301);
and U2950 (N_2950,N_220,N_957);
nor U2951 (N_2951,N_490,N_121);
xor U2952 (N_2952,N_151,N_546);
and U2953 (N_2953,N_1329,N_1230);
nand U2954 (N_2954,N_637,N_813);
xor U2955 (N_2955,N_1149,N_1271);
or U2956 (N_2956,N_990,N_640);
nor U2957 (N_2957,N_707,N_407);
or U2958 (N_2958,N_743,N_1462);
or U2959 (N_2959,N_488,N_290);
or U2960 (N_2960,N_569,N_585);
nand U2961 (N_2961,N_1351,N_384);
and U2962 (N_2962,N_964,N_605);
nor U2963 (N_2963,N_793,N_575);
xor U2964 (N_2964,N_1396,N_388);
nand U2965 (N_2965,N_901,N_15);
xor U2966 (N_2966,N_910,N_1483);
xor U2967 (N_2967,N_591,N_1125);
or U2968 (N_2968,N_471,N_388);
xnor U2969 (N_2969,N_930,N_600);
nor U2970 (N_2970,N_272,N_739);
and U2971 (N_2971,N_119,N_448);
and U2972 (N_2972,N_1034,N_407);
nor U2973 (N_2973,N_710,N_281);
nor U2974 (N_2974,N_368,N_429);
nand U2975 (N_2975,N_1198,N_926);
nand U2976 (N_2976,N_44,N_942);
and U2977 (N_2977,N_1301,N_776);
or U2978 (N_2978,N_779,N_159);
nor U2979 (N_2979,N_207,N_1310);
and U2980 (N_2980,N_1030,N_883);
and U2981 (N_2981,N_1455,N_569);
and U2982 (N_2982,N_1099,N_1116);
nand U2983 (N_2983,N_400,N_228);
xor U2984 (N_2984,N_1376,N_747);
or U2985 (N_2985,N_998,N_252);
xor U2986 (N_2986,N_1213,N_803);
nand U2987 (N_2987,N_483,N_598);
or U2988 (N_2988,N_1059,N_570);
xor U2989 (N_2989,N_1122,N_495);
nor U2990 (N_2990,N_625,N_1093);
or U2991 (N_2991,N_1343,N_22);
nor U2992 (N_2992,N_380,N_1118);
and U2993 (N_2993,N_846,N_415);
xnor U2994 (N_2994,N_379,N_1139);
nand U2995 (N_2995,N_1009,N_1020);
nand U2996 (N_2996,N_596,N_431);
nor U2997 (N_2997,N_1090,N_266);
or U2998 (N_2998,N_1048,N_326);
or U2999 (N_2999,N_1125,N_689);
nor U3000 (N_3000,N_2072,N_2903);
xnor U3001 (N_3001,N_1824,N_2849);
nor U3002 (N_3002,N_1646,N_2214);
and U3003 (N_3003,N_2901,N_2125);
xor U3004 (N_3004,N_2477,N_2334);
and U3005 (N_3005,N_2142,N_2465);
xor U3006 (N_3006,N_1726,N_2019);
nand U3007 (N_3007,N_2170,N_2721);
xor U3008 (N_3008,N_1559,N_2107);
or U3009 (N_3009,N_2825,N_1744);
and U3010 (N_3010,N_1585,N_1718);
xnor U3011 (N_3011,N_1600,N_2470);
nand U3012 (N_3012,N_2444,N_2485);
nor U3013 (N_3013,N_1549,N_2947);
nor U3014 (N_3014,N_2191,N_2434);
and U3015 (N_3015,N_2504,N_2326);
xor U3016 (N_3016,N_1794,N_1916);
nand U3017 (N_3017,N_1759,N_2354);
and U3018 (N_3018,N_2548,N_2871);
nor U3019 (N_3019,N_1776,N_2023);
nand U3020 (N_3020,N_2858,N_1806);
xnor U3021 (N_3021,N_2300,N_2133);
and U3022 (N_3022,N_2843,N_1939);
nand U3023 (N_3023,N_2803,N_2076);
xor U3024 (N_3024,N_1842,N_1567);
nor U3025 (N_3025,N_1708,N_2801);
nor U3026 (N_3026,N_2447,N_1833);
xnor U3027 (N_3027,N_2051,N_2512);
or U3028 (N_3028,N_1642,N_2635);
nand U3029 (N_3029,N_2510,N_2831);
nand U3030 (N_3030,N_2840,N_2994);
xor U3031 (N_3031,N_2507,N_2774);
or U3032 (N_3032,N_2197,N_2511);
and U3033 (N_3033,N_2273,N_1778);
nor U3034 (N_3034,N_2698,N_2140);
or U3035 (N_3035,N_2254,N_1546);
nor U3036 (N_3036,N_2050,N_2755);
xor U3037 (N_3037,N_1922,N_2855);
and U3038 (N_3038,N_2285,N_1754);
nand U3039 (N_3039,N_2523,N_1690);
nor U3040 (N_3040,N_2491,N_1552);
or U3041 (N_3041,N_2976,N_1807);
or U3042 (N_3042,N_2531,N_2919);
xor U3043 (N_3043,N_2058,N_1520);
nor U3044 (N_3044,N_2405,N_2778);
or U3045 (N_3045,N_1563,N_2241);
nor U3046 (N_3046,N_2216,N_2645);
nor U3047 (N_3047,N_2668,N_1623);
and U3048 (N_3048,N_2671,N_2719);
nor U3049 (N_3049,N_2061,N_2094);
nor U3050 (N_3050,N_2652,N_2550);
xnor U3051 (N_3051,N_2717,N_1904);
xor U3052 (N_3052,N_1888,N_2638);
and U3053 (N_3053,N_2852,N_2987);
or U3054 (N_3054,N_2118,N_1606);
or U3055 (N_3055,N_2712,N_2562);
nand U3056 (N_3056,N_2875,N_2618);
nand U3057 (N_3057,N_2088,N_1680);
xor U3058 (N_3058,N_2806,N_1590);
nor U3059 (N_3059,N_2646,N_2603);
nand U3060 (N_3060,N_2406,N_2898);
nor U3061 (N_3061,N_1852,N_2879);
xor U3062 (N_3062,N_2839,N_2126);
xor U3063 (N_3063,N_1630,N_2993);
nand U3064 (N_3064,N_1899,N_1518);
nand U3065 (N_3065,N_2690,N_2832);
xnor U3066 (N_3066,N_2662,N_1709);
nor U3067 (N_3067,N_1535,N_1948);
xnor U3068 (N_3068,N_2538,N_1753);
nand U3069 (N_3069,N_2964,N_2078);
nor U3070 (N_3070,N_2581,N_2663);
xnor U3071 (N_3071,N_2372,N_1737);
or U3072 (N_3072,N_2614,N_2440);
or U3073 (N_3073,N_2678,N_2951);
nand U3074 (N_3074,N_2771,N_1588);
xor U3075 (N_3075,N_2367,N_2127);
nor U3076 (N_3076,N_2394,N_2894);
xor U3077 (N_3077,N_2242,N_2271);
xnor U3078 (N_3078,N_2555,N_2306);
nor U3079 (N_3079,N_1725,N_1942);
nor U3080 (N_3080,N_2817,N_1631);
or U3081 (N_3081,N_2761,N_1715);
or U3082 (N_3082,N_1777,N_1970);
nor U3083 (N_3083,N_2978,N_2457);
nor U3084 (N_3084,N_2380,N_1996);
nand U3085 (N_3085,N_1876,N_2720);
nor U3086 (N_3086,N_2469,N_2694);
xnor U3087 (N_3087,N_1789,N_2233);
or U3088 (N_3088,N_2945,N_1865);
nor U3089 (N_3089,N_1611,N_2033);
nand U3090 (N_3090,N_1637,N_2276);
xnor U3091 (N_3091,N_2456,N_1594);
or U3092 (N_3092,N_2842,N_2924);
or U3093 (N_3093,N_2159,N_2031);
or U3094 (N_3094,N_2569,N_1683);
nor U3095 (N_3095,N_1786,N_1528);
and U3096 (N_3096,N_2965,N_2734);
nand U3097 (N_3097,N_2578,N_2607);
nor U3098 (N_3098,N_1826,N_1873);
nor U3099 (N_3099,N_1539,N_2525);
xnor U3100 (N_3100,N_2151,N_2021);
or U3101 (N_3101,N_2350,N_2794);
or U3102 (N_3102,N_2356,N_2412);
or U3103 (N_3103,N_2480,N_1882);
nand U3104 (N_3104,N_1721,N_1908);
xor U3105 (N_3105,N_2907,N_2174);
nor U3106 (N_3106,N_1799,N_2290);
xnor U3107 (N_3107,N_2878,N_1943);
nor U3108 (N_3108,N_1764,N_2361);
xnor U3109 (N_3109,N_1858,N_2579);
nand U3110 (N_3110,N_2168,N_2758);
nand U3111 (N_3111,N_2837,N_1796);
nor U3112 (N_3112,N_1974,N_2410);
nor U3113 (N_3113,N_1868,N_1879);
and U3114 (N_3114,N_1657,N_2341);
nor U3115 (N_3115,N_1573,N_2561);
and U3116 (N_3116,N_2183,N_2181);
xnor U3117 (N_3117,N_2973,N_2369);
and U3118 (N_3118,N_2443,N_2235);
and U3119 (N_3119,N_2130,N_2592);
or U3120 (N_3120,N_2733,N_2606);
nor U3121 (N_3121,N_1790,N_1607);
and U3122 (N_3122,N_2495,N_2532);
nor U3123 (N_3123,N_1927,N_2808);
nor U3124 (N_3124,N_1689,N_2303);
and U3125 (N_3125,N_1719,N_2139);
xnor U3126 (N_3126,N_1638,N_2153);
nand U3127 (N_3127,N_2672,N_2725);
xor U3128 (N_3128,N_1554,N_1618);
nand U3129 (N_3129,N_2913,N_1728);
nor U3130 (N_3130,N_2805,N_2420);
xnor U3131 (N_3131,N_2403,N_1787);
nand U3132 (N_3132,N_2238,N_1906);
xor U3133 (N_3133,N_2368,N_2591);
nor U3134 (N_3134,N_1816,N_2529);
xnor U3135 (N_3135,N_2508,N_2650);
nand U3136 (N_3136,N_1811,N_2330);
nor U3137 (N_3137,N_2884,N_2038);
xnor U3138 (N_3138,N_2080,N_1932);
xor U3139 (N_3139,N_1980,N_1781);
nand U3140 (N_3140,N_2514,N_2902);
xor U3141 (N_3141,N_2689,N_2043);
nor U3142 (N_3142,N_2194,N_1757);
nand U3143 (N_3143,N_2188,N_2764);
and U3144 (N_3144,N_2044,N_2010);
nor U3145 (N_3145,N_2223,N_2685);
or U3146 (N_3146,N_2893,N_1964);
nand U3147 (N_3147,N_1902,N_2835);
and U3148 (N_3148,N_2732,N_2500);
and U3149 (N_3149,N_2066,N_1592);
nor U3150 (N_3150,N_1930,N_1666);
nand U3151 (N_3151,N_2353,N_1878);
nor U3152 (N_3152,N_2870,N_1752);
or U3153 (N_3153,N_1571,N_2693);
and U3154 (N_3154,N_1771,N_1991);
nand U3155 (N_3155,N_2282,N_1792);
xnor U3156 (N_3156,N_2718,N_2172);
nor U3157 (N_3157,N_2857,N_1524);
xor U3158 (N_3158,N_1541,N_2660);
nand U3159 (N_3159,N_1517,N_2397);
nor U3160 (N_3160,N_2200,N_2014);
or U3161 (N_3161,N_2929,N_2011);
xor U3162 (N_3162,N_2847,N_2438);
nor U3163 (N_3163,N_1863,N_1513);
xnor U3164 (N_3164,N_2358,N_2318);
xor U3165 (N_3165,N_1817,N_1534);
or U3166 (N_3166,N_2383,N_1733);
nor U3167 (N_3167,N_1751,N_1647);
xnor U3168 (N_3168,N_2583,N_2620);
or U3169 (N_3169,N_1820,N_2648);
or U3170 (N_3170,N_2070,N_1619);
and U3171 (N_3171,N_2983,N_1847);
and U3172 (N_3172,N_1921,N_1841);
xnor U3173 (N_3173,N_2960,N_2083);
or U3174 (N_3174,N_2441,N_2921);
or U3175 (N_3175,N_1783,N_2996);
nor U3176 (N_3176,N_2240,N_1960);
nor U3177 (N_3177,N_1562,N_2787);
xor U3178 (N_3178,N_1626,N_1971);
and U3179 (N_3179,N_2427,N_1660);
nand U3180 (N_3180,N_1707,N_2752);
and U3181 (N_3181,N_1935,N_2209);
nor U3182 (N_3182,N_2641,N_2486);
nor U3183 (N_3183,N_2656,N_2262);
and U3184 (N_3184,N_1953,N_2556);
or U3185 (N_3185,N_2553,N_2189);
or U3186 (N_3186,N_2888,N_2112);
or U3187 (N_3187,N_2811,N_1859);
nor U3188 (N_3188,N_2844,N_1684);
or U3189 (N_3189,N_2199,N_1749);
nand U3190 (N_3190,N_2498,N_2281);
and U3191 (N_3191,N_1890,N_1760);
xor U3192 (N_3192,N_1681,N_2552);
and U3193 (N_3193,N_2171,N_2476);
or U3194 (N_3194,N_2742,N_2756);
nand U3195 (N_3195,N_2782,N_2715);
or U3196 (N_3196,N_1654,N_1742);
or U3197 (N_3197,N_2325,N_2362);
nand U3198 (N_3198,N_2055,N_2777);
nand U3199 (N_3199,N_2316,N_2413);
or U3200 (N_3200,N_1695,N_2541);
and U3201 (N_3201,N_2751,N_1838);
nand U3202 (N_3202,N_2845,N_2925);
nand U3203 (N_3203,N_2331,N_1871);
and U3204 (N_3204,N_1987,N_2302);
xnor U3205 (N_3205,N_1941,N_1886);
xor U3206 (N_3206,N_2338,N_1913);
and U3207 (N_3207,N_2814,N_1765);
and U3208 (N_3208,N_1779,N_2201);
and U3209 (N_3209,N_2428,N_2882);
xnor U3210 (N_3210,N_1894,N_2270);
xor U3211 (N_3211,N_2539,N_2727);
or U3212 (N_3212,N_1636,N_2366);
nand U3213 (N_3213,N_2939,N_1505);
nor U3214 (N_3214,N_2386,N_2796);
nor U3215 (N_3215,N_2767,N_1625);
or U3216 (N_3216,N_1530,N_2248);
nand U3217 (N_3217,N_1989,N_2639);
xnor U3218 (N_3218,N_2624,N_2230);
xnor U3219 (N_3219,N_2816,N_2113);
nor U3220 (N_3220,N_2385,N_1555);
nand U3221 (N_3221,N_2173,N_2239);
or U3222 (N_3222,N_2997,N_2069);
nor U3223 (N_3223,N_2377,N_2398);
xnor U3224 (N_3224,N_1575,N_2838);
nand U3225 (N_3225,N_2545,N_2266);
or U3226 (N_3226,N_2707,N_2595);
xor U3227 (N_3227,N_1667,N_1724);
xnor U3228 (N_3228,N_2653,N_1810);
xnor U3229 (N_3229,N_2101,N_2243);
or U3230 (N_3230,N_2382,N_2518);
nor U3231 (N_3231,N_2169,N_2612);
nand U3232 (N_3232,N_2100,N_1525);
nand U3233 (N_3233,N_1761,N_2560);
xnor U3234 (N_3234,N_2793,N_1983);
xor U3235 (N_3235,N_2229,N_2609);
xor U3236 (N_3236,N_2926,N_1803);
or U3237 (N_3237,N_1542,N_2389);
or U3238 (N_3238,N_2096,N_2522);
and U3239 (N_3239,N_1584,N_2745);
nor U3240 (N_3240,N_2513,N_1531);
and U3241 (N_3241,N_1920,N_2575);
nand U3242 (N_3242,N_2679,N_1714);
nor U3243 (N_3243,N_2081,N_1540);
nor U3244 (N_3244,N_2880,N_2779);
xor U3245 (N_3245,N_2820,N_2889);
and U3246 (N_3246,N_1957,N_2472);
xnor U3247 (N_3247,N_1849,N_2952);
xor U3248 (N_3248,N_2824,N_2749);
nor U3249 (N_3249,N_2587,N_2310);
nor U3250 (N_3250,N_2809,N_1972);
and U3251 (N_3251,N_1992,N_1804);
nor U3252 (N_3252,N_2654,N_2846);
or U3253 (N_3253,N_2768,N_1523);
and U3254 (N_3254,N_2900,N_2259);
xnor U3255 (N_3255,N_2800,N_2706);
and U3256 (N_3256,N_2905,N_2527);
nand U3257 (N_3257,N_2815,N_1907);
xor U3258 (N_3258,N_2616,N_2766);
nand U3259 (N_3259,N_1832,N_1954);
and U3260 (N_3260,N_1627,N_2321);
and U3261 (N_3261,N_2705,N_1857);
xnor U3262 (N_3262,N_2425,N_2760);
xor U3263 (N_3263,N_2162,N_2798);
nor U3264 (N_3264,N_2322,N_2002);
nand U3265 (N_3265,N_1617,N_2821);
or U3266 (N_3266,N_2309,N_1526);
nand U3267 (N_3267,N_2328,N_2572);
xor U3268 (N_3268,N_2286,N_2417);
xor U3269 (N_3269,N_2301,N_2134);
xnor U3270 (N_3270,N_2292,N_2899);
and U3271 (N_3271,N_2505,N_2786);
and U3272 (N_3272,N_1864,N_2828);
and U3273 (N_3273,N_1880,N_1655);
or U3274 (N_3274,N_1984,N_2488);
and U3275 (N_3275,N_2812,N_2521);
and U3276 (N_3276,N_2936,N_1867);
xor U3277 (N_3277,N_2941,N_2267);
nand U3278 (N_3278,N_2883,N_2730);
and U3279 (N_3279,N_2818,N_2461);
or U3280 (N_3280,N_2559,N_2625);
xor U3281 (N_3281,N_2391,N_2454);
xor U3282 (N_3282,N_2458,N_2526);
nor U3283 (N_3283,N_1877,N_1965);
nand U3284 (N_3284,N_2891,N_1640);
or U3285 (N_3285,N_2208,N_2776);
xnor U3286 (N_3286,N_2601,N_1769);
and U3287 (N_3287,N_2493,N_1947);
xor U3288 (N_3288,N_2853,N_1860);
nand U3289 (N_3289,N_2363,N_1766);
xor U3290 (N_3290,N_2932,N_1755);
and U3291 (N_3291,N_2378,N_2017);
nand U3292 (N_3292,N_2365,N_1572);
nand U3293 (N_3293,N_2848,N_2633);
xor U3294 (N_3294,N_2288,N_2347);
nor U3295 (N_3295,N_2865,N_2789);
nand U3296 (N_3296,N_1767,N_1919);
nand U3297 (N_3297,N_1529,N_2258);
nand U3298 (N_3298,N_2748,N_2667);
or U3299 (N_3299,N_1918,N_2860);
nor U3300 (N_3300,N_2263,N_2364);
nand U3301 (N_3301,N_2851,N_1537);
nor U3302 (N_3302,N_1897,N_2664);
nor U3303 (N_3303,N_2773,N_2294);
xnor U3304 (N_3304,N_2205,N_2691);
xor U3305 (N_3305,N_2795,N_1874);
nand U3306 (N_3306,N_2016,N_1649);
or U3307 (N_3307,N_1967,N_1866);
nand U3308 (N_3308,N_2744,N_2215);
nor U3309 (N_3309,N_2497,N_2426);
nor U3310 (N_3310,N_2109,N_1604);
nand U3311 (N_3311,N_1955,N_1981);
xor U3312 (N_3312,N_2841,N_2203);
xnor U3313 (N_3313,N_2704,N_2605);
and U3314 (N_3314,N_1774,N_2154);
xor U3315 (N_3315,N_2179,N_2881);
or U3316 (N_3316,N_2830,N_2621);
nor U3317 (N_3317,N_1598,N_2103);
nor U3318 (N_3318,N_1521,N_2762);
xor U3319 (N_3319,N_1901,N_2807);
nand U3320 (N_3320,N_2953,N_1872);
nand U3321 (N_3321,N_2519,N_2687);
nand U3322 (N_3322,N_2264,N_2349);
or U3323 (N_3323,N_2178,N_2298);
or U3324 (N_3324,N_2990,N_1656);
nor U3325 (N_3325,N_2610,N_2731);
or U3326 (N_3326,N_1716,N_2079);
or U3327 (N_3327,N_2392,N_1973);
and U3328 (N_3328,N_2757,N_2729);
and U3329 (N_3329,N_1736,N_2192);
nand U3330 (N_3330,N_2770,N_2297);
nor U3331 (N_3331,N_1608,N_2797);
nand U3332 (N_3332,N_1925,N_1997);
nand U3333 (N_3333,N_2708,N_1545);
xnor U3334 (N_3334,N_2516,N_1602);
nor U3335 (N_3335,N_2063,N_2765);
and U3336 (N_3336,N_2743,N_2198);
nand U3337 (N_3337,N_1664,N_2145);
or U3338 (N_3338,N_1988,N_1805);
nand U3339 (N_3339,N_2370,N_2374);
xor U3340 (N_3340,N_2535,N_1976);
xnor U3341 (N_3341,N_2095,N_1732);
nor U3342 (N_3342,N_2916,N_2528);
xor U3343 (N_3343,N_2670,N_2437);
nor U3344 (N_3344,N_2152,N_2400);
nor U3345 (N_3345,N_1931,N_2041);
nor U3346 (N_3346,N_2682,N_2123);
nor U3347 (N_3347,N_2869,N_2092);
or U3348 (N_3348,N_1504,N_1565);
nor U3349 (N_3349,N_2904,N_2630);
nand U3350 (N_3350,N_1543,N_2336);
and U3351 (N_3351,N_2897,N_1959);
nor U3352 (N_3352,N_1924,N_1712);
xnor U3353 (N_3353,N_2661,N_2138);
nor U3354 (N_3354,N_2613,N_1854);
and U3355 (N_3355,N_2295,N_2911);
or U3356 (N_3356,N_2750,N_2564);
and U3357 (N_3357,N_1648,N_2928);
xnor U3358 (N_3358,N_2039,N_2132);
xor U3359 (N_3359,N_2335,N_1688);
xnor U3360 (N_3360,N_2826,N_1614);
or U3361 (N_3361,N_1516,N_1502);
nor U3362 (N_3362,N_2307,N_2804);
nand U3363 (N_3363,N_2915,N_2588);
nand U3364 (N_3364,N_1784,N_1853);
and U3365 (N_3365,N_1665,N_2675);
and U3366 (N_3366,N_2381,N_2022);
or U3367 (N_3367,N_2989,N_2008);
xor U3368 (N_3368,N_2917,N_2584);
and U3369 (N_3369,N_1809,N_2582);
and U3370 (N_3370,N_1962,N_2567);
xor U3371 (N_3371,N_2467,N_2332);
nand U3372 (N_3372,N_2702,N_2337);
or U3373 (N_3373,N_2202,N_1963);
nor U3374 (N_3374,N_2359,N_2542);
nor U3375 (N_3375,N_2728,N_2261);
and U3376 (N_3376,N_2455,N_2163);
or U3377 (N_3377,N_1578,N_2269);
nand U3378 (N_3378,N_1917,N_2868);
nor U3379 (N_3379,N_2981,N_1603);
nor U3380 (N_3380,N_2466,N_1861);
or U3381 (N_3381,N_2740,N_1643);
or U3382 (N_3382,N_2543,N_1933);
nand U3383 (N_3383,N_1912,N_2234);
or U3384 (N_3384,N_1591,N_2644);
and U3385 (N_3385,N_2020,N_2025);
xnor U3386 (N_3386,N_2217,N_2343);
nand U3387 (N_3387,N_2463,N_2950);
nand U3388 (N_3388,N_2390,N_1609);
nor U3389 (N_3389,N_2085,N_2040);
nor U3390 (N_3390,N_2655,N_2558);
and U3391 (N_3391,N_2714,N_2874);
xnor U3392 (N_3392,N_1628,N_2608);
and U3393 (N_3393,N_2348,N_2255);
xnor U3394 (N_3394,N_2710,N_2135);
and U3395 (N_3395,N_2352,N_2617);
xor U3396 (N_3396,N_1711,N_1685);
xnor U3397 (N_3397,N_2479,N_2090);
xor U3398 (N_3398,N_2161,N_2503);
and U3399 (N_3399,N_2864,N_1605);
nor U3400 (N_3400,N_1895,N_1507);
and U3401 (N_3401,N_2867,N_2697);
nor U3402 (N_3402,N_1610,N_1949);
xor U3403 (N_3403,N_2833,N_2036);
nand U3404 (N_3404,N_2231,N_2175);
xnor U3405 (N_3405,N_2885,N_1900);
and U3406 (N_3406,N_2464,N_2053);
and U3407 (N_3407,N_1560,N_2252);
xnor U3408 (N_3408,N_2696,N_2634);
or U3409 (N_3409,N_2411,N_2150);
nand U3410 (N_3410,N_2206,N_2204);
or U3411 (N_3411,N_1672,N_2184);
or U3412 (N_3412,N_1827,N_1893);
or U3413 (N_3413,N_1687,N_2896);
or U3414 (N_3414,N_1501,N_2709);
and U3415 (N_3415,N_2876,N_1550);
nor U3416 (N_3416,N_1652,N_2097);
nand U3417 (N_3417,N_2586,N_1936);
and U3418 (N_3418,N_2221,N_1875);
nand U3419 (N_3419,N_1999,N_2763);
or U3420 (N_3420,N_1812,N_1547);
nor U3421 (N_3421,N_1819,N_2923);
nand U3422 (N_3422,N_2753,N_2423);
or U3423 (N_3423,N_2345,N_2082);
and U3424 (N_3424,N_2439,N_2029);
xnor U3425 (N_3425,N_2738,N_2433);
or U3426 (N_3426,N_2278,N_2914);
and U3427 (N_3427,N_2086,N_1836);
xnor U3428 (N_3428,N_2813,N_1659);
xnor U3429 (N_3429,N_2665,N_1519);
nand U3430 (N_3430,N_1745,N_1994);
nand U3431 (N_3431,N_2546,N_1579);
and U3432 (N_3432,N_2388,N_2958);
nand U3433 (N_3433,N_2746,N_1596);
or U3434 (N_3434,N_2399,N_2959);
or U3435 (N_3435,N_2000,N_2317);
xnor U3436 (N_3436,N_2272,N_1883);
or U3437 (N_3437,N_1862,N_1693);
nand U3438 (N_3438,N_1780,N_2148);
xor U3439 (N_3439,N_1788,N_2449);
or U3440 (N_3440,N_1844,N_2596);
or U3441 (N_3441,N_2934,N_2442);
xnor U3442 (N_3442,N_2429,N_2649);
or U3443 (N_3443,N_2566,N_2030);
nor U3444 (N_3444,N_1723,N_1797);
and U3445 (N_3445,N_2260,N_1785);
xor U3446 (N_3446,N_2222,N_1775);
nand U3447 (N_3447,N_2157,N_2604);
nor U3448 (N_3448,N_2975,N_2481);
xnor U3449 (N_3449,N_2314,N_2320);
or U3450 (N_3450,N_2979,N_2384);
and U3451 (N_3451,N_2623,N_1696);
xnor U3452 (N_3452,N_1772,N_2506);
or U3453 (N_3453,N_2890,N_2501);
nand U3454 (N_3454,N_2339,N_2268);
or U3455 (N_3455,N_2071,N_2573);
xor U3456 (N_3456,N_1639,N_2593);
or U3457 (N_3457,N_2329,N_1599);
or U3458 (N_3458,N_1923,N_1892);
nand U3459 (N_3459,N_2909,N_2167);
xnor U3460 (N_3460,N_2013,N_2111);
or U3461 (N_3461,N_1944,N_2210);
nor U3462 (N_3462,N_2802,N_2279);
nand U3463 (N_3463,N_1750,N_1905);
xnor U3464 (N_3464,N_1977,N_1650);
nand U3465 (N_3465,N_1586,N_2473);
nor U3466 (N_3466,N_2699,N_1837);
and U3467 (N_3467,N_2676,N_1704);
and U3468 (N_3468,N_2557,N_1669);
and U3469 (N_3469,N_1583,N_2459);
xnor U3470 (N_3470,N_2783,N_2629);
nand U3471 (N_3471,N_2468,N_2536);
xnor U3472 (N_3472,N_1741,N_2483);
and U3473 (N_3473,N_1589,N_1632);
or U3474 (N_3474,N_1710,N_2120);
and U3475 (N_3475,N_1850,N_1763);
xor U3476 (N_3476,N_2251,N_2220);
and U3477 (N_3477,N_1705,N_1670);
nor U3478 (N_3478,N_2971,N_2948);
nor U3479 (N_3479,N_2462,N_1938);
or U3480 (N_3480,N_1722,N_2819);
xor U3481 (N_3481,N_2275,N_1730);
and U3482 (N_3482,N_2283,N_1522);
nor U3483 (N_3483,N_1979,N_2683);
or U3484 (N_3484,N_1808,N_2957);
and U3485 (N_3485,N_1674,N_2052);
nor U3486 (N_3486,N_2930,N_2432);
xnor U3487 (N_3487,N_2619,N_1958);
nor U3488 (N_3488,N_1597,N_2540);
or U3489 (N_3489,N_2492,N_2626);
and U3490 (N_3490,N_2908,N_1995);
nor U3491 (N_3491,N_2227,N_1851);
nor U3492 (N_3492,N_2961,N_2946);
or U3493 (N_3493,N_2128,N_2421);
nor U3494 (N_3494,N_1773,N_2657);
and U3495 (N_3495,N_2344,N_2747);
nor U3496 (N_3496,N_2435,N_2677);
or U3497 (N_3497,N_2713,N_2045);
and U3498 (N_3498,N_2057,N_2155);
nor U3499 (N_3499,N_1569,N_2077);
xor U3500 (N_3500,N_2450,N_2311);
and U3501 (N_3501,N_2219,N_2966);
or U3502 (N_3502,N_2108,N_2313);
nor U3503 (N_3503,N_2861,N_1830);
nand U3504 (N_3504,N_2622,N_2659);
or U3505 (N_3505,N_2549,N_1633);
nand U3506 (N_3506,N_1653,N_2954);
and U3507 (N_3507,N_2424,N_2177);
nor U3508 (N_3508,N_1701,N_1903);
nand U3509 (N_3509,N_1969,N_2315);
nand U3510 (N_3510,N_2631,N_2985);
nor U3511 (N_3511,N_2156,N_2115);
nand U3512 (N_3512,N_2247,N_2106);
and U3513 (N_3513,N_2299,N_1729);
xor U3514 (N_3514,N_1956,N_2565);
xor U3515 (N_3515,N_1746,N_2597);
xor U3516 (N_3516,N_2628,N_2418);
and U3517 (N_3517,N_2274,N_2093);
nand U3518 (N_3518,N_2680,N_2060);
nand U3519 (N_3519,N_2068,N_2836);
nand U3520 (N_3520,N_1740,N_2866);
or U3521 (N_3521,N_2212,N_2700);
nand U3522 (N_3522,N_1770,N_2143);
nand U3523 (N_3523,N_2207,N_1990);
nor U3524 (N_3524,N_1682,N_2489);
xor U3525 (N_3525,N_2598,N_1727);
nor U3526 (N_3526,N_2754,N_1511);
or U3527 (N_3527,N_2146,N_2974);
nor U3528 (N_3528,N_2387,N_1748);
or U3529 (N_3529,N_2688,N_2568);
nand U3530 (N_3530,N_1613,N_1512);
nor U3531 (N_3531,N_2674,N_2166);
xor U3532 (N_3532,N_2873,N_2006);
and U3533 (N_3533,N_1668,N_2360);
xor U3534 (N_3534,N_2788,N_1839);
nand U3535 (N_3535,N_2478,N_2373);
or U3536 (N_3536,N_1676,N_2007);
nand U3537 (N_3537,N_2415,N_1697);
nand U3538 (N_3538,N_2284,N_2375);
xor U3539 (N_3539,N_1885,N_2580);
and U3540 (N_3540,N_2600,N_1678);
nor U3541 (N_3541,N_2327,N_2611);
nand U3542 (N_3542,N_2533,N_2005);
and U3543 (N_3543,N_1782,N_1629);
nand U3544 (N_3544,N_1548,N_2594);
nor U3545 (N_3545,N_1574,N_2099);
xnor U3546 (N_3546,N_1926,N_2193);
nor U3547 (N_3547,N_2636,N_1961);
nand U3548 (N_3548,N_2723,N_2590);
nand U3549 (N_3549,N_2232,N_2445);
xnor U3550 (N_3550,N_2408,N_1570);
and U3551 (N_3551,N_2955,N_1762);
xnor U3552 (N_3552,N_1644,N_2371);
or U3553 (N_3553,N_2577,N_2035);
nor U3554 (N_3554,N_1793,N_1658);
xnor U3555 (N_3555,N_2969,N_2436);
nor U3556 (N_3556,N_2933,N_1679);
nand U3557 (N_3557,N_2859,N_2131);
nand U3558 (N_3558,N_2431,N_2158);
and U3559 (N_3559,N_1993,N_2346);
xnor U3560 (N_3560,N_2850,N_2182);
and U3561 (N_3561,N_2047,N_1692);
nand U3562 (N_3562,N_1595,N_2073);
xor U3563 (N_3563,N_2237,N_1536);
or U3564 (N_3564,N_1914,N_1580);
nor U3565 (N_3565,N_1934,N_1870);
or U3566 (N_3566,N_2487,N_2922);
nor U3567 (N_3567,N_1825,N_1673);
and U3568 (N_3568,N_2324,N_1896);
and U3569 (N_3569,N_2149,N_2213);
xor U3570 (N_3570,N_1587,N_2245);
nor U3571 (N_3571,N_2446,N_2340);
nand U3572 (N_3572,N_2810,N_1635);
nand U3573 (N_3573,N_1831,N_1663);
nand U3574 (N_3574,N_2342,N_1713);
xor U3575 (N_3575,N_1966,N_1514);
nor U3576 (N_3576,N_2827,N_2414);
and U3577 (N_3577,N_1564,N_2121);
nand U3578 (N_3578,N_2333,N_2416);
xnor U3579 (N_3579,N_2822,N_1508);
nand U3580 (N_3580,N_2669,N_1986);
xor U3581 (N_3581,N_1677,N_2854);
xnor U3582 (N_3582,N_1843,N_1577);
and U3583 (N_3583,N_2530,N_1702);
xor U3584 (N_3584,N_2164,N_2992);
or U3585 (N_3585,N_1940,N_2970);
and U3586 (N_3586,N_2906,N_2940);
xnor U3587 (N_3587,N_1978,N_2726);
xnor U3588 (N_3588,N_2910,N_2256);
xor U3589 (N_3589,N_2967,N_2912);
and U3590 (N_3590,N_1566,N_2576);
nand U3591 (N_3591,N_2895,N_2585);
or U3592 (N_3592,N_2537,N_1675);
xor U3593 (N_3593,N_1731,N_2640);
nor U3594 (N_3594,N_2091,N_2064);
and U3595 (N_3595,N_1510,N_1915);
or U3596 (N_3596,N_1945,N_1869);
xnor U3597 (N_3597,N_2937,N_1662);
xor U3598 (N_3598,N_2862,N_2666);
or U3599 (N_3599,N_2393,N_2872);
nand U3600 (N_3600,N_2737,N_1829);
and U3601 (N_3601,N_1509,N_1982);
or U3602 (N_3602,N_2037,N_2474);
xor U3603 (N_3603,N_2938,N_2376);
and U3604 (N_3604,N_1814,N_2059);
or U3605 (N_3605,N_2034,N_2351);
xnor U3606 (N_3606,N_1848,N_2571);
nand U3607 (N_3607,N_2032,N_2995);
and U3608 (N_3608,N_2551,N_1576);
or U3609 (N_3609,N_1985,N_1641);
or U3610 (N_3610,N_2949,N_2249);
or U3611 (N_3611,N_1756,N_2105);
or U3612 (N_3612,N_1700,N_2716);
nor U3613 (N_3613,N_2942,N_2141);
nand U3614 (N_3614,N_2599,N_1855);
xnor U3615 (N_3615,N_2520,N_2003);
and U3616 (N_3616,N_2863,N_1717);
nand U3617 (N_3617,N_2308,N_2102);
xnor U3618 (N_3618,N_2496,N_1691);
nand U3619 (N_3619,N_2026,N_2015);
nor U3620 (N_3620,N_2452,N_1568);
and U3621 (N_3621,N_2291,N_1634);
and U3622 (N_3622,N_2602,N_2956);
or U3623 (N_3623,N_2736,N_2253);
xor U3624 (N_3624,N_1840,N_2739);
or U3625 (N_3625,N_1558,N_1735);
xnor U3626 (N_3626,N_1800,N_1821);
nor U3627 (N_3627,N_2190,N_1557);
nand U3628 (N_3628,N_2165,N_2293);
xnor U3629 (N_3629,N_1527,N_1823);
nand U3630 (N_3630,N_2877,N_2554);
and U3631 (N_3631,N_2935,N_2658);
nor U3632 (N_3632,N_2475,N_2196);
nand U3633 (N_3633,N_2228,N_1845);
nor U3634 (N_3634,N_1612,N_2892);
or U3635 (N_3635,N_2048,N_2074);
nand U3636 (N_3636,N_2009,N_2104);
or U3637 (N_3637,N_2185,N_1891);
nand U3638 (N_3638,N_2963,N_2430);
and U3639 (N_3639,N_2018,N_1556);
nand U3640 (N_3640,N_1856,N_2695);
and U3641 (N_3641,N_1616,N_1881);
nand U3642 (N_3642,N_2004,N_1835);
or U3643 (N_3643,N_1544,N_2117);
nor U3644 (N_3644,N_1515,N_1791);
or U3645 (N_3645,N_2401,N_2065);
nor U3646 (N_3646,N_2887,N_2116);
nor U3647 (N_3647,N_2986,N_2790);
nor U3648 (N_3648,N_2920,N_2280);
nand U3649 (N_3649,N_2570,N_2110);
nor U3650 (N_3650,N_2490,N_1828);
nand U3651 (N_3651,N_2049,N_1738);
nor U3652 (N_3652,N_2012,N_2927);
nand U3653 (N_3653,N_1889,N_1929);
and U3654 (N_3654,N_2067,N_2195);
and U3655 (N_3655,N_1706,N_2775);
xor U3656 (N_3656,N_1551,N_2277);
xor U3657 (N_3657,N_2451,N_2544);
nor U3658 (N_3658,N_2673,N_2176);
xnor U3659 (N_3659,N_2834,N_2792);
and U3660 (N_3660,N_2323,N_2651);
xnor U3661 (N_3661,N_2265,N_1952);
nor U3662 (N_3662,N_2524,N_1975);
nor U3663 (N_3663,N_1822,N_2692);
or U3664 (N_3664,N_1911,N_1743);
nand U3665 (N_3665,N_2943,N_2799);
nor U3666 (N_3666,N_2056,N_1801);
xor U3667 (N_3667,N_2124,N_2735);
xor U3668 (N_3668,N_2711,N_2484);
nor U3669 (N_3669,N_2647,N_2147);
nor U3670 (N_3670,N_1802,N_2257);
nand U3671 (N_3671,N_1720,N_1834);
or U3672 (N_3672,N_2547,N_2046);
nor U3673 (N_3673,N_2098,N_1968);
or U3674 (N_3674,N_2991,N_1818);
nor U3675 (N_3675,N_2759,N_1694);
nor U3676 (N_3676,N_2615,N_2589);
or U3677 (N_3677,N_2225,N_1532);
nand U3678 (N_3678,N_1699,N_2296);
and U3679 (N_3679,N_1651,N_1898);
or U3680 (N_3680,N_2988,N_2355);
or U3681 (N_3681,N_2681,N_2144);
or U3682 (N_3682,N_2114,N_1621);
and U3683 (N_3683,N_1703,N_2305);
nor U3684 (N_3684,N_2319,N_2471);
xnor U3685 (N_3685,N_1937,N_2534);
and U3686 (N_3686,N_2407,N_2042);
or U3687 (N_3687,N_1661,N_2404);
nor U3688 (N_3688,N_1910,N_1500);
nand U3689 (N_3689,N_2419,N_1946);
nand U3690 (N_3690,N_1561,N_2395);
nand U3691 (N_3691,N_2001,N_2998);
nor U3692 (N_3692,N_2509,N_1795);
xnor U3693 (N_3693,N_2244,N_2304);
and U3694 (N_3694,N_1645,N_1747);
nor U3695 (N_3695,N_1768,N_2823);
nor U3696 (N_3696,N_2999,N_1739);
nor U3697 (N_3697,N_2980,N_2062);
and U3698 (N_3698,N_1686,N_1593);
nor U3699 (N_3699,N_1758,N_2722);
xor U3700 (N_3700,N_2396,N_2218);
nor U3701 (N_3701,N_1533,N_2944);
nand U3702 (N_3702,N_2517,N_2226);
xor U3703 (N_3703,N_2856,N_1951);
nor U3704 (N_3704,N_1622,N_2287);
nand U3705 (N_3705,N_1601,N_2357);
and U3706 (N_3706,N_2637,N_2977);
or U3707 (N_3707,N_1813,N_1998);
or U3708 (N_3708,N_1909,N_1581);
or U3709 (N_3709,N_1798,N_2027);
nand U3710 (N_3710,N_2499,N_2563);
or U3711 (N_3711,N_2701,N_2502);
nor U3712 (N_3712,N_2482,N_1615);
and U3713 (N_3713,N_2780,N_1884);
or U3714 (N_3714,N_1928,N_2643);
nor U3715 (N_3715,N_2180,N_2187);
xor U3716 (N_3716,N_2236,N_1620);
or U3717 (N_3717,N_2186,N_2289);
or U3718 (N_3718,N_2379,N_2984);
nor U3719 (N_3719,N_2402,N_2028);
or U3720 (N_3720,N_1698,N_2211);
nor U3721 (N_3721,N_2972,N_2409);
nand U3722 (N_3722,N_2224,N_1815);
xor U3723 (N_3723,N_2460,N_1503);
or U3724 (N_3724,N_1553,N_2246);
nor U3725 (N_3725,N_2087,N_2024);
nand U3726 (N_3726,N_2772,N_2129);
nor U3727 (N_3727,N_2075,N_2724);
and U3728 (N_3728,N_2741,N_2119);
nand U3729 (N_3729,N_1734,N_1887);
or U3730 (N_3730,N_1624,N_2084);
or U3731 (N_3731,N_2791,N_2137);
nor U3732 (N_3732,N_2632,N_2684);
or U3733 (N_3733,N_1846,N_2886);
nand U3734 (N_3734,N_2250,N_2781);
or U3735 (N_3735,N_2160,N_2122);
or U3736 (N_3736,N_2982,N_2769);
xnor U3737 (N_3737,N_2054,N_2784);
and U3738 (N_3738,N_2642,N_1506);
xnor U3739 (N_3739,N_2785,N_2627);
xor U3740 (N_3740,N_2136,N_1582);
nor U3741 (N_3741,N_2494,N_2453);
or U3742 (N_3742,N_1950,N_2312);
or U3743 (N_3743,N_2968,N_2703);
nor U3744 (N_3744,N_2918,N_2931);
xnor U3745 (N_3745,N_2574,N_2686);
xor U3746 (N_3746,N_2089,N_1538);
xor U3747 (N_3747,N_1671,N_2515);
and U3748 (N_3748,N_2829,N_2962);
xnor U3749 (N_3749,N_2448,N_2422);
or U3750 (N_3750,N_1516,N_2289);
or U3751 (N_3751,N_1953,N_1660);
nor U3752 (N_3752,N_1590,N_2226);
xnor U3753 (N_3753,N_2553,N_1562);
nor U3754 (N_3754,N_2868,N_2227);
nand U3755 (N_3755,N_2931,N_2464);
or U3756 (N_3756,N_1831,N_2308);
and U3757 (N_3757,N_1515,N_2857);
and U3758 (N_3758,N_2305,N_1581);
and U3759 (N_3759,N_1813,N_2011);
nor U3760 (N_3760,N_1543,N_1629);
and U3761 (N_3761,N_2660,N_2530);
nor U3762 (N_3762,N_2720,N_2385);
nand U3763 (N_3763,N_2132,N_2550);
nand U3764 (N_3764,N_1654,N_2703);
nand U3765 (N_3765,N_2024,N_2914);
nor U3766 (N_3766,N_1648,N_2734);
or U3767 (N_3767,N_2653,N_2790);
nor U3768 (N_3768,N_2051,N_1618);
nand U3769 (N_3769,N_2555,N_1800);
nand U3770 (N_3770,N_2494,N_2052);
or U3771 (N_3771,N_1734,N_2211);
nor U3772 (N_3772,N_1716,N_1626);
and U3773 (N_3773,N_1865,N_1633);
nor U3774 (N_3774,N_2281,N_2670);
or U3775 (N_3775,N_1867,N_2569);
xor U3776 (N_3776,N_2572,N_1529);
nor U3777 (N_3777,N_2926,N_2734);
and U3778 (N_3778,N_2605,N_2275);
xor U3779 (N_3779,N_2437,N_2355);
nor U3780 (N_3780,N_1666,N_2954);
nor U3781 (N_3781,N_2644,N_2327);
nor U3782 (N_3782,N_2106,N_1880);
nand U3783 (N_3783,N_2708,N_2340);
or U3784 (N_3784,N_1669,N_2842);
and U3785 (N_3785,N_2881,N_2060);
nand U3786 (N_3786,N_2351,N_2186);
or U3787 (N_3787,N_2351,N_2867);
or U3788 (N_3788,N_2920,N_2864);
and U3789 (N_3789,N_2450,N_2613);
xnor U3790 (N_3790,N_2729,N_2538);
and U3791 (N_3791,N_1855,N_2861);
nor U3792 (N_3792,N_1917,N_2891);
nor U3793 (N_3793,N_2642,N_2626);
or U3794 (N_3794,N_2519,N_2791);
nand U3795 (N_3795,N_1785,N_2943);
nand U3796 (N_3796,N_1577,N_2021);
and U3797 (N_3797,N_2124,N_2650);
nor U3798 (N_3798,N_2443,N_2699);
nor U3799 (N_3799,N_2193,N_1955);
and U3800 (N_3800,N_2676,N_2442);
xnor U3801 (N_3801,N_2029,N_1963);
xnor U3802 (N_3802,N_2664,N_2650);
nor U3803 (N_3803,N_1970,N_2868);
or U3804 (N_3804,N_1607,N_2311);
or U3805 (N_3805,N_1978,N_2519);
nor U3806 (N_3806,N_1731,N_2886);
nor U3807 (N_3807,N_2320,N_1778);
or U3808 (N_3808,N_1522,N_1520);
and U3809 (N_3809,N_1896,N_2831);
nand U3810 (N_3810,N_2959,N_2552);
and U3811 (N_3811,N_2071,N_2186);
and U3812 (N_3812,N_1948,N_1566);
or U3813 (N_3813,N_2905,N_2501);
xor U3814 (N_3814,N_2895,N_2315);
nor U3815 (N_3815,N_2017,N_1788);
xor U3816 (N_3816,N_2643,N_1887);
and U3817 (N_3817,N_1857,N_2819);
or U3818 (N_3818,N_2802,N_1915);
xor U3819 (N_3819,N_2243,N_2190);
and U3820 (N_3820,N_2623,N_2288);
or U3821 (N_3821,N_1861,N_1707);
nand U3822 (N_3822,N_1820,N_2791);
nor U3823 (N_3823,N_2627,N_1838);
or U3824 (N_3824,N_2302,N_2819);
and U3825 (N_3825,N_2005,N_2210);
nand U3826 (N_3826,N_2791,N_2439);
and U3827 (N_3827,N_1601,N_2419);
nor U3828 (N_3828,N_2023,N_2770);
or U3829 (N_3829,N_1677,N_2721);
or U3830 (N_3830,N_1661,N_2839);
nor U3831 (N_3831,N_2195,N_2644);
nor U3832 (N_3832,N_2904,N_1833);
nor U3833 (N_3833,N_2213,N_2828);
nand U3834 (N_3834,N_2440,N_1745);
or U3835 (N_3835,N_2897,N_2240);
nand U3836 (N_3836,N_2036,N_1540);
nand U3837 (N_3837,N_2381,N_1681);
and U3838 (N_3838,N_2584,N_2225);
or U3839 (N_3839,N_1681,N_2104);
or U3840 (N_3840,N_1952,N_2284);
and U3841 (N_3841,N_2375,N_1792);
and U3842 (N_3842,N_2621,N_2398);
or U3843 (N_3843,N_2791,N_2598);
or U3844 (N_3844,N_1610,N_2479);
nor U3845 (N_3845,N_2694,N_1633);
nand U3846 (N_3846,N_1620,N_2518);
nor U3847 (N_3847,N_2961,N_2872);
and U3848 (N_3848,N_2071,N_1859);
nor U3849 (N_3849,N_2674,N_1850);
nor U3850 (N_3850,N_2918,N_2350);
nand U3851 (N_3851,N_2323,N_2372);
and U3852 (N_3852,N_2388,N_2031);
or U3853 (N_3853,N_1574,N_2926);
and U3854 (N_3854,N_2030,N_2023);
nand U3855 (N_3855,N_2415,N_1708);
nand U3856 (N_3856,N_1802,N_2093);
nand U3857 (N_3857,N_1872,N_1979);
nor U3858 (N_3858,N_2496,N_2610);
and U3859 (N_3859,N_2542,N_2404);
xor U3860 (N_3860,N_2267,N_2920);
and U3861 (N_3861,N_2069,N_2775);
nor U3862 (N_3862,N_1825,N_2491);
xnor U3863 (N_3863,N_2463,N_2792);
or U3864 (N_3864,N_2612,N_1726);
xnor U3865 (N_3865,N_1597,N_2463);
nand U3866 (N_3866,N_2364,N_2994);
xor U3867 (N_3867,N_2330,N_2045);
nor U3868 (N_3868,N_2305,N_1898);
xnor U3869 (N_3869,N_1695,N_2333);
nor U3870 (N_3870,N_2177,N_1870);
and U3871 (N_3871,N_2961,N_1611);
xor U3872 (N_3872,N_2170,N_2473);
xnor U3873 (N_3873,N_1966,N_2107);
nor U3874 (N_3874,N_1915,N_1566);
xnor U3875 (N_3875,N_1732,N_2066);
xnor U3876 (N_3876,N_2403,N_1682);
or U3877 (N_3877,N_2642,N_2023);
nand U3878 (N_3878,N_1900,N_2673);
nor U3879 (N_3879,N_2494,N_1968);
nor U3880 (N_3880,N_2654,N_2590);
xor U3881 (N_3881,N_2536,N_1904);
nor U3882 (N_3882,N_1879,N_2250);
xor U3883 (N_3883,N_2182,N_1623);
nor U3884 (N_3884,N_2806,N_2040);
or U3885 (N_3885,N_1519,N_2426);
nor U3886 (N_3886,N_2503,N_2382);
nand U3887 (N_3887,N_2017,N_2996);
xor U3888 (N_3888,N_2094,N_2458);
and U3889 (N_3889,N_2352,N_1694);
or U3890 (N_3890,N_2510,N_1519);
xor U3891 (N_3891,N_2041,N_2211);
nor U3892 (N_3892,N_2894,N_2296);
and U3893 (N_3893,N_2099,N_2124);
nand U3894 (N_3894,N_1969,N_2277);
and U3895 (N_3895,N_2876,N_2552);
nand U3896 (N_3896,N_1864,N_2176);
nor U3897 (N_3897,N_2688,N_2146);
nand U3898 (N_3898,N_1977,N_1717);
xnor U3899 (N_3899,N_1627,N_2206);
or U3900 (N_3900,N_2471,N_2796);
xnor U3901 (N_3901,N_2686,N_2301);
nand U3902 (N_3902,N_2660,N_2439);
nand U3903 (N_3903,N_1573,N_2485);
or U3904 (N_3904,N_2687,N_2444);
nor U3905 (N_3905,N_1808,N_2230);
xnor U3906 (N_3906,N_2137,N_1679);
or U3907 (N_3907,N_2926,N_1794);
or U3908 (N_3908,N_2272,N_1645);
nor U3909 (N_3909,N_1659,N_2587);
or U3910 (N_3910,N_1729,N_1536);
nand U3911 (N_3911,N_2702,N_2517);
nor U3912 (N_3912,N_1528,N_2486);
nand U3913 (N_3913,N_2658,N_1863);
nand U3914 (N_3914,N_2074,N_2521);
and U3915 (N_3915,N_1949,N_2400);
xnor U3916 (N_3916,N_1796,N_1928);
or U3917 (N_3917,N_1512,N_2068);
xnor U3918 (N_3918,N_1557,N_1977);
or U3919 (N_3919,N_2584,N_2386);
nand U3920 (N_3920,N_1505,N_1543);
nor U3921 (N_3921,N_2283,N_2692);
or U3922 (N_3922,N_2636,N_2501);
and U3923 (N_3923,N_1832,N_2637);
and U3924 (N_3924,N_2422,N_2263);
or U3925 (N_3925,N_2778,N_2874);
and U3926 (N_3926,N_2233,N_1794);
and U3927 (N_3927,N_2102,N_1775);
and U3928 (N_3928,N_2608,N_2459);
nand U3929 (N_3929,N_1717,N_2700);
xor U3930 (N_3930,N_1883,N_2108);
nand U3931 (N_3931,N_1764,N_2516);
or U3932 (N_3932,N_2410,N_1534);
xnor U3933 (N_3933,N_2898,N_1794);
nand U3934 (N_3934,N_2187,N_1612);
and U3935 (N_3935,N_2769,N_2570);
or U3936 (N_3936,N_2462,N_2878);
or U3937 (N_3937,N_2952,N_2116);
xor U3938 (N_3938,N_2075,N_2828);
nor U3939 (N_3939,N_2128,N_1579);
xnor U3940 (N_3940,N_1522,N_2643);
or U3941 (N_3941,N_2817,N_2057);
nor U3942 (N_3942,N_2832,N_2109);
and U3943 (N_3943,N_1894,N_2937);
and U3944 (N_3944,N_2434,N_2285);
or U3945 (N_3945,N_2174,N_2570);
or U3946 (N_3946,N_2033,N_2042);
xor U3947 (N_3947,N_2302,N_2728);
nand U3948 (N_3948,N_1734,N_2832);
and U3949 (N_3949,N_1501,N_2954);
nor U3950 (N_3950,N_2064,N_2003);
or U3951 (N_3951,N_2244,N_1989);
and U3952 (N_3952,N_2143,N_2519);
and U3953 (N_3953,N_2294,N_2965);
nand U3954 (N_3954,N_1687,N_1604);
nor U3955 (N_3955,N_1852,N_1803);
xor U3956 (N_3956,N_1825,N_2321);
nand U3957 (N_3957,N_2482,N_2286);
and U3958 (N_3958,N_2781,N_2979);
or U3959 (N_3959,N_2254,N_2571);
nand U3960 (N_3960,N_2361,N_2433);
nor U3961 (N_3961,N_2294,N_2680);
or U3962 (N_3962,N_2955,N_2633);
and U3963 (N_3963,N_1619,N_1729);
nand U3964 (N_3964,N_2124,N_1954);
or U3965 (N_3965,N_1862,N_2731);
xnor U3966 (N_3966,N_1713,N_1867);
and U3967 (N_3967,N_2316,N_2305);
nand U3968 (N_3968,N_2472,N_1793);
nand U3969 (N_3969,N_2901,N_1707);
xor U3970 (N_3970,N_2333,N_2122);
xnor U3971 (N_3971,N_1550,N_2840);
xor U3972 (N_3972,N_2850,N_2666);
nor U3973 (N_3973,N_2517,N_2532);
or U3974 (N_3974,N_1593,N_1699);
nand U3975 (N_3975,N_2800,N_2709);
nand U3976 (N_3976,N_2899,N_2192);
nand U3977 (N_3977,N_1922,N_1652);
and U3978 (N_3978,N_1789,N_1559);
or U3979 (N_3979,N_2073,N_2825);
or U3980 (N_3980,N_2533,N_2389);
and U3981 (N_3981,N_1666,N_2811);
xnor U3982 (N_3982,N_2009,N_2560);
nor U3983 (N_3983,N_2848,N_1532);
and U3984 (N_3984,N_1871,N_2530);
xor U3985 (N_3985,N_2804,N_1648);
nand U3986 (N_3986,N_2267,N_2355);
or U3987 (N_3987,N_1694,N_1730);
or U3988 (N_3988,N_2226,N_2912);
xnor U3989 (N_3989,N_2930,N_2080);
xor U3990 (N_3990,N_2351,N_2072);
and U3991 (N_3991,N_2154,N_1764);
or U3992 (N_3992,N_2235,N_2157);
and U3993 (N_3993,N_2796,N_2887);
or U3994 (N_3994,N_2852,N_2285);
nand U3995 (N_3995,N_2125,N_1534);
xnor U3996 (N_3996,N_1804,N_2972);
and U3997 (N_3997,N_2958,N_1995);
nor U3998 (N_3998,N_1898,N_1710);
or U3999 (N_3999,N_2154,N_1629);
xnor U4000 (N_4000,N_1682,N_2945);
or U4001 (N_4001,N_2306,N_2726);
nor U4002 (N_4002,N_2687,N_2955);
nor U4003 (N_4003,N_1554,N_1936);
or U4004 (N_4004,N_2428,N_2904);
and U4005 (N_4005,N_1642,N_2543);
xnor U4006 (N_4006,N_2704,N_2033);
and U4007 (N_4007,N_2722,N_1850);
xnor U4008 (N_4008,N_1581,N_2749);
or U4009 (N_4009,N_1829,N_2850);
xnor U4010 (N_4010,N_2895,N_2829);
and U4011 (N_4011,N_1884,N_1948);
and U4012 (N_4012,N_1743,N_1900);
or U4013 (N_4013,N_1823,N_2915);
xor U4014 (N_4014,N_2713,N_2913);
xor U4015 (N_4015,N_2325,N_1568);
nand U4016 (N_4016,N_2708,N_1566);
or U4017 (N_4017,N_2406,N_2271);
and U4018 (N_4018,N_2725,N_2796);
nand U4019 (N_4019,N_2049,N_1501);
nand U4020 (N_4020,N_1737,N_1640);
nor U4021 (N_4021,N_2591,N_2704);
nand U4022 (N_4022,N_2024,N_2012);
xnor U4023 (N_4023,N_1992,N_1502);
or U4024 (N_4024,N_1613,N_2413);
xnor U4025 (N_4025,N_2859,N_1710);
nor U4026 (N_4026,N_2960,N_2670);
or U4027 (N_4027,N_2124,N_2036);
nand U4028 (N_4028,N_2256,N_2329);
or U4029 (N_4029,N_1934,N_1542);
and U4030 (N_4030,N_2641,N_2724);
xnor U4031 (N_4031,N_2637,N_2117);
xor U4032 (N_4032,N_2249,N_1931);
xnor U4033 (N_4033,N_2980,N_2349);
nor U4034 (N_4034,N_2097,N_2045);
xor U4035 (N_4035,N_1812,N_2124);
nand U4036 (N_4036,N_2477,N_2044);
xor U4037 (N_4037,N_2945,N_2038);
xor U4038 (N_4038,N_2961,N_1708);
or U4039 (N_4039,N_2042,N_2726);
nand U4040 (N_4040,N_1683,N_2307);
or U4041 (N_4041,N_2671,N_2411);
and U4042 (N_4042,N_2046,N_1503);
xor U4043 (N_4043,N_2497,N_2223);
nor U4044 (N_4044,N_2157,N_2998);
nand U4045 (N_4045,N_1551,N_2330);
nor U4046 (N_4046,N_2700,N_2997);
and U4047 (N_4047,N_2701,N_1683);
xor U4048 (N_4048,N_1987,N_1661);
and U4049 (N_4049,N_2258,N_2007);
and U4050 (N_4050,N_1863,N_2963);
xor U4051 (N_4051,N_2012,N_1507);
nand U4052 (N_4052,N_2712,N_2804);
nor U4053 (N_4053,N_2345,N_2063);
and U4054 (N_4054,N_1973,N_1919);
or U4055 (N_4055,N_2386,N_2432);
nand U4056 (N_4056,N_1687,N_2190);
and U4057 (N_4057,N_2418,N_2292);
nand U4058 (N_4058,N_1599,N_1538);
and U4059 (N_4059,N_1875,N_2395);
nand U4060 (N_4060,N_2243,N_1798);
nor U4061 (N_4061,N_2534,N_2624);
nor U4062 (N_4062,N_1903,N_1583);
or U4063 (N_4063,N_1579,N_1882);
nor U4064 (N_4064,N_2920,N_2873);
and U4065 (N_4065,N_2878,N_1649);
nor U4066 (N_4066,N_2619,N_2280);
nand U4067 (N_4067,N_1968,N_1636);
xnor U4068 (N_4068,N_1789,N_2854);
nand U4069 (N_4069,N_1691,N_2439);
nand U4070 (N_4070,N_1572,N_1801);
and U4071 (N_4071,N_2107,N_2928);
or U4072 (N_4072,N_1593,N_2901);
or U4073 (N_4073,N_2238,N_2122);
nand U4074 (N_4074,N_2188,N_1833);
or U4075 (N_4075,N_2288,N_2837);
xor U4076 (N_4076,N_2465,N_2451);
and U4077 (N_4077,N_1548,N_1757);
or U4078 (N_4078,N_2101,N_1730);
and U4079 (N_4079,N_2809,N_2345);
and U4080 (N_4080,N_2845,N_2318);
xnor U4081 (N_4081,N_1669,N_2569);
nor U4082 (N_4082,N_1935,N_2046);
xor U4083 (N_4083,N_1647,N_1771);
nor U4084 (N_4084,N_2217,N_2766);
nor U4085 (N_4085,N_2850,N_1822);
nand U4086 (N_4086,N_2187,N_2897);
xnor U4087 (N_4087,N_2800,N_2757);
nor U4088 (N_4088,N_1625,N_2480);
and U4089 (N_4089,N_2875,N_2003);
xnor U4090 (N_4090,N_1603,N_2150);
or U4091 (N_4091,N_2454,N_1908);
or U4092 (N_4092,N_2965,N_1575);
nor U4093 (N_4093,N_2005,N_2539);
xor U4094 (N_4094,N_1912,N_2188);
xnor U4095 (N_4095,N_1948,N_2853);
or U4096 (N_4096,N_1591,N_2276);
nand U4097 (N_4097,N_2654,N_2796);
and U4098 (N_4098,N_1583,N_2980);
nand U4099 (N_4099,N_1609,N_2309);
and U4100 (N_4100,N_1784,N_2829);
nor U4101 (N_4101,N_2907,N_2531);
xnor U4102 (N_4102,N_1525,N_1839);
nor U4103 (N_4103,N_2804,N_2736);
xnor U4104 (N_4104,N_1633,N_2011);
nor U4105 (N_4105,N_2060,N_1645);
or U4106 (N_4106,N_1795,N_1530);
and U4107 (N_4107,N_2675,N_2608);
or U4108 (N_4108,N_2030,N_1852);
or U4109 (N_4109,N_1976,N_1784);
or U4110 (N_4110,N_1756,N_2637);
nand U4111 (N_4111,N_1832,N_2938);
and U4112 (N_4112,N_2984,N_2736);
xor U4113 (N_4113,N_2226,N_2086);
xor U4114 (N_4114,N_1896,N_2047);
and U4115 (N_4115,N_2247,N_1535);
and U4116 (N_4116,N_1913,N_1919);
nor U4117 (N_4117,N_2557,N_1663);
or U4118 (N_4118,N_2657,N_1980);
xor U4119 (N_4119,N_2287,N_2521);
xor U4120 (N_4120,N_1885,N_1585);
or U4121 (N_4121,N_2689,N_2433);
and U4122 (N_4122,N_2569,N_1890);
xor U4123 (N_4123,N_2213,N_2559);
or U4124 (N_4124,N_1936,N_1730);
and U4125 (N_4125,N_2034,N_2804);
and U4126 (N_4126,N_2356,N_1622);
nand U4127 (N_4127,N_2692,N_2107);
and U4128 (N_4128,N_2793,N_2217);
or U4129 (N_4129,N_2448,N_1618);
nor U4130 (N_4130,N_2735,N_2447);
and U4131 (N_4131,N_2603,N_2472);
nor U4132 (N_4132,N_1886,N_2254);
xnor U4133 (N_4133,N_2598,N_2465);
nand U4134 (N_4134,N_1907,N_2269);
or U4135 (N_4135,N_2037,N_2306);
or U4136 (N_4136,N_1736,N_2518);
nor U4137 (N_4137,N_1722,N_2599);
nand U4138 (N_4138,N_2116,N_2257);
or U4139 (N_4139,N_1914,N_1984);
nand U4140 (N_4140,N_2190,N_2567);
or U4141 (N_4141,N_2307,N_2211);
nor U4142 (N_4142,N_2818,N_1513);
or U4143 (N_4143,N_2562,N_2667);
nand U4144 (N_4144,N_1566,N_1826);
or U4145 (N_4145,N_2668,N_2506);
and U4146 (N_4146,N_2342,N_2742);
xnor U4147 (N_4147,N_2447,N_2928);
or U4148 (N_4148,N_2786,N_1821);
or U4149 (N_4149,N_2743,N_1680);
and U4150 (N_4150,N_2949,N_2783);
xnor U4151 (N_4151,N_2814,N_1843);
or U4152 (N_4152,N_2136,N_2370);
or U4153 (N_4153,N_2974,N_2654);
and U4154 (N_4154,N_2466,N_1908);
nor U4155 (N_4155,N_2317,N_2090);
nand U4156 (N_4156,N_1674,N_1869);
xnor U4157 (N_4157,N_1821,N_2629);
nor U4158 (N_4158,N_2813,N_2245);
or U4159 (N_4159,N_1517,N_1614);
or U4160 (N_4160,N_2356,N_2929);
xor U4161 (N_4161,N_2383,N_2254);
nor U4162 (N_4162,N_2062,N_2197);
nand U4163 (N_4163,N_2050,N_2859);
nand U4164 (N_4164,N_2037,N_1864);
nand U4165 (N_4165,N_1922,N_2982);
nor U4166 (N_4166,N_2935,N_2359);
or U4167 (N_4167,N_1641,N_2898);
or U4168 (N_4168,N_2968,N_2985);
xnor U4169 (N_4169,N_2794,N_2416);
xnor U4170 (N_4170,N_2999,N_1724);
nor U4171 (N_4171,N_2344,N_1980);
or U4172 (N_4172,N_2646,N_1612);
and U4173 (N_4173,N_1834,N_2121);
nand U4174 (N_4174,N_2694,N_2887);
nand U4175 (N_4175,N_2920,N_2991);
or U4176 (N_4176,N_2557,N_1598);
nor U4177 (N_4177,N_2396,N_2569);
and U4178 (N_4178,N_2790,N_1513);
nand U4179 (N_4179,N_1909,N_1583);
xor U4180 (N_4180,N_2322,N_2042);
or U4181 (N_4181,N_1570,N_2325);
or U4182 (N_4182,N_2821,N_2425);
xor U4183 (N_4183,N_2453,N_2911);
nor U4184 (N_4184,N_1995,N_2856);
nand U4185 (N_4185,N_2396,N_2308);
nand U4186 (N_4186,N_1684,N_1930);
or U4187 (N_4187,N_2447,N_1584);
nand U4188 (N_4188,N_2196,N_2182);
nand U4189 (N_4189,N_2047,N_2736);
xor U4190 (N_4190,N_2051,N_2632);
or U4191 (N_4191,N_2317,N_1912);
nor U4192 (N_4192,N_2929,N_2180);
and U4193 (N_4193,N_2026,N_2195);
nor U4194 (N_4194,N_1713,N_2756);
and U4195 (N_4195,N_2514,N_2326);
nor U4196 (N_4196,N_2575,N_1825);
nor U4197 (N_4197,N_1792,N_2657);
nand U4198 (N_4198,N_2633,N_2403);
nor U4199 (N_4199,N_2167,N_2223);
nand U4200 (N_4200,N_2118,N_1664);
xnor U4201 (N_4201,N_1628,N_2784);
and U4202 (N_4202,N_2766,N_1692);
or U4203 (N_4203,N_2729,N_1899);
or U4204 (N_4204,N_1721,N_1529);
and U4205 (N_4205,N_2439,N_2540);
and U4206 (N_4206,N_2041,N_1769);
nor U4207 (N_4207,N_2750,N_1954);
nor U4208 (N_4208,N_1916,N_1829);
xor U4209 (N_4209,N_1678,N_2771);
nor U4210 (N_4210,N_1535,N_2405);
or U4211 (N_4211,N_2649,N_2189);
nor U4212 (N_4212,N_1614,N_2751);
or U4213 (N_4213,N_2373,N_2533);
or U4214 (N_4214,N_1723,N_1660);
and U4215 (N_4215,N_1521,N_2995);
xor U4216 (N_4216,N_1798,N_2240);
and U4217 (N_4217,N_2675,N_2876);
or U4218 (N_4218,N_2740,N_2797);
xor U4219 (N_4219,N_2047,N_1983);
or U4220 (N_4220,N_2121,N_1981);
xor U4221 (N_4221,N_1883,N_2658);
nand U4222 (N_4222,N_1879,N_2470);
or U4223 (N_4223,N_2509,N_2018);
xnor U4224 (N_4224,N_1505,N_2883);
xor U4225 (N_4225,N_1567,N_1501);
and U4226 (N_4226,N_1910,N_1647);
nor U4227 (N_4227,N_1921,N_1900);
or U4228 (N_4228,N_2165,N_2191);
and U4229 (N_4229,N_2265,N_2519);
nand U4230 (N_4230,N_1974,N_2352);
nand U4231 (N_4231,N_2572,N_1869);
and U4232 (N_4232,N_2258,N_1614);
or U4233 (N_4233,N_2805,N_1543);
nand U4234 (N_4234,N_2926,N_2657);
or U4235 (N_4235,N_1868,N_1705);
and U4236 (N_4236,N_2739,N_2047);
xnor U4237 (N_4237,N_2988,N_2091);
xnor U4238 (N_4238,N_2325,N_2515);
and U4239 (N_4239,N_2743,N_2350);
nor U4240 (N_4240,N_2758,N_2728);
nor U4241 (N_4241,N_1672,N_2923);
xnor U4242 (N_4242,N_1686,N_1589);
nand U4243 (N_4243,N_2017,N_2447);
and U4244 (N_4244,N_1729,N_1995);
and U4245 (N_4245,N_2175,N_1533);
nand U4246 (N_4246,N_1864,N_2476);
nand U4247 (N_4247,N_2376,N_2472);
nand U4248 (N_4248,N_2216,N_2571);
nand U4249 (N_4249,N_1835,N_2432);
xor U4250 (N_4250,N_1822,N_2917);
or U4251 (N_4251,N_2218,N_1893);
and U4252 (N_4252,N_2934,N_2579);
or U4253 (N_4253,N_1706,N_2201);
xor U4254 (N_4254,N_2721,N_2625);
xor U4255 (N_4255,N_2987,N_2326);
xnor U4256 (N_4256,N_2305,N_2704);
and U4257 (N_4257,N_2710,N_2864);
and U4258 (N_4258,N_2724,N_2439);
and U4259 (N_4259,N_1913,N_2161);
nor U4260 (N_4260,N_1972,N_2474);
xor U4261 (N_4261,N_2136,N_2042);
nand U4262 (N_4262,N_2227,N_2670);
nand U4263 (N_4263,N_2332,N_1768);
nor U4264 (N_4264,N_2065,N_1785);
nor U4265 (N_4265,N_2212,N_1776);
or U4266 (N_4266,N_1837,N_2229);
nand U4267 (N_4267,N_1957,N_2886);
nor U4268 (N_4268,N_2070,N_2207);
and U4269 (N_4269,N_2175,N_1821);
and U4270 (N_4270,N_1529,N_2748);
nand U4271 (N_4271,N_2763,N_2191);
nand U4272 (N_4272,N_2188,N_1688);
or U4273 (N_4273,N_1944,N_2508);
or U4274 (N_4274,N_2716,N_2611);
xnor U4275 (N_4275,N_1711,N_1876);
nor U4276 (N_4276,N_1628,N_2536);
or U4277 (N_4277,N_1583,N_1983);
xnor U4278 (N_4278,N_2110,N_2290);
xor U4279 (N_4279,N_2908,N_2924);
xnor U4280 (N_4280,N_2447,N_1508);
xor U4281 (N_4281,N_2626,N_2025);
and U4282 (N_4282,N_2707,N_1836);
nor U4283 (N_4283,N_2087,N_1647);
and U4284 (N_4284,N_1887,N_1878);
nand U4285 (N_4285,N_2528,N_2853);
or U4286 (N_4286,N_2464,N_2101);
xor U4287 (N_4287,N_2658,N_2495);
or U4288 (N_4288,N_1781,N_1782);
nor U4289 (N_4289,N_1872,N_2560);
and U4290 (N_4290,N_2976,N_1986);
xor U4291 (N_4291,N_2873,N_1650);
or U4292 (N_4292,N_2221,N_2409);
nand U4293 (N_4293,N_2583,N_1537);
or U4294 (N_4294,N_1722,N_1791);
nor U4295 (N_4295,N_2719,N_2334);
nand U4296 (N_4296,N_2812,N_2546);
or U4297 (N_4297,N_2165,N_2443);
or U4298 (N_4298,N_1952,N_2723);
nand U4299 (N_4299,N_2654,N_2456);
or U4300 (N_4300,N_2812,N_2866);
xnor U4301 (N_4301,N_2225,N_2132);
xor U4302 (N_4302,N_2577,N_2897);
nand U4303 (N_4303,N_1993,N_2265);
xnor U4304 (N_4304,N_1791,N_2608);
or U4305 (N_4305,N_2475,N_2083);
and U4306 (N_4306,N_2728,N_1566);
nand U4307 (N_4307,N_1724,N_2314);
and U4308 (N_4308,N_1931,N_2780);
xnor U4309 (N_4309,N_2187,N_2758);
xnor U4310 (N_4310,N_2909,N_1573);
nand U4311 (N_4311,N_2707,N_2797);
or U4312 (N_4312,N_2525,N_2698);
nand U4313 (N_4313,N_2088,N_1903);
nor U4314 (N_4314,N_2160,N_2599);
xnor U4315 (N_4315,N_2662,N_2724);
nor U4316 (N_4316,N_1944,N_2353);
and U4317 (N_4317,N_2000,N_2112);
and U4318 (N_4318,N_1646,N_2622);
xnor U4319 (N_4319,N_2285,N_1755);
or U4320 (N_4320,N_2888,N_2363);
nor U4321 (N_4321,N_2227,N_1962);
and U4322 (N_4322,N_2680,N_2195);
nor U4323 (N_4323,N_1969,N_1832);
xnor U4324 (N_4324,N_2353,N_2986);
xor U4325 (N_4325,N_1724,N_2921);
and U4326 (N_4326,N_2657,N_1561);
xor U4327 (N_4327,N_1902,N_2952);
xnor U4328 (N_4328,N_2264,N_1931);
and U4329 (N_4329,N_1862,N_1769);
xor U4330 (N_4330,N_2933,N_1597);
xor U4331 (N_4331,N_1656,N_1636);
and U4332 (N_4332,N_1574,N_2708);
nand U4333 (N_4333,N_2526,N_2878);
or U4334 (N_4334,N_2561,N_1544);
and U4335 (N_4335,N_1597,N_2021);
nand U4336 (N_4336,N_2005,N_2087);
nor U4337 (N_4337,N_2091,N_2677);
or U4338 (N_4338,N_2245,N_1854);
xor U4339 (N_4339,N_1702,N_1746);
nand U4340 (N_4340,N_2132,N_2400);
nor U4341 (N_4341,N_2036,N_1880);
nand U4342 (N_4342,N_2258,N_1709);
nand U4343 (N_4343,N_1851,N_1530);
nor U4344 (N_4344,N_1552,N_1753);
xnor U4345 (N_4345,N_2310,N_2824);
and U4346 (N_4346,N_2212,N_2034);
or U4347 (N_4347,N_2966,N_2845);
nor U4348 (N_4348,N_2096,N_2587);
or U4349 (N_4349,N_2276,N_2017);
xor U4350 (N_4350,N_1554,N_1565);
nand U4351 (N_4351,N_1683,N_2571);
xor U4352 (N_4352,N_2319,N_1595);
xor U4353 (N_4353,N_1755,N_2401);
xnor U4354 (N_4354,N_2940,N_1693);
and U4355 (N_4355,N_2976,N_1781);
xor U4356 (N_4356,N_1767,N_2475);
xnor U4357 (N_4357,N_2024,N_1748);
and U4358 (N_4358,N_1735,N_2331);
nor U4359 (N_4359,N_2274,N_2534);
nand U4360 (N_4360,N_1605,N_1915);
xor U4361 (N_4361,N_1970,N_2948);
nand U4362 (N_4362,N_2701,N_1513);
nand U4363 (N_4363,N_2173,N_2692);
or U4364 (N_4364,N_1795,N_2085);
or U4365 (N_4365,N_2491,N_2886);
and U4366 (N_4366,N_2959,N_2810);
nand U4367 (N_4367,N_2335,N_2152);
and U4368 (N_4368,N_2084,N_2050);
nand U4369 (N_4369,N_2098,N_1583);
or U4370 (N_4370,N_2825,N_2145);
xnor U4371 (N_4371,N_2843,N_2767);
nor U4372 (N_4372,N_2529,N_1753);
nor U4373 (N_4373,N_2151,N_1657);
and U4374 (N_4374,N_2156,N_2075);
nor U4375 (N_4375,N_2389,N_1777);
nor U4376 (N_4376,N_2541,N_1748);
and U4377 (N_4377,N_1833,N_2516);
or U4378 (N_4378,N_1994,N_2189);
nand U4379 (N_4379,N_2749,N_2105);
xnor U4380 (N_4380,N_1846,N_2630);
and U4381 (N_4381,N_1891,N_2171);
xnor U4382 (N_4382,N_2351,N_2097);
nand U4383 (N_4383,N_2283,N_2993);
and U4384 (N_4384,N_2995,N_2286);
xnor U4385 (N_4385,N_1829,N_1670);
nor U4386 (N_4386,N_2105,N_2730);
or U4387 (N_4387,N_2459,N_2235);
or U4388 (N_4388,N_1502,N_2454);
nand U4389 (N_4389,N_2967,N_1947);
xnor U4390 (N_4390,N_1928,N_2398);
and U4391 (N_4391,N_2060,N_1961);
nand U4392 (N_4392,N_2551,N_1611);
xor U4393 (N_4393,N_1784,N_1824);
nand U4394 (N_4394,N_1753,N_2833);
xor U4395 (N_4395,N_1632,N_2982);
or U4396 (N_4396,N_2863,N_1668);
nor U4397 (N_4397,N_1526,N_1840);
and U4398 (N_4398,N_2234,N_2089);
and U4399 (N_4399,N_2332,N_2412);
nor U4400 (N_4400,N_2950,N_2127);
and U4401 (N_4401,N_1584,N_2464);
xnor U4402 (N_4402,N_1845,N_1630);
and U4403 (N_4403,N_1901,N_1520);
and U4404 (N_4404,N_2974,N_2855);
or U4405 (N_4405,N_2814,N_1938);
nor U4406 (N_4406,N_2675,N_2163);
nand U4407 (N_4407,N_2370,N_1681);
nand U4408 (N_4408,N_2229,N_2271);
or U4409 (N_4409,N_2038,N_2521);
nor U4410 (N_4410,N_2905,N_1809);
xor U4411 (N_4411,N_2035,N_2547);
nor U4412 (N_4412,N_1759,N_2714);
and U4413 (N_4413,N_1862,N_2192);
xnor U4414 (N_4414,N_2394,N_2461);
nor U4415 (N_4415,N_2221,N_2602);
and U4416 (N_4416,N_2136,N_1795);
xnor U4417 (N_4417,N_1662,N_2366);
xor U4418 (N_4418,N_1529,N_2028);
nor U4419 (N_4419,N_2315,N_1648);
nor U4420 (N_4420,N_2332,N_2078);
and U4421 (N_4421,N_1856,N_2514);
nand U4422 (N_4422,N_2713,N_2184);
nor U4423 (N_4423,N_1814,N_2233);
nand U4424 (N_4424,N_2378,N_2140);
nor U4425 (N_4425,N_2131,N_1748);
or U4426 (N_4426,N_2521,N_2791);
nand U4427 (N_4427,N_2778,N_1731);
nor U4428 (N_4428,N_2019,N_2785);
or U4429 (N_4429,N_2288,N_1529);
or U4430 (N_4430,N_2459,N_1783);
nor U4431 (N_4431,N_2212,N_2924);
xor U4432 (N_4432,N_2976,N_2323);
nand U4433 (N_4433,N_2059,N_1959);
nor U4434 (N_4434,N_2709,N_1681);
nand U4435 (N_4435,N_2272,N_1815);
nand U4436 (N_4436,N_2645,N_2984);
xnor U4437 (N_4437,N_2744,N_1636);
and U4438 (N_4438,N_1847,N_2565);
and U4439 (N_4439,N_2803,N_1965);
and U4440 (N_4440,N_2975,N_2582);
nor U4441 (N_4441,N_2040,N_2940);
nor U4442 (N_4442,N_2908,N_2004);
nand U4443 (N_4443,N_1708,N_1663);
nor U4444 (N_4444,N_2476,N_2397);
or U4445 (N_4445,N_2473,N_1995);
nand U4446 (N_4446,N_2258,N_1587);
nand U4447 (N_4447,N_1582,N_2988);
and U4448 (N_4448,N_2970,N_1651);
and U4449 (N_4449,N_1726,N_1942);
nand U4450 (N_4450,N_2749,N_2909);
xor U4451 (N_4451,N_2456,N_2007);
nand U4452 (N_4452,N_1605,N_2786);
and U4453 (N_4453,N_2590,N_2738);
xor U4454 (N_4454,N_2232,N_2214);
xnor U4455 (N_4455,N_2933,N_2842);
nand U4456 (N_4456,N_2907,N_1917);
nor U4457 (N_4457,N_1874,N_1546);
or U4458 (N_4458,N_2763,N_2627);
nor U4459 (N_4459,N_2322,N_1576);
nand U4460 (N_4460,N_2708,N_1794);
or U4461 (N_4461,N_2215,N_2000);
or U4462 (N_4462,N_2092,N_2754);
or U4463 (N_4463,N_1939,N_2196);
xor U4464 (N_4464,N_1998,N_1994);
or U4465 (N_4465,N_1603,N_2707);
and U4466 (N_4466,N_2174,N_2408);
and U4467 (N_4467,N_2195,N_2309);
xor U4468 (N_4468,N_1830,N_1882);
xnor U4469 (N_4469,N_2156,N_2082);
and U4470 (N_4470,N_2817,N_2337);
or U4471 (N_4471,N_2281,N_1979);
and U4472 (N_4472,N_1654,N_2371);
xor U4473 (N_4473,N_2458,N_1920);
and U4474 (N_4474,N_2313,N_2551);
nor U4475 (N_4475,N_2559,N_2016);
or U4476 (N_4476,N_2844,N_2828);
and U4477 (N_4477,N_1871,N_2168);
or U4478 (N_4478,N_2895,N_2057);
and U4479 (N_4479,N_2703,N_1829);
and U4480 (N_4480,N_1595,N_1942);
nor U4481 (N_4481,N_2564,N_2098);
or U4482 (N_4482,N_2525,N_2248);
nand U4483 (N_4483,N_1537,N_1980);
nand U4484 (N_4484,N_2548,N_1687);
nand U4485 (N_4485,N_2432,N_2365);
nor U4486 (N_4486,N_2901,N_2500);
or U4487 (N_4487,N_2373,N_1620);
or U4488 (N_4488,N_2292,N_2805);
and U4489 (N_4489,N_1938,N_2597);
or U4490 (N_4490,N_1753,N_2294);
nor U4491 (N_4491,N_1950,N_2811);
or U4492 (N_4492,N_1982,N_1888);
or U4493 (N_4493,N_1813,N_2585);
nor U4494 (N_4494,N_1693,N_2252);
xor U4495 (N_4495,N_1939,N_2879);
or U4496 (N_4496,N_2452,N_1793);
nor U4497 (N_4497,N_2868,N_1877);
or U4498 (N_4498,N_2370,N_1943);
or U4499 (N_4499,N_1910,N_2701);
and U4500 (N_4500,N_3833,N_3306);
or U4501 (N_4501,N_3473,N_3603);
nor U4502 (N_4502,N_4481,N_4362);
nor U4503 (N_4503,N_3291,N_3887);
or U4504 (N_4504,N_3043,N_3038);
nand U4505 (N_4505,N_3791,N_4143);
and U4506 (N_4506,N_3104,N_4389);
and U4507 (N_4507,N_3027,N_3072);
and U4508 (N_4508,N_3957,N_3383);
xor U4509 (N_4509,N_3434,N_4117);
xnor U4510 (N_4510,N_4409,N_4152);
or U4511 (N_4511,N_3889,N_3784);
and U4512 (N_4512,N_3377,N_4249);
nor U4513 (N_4513,N_4209,N_3412);
or U4514 (N_4514,N_3663,N_3790);
nand U4515 (N_4515,N_3276,N_4078);
xor U4516 (N_4516,N_3742,N_3367);
xor U4517 (N_4517,N_3189,N_3334);
or U4518 (N_4518,N_3193,N_3696);
and U4519 (N_4519,N_3135,N_3360);
or U4520 (N_4520,N_3551,N_3998);
or U4521 (N_4521,N_4057,N_3967);
and U4522 (N_4522,N_3654,N_3853);
nor U4523 (N_4523,N_3869,N_3927);
or U4524 (N_4524,N_3908,N_4102);
and U4525 (N_4525,N_4482,N_3681);
or U4526 (N_4526,N_4134,N_4111);
and U4527 (N_4527,N_4180,N_3323);
and U4528 (N_4528,N_3392,N_4181);
and U4529 (N_4529,N_3870,N_3232);
nand U4530 (N_4530,N_3764,N_4464);
nand U4531 (N_4531,N_3425,N_4351);
xor U4532 (N_4532,N_3959,N_4088);
and U4533 (N_4533,N_3989,N_3021);
nor U4534 (N_4534,N_3263,N_3670);
xor U4535 (N_4535,N_4240,N_4420);
nand U4536 (N_4536,N_3865,N_3147);
nor U4537 (N_4537,N_3910,N_3627);
nor U4538 (N_4538,N_3036,N_4321);
nand U4539 (N_4539,N_4026,N_4113);
or U4540 (N_4540,N_3535,N_4148);
and U4541 (N_4541,N_3279,N_3732);
or U4542 (N_4542,N_4040,N_3210);
and U4543 (N_4543,N_3891,N_4319);
nor U4544 (N_4544,N_3126,N_3305);
nand U4545 (N_4545,N_4301,N_3186);
nand U4546 (N_4546,N_4374,N_3589);
and U4547 (N_4547,N_3299,N_4480);
xor U4548 (N_4548,N_4202,N_3413);
and U4549 (N_4549,N_4170,N_3288);
and U4550 (N_4550,N_3559,N_3924);
nor U4551 (N_4551,N_3131,N_3475);
and U4552 (N_4552,N_3289,N_3039);
xor U4553 (N_4553,N_3754,N_4386);
xnor U4554 (N_4554,N_3648,N_4214);
and U4555 (N_4555,N_3084,N_3350);
or U4556 (N_4556,N_3612,N_3786);
xnor U4557 (N_4557,N_3270,N_3164);
nor U4558 (N_4558,N_4410,N_3639);
or U4559 (N_4559,N_4444,N_3173);
xnor U4560 (N_4560,N_3493,N_3757);
nor U4561 (N_4561,N_3642,N_3448);
or U4562 (N_4562,N_4108,N_3222);
xor U4563 (N_4563,N_3883,N_4097);
nor U4564 (N_4564,N_4109,N_3057);
and U4565 (N_4565,N_4281,N_3258);
or U4566 (N_4566,N_3008,N_3911);
xor U4567 (N_4567,N_3205,N_4032);
or U4568 (N_4568,N_4167,N_3484);
nand U4569 (N_4569,N_3093,N_3481);
xor U4570 (N_4570,N_3549,N_3874);
xnor U4571 (N_4571,N_3525,N_4082);
xnor U4572 (N_4572,N_3649,N_3191);
nand U4573 (N_4573,N_4245,N_3864);
xor U4574 (N_4574,N_4408,N_3725);
and U4575 (N_4575,N_3937,N_3406);
or U4576 (N_4576,N_3029,N_3839);
nor U4577 (N_4577,N_3515,N_3999);
or U4578 (N_4578,N_4308,N_4264);
xnor U4579 (N_4579,N_3547,N_3563);
and U4580 (N_4580,N_4018,N_3932);
xor U4581 (N_4581,N_3153,N_4427);
and U4582 (N_4582,N_4135,N_4165);
nor U4583 (N_4583,N_4411,N_3097);
or U4584 (N_4584,N_3092,N_3058);
or U4585 (N_4585,N_4008,N_4471);
or U4586 (N_4586,N_3068,N_3200);
or U4587 (N_4587,N_3028,N_3693);
xor U4588 (N_4588,N_3139,N_3965);
nor U4589 (N_4589,N_3235,N_3509);
and U4590 (N_4590,N_4207,N_4350);
nor U4591 (N_4591,N_3255,N_4277);
nor U4592 (N_4592,N_4392,N_3183);
xnor U4593 (N_4593,N_4388,N_3431);
or U4594 (N_4594,N_3492,N_3777);
nor U4595 (N_4595,N_3437,N_3984);
xnor U4596 (N_4596,N_3803,N_4403);
or U4597 (N_4597,N_4068,N_3992);
nand U4598 (N_4598,N_4052,N_4022);
nand U4599 (N_4599,N_3469,N_4150);
nor U4600 (N_4600,N_3579,N_3768);
xor U4601 (N_4601,N_4270,N_4356);
xnor U4602 (N_4602,N_3931,N_4456);
nand U4603 (N_4603,N_4428,N_3441);
xor U4604 (N_4604,N_3944,N_3562);
xnor U4605 (N_4605,N_3101,N_3909);
xnor U4606 (N_4606,N_4103,N_4033);
nor U4607 (N_4607,N_3792,N_4457);
xnor U4608 (N_4608,N_3672,N_4314);
xor U4609 (N_4609,N_4125,N_3209);
xor U4610 (N_4610,N_3960,N_3476);
xor U4611 (N_4611,N_3928,N_4404);
and U4612 (N_4612,N_3733,N_3806);
xor U4613 (N_4613,N_3304,N_4426);
nor U4614 (N_4614,N_3505,N_3665);
nor U4615 (N_4615,N_3320,N_4476);
and U4616 (N_4616,N_4062,N_3682);
xor U4617 (N_4617,N_3148,N_3100);
nor U4618 (N_4618,N_3180,N_3022);
nor U4619 (N_4619,N_3014,N_3716);
and U4620 (N_4620,N_3391,N_3423);
nor U4621 (N_4621,N_3686,N_3502);
xor U4622 (N_4622,N_3026,N_3385);
xnor U4623 (N_4623,N_4415,N_3961);
and U4624 (N_4624,N_3185,N_4038);
nor U4625 (N_4625,N_4246,N_3694);
nor U4626 (N_4626,N_3607,N_4247);
or U4627 (N_4627,N_4244,N_3794);
or U4628 (N_4628,N_3948,N_3284);
nor U4629 (N_4629,N_4210,N_3583);
nor U4630 (N_4630,N_4071,N_4373);
or U4631 (N_4631,N_4161,N_4394);
and U4632 (N_4632,N_3763,N_3424);
nor U4633 (N_4633,N_3459,N_3328);
and U4634 (N_4634,N_3988,N_3608);
nor U4635 (N_4635,N_3950,N_3503);
and U4636 (N_4636,N_3368,N_3482);
xnor U4637 (N_4637,N_4405,N_3138);
nand U4638 (N_4638,N_3979,N_4274);
nand U4639 (N_4639,N_4442,N_3062);
and U4640 (N_4640,N_3737,N_3049);
nor U4641 (N_4641,N_3478,N_4304);
or U4642 (N_4642,N_3526,N_3146);
nand U4643 (N_4643,N_4424,N_3894);
xor U4644 (N_4644,N_4174,N_4208);
nor U4645 (N_4645,N_4498,N_3316);
and U4646 (N_4646,N_4090,N_3685);
xnor U4647 (N_4647,N_4357,N_4486);
nand U4648 (N_4648,N_3850,N_4275);
or U4649 (N_4649,N_4056,N_4188);
or U4650 (N_4650,N_4029,N_3662);
nand U4651 (N_4651,N_4300,N_3176);
nor U4652 (N_4652,N_4230,N_3644);
xnor U4653 (N_4653,N_3201,N_3252);
nor U4654 (N_4654,N_3647,N_3743);
nor U4655 (N_4655,N_3674,N_4043);
nand U4656 (N_4656,N_3370,N_4064);
xor U4657 (N_4657,N_3310,N_4422);
or U4658 (N_4658,N_4348,N_3512);
xnor U4659 (N_4659,N_4127,N_4273);
nor U4660 (N_4660,N_3472,N_3553);
nand U4661 (N_4661,N_4157,N_3446);
nor U4662 (N_4662,N_4067,N_3913);
nor U4663 (N_4663,N_3426,N_3409);
nor U4664 (N_4664,N_4081,N_3699);
nor U4665 (N_4665,N_4168,N_3567);
nor U4666 (N_4666,N_3531,N_3326);
xor U4667 (N_4667,N_3366,N_3861);
and U4668 (N_4668,N_4325,N_3449);
and U4669 (N_4669,N_3812,N_4401);
nor U4670 (N_4670,N_4002,N_4126);
xnor U4671 (N_4671,N_3397,N_4285);
nor U4672 (N_4672,N_3394,N_3741);
or U4673 (N_4673,N_3797,N_3919);
and U4674 (N_4674,N_3990,N_3041);
or U4675 (N_4675,N_3046,N_3402);
and U4676 (N_4676,N_4490,N_3108);
nand U4677 (N_4677,N_4298,N_4179);
nor U4678 (N_4678,N_4009,N_4139);
xnor U4679 (N_4679,N_3691,N_3332);
nand U4680 (N_4680,N_3116,N_4192);
or U4681 (N_4681,N_3762,N_4027);
nand U4682 (N_4682,N_3165,N_4254);
or U4683 (N_4683,N_3712,N_3067);
nor U4684 (N_4684,N_3309,N_4162);
or U4685 (N_4685,N_4204,N_3617);
xnor U4686 (N_4686,N_3892,N_4235);
nor U4687 (N_4687,N_3697,N_3985);
nand U4688 (N_4688,N_4006,N_3817);
and U4689 (N_4689,N_3707,N_3430);
or U4690 (N_4690,N_3411,N_3554);
nand U4691 (N_4691,N_3187,N_4058);
and U4692 (N_4692,N_4084,N_4454);
or U4693 (N_4693,N_4294,N_3669);
nand U4694 (N_4694,N_4114,N_3088);
nor U4695 (N_4695,N_3233,N_3467);
nor U4696 (N_4696,N_3523,N_3219);
or U4697 (N_4697,N_3064,N_3011);
xor U4698 (N_4698,N_3157,N_4474);
xnor U4699 (N_4699,N_3390,N_3372);
and U4700 (N_4700,N_4098,N_3254);
and U4701 (N_4701,N_3888,N_3800);
xnor U4702 (N_4702,N_4198,N_4320);
xnor U4703 (N_4703,N_3398,N_4359);
xor U4704 (N_4704,N_3900,N_3646);
xnor U4705 (N_4705,N_3516,N_3970);
and U4706 (N_4706,N_3890,N_3635);
nand U4707 (N_4707,N_3816,N_3872);
xor U4708 (N_4708,N_3442,N_3977);
nand U4709 (N_4709,N_3722,N_3436);
nor U4710 (N_4710,N_4289,N_4226);
nand U4711 (N_4711,N_4039,N_3375);
nor U4712 (N_4712,N_4129,N_3296);
and U4713 (N_4713,N_4242,N_3374);
nand U4714 (N_4714,N_3103,N_4451);
nor U4715 (N_4715,N_3450,N_3899);
or U4716 (N_4716,N_4305,N_3204);
xnor U4717 (N_4717,N_3798,N_4154);
and U4718 (N_4718,N_3259,N_3843);
nand U4719 (N_4719,N_4206,N_3528);
or U4720 (N_4720,N_4104,N_3115);
xnor U4721 (N_4721,N_4333,N_3618);
and U4722 (N_4722,N_3756,N_3271);
or U4723 (N_4723,N_4407,N_4203);
xnor U4724 (N_4724,N_4326,N_4074);
or U4725 (N_4725,N_4217,N_4335);
xnor U4726 (N_4726,N_3852,N_4156);
nand U4727 (N_4727,N_4155,N_4286);
or U4728 (N_4728,N_4019,N_4434);
or U4729 (N_4729,N_4296,N_3128);
and U4730 (N_4730,N_3904,N_3506);
nor U4731 (N_4731,N_3595,N_3190);
nand U4732 (N_4732,N_3749,N_3215);
nor U4733 (N_4733,N_3020,N_3381);
or U4734 (N_4734,N_4121,N_4462);
and U4735 (N_4735,N_4073,N_4306);
xnor U4736 (N_4736,N_4193,N_3250);
and U4737 (N_4737,N_3161,N_4160);
nor U4738 (N_4738,N_3311,N_3519);
and U4739 (N_4739,N_4372,N_3956);
and U4740 (N_4740,N_3621,N_3227);
nand U4741 (N_4741,N_4382,N_4412);
or U4742 (N_4742,N_3421,N_3314);
or U4743 (N_4743,N_3991,N_3659);
and U4744 (N_4744,N_3018,N_3051);
nor U4745 (N_4745,N_4460,N_3238);
and U4746 (N_4746,N_3748,N_4238);
and U4747 (N_4747,N_3923,N_3983);
and U4748 (N_4748,N_3091,N_3281);
xor U4749 (N_4749,N_3844,N_4353);
or U4750 (N_4750,N_3212,N_4363);
nand U4751 (N_4751,N_4086,N_4263);
or U4752 (N_4752,N_3521,N_3119);
xor U4753 (N_4753,N_3594,N_4429);
and U4754 (N_4754,N_3941,N_3156);
nand U4755 (N_4755,N_3832,N_3224);
nand U4756 (N_4756,N_3075,N_4438);
nor U4757 (N_4757,N_3601,N_4303);
nor U4758 (N_4758,N_3973,N_3445);
nand U4759 (N_4759,N_4091,N_3327);
or U4760 (N_4760,N_3572,N_3282);
xor U4761 (N_4761,N_3795,N_3925);
nand U4762 (N_4762,N_3129,N_3048);
nor U4763 (N_4763,N_3074,N_3407);
or U4764 (N_4764,N_4145,N_4315);
xnor U4765 (N_4765,N_3231,N_4488);
or U4766 (N_4766,N_3930,N_3929);
and U4767 (N_4767,N_4371,N_3468);
or U4768 (N_4768,N_3125,N_4259);
and U4769 (N_4769,N_3982,N_3471);
nor U4770 (N_4770,N_4099,N_3102);
or U4771 (N_4771,N_3596,N_3590);
or U4772 (N_4772,N_3568,N_4378);
nand U4773 (N_4773,N_3836,N_3804);
and U4774 (N_4774,N_3172,N_4096);
xor U4775 (N_4775,N_3246,N_4045);
nor U4776 (N_4776,N_4177,N_3599);
nor U4777 (N_4777,N_4212,N_3474);
nand U4778 (N_4778,N_3822,N_3401);
or U4779 (N_4779,N_4331,N_3477);
and U4780 (N_4780,N_4484,N_4499);
and U4781 (N_4781,N_3671,N_3280);
nor U4782 (N_4782,N_3962,N_4037);
xnor U4783 (N_4783,N_3915,N_4385);
nand U4784 (N_4784,N_3229,N_3490);
nor U4785 (N_4785,N_3295,N_4122);
and U4786 (N_4786,N_3858,N_3239);
or U4787 (N_4787,N_3054,N_3220);
or U4788 (N_4788,N_4302,N_3945);
and U4789 (N_4789,N_3428,N_3464);
and U4790 (N_4790,N_3668,N_3609);
nor U4791 (N_4791,N_3859,N_4169);
nand U4792 (N_4792,N_4178,N_3420);
nand U4793 (N_4793,N_4199,N_3855);
or U4794 (N_4794,N_4219,N_4358);
xnor U4795 (N_4795,N_3237,N_3511);
and U4796 (N_4796,N_3631,N_3604);
or U4797 (N_4797,N_3082,N_4376);
and U4798 (N_4798,N_3522,N_3630);
and U4799 (N_4799,N_3629,N_4465);
or U4800 (N_4800,N_3767,N_3292);
xnor U4801 (N_4801,N_3574,N_4477);
and U4802 (N_4802,N_4345,N_3706);
nor U4803 (N_4803,N_4398,N_4231);
and U4804 (N_4804,N_3234,N_3285);
nor U4805 (N_4805,N_4436,N_3868);
or U4806 (N_4806,N_3110,N_3069);
nand U4807 (N_4807,N_3435,N_3010);
or U4808 (N_4808,N_4468,N_3071);
nand U4809 (N_4809,N_3178,N_4232);
nor U4810 (N_4810,N_4370,N_3337);
and U4811 (N_4811,N_3249,N_3779);
nor U4812 (N_4812,N_3939,N_4241);
or U4813 (N_4813,N_3688,N_4280);
and U4814 (N_4814,N_3841,N_4375);
or U4815 (N_4815,N_3247,N_3753);
and U4816 (N_4816,N_3121,N_3333);
xnor U4817 (N_4817,N_3486,N_3650);
xnor U4818 (N_4818,N_3901,N_4307);
nand U4819 (N_4819,N_4228,N_3940);
nand U4820 (N_4820,N_3953,N_3162);
or U4821 (N_4821,N_3163,N_4458);
nand U4822 (N_4822,N_4138,N_3065);
or U4823 (N_4823,N_3345,N_3721);
or U4824 (N_4824,N_3628,N_4418);
and U4825 (N_4825,N_3277,N_4431);
and U4826 (N_4826,N_3954,N_3731);
xnor U4827 (N_4827,N_3873,N_3702);
and U4828 (N_4828,N_3854,N_3943);
and U4829 (N_4829,N_4028,N_3564);
xnor U4830 (N_4830,N_3632,N_4175);
or U4831 (N_4831,N_3565,N_4459);
and U4832 (N_4832,N_3458,N_3545);
nand U4833 (N_4833,N_3417,N_3349);
nor U4834 (N_4834,N_3501,N_3329);
nor U4835 (N_4835,N_3826,N_3689);
nor U4836 (N_4836,N_4128,N_4316);
and U4837 (N_4837,N_4092,N_3499);
xnor U4838 (N_4838,N_3881,N_4447);
xnor U4839 (N_4839,N_3199,N_3061);
and U4840 (N_4840,N_3044,N_3677);
nor U4841 (N_4841,N_3035,N_3997);
nor U4842 (N_4842,N_3443,N_3776);
xnor U4843 (N_4843,N_3532,N_3801);
and U4844 (N_4844,N_4191,N_3585);
nor U4845 (N_4845,N_3969,N_4318);
nand U4846 (N_4846,N_4110,N_3256);
xor U4847 (N_4847,N_4144,N_3266);
and U4848 (N_4848,N_3321,N_4284);
xnor U4849 (N_4849,N_3815,N_3752);
and U4850 (N_4850,N_3419,N_3507);
xor U4851 (N_4851,N_4227,N_3358);
xnor U4852 (N_4852,N_3060,N_4417);
nand U4853 (N_4853,N_3660,N_3695);
or U4854 (N_4854,N_4149,N_3085);
or U4855 (N_4855,N_3454,N_4140);
and U4856 (N_4856,N_3758,N_4196);
nor U4857 (N_4857,N_4063,N_3009);
nor U4858 (N_4858,N_4347,N_3771);
nand U4859 (N_4859,N_4051,N_3313);
and U4860 (N_4860,N_4224,N_4133);
xor U4861 (N_4861,N_3346,N_3253);
and U4862 (N_4862,N_3228,N_4124);
and U4863 (N_4863,N_3095,N_3203);
xor U4864 (N_4864,N_3302,N_4059);
nor U4865 (N_4865,N_3016,N_3557);
or U4866 (N_4866,N_4147,N_3746);
or U4867 (N_4867,N_3917,N_3181);
nor U4868 (N_4868,N_3750,N_3877);
xnor U4869 (N_4869,N_4171,N_4479);
xnor U4870 (N_4870,N_4036,N_3500);
nor U4871 (N_4871,N_4271,N_3405);
xnor U4872 (N_4872,N_3614,N_4349);
nand U4873 (N_4873,N_3623,N_4257);
and U4874 (N_4874,N_3141,N_3684);
nand U4875 (N_4875,N_3013,N_3728);
or U4876 (N_4876,N_4066,N_3529);
or U4877 (N_4877,N_3453,N_3542);
nor U4878 (N_4878,N_4268,N_3037);
nor U4879 (N_4879,N_3335,N_3462);
xor U4880 (N_4880,N_3533,N_3031);
nand U4881 (N_4881,N_3343,N_4360);
nand U4882 (N_4882,N_4163,N_4260);
nor U4883 (N_4883,N_4183,N_4317);
and U4884 (N_4884,N_3679,N_3903);
nor U4885 (N_4885,N_3396,N_3971);
xor U4886 (N_4886,N_4361,N_3655);
nand U4887 (N_4887,N_4119,N_4288);
nor U4888 (N_4888,N_4000,N_3914);
or U4889 (N_4889,N_4323,N_3560);
or U4890 (N_4890,N_3602,N_3633);
nor U4891 (N_4891,N_4072,N_3575);
nor U4892 (N_4892,N_3303,N_3106);
nand U4893 (N_4893,N_4322,N_4186);
and U4894 (N_4894,N_3179,N_3298);
and U4895 (N_4895,N_4369,N_3624);
or U4896 (N_4896,N_3745,N_4076);
xnor U4897 (N_4897,N_3625,N_3720);
nand U4898 (N_4898,N_3050,N_3678);
xor U4899 (N_4899,N_3317,N_4237);
xnor U4900 (N_4900,N_3751,N_4282);
nand U4901 (N_4901,N_4223,N_3325);
nor U4902 (N_4902,N_3034,N_3840);
nor U4903 (N_4903,N_3494,N_3498);
nor U4904 (N_4904,N_4310,N_3824);
nor U4905 (N_4905,N_3196,N_4469);
and U4906 (N_4906,N_3033,N_3393);
and U4907 (N_4907,N_3637,N_3548);
and U4908 (N_4908,N_3895,N_4450);
nand U4909 (N_4909,N_3882,N_3087);
nor U4910 (N_4910,N_4011,N_4205);
or U4911 (N_4911,N_4010,N_3024);
or U4912 (N_4912,N_3319,N_3336);
nand U4913 (N_4913,N_3922,N_3142);
nor U4914 (N_4914,N_4251,N_3269);
or U4915 (N_4915,N_3827,N_3318);
nand U4916 (N_4916,N_4485,N_4159);
or U4917 (N_4917,N_3508,N_3112);
nor U4918 (N_4918,N_4266,N_3056);
nor U4919 (N_4919,N_3415,N_3759);
xnor U4920 (N_4920,N_4107,N_3080);
xor U4921 (N_4921,N_4297,N_3105);
nor U4922 (N_4922,N_3986,N_4213);
nand U4923 (N_4923,N_3818,N_4399);
or U4924 (N_4924,N_4055,N_3152);
and U4925 (N_4925,N_4070,N_4229);
nand U4926 (N_4926,N_3000,N_4041);
and U4927 (N_4927,N_4402,N_3831);
nor U4928 (N_4928,N_3566,N_3182);
xnor U4929 (N_4929,N_3395,N_3550);
nor U4930 (N_4930,N_3879,N_3359);
xnor U4931 (N_4931,N_4478,N_3862);
and U4932 (N_4932,N_3847,N_3369);
or U4933 (N_4933,N_3781,N_4397);
xor U4934 (N_4934,N_3729,N_4467);
and U4935 (N_4935,N_3513,N_4466);
nand U4936 (N_4936,N_3651,N_4118);
xor U4937 (N_4937,N_4441,N_3848);
and U4938 (N_4938,N_3086,N_4433);
xor U4939 (N_4939,N_3120,N_4283);
and U4940 (N_4940,N_3495,N_4137);
and U4941 (N_4941,N_3171,N_3719);
nand U4942 (N_4942,N_4042,N_4220);
or U4943 (N_4943,N_3213,N_3963);
and U4944 (N_4944,N_3667,N_3740);
or U4945 (N_4945,N_3145,N_4406);
xnor U4946 (N_4946,N_3261,N_3378);
and U4947 (N_4947,N_3243,N_3144);
and U4948 (N_4948,N_3921,N_4425);
xor U4949 (N_4949,N_3993,N_3480);
nor U4950 (N_4950,N_3275,N_4496);
and U4951 (N_4951,N_3709,N_3636);
or U4952 (N_4952,N_3040,N_3598);
or U4953 (N_4953,N_3287,N_3555);
or U4954 (N_4954,N_3273,N_3202);
and U4955 (N_4955,N_4158,N_3114);
nor U4956 (N_4956,N_4190,N_3324);
or U4957 (N_4957,N_3004,N_3355);
nand U4958 (N_4958,N_3537,N_3496);
or U4959 (N_4959,N_3770,N_3137);
or U4960 (N_4960,N_4034,N_3880);
nand U4961 (N_4961,N_4390,N_3134);
and U4962 (N_4962,N_3638,N_3342);
or U4963 (N_4963,N_3726,N_3704);
nor U4964 (N_4964,N_3174,N_3641);
or U4965 (N_4965,N_3825,N_4030);
and U4966 (N_4966,N_3077,N_3030);
nor U4967 (N_4967,N_3207,N_4377);
or U4968 (N_4968,N_3404,N_3714);
and U4969 (N_4969,N_4354,N_4341);
nor U4970 (N_4970,N_3440,N_4222);
nor U4971 (N_4971,N_3055,N_4387);
nor U4972 (N_4972,N_4211,N_3775);
and U4973 (N_4973,N_3788,N_3301);
nand U4974 (N_4974,N_4012,N_3221);
nor U4975 (N_4975,N_3580,N_3738);
or U4976 (N_4976,N_4430,N_3130);
xnor U4977 (N_4977,N_3081,N_4435);
nand U4978 (N_4978,N_3416,N_3339);
and U4979 (N_4979,N_3208,N_3687);
xor U4980 (N_4980,N_4024,N_3123);
nor U4981 (N_4981,N_3673,N_4336);
or U4982 (N_4982,N_3322,N_4250);
or U4983 (N_4983,N_3257,N_3347);
and U4984 (N_4984,N_3514,N_3968);
nor U4985 (N_4985,N_3573,N_3111);
xnor U4986 (N_4986,N_3666,N_3782);
and U4987 (N_4987,N_4355,N_4414);
or U4988 (N_4988,N_4001,N_4287);
and U4989 (N_4989,N_4120,N_4381);
nor U4990 (N_4990,N_3427,N_3810);
nor U4991 (N_4991,N_3588,N_3331);
and U4992 (N_4992,N_3373,N_3422);
nand U4993 (N_4993,N_3994,N_3197);
or U4994 (N_4994,N_3546,N_4342);
nor U4995 (N_4995,N_3225,N_3947);
nand U4996 (N_4996,N_4101,N_3878);
xor U4997 (N_4997,N_3774,N_3244);
or U4998 (N_4998,N_3905,N_4077);
and U4999 (N_4999,N_3400,N_4324);
xor U5000 (N_5000,N_3151,N_3063);
and U5001 (N_5001,N_3705,N_3444);
nor U5002 (N_5002,N_3032,N_4233);
nand U5003 (N_5003,N_3076,N_3015);
and U5004 (N_5004,N_3701,N_3823);
xor U5005 (N_5005,N_3543,N_4334);
and U5006 (N_5006,N_3047,N_4366);
nand U5007 (N_5007,N_3799,N_3098);
xor U5008 (N_5008,N_3113,N_3133);
nand U5009 (N_5009,N_3059,N_4164);
and U5010 (N_5010,N_3886,N_3274);
xnor U5011 (N_5011,N_3168,N_4020);
xnor U5012 (N_5012,N_3278,N_4236);
nand U5013 (N_5013,N_3561,N_3184);
nand U5014 (N_5014,N_3727,N_3976);
or U5015 (N_5015,N_3294,N_4146);
nor U5016 (N_5016,N_4329,N_3361);
nor U5017 (N_5017,N_3264,N_4080);
nor U5018 (N_5018,N_4053,N_3558);
and U5019 (N_5019,N_3734,N_4075);
or U5020 (N_5020,N_3690,N_4089);
and U5021 (N_5021,N_3338,N_3211);
or U5022 (N_5022,N_4437,N_3357);
nand U5023 (N_5023,N_3620,N_3592);
or U5024 (N_5024,N_3109,N_3127);
nand U5025 (N_5025,N_3613,N_3723);
or U5026 (N_5026,N_4194,N_3692);
or U5027 (N_5027,N_4115,N_3089);
and U5028 (N_5028,N_3830,N_3388);
and U5029 (N_5029,N_4166,N_3491);
nand U5030 (N_5030,N_3597,N_3918);
nand U5031 (N_5031,N_3083,N_3297);
nor U5032 (N_5032,N_3610,N_3814);
nand U5033 (N_5033,N_3463,N_4239);
nand U5034 (N_5034,N_3569,N_3805);
nor U5035 (N_5035,N_3094,N_4035);
xor U5036 (N_5036,N_3975,N_3132);
xor U5037 (N_5037,N_4332,N_3414);
or U5038 (N_5038,N_3640,N_3717);
xor U5039 (N_5039,N_4293,N_4031);
or U5040 (N_5040,N_3838,N_4234);
xnor U5041 (N_5041,N_3452,N_3996);
nor U5042 (N_5042,N_3090,N_4094);
and U5043 (N_5043,N_3410,N_4344);
xnor U5044 (N_5044,N_4131,N_3170);
xnor U5045 (N_5045,N_4061,N_3808);
xor U5046 (N_5046,N_3117,N_3140);
xnor U5047 (N_5047,N_4453,N_3150);
or U5048 (N_5048,N_3169,N_3916);
or U5049 (N_5049,N_3926,N_3308);
or U5050 (N_5050,N_3096,N_3736);
nor U5051 (N_5051,N_4495,N_3735);
xor U5052 (N_5052,N_4446,N_3483);
xnor U5053 (N_5053,N_4225,N_3226);
nor U5054 (N_5054,N_3896,N_3821);
and U5055 (N_5055,N_3934,N_4470);
xnor U5056 (N_5056,N_3195,N_3175);
xor U5057 (N_5057,N_3643,N_3787);
or U5058 (N_5058,N_4413,N_3972);
nand U5059 (N_5059,N_4449,N_3122);
or U5060 (N_5060,N_4443,N_3461);
or U5061 (N_5061,N_4278,N_4497);
nor U5062 (N_5062,N_3007,N_4093);
or U5063 (N_5063,N_3286,N_3365);
or U5064 (N_5064,N_4005,N_3661);
nand U5065 (N_5065,N_3765,N_4112);
nor U5066 (N_5066,N_3364,N_4048);
nand U5067 (N_5067,N_3793,N_3517);
nor U5068 (N_5068,N_3760,N_3362);
and U5069 (N_5069,N_4184,N_4328);
or U5070 (N_5070,N_4393,N_3188);
and U5071 (N_5071,N_3813,N_4489);
nand U5072 (N_5072,N_3656,N_3964);
nor U5073 (N_5073,N_4493,N_4364);
nand U5074 (N_5074,N_4049,N_3262);
xnor U5075 (N_5075,N_3363,N_3524);
or U5076 (N_5076,N_3042,N_3019);
or U5077 (N_5077,N_3005,N_3376);
and U5078 (N_5078,N_3330,N_4106);
nand U5079 (N_5079,N_3974,N_3796);
nor U5080 (N_5080,N_3946,N_4279);
nand U5081 (N_5081,N_4153,N_4313);
or U5082 (N_5082,N_3245,N_4365);
nor U5083 (N_5083,N_3809,N_3192);
nor U5084 (N_5084,N_4016,N_4085);
nand U5085 (N_5085,N_4116,N_3920);
and U5086 (N_5086,N_4141,N_4054);
xnor U5087 (N_5087,N_3315,N_3653);
and U5088 (N_5088,N_3807,N_3389);
or U5089 (N_5089,N_3240,N_4383);
and U5090 (N_5090,N_4423,N_3842);
xnor U5091 (N_5091,N_3456,N_3099);
and U5092 (N_5092,N_3341,N_3487);
xor U5093 (N_5093,N_4338,N_3418);
nor U5094 (N_5094,N_4021,N_3846);
and U5095 (N_5095,N_4087,N_4200);
and U5096 (N_5096,N_4023,N_4216);
nand U5097 (N_5097,N_3698,N_3586);
xnor U5098 (N_5098,N_4046,N_3344);
and U5099 (N_5099,N_4017,N_3433);
nand U5100 (N_5100,N_4491,N_3136);
xor U5101 (N_5101,N_3465,N_3070);
or U5102 (N_5102,N_4065,N_3761);
or U5103 (N_5103,N_4197,N_3849);
nand U5104 (N_5104,N_3520,N_3785);
xor U5105 (N_5105,N_3936,N_3576);
xnor U5106 (N_5106,N_4007,N_3616);
xor U5107 (N_5107,N_3143,N_3079);
nor U5108 (N_5108,N_3403,N_3236);
nand U5109 (N_5109,N_3626,N_3206);
xnor U5110 (N_5110,N_4346,N_3871);
nor U5111 (N_5111,N_3587,N_4339);
or U5112 (N_5112,N_3884,N_3149);
xor U5113 (N_5113,N_4142,N_3466);
and U5114 (N_5114,N_3851,N_3382);
and U5115 (N_5115,N_3251,N_3352);
nor U5116 (N_5116,N_3003,N_4421);
and U5117 (N_5117,N_4455,N_3885);
and U5118 (N_5118,N_3893,N_3898);
and U5119 (N_5119,N_3399,N_3724);
or U5120 (N_5120,N_4025,N_3006);
or U5121 (N_5121,N_3439,N_3540);
xor U5122 (N_5122,N_3265,N_3460);
and U5123 (N_5123,N_3897,N_3981);
nand U5124 (N_5124,N_3012,N_4255);
and U5125 (N_5125,N_3160,N_3300);
and U5126 (N_5126,N_3497,N_3447);
xnor U5127 (N_5127,N_3866,N_4123);
nor U5128 (N_5128,N_4187,N_4448);
nand U5129 (N_5129,N_3408,N_4172);
nand U5130 (N_5130,N_3429,N_3538);
and U5131 (N_5131,N_3766,N_4327);
and U5132 (N_5132,N_3744,N_4221);
or U5133 (N_5133,N_4253,N_3718);
xor U5134 (N_5134,N_3708,N_4044);
nor U5135 (N_5135,N_4215,N_3078);
nor U5136 (N_5136,N_4432,N_3657);
and U5137 (N_5137,N_4189,N_3159);
or U5138 (N_5138,N_3223,N_3351);
and U5139 (N_5139,N_4136,N_3107);
nand U5140 (N_5140,N_4050,N_3248);
nand U5141 (N_5141,N_3242,N_3634);
and U5142 (N_5142,N_3755,N_3828);
and U5143 (N_5143,N_3652,N_4100);
nor U5144 (N_5144,N_3124,N_3942);
nor U5145 (N_5145,N_4299,N_3489);
nand U5146 (N_5146,N_4396,N_4130);
xor U5147 (N_5147,N_3214,N_3158);
xor U5148 (N_5148,N_3955,N_3875);
or U5149 (N_5149,N_3952,N_4379);
xnor U5150 (N_5150,N_3380,N_3578);
nand U5151 (N_5151,N_3980,N_3017);
xnor U5152 (N_5152,N_4176,N_4265);
and U5153 (N_5153,N_4473,N_3577);
and U5154 (N_5154,N_4439,N_3530);
xnor U5155 (N_5155,N_3606,N_3780);
or U5156 (N_5156,N_3544,N_3683);
xor U5157 (N_5157,N_3582,N_3611);
nor U5158 (N_5158,N_4440,N_3778);
nand U5159 (N_5159,N_3581,N_4079);
nor U5160 (N_5160,N_4004,N_3739);
xnor U5161 (N_5161,N_3534,N_3676);
and U5162 (N_5162,N_3619,N_4384);
nand U5163 (N_5163,N_3488,N_3710);
nor U5164 (N_5164,N_3622,N_4483);
or U5165 (N_5165,N_3675,N_4400);
and U5166 (N_5166,N_4003,N_3860);
nor U5167 (N_5167,N_3584,N_3384);
nor U5168 (N_5168,N_3177,N_4267);
xnor U5169 (N_5169,N_4218,N_3166);
xnor U5170 (N_5170,N_3591,N_4243);
and U5171 (N_5171,N_4276,N_4487);
xor U5172 (N_5172,N_3680,N_4173);
nand U5173 (N_5173,N_3432,N_3053);
xor U5174 (N_5174,N_3455,N_4182);
nand U5175 (N_5175,N_3527,N_3118);
xnor U5176 (N_5176,N_3906,N_3715);
xor U5177 (N_5177,N_3664,N_3802);
or U5178 (N_5178,N_3935,N_3711);
and U5179 (N_5179,N_4312,N_4494);
nor U5180 (N_5180,N_3353,N_4416);
or U5181 (N_5181,N_4095,N_4291);
or U5182 (N_5182,N_4015,N_3658);
nor U5183 (N_5183,N_4343,N_4185);
and U5184 (N_5184,N_3167,N_3829);
or U5185 (N_5185,N_3700,N_4445);
or U5186 (N_5186,N_3371,N_4083);
nor U5187 (N_5187,N_4261,N_3379);
or U5188 (N_5188,N_4201,N_4256);
nand U5189 (N_5189,N_3856,N_3867);
xor U5190 (N_5190,N_3216,N_4352);
nor U5191 (N_5191,N_3747,N_3820);
nand U5192 (N_5192,N_3556,N_3876);
xnor U5193 (N_5193,N_3834,N_3600);
xnor U5194 (N_5194,N_3539,N_3260);
nor U5195 (N_5195,N_4014,N_4330);
and U5196 (N_5196,N_3541,N_3966);
nor U5197 (N_5197,N_4391,N_4272);
nand U5198 (N_5198,N_4258,N_4269);
nand U5199 (N_5199,N_3987,N_4060);
or U5200 (N_5200,N_3938,N_3845);
xnor U5201 (N_5201,N_3479,N_4492);
xor U5202 (N_5202,N_3268,N_3978);
or U5203 (N_5203,N_3902,N_3837);
and U5204 (N_5204,N_4452,N_3354);
and U5205 (N_5205,N_3552,N_3571);
nand U5206 (N_5206,N_3645,N_3615);
or U5207 (N_5207,N_3789,N_3348);
or U5208 (N_5208,N_3536,N_4419);
nor U5209 (N_5209,N_3857,N_3002);
nand U5210 (N_5210,N_4295,N_3230);
and U5211 (N_5211,N_3356,N_3387);
or U5212 (N_5212,N_4290,N_4472);
and U5213 (N_5213,N_4461,N_3485);
and U5214 (N_5214,N_3504,N_3605);
nor U5215 (N_5215,N_4309,N_4292);
or U5216 (N_5216,N_3073,N_3783);
xnor U5217 (N_5217,N_3518,N_4262);
and U5218 (N_5218,N_3912,N_3835);
xor U5219 (N_5219,N_3052,N_4337);
and U5220 (N_5220,N_3386,N_3001);
and U5221 (N_5221,N_3340,N_3907);
and U5222 (N_5222,N_3863,N_4013);
or U5223 (N_5223,N_3457,N_3995);
or U5224 (N_5224,N_3293,N_3023);
nor U5225 (N_5225,N_4248,N_4195);
nand U5226 (N_5226,N_4475,N_3217);
nand U5227 (N_5227,N_3933,N_3198);
and U5228 (N_5228,N_4340,N_3307);
or U5229 (N_5229,N_3272,N_4311);
nand U5230 (N_5230,N_3570,N_4132);
and U5231 (N_5231,N_3025,N_4105);
and U5232 (N_5232,N_3312,N_3267);
nor U5233 (N_5233,N_4380,N_3290);
nor U5234 (N_5234,N_3241,N_3451);
or U5235 (N_5235,N_3470,N_4463);
or U5236 (N_5236,N_3438,N_3773);
nor U5237 (N_5237,N_4368,N_3593);
and U5238 (N_5238,N_3730,N_3194);
nor U5239 (N_5239,N_4395,N_3819);
and U5240 (N_5240,N_3811,N_3045);
nor U5241 (N_5241,N_4069,N_3769);
nand U5242 (N_5242,N_3951,N_4367);
or U5243 (N_5243,N_3155,N_3510);
nand U5244 (N_5244,N_3066,N_3154);
nand U5245 (N_5245,N_3713,N_3772);
and U5246 (N_5246,N_3283,N_3218);
xnor U5247 (N_5247,N_3958,N_4047);
nor U5248 (N_5248,N_3949,N_4252);
xnor U5249 (N_5249,N_4151,N_3703);
nor U5250 (N_5250,N_3491,N_4176);
nand U5251 (N_5251,N_4171,N_3669);
xnor U5252 (N_5252,N_4009,N_4481);
xor U5253 (N_5253,N_3298,N_4419);
or U5254 (N_5254,N_3542,N_3514);
xnor U5255 (N_5255,N_4020,N_3284);
nand U5256 (N_5256,N_3504,N_3787);
or U5257 (N_5257,N_3924,N_3379);
xnor U5258 (N_5258,N_3459,N_3968);
nand U5259 (N_5259,N_3247,N_4198);
xor U5260 (N_5260,N_3652,N_3859);
nor U5261 (N_5261,N_3012,N_3966);
xnor U5262 (N_5262,N_3947,N_3123);
xnor U5263 (N_5263,N_4184,N_3690);
or U5264 (N_5264,N_3683,N_3371);
nor U5265 (N_5265,N_3323,N_4347);
nor U5266 (N_5266,N_3207,N_4142);
nor U5267 (N_5267,N_3694,N_4238);
and U5268 (N_5268,N_3003,N_3462);
or U5269 (N_5269,N_4345,N_3808);
nor U5270 (N_5270,N_3352,N_4147);
or U5271 (N_5271,N_3943,N_3296);
xor U5272 (N_5272,N_3632,N_3747);
xor U5273 (N_5273,N_4241,N_3505);
nor U5274 (N_5274,N_4358,N_4131);
xnor U5275 (N_5275,N_3846,N_3441);
nand U5276 (N_5276,N_4348,N_3896);
or U5277 (N_5277,N_3729,N_3632);
or U5278 (N_5278,N_3735,N_3415);
or U5279 (N_5279,N_4034,N_3776);
nor U5280 (N_5280,N_3093,N_3604);
nand U5281 (N_5281,N_3704,N_3075);
xnor U5282 (N_5282,N_4082,N_4096);
and U5283 (N_5283,N_3146,N_3399);
and U5284 (N_5284,N_3485,N_4474);
nand U5285 (N_5285,N_3250,N_3587);
xnor U5286 (N_5286,N_3724,N_3937);
nand U5287 (N_5287,N_3673,N_3295);
and U5288 (N_5288,N_3464,N_4211);
or U5289 (N_5289,N_4298,N_4472);
and U5290 (N_5290,N_4448,N_3228);
nand U5291 (N_5291,N_3465,N_3584);
nand U5292 (N_5292,N_3881,N_4061);
nand U5293 (N_5293,N_4419,N_3681);
and U5294 (N_5294,N_3571,N_3819);
nor U5295 (N_5295,N_4099,N_3325);
and U5296 (N_5296,N_4316,N_3958);
nand U5297 (N_5297,N_3018,N_3540);
xor U5298 (N_5298,N_3734,N_3579);
nand U5299 (N_5299,N_4313,N_4095);
or U5300 (N_5300,N_3108,N_4292);
nand U5301 (N_5301,N_3691,N_4377);
nor U5302 (N_5302,N_4017,N_3648);
nor U5303 (N_5303,N_3631,N_3178);
or U5304 (N_5304,N_4080,N_3102);
or U5305 (N_5305,N_3605,N_3395);
nand U5306 (N_5306,N_4200,N_3627);
and U5307 (N_5307,N_4087,N_4212);
nor U5308 (N_5308,N_4208,N_3909);
nor U5309 (N_5309,N_3785,N_3152);
nand U5310 (N_5310,N_3370,N_4332);
xnor U5311 (N_5311,N_3238,N_3688);
nor U5312 (N_5312,N_4026,N_3030);
nor U5313 (N_5313,N_4248,N_3827);
xor U5314 (N_5314,N_3512,N_3039);
xor U5315 (N_5315,N_4342,N_4128);
and U5316 (N_5316,N_4491,N_3574);
nor U5317 (N_5317,N_3501,N_4420);
or U5318 (N_5318,N_4373,N_4451);
nor U5319 (N_5319,N_3574,N_3744);
and U5320 (N_5320,N_3415,N_3187);
nor U5321 (N_5321,N_4271,N_4376);
and U5322 (N_5322,N_3445,N_3708);
and U5323 (N_5323,N_4023,N_3355);
nor U5324 (N_5324,N_3786,N_3438);
xor U5325 (N_5325,N_4221,N_4026);
xor U5326 (N_5326,N_3178,N_3198);
and U5327 (N_5327,N_3454,N_3316);
and U5328 (N_5328,N_3286,N_3075);
nand U5329 (N_5329,N_3869,N_3053);
nor U5330 (N_5330,N_4378,N_3772);
nand U5331 (N_5331,N_4291,N_3665);
nor U5332 (N_5332,N_3679,N_4001);
nor U5333 (N_5333,N_4121,N_3703);
or U5334 (N_5334,N_4346,N_3157);
nor U5335 (N_5335,N_3183,N_3878);
nor U5336 (N_5336,N_3788,N_4293);
nor U5337 (N_5337,N_4427,N_3717);
or U5338 (N_5338,N_3254,N_4370);
xor U5339 (N_5339,N_3364,N_3712);
and U5340 (N_5340,N_4314,N_4003);
xor U5341 (N_5341,N_3306,N_3362);
nor U5342 (N_5342,N_3301,N_3771);
and U5343 (N_5343,N_4435,N_3085);
nand U5344 (N_5344,N_4349,N_4097);
and U5345 (N_5345,N_3760,N_4068);
xnor U5346 (N_5346,N_3237,N_3376);
nor U5347 (N_5347,N_3335,N_4138);
and U5348 (N_5348,N_3930,N_3721);
or U5349 (N_5349,N_3033,N_3942);
xnor U5350 (N_5350,N_3700,N_3973);
xnor U5351 (N_5351,N_3502,N_4049);
or U5352 (N_5352,N_3607,N_3655);
or U5353 (N_5353,N_3963,N_3709);
nor U5354 (N_5354,N_3897,N_3115);
xor U5355 (N_5355,N_3327,N_4367);
nand U5356 (N_5356,N_3292,N_4361);
or U5357 (N_5357,N_4385,N_3757);
nand U5358 (N_5358,N_3757,N_3128);
nor U5359 (N_5359,N_3220,N_4377);
nor U5360 (N_5360,N_3284,N_4309);
xor U5361 (N_5361,N_3201,N_3700);
and U5362 (N_5362,N_4483,N_3535);
nor U5363 (N_5363,N_4186,N_4050);
or U5364 (N_5364,N_3184,N_3363);
nor U5365 (N_5365,N_3910,N_3112);
or U5366 (N_5366,N_3690,N_3090);
xnor U5367 (N_5367,N_3481,N_3684);
nand U5368 (N_5368,N_3475,N_4245);
and U5369 (N_5369,N_3633,N_3073);
nor U5370 (N_5370,N_4494,N_4372);
nor U5371 (N_5371,N_3195,N_3945);
or U5372 (N_5372,N_3457,N_3249);
xnor U5373 (N_5373,N_4085,N_4369);
nand U5374 (N_5374,N_3244,N_4219);
nor U5375 (N_5375,N_3937,N_3426);
or U5376 (N_5376,N_3919,N_3110);
or U5377 (N_5377,N_3574,N_4007);
nor U5378 (N_5378,N_3402,N_3561);
nor U5379 (N_5379,N_3731,N_4186);
or U5380 (N_5380,N_3928,N_3003);
nand U5381 (N_5381,N_4263,N_3062);
and U5382 (N_5382,N_3872,N_4299);
xor U5383 (N_5383,N_3336,N_3509);
nand U5384 (N_5384,N_3396,N_4182);
nor U5385 (N_5385,N_3502,N_4134);
xnor U5386 (N_5386,N_3318,N_3415);
nand U5387 (N_5387,N_3445,N_4194);
nand U5388 (N_5388,N_3811,N_3968);
or U5389 (N_5389,N_3638,N_3966);
or U5390 (N_5390,N_3005,N_3157);
and U5391 (N_5391,N_4436,N_3920);
or U5392 (N_5392,N_4301,N_3722);
nor U5393 (N_5393,N_4485,N_4370);
nand U5394 (N_5394,N_3587,N_3745);
nand U5395 (N_5395,N_4449,N_3696);
and U5396 (N_5396,N_3816,N_3745);
nor U5397 (N_5397,N_3585,N_3517);
and U5398 (N_5398,N_3345,N_3268);
or U5399 (N_5399,N_3016,N_3692);
nand U5400 (N_5400,N_3240,N_3892);
xnor U5401 (N_5401,N_4336,N_3552);
xnor U5402 (N_5402,N_3538,N_3465);
xor U5403 (N_5403,N_3858,N_3318);
and U5404 (N_5404,N_3701,N_3917);
or U5405 (N_5405,N_3349,N_3724);
xor U5406 (N_5406,N_3551,N_3743);
or U5407 (N_5407,N_3482,N_3336);
xnor U5408 (N_5408,N_3874,N_3645);
nor U5409 (N_5409,N_3625,N_4317);
or U5410 (N_5410,N_3510,N_3722);
nand U5411 (N_5411,N_4368,N_3142);
xor U5412 (N_5412,N_3552,N_3726);
nor U5413 (N_5413,N_4492,N_3735);
nor U5414 (N_5414,N_4257,N_4463);
or U5415 (N_5415,N_3357,N_3544);
and U5416 (N_5416,N_4368,N_3041);
nand U5417 (N_5417,N_4312,N_3626);
nand U5418 (N_5418,N_3874,N_3965);
nor U5419 (N_5419,N_3653,N_3841);
and U5420 (N_5420,N_3205,N_3927);
xor U5421 (N_5421,N_4318,N_4450);
nor U5422 (N_5422,N_3064,N_3291);
nand U5423 (N_5423,N_3618,N_3880);
nand U5424 (N_5424,N_4097,N_4414);
nor U5425 (N_5425,N_4344,N_3988);
nand U5426 (N_5426,N_3036,N_4387);
xor U5427 (N_5427,N_4257,N_3844);
and U5428 (N_5428,N_3259,N_3856);
or U5429 (N_5429,N_4436,N_3280);
xor U5430 (N_5430,N_3909,N_3170);
nor U5431 (N_5431,N_3293,N_4212);
or U5432 (N_5432,N_3465,N_4474);
and U5433 (N_5433,N_3500,N_3557);
or U5434 (N_5434,N_3567,N_3186);
xor U5435 (N_5435,N_3274,N_3404);
or U5436 (N_5436,N_4202,N_3175);
nand U5437 (N_5437,N_4336,N_3505);
xnor U5438 (N_5438,N_4032,N_3199);
xor U5439 (N_5439,N_3645,N_3279);
and U5440 (N_5440,N_3651,N_3919);
nand U5441 (N_5441,N_3747,N_3643);
nor U5442 (N_5442,N_3869,N_4443);
and U5443 (N_5443,N_3100,N_3931);
nor U5444 (N_5444,N_3354,N_3936);
nor U5445 (N_5445,N_4201,N_3304);
xnor U5446 (N_5446,N_3479,N_3751);
nor U5447 (N_5447,N_3951,N_3367);
nor U5448 (N_5448,N_3060,N_4132);
xor U5449 (N_5449,N_4443,N_3420);
xor U5450 (N_5450,N_4067,N_4150);
or U5451 (N_5451,N_3557,N_3981);
and U5452 (N_5452,N_4449,N_3019);
nand U5453 (N_5453,N_4334,N_4225);
nand U5454 (N_5454,N_3956,N_4088);
nand U5455 (N_5455,N_4193,N_3669);
or U5456 (N_5456,N_3730,N_3826);
xor U5457 (N_5457,N_3487,N_4101);
nand U5458 (N_5458,N_4356,N_4477);
nor U5459 (N_5459,N_3027,N_3177);
nand U5460 (N_5460,N_4206,N_3902);
and U5461 (N_5461,N_4185,N_4437);
nor U5462 (N_5462,N_3442,N_4209);
xnor U5463 (N_5463,N_3916,N_3526);
or U5464 (N_5464,N_3022,N_4284);
or U5465 (N_5465,N_3174,N_3088);
nand U5466 (N_5466,N_3521,N_3945);
nand U5467 (N_5467,N_3676,N_4253);
and U5468 (N_5468,N_4026,N_4042);
or U5469 (N_5469,N_4426,N_4430);
xor U5470 (N_5470,N_3335,N_3483);
nand U5471 (N_5471,N_3157,N_3419);
nor U5472 (N_5472,N_4455,N_3779);
xnor U5473 (N_5473,N_4478,N_3350);
or U5474 (N_5474,N_4101,N_3647);
or U5475 (N_5475,N_3182,N_3237);
nand U5476 (N_5476,N_3521,N_4446);
xnor U5477 (N_5477,N_3262,N_3881);
nor U5478 (N_5478,N_3063,N_3736);
and U5479 (N_5479,N_3100,N_3435);
xnor U5480 (N_5480,N_3705,N_3978);
nor U5481 (N_5481,N_3366,N_3375);
xnor U5482 (N_5482,N_4345,N_3664);
xor U5483 (N_5483,N_4346,N_4027);
nor U5484 (N_5484,N_4029,N_3952);
xnor U5485 (N_5485,N_4122,N_3007);
or U5486 (N_5486,N_4097,N_3315);
xnor U5487 (N_5487,N_3161,N_4079);
or U5488 (N_5488,N_4430,N_3223);
nor U5489 (N_5489,N_3188,N_3764);
xor U5490 (N_5490,N_3799,N_3537);
xnor U5491 (N_5491,N_3947,N_3250);
and U5492 (N_5492,N_3992,N_3973);
nand U5493 (N_5493,N_4000,N_4450);
nor U5494 (N_5494,N_3753,N_3589);
nor U5495 (N_5495,N_3998,N_3736);
xor U5496 (N_5496,N_4136,N_3733);
nor U5497 (N_5497,N_4364,N_4310);
xor U5498 (N_5498,N_4097,N_3354);
and U5499 (N_5499,N_4252,N_3178);
and U5500 (N_5500,N_4030,N_3843);
and U5501 (N_5501,N_4318,N_3483);
nand U5502 (N_5502,N_3881,N_3663);
nor U5503 (N_5503,N_3973,N_3555);
and U5504 (N_5504,N_4396,N_4028);
and U5505 (N_5505,N_4102,N_4483);
or U5506 (N_5506,N_3966,N_4262);
nor U5507 (N_5507,N_3846,N_3121);
nor U5508 (N_5508,N_4392,N_3146);
or U5509 (N_5509,N_3907,N_3270);
and U5510 (N_5510,N_4349,N_3855);
xor U5511 (N_5511,N_4317,N_3898);
nand U5512 (N_5512,N_3377,N_4133);
and U5513 (N_5513,N_4466,N_3965);
or U5514 (N_5514,N_3197,N_3977);
xnor U5515 (N_5515,N_4375,N_3502);
xor U5516 (N_5516,N_3808,N_3935);
nor U5517 (N_5517,N_3472,N_3678);
nand U5518 (N_5518,N_3931,N_3590);
xnor U5519 (N_5519,N_3977,N_4432);
and U5520 (N_5520,N_3039,N_3548);
nor U5521 (N_5521,N_4279,N_4111);
xor U5522 (N_5522,N_4462,N_3346);
nor U5523 (N_5523,N_4493,N_4289);
xnor U5524 (N_5524,N_3235,N_4393);
xor U5525 (N_5525,N_3094,N_3974);
and U5526 (N_5526,N_4226,N_4350);
or U5527 (N_5527,N_3436,N_3489);
xnor U5528 (N_5528,N_4186,N_3267);
or U5529 (N_5529,N_3950,N_4312);
nor U5530 (N_5530,N_4128,N_3346);
or U5531 (N_5531,N_4164,N_3836);
nand U5532 (N_5532,N_3912,N_4467);
and U5533 (N_5533,N_3975,N_4396);
or U5534 (N_5534,N_4336,N_3950);
xor U5535 (N_5535,N_4234,N_4440);
nand U5536 (N_5536,N_4030,N_4416);
nor U5537 (N_5537,N_3816,N_3957);
nand U5538 (N_5538,N_3782,N_3834);
nor U5539 (N_5539,N_3171,N_4134);
nand U5540 (N_5540,N_3588,N_4446);
xor U5541 (N_5541,N_3722,N_3317);
nor U5542 (N_5542,N_3565,N_3083);
xor U5543 (N_5543,N_3559,N_4374);
or U5544 (N_5544,N_3016,N_3798);
nor U5545 (N_5545,N_3041,N_3474);
nand U5546 (N_5546,N_4235,N_4110);
xor U5547 (N_5547,N_4073,N_4166);
xor U5548 (N_5548,N_3469,N_3084);
or U5549 (N_5549,N_3218,N_3732);
xor U5550 (N_5550,N_3362,N_3428);
nor U5551 (N_5551,N_3150,N_3629);
or U5552 (N_5552,N_3248,N_3580);
or U5553 (N_5553,N_3561,N_3489);
xnor U5554 (N_5554,N_3472,N_4494);
and U5555 (N_5555,N_3246,N_3534);
and U5556 (N_5556,N_3074,N_3103);
nand U5557 (N_5557,N_3819,N_3481);
nor U5558 (N_5558,N_3827,N_3962);
nand U5559 (N_5559,N_3047,N_4433);
and U5560 (N_5560,N_3634,N_3867);
nor U5561 (N_5561,N_4166,N_4212);
and U5562 (N_5562,N_3294,N_4206);
and U5563 (N_5563,N_3716,N_3451);
and U5564 (N_5564,N_3112,N_3401);
and U5565 (N_5565,N_4212,N_3945);
xnor U5566 (N_5566,N_3536,N_3678);
xnor U5567 (N_5567,N_3943,N_4121);
or U5568 (N_5568,N_3296,N_4016);
or U5569 (N_5569,N_4405,N_3589);
nand U5570 (N_5570,N_3725,N_3643);
or U5571 (N_5571,N_4155,N_3313);
xnor U5572 (N_5572,N_3846,N_4107);
nor U5573 (N_5573,N_4098,N_3453);
nor U5574 (N_5574,N_3399,N_4131);
nor U5575 (N_5575,N_3087,N_3277);
nor U5576 (N_5576,N_3290,N_3793);
or U5577 (N_5577,N_3434,N_4310);
nand U5578 (N_5578,N_3727,N_3505);
nand U5579 (N_5579,N_3357,N_3741);
and U5580 (N_5580,N_3665,N_4412);
or U5581 (N_5581,N_3394,N_3307);
nor U5582 (N_5582,N_3085,N_3303);
and U5583 (N_5583,N_4104,N_4270);
or U5584 (N_5584,N_3613,N_3150);
nor U5585 (N_5585,N_3424,N_3531);
and U5586 (N_5586,N_3108,N_3789);
xnor U5587 (N_5587,N_4052,N_3910);
and U5588 (N_5588,N_4464,N_3805);
nand U5589 (N_5589,N_4143,N_4196);
xnor U5590 (N_5590,N_3222,N_4314);
nor U5591 (N_5591,N_3212,N_3323);
and U5592 (N_5592,N_3923,N_4058);
nor U5593 (N_5593,N_3764,N_3399);
and U5594 (N_5594,N_3768,N_3112);
and U5595 (N_5595,N_3914,N_3868);
nand U5596 (N_5596,N_3885,N_3705);
nor U5597 (N_5597,N_3861,N_3954);
nand U5598 (N_5598,N_3017,N_3455);
or U5599 (N_5599,N_3597,N_3749);
or U5600 (N_5600,N_4203,N_4090);
nand U5601 (N_5601,N_3428,N_3014);
nor U5602 (N_5602,N_4441,N_4459);
xor U5603 (N_5603,N_4131,N_3888);
and U5604 (N_5604,N_3828,N_3613);
nor U5605 (N_5605,N_3747,N_3940);
nand U5606 (N_5606,N_3283,N_3458);
xor U5607 (N_5607,N_3454,N_3715);
nor U5608 (N_5608,N_3330,N_4479);
xor U5609 (N_5609,N_3113,N_3439);
nor U5610 (N_5610,N_3196,N_4037);
nor U5611 (N_5611,N_3146,N_3944);
nand U5612 (N_5612,N_3714,N_4033);
xor U5613 (N_5613,N_4482,N_3325);
nor U5614 (N_5614,N_3018,N_3195);
and U5615 (N_5615,N_3059,N_3512);
nand U5616 (N_5616,N_3724,N_3080);
nand U5617 (N_5617,N_3942,N_3821);
and U5618 (N_5618,N_3135,N_3114);
xnor U5619 (N_5619,N_4255,N_3498);
xor U5620 (N_5620,N_3203,N_4415);
nor U5621 (N_5621,N_3420,N_3380);
or U5622 (N_5622,N_4212,N_4285);
nor U5623 (N_5623,N_3460,N_3005);
nand U5624 (N_5624,N_4368,N_4189);
nand U5625 (N_5625,N_4316,N_3590);
and U5626 (N_5626,N_3716,N_3437);
nor U5627 (N_5627,N_4297,N_3615);
or U5628 (N_5628,N_4390,N_4166);
xor U5629 (N_5629,N_4352,N_4475);
and U5630 (N_5630,N_3724,N_3452);
and U5631 (N_5631,N_3769,N_3344);
or U5632 (N_5632,N_3885,N_3259);
and U5633 (N_5633,N_4130,N_3172);
nor U5634 (N_5634,N_3712,N_3041);
xor U5635 (N_5635,N_3231,N_3901);
nor U5636 (N_5636,N_4058,N_3373);
or U5637 (N_5637,N_4365,N_3286);
xnor U5638 (N_5638,N_4462,N_4413);
xnor U5639 (N_5639,N_3647,N_3618);
nor U5640 (N_5640,N_3731,N_4335);
xnor U5641 (N_5641,N_4237,N_3406);
nand U5642 (N_5642,N_4373,N_3740);
and U5643 (N_5643,N_4215,N_3873);
nor U5644 (N_5644,N_3110,N_3703);
xor U5645 (N_5645,N_4276,N_4052);
and U5646 (N_5646,N_3311,N_4140);
xnor U5647 (N_5647,N_3895,N_3109);
xor U5648 (N_5648,N_4000,N_3560);
nor U5649 (N_5649,N_3319,N_3470);
or U5650 (N_5650,N_4324,N_3491);
xor U5651 (N_5651,N_3038,N_4105);
or U5652 (N_5652,N_3361,N_4174);
nor U5653 (N_5653,N_3213,N_3697);
or U5654 (N_5654,N_3794,N_4403);
or U5655 (N_5655,N_4332,N_3930);
or U5656 (N_5656,N_4304,N_3665);
xor U5657 (N_5657,N_3054,N_3356);
and U5658 (N_5658,N_4104,N_3735);
and U5659 (N_5659,N_3664,N_3696);
nand U5660 (N_5660,N_3657,N_4013);
and U5661 (N_5661,N_3284,N_4429);
xnor U5662 (N_5662,N_3524,N_4356);
xnor U5663 (N_5663,N_4161,N_3325);
and U5664 (N_5664,N_3451,N_3384);
nand U5665 (N_5665,N_3760,N_3764);
nor U5666 (N_5666,N_4188,N_3021);
xnor U5667 (N_5667,N_3866,N_3037);
and U5668 (N_5668,N_4008,N_4078);
or U5669 (N_5669,N_4060,N_3937);
or U5670 (N_5670,N_3514,N_4020);
and U5671 (N_5671,N_4186,N_4118);
nor U5672 (N_5672,N_3400,N_4379);
xor U5673 (N_5673,N_3689,N_3616);
and U5674 (N_5674,N_3681,N_3721);
xnor U5675 (N_5675,N_4127,N_4122);
xor U5676 (N_5676,N_3460,N_3349);
nor U5677 (N_5677,N_3536,N_3763);
nand U5678 (N_5678,N_4446,N_3310);
xor U5679 (N_5679,N_3449,N_3528);
xor U5680 (N_5680,N_4068,N_4405);
and U5681 (N_5681,N_3064,N_3101);
or U5682 (N_5682,N_3074,N_4127);
xnor U5683 (N_5683,N_3948,N_3333);
nor U5684 (N_5684,N_3661,N_4432);
or U5685 (N_5685,N_3224,N_3522);
nand U5686 (N_5686,N_3896,N_4208);
nand U5687 (N_5687,N_3926,N_4410);
xor U5688 (N_5688,N_3664,N_3820);
nand U5689 (N_5689,N_3309,N_3426);
or U5690 (N_5690,N_4347,N_4390);
or U5691 (N_5691,N_3807,N_4190);
xnor U5692 (N_5692,N_4413,N_4294);
and U5693 (N_5693,N_3669,N_3277);
nand U5694 (N_5694,N_3709,N_3300);
xor U5695 (N_5695,N_4277,N_3969);
or U5696 (N_5696,N_3070,N_4271);
or U5697 (N_5697,N_3596,N_4225);
and U5698 (N_5698,N_3870,N_3459);
or U5699 (N_5699,N_4426,N_4298);
nor U5700 (N_5700,N_3931,N_3153);
or U5701 (N_5701,N_4042,N_3323);
and U5702 (N_5702,N_3434,N_4107);
nor U5703 (N_5703,N_3795,N_3617);
xnor U5704 (N_5704,N_4494,N_3591);
nor U5705 (N_5705,N_3606,N_4226);
nor U5706 (N_5706,N_4185,N_3151);
nand U5707 (N_5707,N_4396,N_3877);
nor U5708 (N_5708,N_3154,N_4420);
nand U5709 (N_5709,N_3430,N_3105);
and U5710 (N_5710,N_3427,N_3658);
or U5711 (N_5711,N_4149,N_3183);
and U5712 (N_5712,N_3255,N_3239);
or U5713 (N_5713,N_3460,N_3687);
xor U5714 (N_5714,N_3972,N_3610);
nand U5715 (N_5715,N_3631,N_3435);
xnor U5716 (N_5716,N_3926,N_3469);
nand U5717 (N_5717,N_4184,N_3013);
nor U5718 (N_5718,N_3569,N_3299);
and U5719 (N_5719,N_4281,N_3786);
xor U5720 (N_5720,N_3972,N_3197);
nand U5721 (N_5721,N_4126,N_4483);
and U5722 (N_5722,N_4223,N_3365);
and U5723 (N_5723,N_3048,N_4285);
or U5724 (N_5724,N_3245,N_3118);
xor U5725 (N_5725,N_3647,N_4072);
and U5726 (N_5726,N_3070,N_3327);
nand U5727 (N_5727,N_4139,N_3308);
and U5728 (N_5728,N_3268,N_3829);
nand U5729 (N_5729,N_3783,N_3403);
or U5730 (N_5730,N_3139,N_4084);
nor U5731 (N_5731,N_4157,N_4450);
and U5732 (N_5732,N_3410,N_3419);
xor U5733 (N_5733,N_3293,N_3973);
nor U5734 (N_5734,N_3912,N_3326);
xor U5735 (N_5735,N_3552,N_3646);
and U5736 (N_5736,N_3915,N_3738);
xnor U5737 (N_5737,N_3011,N_3838);
or U5738 (N_5738,N_3166,N_3629);
xor U5739 (N_5739,N_3710,N_3098);
nand U5740 (N_5740,N_3975,N_3569);
nor U5741 (N_5741,N_3066,N_3055);
or U5742 (N_5742,N_4207,N_3215);
nor U5743 (N_5743,N_3536,N_3413);
xnor U5744 (N_5744,N_4358,N_4034);
nor U5745 (N_5745,N_3122,N_3079);
and U5746 (N_5746,N_4052,N_3059);
nand U5747 (N_5747,N_3253,N_3855);
or U5748 (N_5748,N_3338,N_3652);
nor U5749 (N_5749,N_4068,N_3033);
and U5750 (N_5750,N_3383,N_3189);
xor U5751 (N_5751,N_3522,N_3475);
or U5752 (N_5752,N_3298,N_3611);
nor U5753 (N_5753,N_3595,N_3981);
nand U5754 (N_5754,N_3799,N_4351);
nand U5755 (N_5755,N_4468,N_3327);
or U5756 (N_5756,N_3834,N_3039);
and U5757 (N_5757,N_4090,N_3002);
and U5758 (N_5758,N_3955,N_3583);
xnor U5759 (N_5759,N_3233,N_3400);
or U5760 (N_5760,N_4338,N_4479);
xnor U5761 (N_5761,N_3896,N_3027);
xnor U5762 (N_5762,N_4387,N_4325);
and U5763 (N_5763,N_4473,N_4318);
nor U5764 (N_5764,N_3264,N_4348);
nand U5765 (N_5765,N_3983,N_4134);
and U5766 (N_5766,N_3215,N_4266);
nand U5767 (N_5767,N_4394,N_3970);
xnor U5768 (N_5768,N_4266,N_4187);
nor U5769 (N_5769,N_3386,N_3797);
nand U5770 (N_5770,N_3886,N_4379);
nand U5771 (N_5771,N_4090,N_4372);
or U5772 (N_5772,N_3521,N_3273);
xor U5773 (N_5773,N_3374,N_3876);
nand U5774 (N_5774,N_3831,N_3122);
and U5775 (N_5775,N_4119,N_3382);
nand U5776 (N_5776,N_3778,N_3469);
and U5777 (N_5777,N_3235,N_4156);
nor U5778 (N_5778,N_4149,N_4462);
nand U5779 (N_5779,N_4221,N_3378);
nand U5780 (N_5780,N_3763,N_4120);
or U5781 (N_5781,N_3622,N_3614);
or U5782 (N_5782,N_3293,N_3743);
xor U5783 (N_5783,N_3277,N_3208);
xnor U5784 (N_5784,N_3192,N_4218);
xnor U5785 (N_5785,N_3182,N_3353);
or U5786 (N_5786,N_3206,N_4382);
nand U5787 (N_5787,N_3980,N_4023);
xor U5788 (N_5788,N_3586,N_3142);
nand U5789 (N_5789,N_3320,N_3591);
and U5790 (N_5790,N_3695,N_3100);
xor U5791 (N_5791,N_3063,N_4073);
or U5792 (N_5792,N_4320,N_3522);
or U5793 (N_5793,N_4462,N_3162);
xor U5794 (N_5794,N_3992,N_3656);
and U5795 (N_5795,N_4049,N_3028);
nand U5796 (N_5796,N_3768,N_3853);
and U5797 (N_5797,N_3146,N_3696);
nand U5798 (N_5798,N_4485,N_4251);
or U5799 (N_5799,N_4484,N_4183);
nand U5800 (N_5800,N_4493,N_3109);
nand U5801 (N_5801,N_3542,N_3084);
nor U5802 (N_5802,N_3357,N_4493);
nand U5803 (N_5803,N_3035,N_3554);
or U5804 (N_5804,N_4029,N_3370);
nor U5805 (N_5805,N_4477,N_3186);
xor U5806 (N_5806,N_3464,N_3260);
nand U5807 (N_5807,N_3646,N_3899);
or U5808 (N_5808,N_3162,N_3298);
or U5809 (N_5809,N_4327,N_3747);
and U5810 (N_5810,N_3530,N_3801);
nand U5811 (N_5811,N_4465,N_4225);
nand U5812 (N_5812,N_4200,N_3916);
nor U5813 (N_5813,N_3933,N_4262);
or U5814 (N_5814,N_4155,N_3377);
nand U5815 (N_5815,N_3377,N_3044);
nand U5816 (N_5816,N_4105,N_4408);
xnor U5817 (N_5817,N_4167,N_3933);
nand U5818 (N_5818,N_3346,N_4488);
xor U5819 (N_5819,N_3848,N_4280);
nand U5820 (N_5820,N_3009,N_4014);
nand U5821 (N_5821,N_3618,N_3609);
nand U5822 (N_5822,N_3368,N_4018);
and U5823 (N_5823,N_4061,N_3323);
nor U5824 (N_5824,N_3746,N_3339);
and U5825 (N_5825,N_3869,N_3921);
xor U5826 (N_5826,N_3834,N_4425);
and U5827 (N_5827,N_3252,N_3159);
xnor U5828 (N_5828,N_4000,N_4311);
xnor U5829 (N_5829,N_3574,N_4004);
nand U5830 (N_5830,N_3081,N_4087);
xor U5831 (N_5831,N_3970,N_4466);
nor U5832 (N_5832,N_3804,N_3019);
and U5833 (N_5833,N_4106,N_4287);
xor U5834 (N_5834,N_4196,N_3068);
xor U5835 (N_5835,N_4408,N_3055);
or U5836 (N_5836,N_4424,N_3149);
xor U5837 (N_5837,N_3642,N_3078);
and U5838 (N_5838,N_3865,N_4097);
xor U5839 (N_5839,N_3695,N_3450);
nand U5840 (N_5840,N_4002,N_4086);
xor U5841 (N_5841,N_3233,N_3718);
and U5842 (N_5842,N_3365,N_3069);
xnor U5843 (N_5843,N_4440,N_4212);
nand U5844 (N_5844,N_3217,N_3390);
or U5845 (N_5845,N_3829,N_3208);
xor U5846 (N_5846,N_4092,N_4463);
xor U5847 (N_5847,N_3567,N_4388);
and U5848 (N_5848,N_3277,N_3657);
nand U5849 (N_5849,N_4003,N_4445);
nor U5850 (N_5850,N_3104,N_4236);
nand U5851 (N_5851,N_3177,N_3299);
and U5852 (N_5852,N_3226,N_4012);
and U5853 (N_5853,N_3874,N_3608);
or U5854 (N_5854,N_3423,N_3814);
nand U5855 (N_5855,N_3755,N_4446);
or U5856 (N_5856,N_3079,N_4130);
or U5857 (N_5857,N_3379,N_3760);
nand U5858 (N_5858,N_3193,N_3150);
and U5859 (N_5859,N_4250,N_3697);
or U5860 (N_5860,N_3268,N_4488);
and U5861 (N_5861,N_3119,N_3858);
or U5862 (N_5862,N_4307,N_4240);
or U5863 (N_5863,N_4099,N_3018);
and U5864 (N_5864,N_4473,N_3621);
nand U5865 (N_5865,N_3933,N_3265);
nor U5866 (N_5866,N_3435,N_4320);
xor U5867 (N_5867,N_3034,N_3674);
and U5868 (N_5868,N_4170,N_4096);
and U5869 (N_5869,N_3421,N_3255);
and U5870 (N_5870,N_3019,N_4297);
or U5871 (N_5871,N_3330,N_3370);
or U5872 (N_5872,N_4187,N_3262);
nor U5873 (N_5873,N_3804,N_3891);
nor U5874 (N_5874,N_3668,N_3042);
xnor U5875 (N_5875,N_3900,N_3467);
and U5876 (N_5876,N_3076,N_3795);
or U5877 (N_5877,N_3617,N_4076);
xor U5878 (N_5878,N_3858,N_4164);
or U5879 (N_5879,N_4310,N_3484);
or U5880 (N_5880,N_3017,N_4440);
nand U5881 (N_5881,N_3723,N_4391);
xor U5882 (N_5882,N_3036,N_4482);
xor U5883 (N_5883,N_3370,N_3719);
or U5884 (N_5884,N_3372,N_4022);
xor U5885 (N_5885,N_3909,N_4144);
xor U5886 (N_5886,N_4209,N_3451);
nor U5887 (N_5887,N_3777,N_3372);
and U5888 (N_5888,N_4475,N_3391);
nor U5889 (N_5889,N_4428,N_4380);
or U5890 (N_5890,N_3343,N_4213);
or U5891 (N_5891,N_3608,N_3135);
xnor U5892 (N_5892,N_3511,N_3615);
nand U5893 (N_5893,N_4187,N_3955);
nor U5894 (N_5894,N_3025,N_3125);
nand U5895 (N_5895,N_3853,N_4300);
xor U5896 (N_5896,N_3456,N_3448);
or U5897 (N_5897,N_3147,N_3870);
and U5898 (N_5898,N_3282,N_3859);
nor U5899 (N_5899,N_3529,N_3711);
and U5900 (N_5900,N_3393,N_3570);
and U5901 (N_5901,N_3530,N_3714);
nand U5902 (N_5902,N_3509,N_4146);
xnor U5903 (N_5903,N_3237,N_3624);
xor U5904 (N_5904,N_3866,N_4474);
and U5905 (N_5905,N_3770,N_3073);
and U5906 (N_5906,N_3728,N_3960);
nor U5907 (N_5907,N_3642,N_4466);
or U5908 (N_5908,N_3469,N_4200);
and U5909 (N_5909,N_4348,N_4093);
and U5910 (N_5910,N_3716,N_4199);
nand U5911 (N_5911,N_4305,N_3666);
and U5912 (N_5912,N_4458,N_3770);
xor U5913 (N_5913,N_3414,N_3659);
and U5914 (N_5914,N_3390,N_3967);
and U5915 (N_5915,N_4051,N_4048);
or U5916 (N_5916,N_4065,N_3052);
nor U5917 (N_5917,N_3812,N_3428);
and U5918 (N_5918,N_3881,N_4263);
nor U5919 (N_5919,N_4019,N_4097);
and U5920 (N_5920,N_3251,N_4054);
xnor U5921 (N_5921,N_3667,N_3593);
nand U5922 (N_5922,N_3548,N_4425);
nor U5923 (N_5923,N_3575,N_4262);
nand U5924 (N_5924,N_3584,N_3835);
or U5925 (N_5925,N_3916,N_3847);
nand U5926 (N_5926,N_4285,N_4439);
nor U5927 (N_5927,N_3616,N_3348);
or U5928 (N_5928,N_3777,N_3431);
nand U5929 (N_5929,N_4305,N_4136);
or U5930 (N_5930,N_3540,N_4182);
and U5931 (N_5931,N_3287,N_3101);
xnor U5932 (N_5932,N_3925,N_4113);
and U5933 (N_5933,N_3371,N_4174);
nand U5934 (N_5934,N_4088,N_4403);
or U5935 (N_5935,N_3459,N_3491);
nor U5936 (N_5936,N_3389,N_3226);
or U5937 (N_5937,N_4114,N_3484);
and U5938 (N_5938,N_3826,N_3934);
and U5939 (N_5939,N_3235,N_4175);
and U5940 (N_5940,N_3762,N_4133);
nor U5941 (N_5941,N_4331,N_4123);
or U5942 (N_5942,N_3414,N_3916);
xor U5943 (N_5943,N_3610,N_4128);
nor U5944 (N_5944,N_3043,N_3303);
nand U5945 (N_5945,N_3213,N_3955);
nor U5946 (N_5946,N_3760,N_4209);
nor U5947 (N_5947,N_3162,N_3904);
nor U5948 (N_5948,N_3202,N_4422);
or U5949 (N_5949,N_3382,N_3621);
or U5950 (N_5950,N_4440,N_4134);
or U5951 (N_5951,N_3554,N_3923);
and U5952 (N_5952,N_4159,N_3664);
and U5953 (N_5953,N_3972,N_3335);
xor U5954 (N_5954,N_3175,N_4377);
and U5955 (N_5955,N_4150,N_3608);
and U5956 (N_5956,N_4119,N_4418);
xor U5957 (N_5957,N_4270,N_4331);
and U5958 (N_5958,N_3237,N_4189);
or U5959 (N_5959,N_4381,N_3789);
xor U5960 (N_5960,N_3913,N_3450);
nand U5961 (N_5961,N_4053,N_4055);
nor U5962 (N_5962,N_4030,N_3612);
or U5963 (N_5963,N_4070,N_4473);
and U5964 (N_5964,N_4247,N_4034);
nor U5965 (N_5965,N_4132,N_3593);
nor U5966 (N_5966,N_3340,N_4236);
xor U5967 (N_5967,N_3257,N_3415);
nor U5968 (N_5968,N_4139,N_3765);
or U5969 (N_5969,N_4477,N_3214);
or U5970 (N_5970,N_3227,N_3584);
and U5971 (N_5971,N_4357,N_3317);
nor U5972 (N_5972,N_3221,N_4090);
nand U5973 (N_5973,N_3219,N_3819);
or U5974 (N_5974,N_3423,N_3782);
nand U5975 (N_5975,N_3658,N_3278);
nand U5976 (N_5976,N_4394,N_3408);
and U5977 (N_5977,N_3179,N_3808);
xor U5978 (N_5978,N_4122,N_3873);
and U5979 (N_5979,N_4316,N_3021);
nand U5980 (N_5980,N_3859,N_4348);
and U5981 (N_5981,N_3929,N_3308);
xnor U5982 (N_5982,N_3153,N_3094);
or U5983 (N_5983,N_3508,N_3545);
nor U5984 (N_5984,N_3923,N_3143);
nand U5985 (N_5985,N_3900,N_3558);
nand U5986 (N_5986,N_3742,N_3171);
xnor U5987 (N_5987,N_3726,N_3738);
xor U5988 (N_5988,N_3909,N_4462);
nand U5989 (N_5989,N_3674,N_4435);
or U5990 (N_5990,N_4423,N_4076);
nand U5991 (N_5991,N_3732,N_3848);
nor U5992 (N_5992,N_3903,N_3554);
or U5993 (N_5993,N_4181,N_4357);
nand U5994 (N_5994,N_3725,N_3618);
nand U5995 (N_5995,N_3353,N_4017);
nand U5996 (N_5996,N_3737,N_3258);
nor U5997 (N_5997,N_3010,N_4448);
or U5998 (N_5998,N_3149,N_3668);
or U5999 (N_5999,N_4406,N_3013);
nor U6000 (N_6000,N_5407,N_5536);
and U6001 (N_6001,N_5383,N_5488);
xor U6002 (N_6002,N_4967,N_4956);
xor U6003 (N_6003,N_5323,N_4861);
nand U6004 (N_6004,N_4917,N_4675);
nor U6005 (N_6005,N_4634,N_5212);
nand U6006 (N_6006,N_5576,N_5505);
nand U6007 (N_6007,N_5503,N_5763);
and U6008 (N_6008,N_5250,N_5298);
or U6009 (N_6009,N_5568,N_5064);
and U6010 (N_6010,N_5710,N_4929);
or U6011 (N_6011,N_4742,N_5045);
xnor U6012 (N_6012,N_5947,N_5902);
nor U6013 (N_6013,N_5377,N_4782);
or U6014 (N_6014,N_5873,N_5297);
or U6015 (N_6015,N_4893,N_4804);
nand U6016 (N_6016,N_4565,N_5230);
and U6017 (N_6017,N_4984,N_4784);
or U6018 (N_6018,N_5210,N_5721);
nand U6019 (N_6019,N_5700,N_4641);
and U6020 (N_6020,N_4875,N_4775);
and U6021 (N_6021,N_4665,N_5268);
or U6022 (N_6022,N_5941,N_5487);
nor U6023 (N_6023,N_5078,N_5754);
or U6024 (N_6024,N_5222,N_5807);
or U6025 (N_6025,N_5997,N_5107);
or U6026 (N_6026,N_5269,N_5110);
or U6027 (N_6027,N_4791,N_5315);
nand U6028 (N_6028,N_5467,N_4723);
nand U6029 (N_6029,N_4809,N_5002);
and U6030 (N_6030,N_4643,N_5195);
xor U6031 (N_6031,N_5314,N_4805);
nand U6032 (N_6032,N_4844,N_5845);
nor U6033 (N_6033,N_5897,N_5157);
nor U6034 (N_6034,N_5284,N_4683);
nor U6035 (N_6035,N_4873,N_4567);
xnor U6036 (N_6036,N_4661,N_4704);
nor U6037 (N_6037,N_4635,N_5464);
nor U6038 (N_6038,N_5272,N_5875);
and U6039 (N_6039,N_5402,N_5975);
and U6040 (N_6040,N_5019,N_4583);
or U6041 (N_6041,N_5563,N_5066);
nand U6042 (N_6042,N_5816,N_5933);
and U6043 (N_6043,N_5567,N_5709);
nand U6044 (N_6044,N_5663,N_4772);
xnor U6045 (N_6045,N_4667,N_5055);
nand U6046 (N_6046,N_5234,N_4858);
nand U6047 (N_6047,N_5499,N_4989);
nor U6048 (N_6048,N_4876,N_4783);
and U6049 (N_6049,N_4953,N_5137);
nor U6050 (N_6050,N_5634,N_5651);
nand U6051 (N_6051,N_5231,N_4644);
nor U6052 (N_6052,N_4934,N_4759);
nor U6053 (N_6053,N_5398,N_5028);
nand U6054 (N_6054,N_4773,N_5923);
nor U6055 (N_6055,N_4740,N_5591);
xor U6056 (N_6056,N_5860,N_4849);
nor U6057 (N_6057,N_5547,N_4733);
nor U6058 (N_6058,N_4698,N_5711);
xor U6059 (N_6059,N_5867,N_4749);
or U6060 (N_6060,N_4509,N_5207);
xor U6061 (N_6061,N_5558,N_4652);
and U6062 (N_6062,N_5176,N_4766);
nor U6063 (N_6063,N_4600,N_4793);
or U6064 (N_6064,N_5452,N_4883);
and U6065 (N_6065,N_5540,N_5043);
xor U6066 (N_6066,N_5332,N_5989);
and U6067 (N_6067,N_5804,N_4975);
nand U6068 (N_6068,N_5057,N_5512);
nand U6069 (N_6069,N_4713,N_4633);
nand U6070 (N_6070,N_4913,N_5324);
nor U6071 (N_6071,N_5815,N_5713);
nor U6072 (N_6072,N_5723,N_5824);
or U6073 (N_6073,N_4769,N_5500);
or U6074 (N_6074,N_5904,N_4719);
xnor U6075 (N_6075,N_5380,N_5492);
nor U6076 (N_6076,N_5665,N_5349);
nand U6077 (N_6077,N_5929,N_4886);
xnor U6078 (N_6078,N_5701,N_5001);
xor U6079 (N_6079,N_5186,N_5042);
or U6080 (N_6080,N_5498,N_5173);
nor U6081 (N_6081,N_5656,N_5046);
xnor U6082 (N_6082,N_5388,N_5906);
xor U6083 (N_6083,N_5917,N_5140);
and U6084 (N_6084,N_4559,N_4538);
or U6085 (N_6085,N_5138,N_4928);
xor U6086 (N_6086,N_5326,N_5361);
xor U6087 (N_6087,N_4959,N_4711);
or U6088 (N_6088,N_5616,N_4785);
xnor U6089 (N_6089,N_5310,N_5257);
and U6090 (N_6090,N_5708,N_5649);
nor U6091 (N_6091,N_5330,N_5992);
nand U6092 (N_6092,N_5356,N_5530);
or U6093 (N_6093,N_5574,N_5657);
and U6094 (N_6094,N_5116,N_5986);
or U6095 (N_6095,N_4828,N_5965);
and U6096 (N_6096,N_5539,N_5187);
xor U6097 (N_6097,N_5014,N_5274);
and U6098 (N_6098,N_4827,N_5910);
xor U6099 (N_6099,N_4799,N_5239);
nand U6100 (N_6100,N_5534,N_5853);
nor U6101 (N_6101,N_4969,N_5661);
or U6102 (N_6102,N_5320,N_5504);
nand U6103 (N_6103,N_4838,N_5171);
xor U6104 (N_6104,N_5757,N_5911);
nor U6105 (N_6105,N_5739,N_5892);
nand U6106 (N_6106,N_4700,N_5783);
and U6107 (N_6107,N_5821,N_5003);
xor U6108 (N_6108,N_5172,N_5448);
nor U6109 (N_6109,N_5866,N_4765);
or U6110 (N_6110,N_5553,N_5333);
xor U6111 (N_6111,N_4527,N_5637);
nor U6112 (N_6112,N_5981,N_5618);
or U6113 (N_6113,N_5404,N_4763);
xnor U6114 (N_6114,N_5000,N_5350);
or U6115 (N_6115,N_5516,N_5608);
and U6116 (N_6116,N_5973,N_4800);
or U6117 (N_6117,N_5409,N_4671);
and U6118 (N_6118,N_5422,N_4682);
xor U6119 (N_6119,N_5309,N_5327);
nor U6120 (N_6120,N_4914,N_4560);
nor U6121 (N_6121,N_4825,N_5061);
or U6122 (N_6122,N_5316,N_5146);
nor U6123 (N_6123,N_5185,N_5513);
and U6124 (N_6124,N_4903,N_4691);
nor U6125 (N_6125,N_5428,N_4856);
or U6126 (N_6126,N_4790,N_4576);
and U6127 (N_6127,N_5286,N_5972);
nor U6128 (N_6128,N_4689,N_5340);
or U6129 (N_6129,N_4970,N_4907);
nor U6130 (N_6130,N_5677,N_5366);
or U6131 (N_6131,N_5605,N_5680);
xnor U6132 (N_6132,N_4614,N_5205);
nor U6133 (N_6133,N_5961,N_4568);
nor U6134 (N_6134,N_5996,N_4620);
or U6135 (N_6135,N_4788,N_5664);
or U6136 (N_6136,N_4517,N_4736);
and U6137 (N_6137,N_5432,N_5518);
or U6138 (N_6138,N_5450,N_5347);
xnor U6139 (N_6139,N_5926,N_5049);
nor U6140 (N_6140,N_5510,N_5063);
nand U6141 (N_6141,N_5255,N_4944);
or U6142 (N_6142,N_4938,N_5672);
xnor U6143 (N_6143,N_5589,N_5753);
or U6144 (N_6144,N_5982,N_5397);
and U6145 (N_6145,N_5495,N_5208);
nor U6146 (N_6146,N_5979,N_5312);
nor U6147 (N_6147,N_4549,N_4915);
and U6148 (N_6148,N_4995,N_4728);
nand U6149 (N_6149,N_5174,N_4627);
or U6150 (N_6150,N_4982,N_4958);
nand U6151 (N_6151,N_4658,N_5582);
xor U6152 (N_6152,N_4739,N_5266);
and U6153 (N_6153,N_5264,N_4647);
and U6154 (N_6154,N_4555,N_4850);
and U6155 (N_6155,N_5123,N_4696);
and U6156 (N_6156,N_5431,N_5722);
nor U6157 (N_6157,N_5854,N_5196);
nor U6158 (N_6158,N_4690,N_5581);
and U6159 (N_6159,N_5957,N_5977);
nor U6160 (N_6160,N_4878,N_5502);
xnor U6161 (N_6161,N_4976,N_5937);
nand U6162 (N_6162,N_4720,N_5375);
and U6163 (N_6163,N_4891,N_4919);
and U6164 (N_6164,N_4801,N_4911);
and U6165 (N_6165,N_4706,N_4843);
nand U6166 (N_6166,N_5494,N_5777);
xor U6167 (N_6167,N_5802,N_4553);
or U6168 (N_6168,N_5344,N_5449);
and U6169 (N_6169,N_5561,N_5717);
nor U6170 (N_6170,N_5141,N_5243);
nor U6171 (N_6171,N_4566,N_5592);
xor U6172 (N_6172,N_5299,N_4610);
or U6173 (N_6173,N_5496,N_5552);
nor U6174 (N_6174,N_5016,N_4859);
xor U6175 (N_6175,N_4522,N_5348);
or U6176 (N_6176,N_5408,N_5541);
xor U6177 (N_6177,N_5863,N_4797);
nand U6178 (N_6178,N_5912,N_5287);
xnor U6179 (N_6179,N_5859,N_5376);
and U6180 (N_6180,N_5679,N_5006);
or U6181 (N_6181,N_4852,N_5158);
or U6182 (N_6182,N_4892,N_5412);
nand U6183 (N_6183,N_4653,N_5810);
and U6184 (N_6184,N_5068,N_5844);
xor U6185 (N_6185,N_5511,N_4776);
nand U6186 (N_6186,N_5319,N_4974);
xnor U6187 (N_6187,N_5650,N_4879);
and U6188 (N_6188,N_5420,N_5341);
or U6189 (N_6189,N_4694,N_5065);
nor U6190 (N_6190,N_5600,N_4676);
nand U6191 (N_6191,N_5751,N_5690);
nor U6192 (N_6192,N_5067,N_4586);
nand U6193 (N_6193,N_4543,N_5745);
and U6194 (N_6194,N_5771,N_5814);
or U6195 (N_6195,N_5719,N_5833);
xnor U6196 (N_6196,N_5900,N_4884);
and U6197 (N_6197,N_4507,N_4983);
xor U6198 (N_6198,N_5267,N_5152);
nand U6199 (N_6199,N_5085,N_5392);
or U6200 (N_6200,N_4999,N_4585);
nor U6201 (N_6201,N_5443,N_5405);
nor U6202 (N_6202,N_5183,N_4758);
nor U6203 (N_6203,N_5129,N_5162);
nand U6204 (N_6204,N_5092,N_5059);
xor U6205 (N_6205,N_5285,N_5189);
or U6206 (N_6206,N_5683,N_5275);
or U6207 (N_6207,N_4991,N_4598);
or U6208 (N_6208,N_5098,N_5079);
nand U6209 (N_6209,N_5096,N_5857);
or U6210 (N_6210,N_5031,N_5134);
and U6211 (N_6211,N_5336,N_5281);
nor U6212 (N_6212,N_5217,N_4881);
nor U6213 (N_6213,N_5778,N_4869);
or U6214 (N_6214,N_4823,N_5072);
xnor U6215 (N_6215,N_4607,N_5569);
xor U6216 (N_6216,N_4954,N_5038);
or U6217 (N_6217,N_4812,N_5242);
and U6218 (N_6218,N_5458,N_5696);
xor U6219 (N_6219,N_4948,N_4853);
or U6220 (N_6220,N_5232,N_4596);
and U6221 (N_6221,N_4997,N_5627);
nor U6222 (N_6222,N_4744,N_5945);
xnor U6223 (N_6223,N_4898,N_4557);
or U6224 (N_6224,N_5220,N_5542);
and U6225 (N_6225,N_5877,N_5226);
nand U6226 (N_6226,N_5258,N_5644);
and U6227 (N_6227,N_5070,N_4525);
nor U6228 (N_6228,N_5703,N_5288);
xnor U6229 (N_6229,N_4807,N_5642);
and U6230 (N_6230,N_4714,N_5638);
and U6231 (N_6231,N_5507,N_4539);
nand U6232 (N_6232,N_5084,N_5653);
nand U6233 (N_6233,N_5543,N_5612);
and U6234 (N_6234,N_4552,N_5521);
or U6235 (N_6235,N_4792,N_5074);
or U6236 (N_6236,N_5523,N_4837);
nor U6237 (N_6237,N_4702,N_5546);
and U6238 (N_6238,N_4924,N_5842);
xor U6239 (N_6239,N_5209,N_5290);
xnor U6240 (N_6240,N_5983,N_4636);
nor U6241 (N_6241,N_5675,N_5876);
or U6242 (N_6242,N_5473,N_5936);
xor U6243 (N_6243,N_4645,N_5856);
nand U6244 (N_6244,N_4528,N_4973);
xor U6245 (N_6245,N_5924,N_5953);
nand U6246 (N_6246,N_5741,N_5871);
and U6247 (N_6247,N_5378,N_5273);
nor U6248 (N_6248,N_4669,N_5598);
or U6249 (N_6249,N_5437,N_5706);
xnor U6250 (N_6250,N_4582,N_5594);
nand U6251 (N_6251,N_5832,N_5508);
xnor U6252 (N_6252,N_5619,N_4868);
and U6253 (N_6253,N_4612,N_5988);
xnor U6254 (N_6254,N_4595,N_4951);
nor U6255 (N_6255,N_5839,N_5565);
nor U6256 (N_6256,N_5426,N_5687);
and U6257 (N_6257,N_4615,N_5401);
nand U6258 (N_6258,N_5386,N_5438);
xnor U6259 (N_6259,N_5115,N_5825);
or U6260 (N_6260,N_5837,N_4960);
nor U6261 (N_6261,N_5396,N_5725);
or U6262 (N_6262,N_4544,N_5762);
xor U6263 (N_6263,N_5993,N_4685);
nor U6264 (N_6264,N_4894,N_5476);
xor U6265 (N_6265,N_5971,N_4777);
nor U6266 (N_6266,N_5237,N_5313);
nor U6267 (N_6267,N_5538,N_5203);
nor U6268 (N_6268,N_5305,N_5279);
or U6269 (N_6269,N_5303,N_4655);
or U6270 (N_6270,N_5629,N_4977);
and U6271 (N_6271,N_5168,N_5497);
and U6272 (N_6272,N_5724,N_5654);
and U6273 (N_6273,N_5640,N_4754);
nand U6274 (N_6274,N_5682,N_5781);
nor U6275 (N_6275,N_5260,N_5277);
xor U6276 (N_6276,N_5609,N_5236);
and U6277 (N_6277,N_5430,N_5101);
or U6278 (N_6278,N_5916,N_5836);
or U6279 (N_6279,N_5673,N_5932);
or U6280 (N_6280,N_4651,N_4889);
xnor U6281 (N_6281,N_5572,N_4523);
or U6282 (N_6282,N_5951,N_5009);
nand U6283 (N_6283,N_5840,N_5088);
xor U6284 (N_6284,N_5143,N_4591);
and U6285 (N_6285,N_4729,N_5238);
nand U6286 (N_6286,N_5485,N_4926);
xnor U6287 (N_6287,N_4734,N_4811);
and U6288 (N_6288,N_5968,N_4516);
nor U6289 (N_6289,N_5394,N_5354);
or U6290 (N_6290,N_5159,N_4540);
xnor U6291 (N_6291,N_4945,N_5628);
nand U6292 (N_6292,N_4980,N_5051);
nand U6293 (N_6293,N_4795,N_5881);
nor U6294 (N_6294,N_5610,N_5228);
or U6295 (N_6295,N_5446,N_4978);
and U6296 (N_6296,N_5121,N_5280);
nand U6297 (N_6297,N_5834,N_5630);
nor U6298 (N_6298,N_5381,N_4745);
and U6299 (N_6299,N_5334,N_4841);
nand U6300 (N_6300,N_5410,N_5964);
or U6301 (N_6301,N_5588,N_4677);
xnor U6302 (N_6302,N_5052,N_5603);
or U6303 (N_6303,N_5517,N_5761);
nor U6304 (N_6304,N_5075,N_5111);
and U6305 (N_6305,N_5604,N_5077);
xnor U6306 (N_6306,N_5577,N_5584);
nor U6307 (N_6307,N_4504,N_4864);
xnor U6308 (N_6308,N_5477,N_4818);
nand U6309 (N_6309,N_5202,N_4588);
or U6310 (N_6310,N_5128,N_4916);
or U6311 (N_6311,N_5817,N_5966);
nand U6312 (N_6312,N_5960,N_5669);
xnor U6313 (N_6313,N_5958,N_5671);
nand U6314 (N_6314,N_5774,N_5252);
nand U6315 (N_6315,N_5794,N_4966);
and U6316 (N_6316,N_4630,N_5328);
and U6317 (N_6317,N_4510,N_4931);
and U6318 (N_6318,N_5922,N_5411);
nand U6319 (N_6319,N_5304,N_4707);
nand U6320 (N_6320,N_5602,N_5613);
nand U6321 (N_6321,N_5740,N_5165);
nor U6322 (N_6322,N_4832,N_5639);
nand U6323 (N_6323,N_5345,N_5225);
xnor U6324 (N_6324,N_4985,N_5828);
and U6325 (N_6325,N_5155,N_4981);
and U6326 (N_6326,N_5484,N_5192);
nor U6327 (N_6327,N_5076,N_5124);
xnor U6328 (N_6328,N_4762,N_4617);
xor U6329 (N_6329,N_5200,N_4952);
xor U6330 (N_6330,N_4554,N_4697);
nor U6331 (N_6331,N_4955,N_5685);
or U6332 (N_6332,N_5890,N_5413);
nor U6333 (N_6333,N_4501,N_5224);
xor U6334 (N_6334,N_4962,N_5823);
nand U6335 (N_6335,N_4836,N_5718);
and U6336 (N_6336,N_5213,N_5712);
nand U6337 (N_6337,N_5573,N_5535);
xnor U6338 (N_6338,N_5697,N_4608);
or U6339 (N_6339,N_5417,N_5033);
xor U6340 (N_6340,N_4663,N_5219);
nor U6341 (N_6341,N_5080,N_5767);
or U6342 (N_6342,N_5611,N_4904);
and U6343 (N_6343,N_5191,N_5453);
or U6344 (N_6344,N_5465,N_5083);
nand U6345 (N_6345,N_5199,N_4609);
xnor U6346 (N_6346,N_5974,N_5005);
or U6347 (N_6347,N_5151,N_4724);
nand U6348 (N_6348,N_4672,N_5564);
xor U6349 (N_6349,N_4863,N_4918);
nor U6350 (N_6350,N_5419,N_4551);
and U6351 (N_6351,N_5743,N_5515);
or U6352 (N_6352,N_5704,N_5976);
nand U6353 (N_6353,N_5647,N_5100);
nor U6354 (N_6354,N_5551,N_5583);
or U6355 (N_6355,N_4834,N_5062);
nor U6356 (N_6356,N_5197,N_5013);
nand U6357 (N_6357,N_5154,N_4871);
nand U6358 (N_6358,N_5265,N_4885);
nand U6359 (N_6359,N_5468,N_5635);
xnor U6360 (N_6360,N_5166,N_5908);
or U6361 (N_6361,N_4753,N_5931);
nor U6362 (N_6362,N_5896,N_4870);
and U6363 (N_6363,N_4575,N_4637);
nor U6364 (N_6364,N_4752,N_5729);
nor U6365 (N_6365,N_5011,N_4535);
nand U6366 (N_6366,N_5241,N_5820);
and U6367 (N_6367,N_5302,N_4840);
xor U6368 (N_6368,N_5474,N_5689);
or U6369 (N_6369,N_5811,N_5012);
or U6370 (N_6370,N_4822,N_5784);
or U6371 (N_6371,N_5714,N_5081);
nand U6372 (N_6372,N_5841,N_4578);
or U6373 (N_6373,N_4987,N_4988);
xnor U6374 (N_6374,N_5869,N_5984);
or U6375 (N_6375,N_5755,N_5956);
and U6376 (N_6376,N_5670,N_4761);
or U6377 (N_6377,N_4896,N_5668);
and U6378 (N_6378,N_4530,N_5032);
nor U6379 (N_6379,N_5481,N_5803);
nor U6380 (N_6380,N_4709,N_5749);
xor U6381 (N_6381,N_5733,N_5575);
xnor U6382 (N_6382,N_5434,N_5899);
or U6383 (N_6383,N_5439,N_5261);
or U6384 (N_6384,N_5695,N_4648);
nor U6385 (N_6385,N_5416,N_4780);
and U6386 (N_6386,N_5442,N_4848);
or U6387 (N_6387,N_5099,N_5015);
or U6388 (N_6388,N_4851,N_5940);
nand U6389 (N_6389,N_5934,N_4593);
nand U6390 (N_6390,N_4756,N_5660);
nand U6391 (N_6391,N_5469,N_5486);
nor U6392 (N_6392,N_4865,N_5295);
and U6393 (N_6393,N_5136,N_5533);
or U6394 (N_6394,N_5991,N_5395);
nor U6395 (N_6395,N_5570,N_5292);
nand U6396 (N_6396,N_4562,N_4943);
xor U6397 (N_6397,N_5526,N_5631);
nand U6398 (N_6398,N_4536,N_5607);
nand U6399 (N_6399,N_5698,N_5893);
xor U6400 (N_6400,N_5097,N_4748);
nor U6401 (N_6401,N_4664,N_5221);
nor U6402 (N_6402,N_5980,N_5694);
nor U6403 (N_6403,N_5296,N_5091);
nand U6404 (N_6404,N_4695,N_4547);
nand U6405 (N_6405,N_5636,N_4855);
nand U6406 (N_6406,N_5278,N_4680);
and U6407 (N_6407,N_5532,N_5247);
nor U6408 (N_6408,N_5978,N_5962);
nor U6409 (N_6409,N_4511,N_4558);
xnor U6410 (N_6410,N_4899,N_5994);
nor U6411 (N_6411,N_4550,N_5367);
nand U6412 (N_6412,N_4601,N_5331);
and U6413 (N_6413,N_5970,N_4626);
xor U6414 (N_6414,N_5374,N_5240);
nand U6415 (N_6415,N_5145,N_4806);
xnor U6416 (N_6416,N_5480,N_5579);
or U6417 (N_6417,N_5999,N_5773);
nor U6418 (N_6418,N_4571,N_5479);
or U6419 (N_6419,N_4887,N_4721);
nand U6420 (N_6420,N_4725,N_5418);
xnor U6421 (N_6421,N_5891,N_5321);
nand U6422 (N_6422,N_5641,N_5692);
and U6423 (N_6423,N_5271,N_5435);
nand U6424 (N_6424,N_5263,N_4692);
and U6425 (N_6425,N_5593,N_5809);
xor U6426 (N_6426,N_5335,N_5625);
nand U6427 (N_6427,N_5525,N_5294);
nand U6428 (N_6428,N_4814,N_4660);
xnor U6429 (N_6429,N_4673,N_5193);
or U6430 (N_6430,N_5399,N_5370);
xor U6431 (N_6431,N_4992,N_5843);
or U6432 (N_6432,N_4674,N_4802);
or U6433 (N_6433,N_5786,N_5522);
nor U6434 (N_6434,N_5805,N_4526);
and U6435 (N_6435,N_4556,N_4574);
xor U6436 (N_6436,N_5427,N_5788);
nor U6437 (N_6437,N_5029,N_5944);
and U6438 (N_6438,N_5880,N_4681);
nand U6439 (N_6439,N_5126,N_4813);
and U6440 (N_6440,N_5519,N_4606);
and U6441 (N_6441,N_5177,N_4909);
nand U6442 (N_6442,N_5681,N_5585);
nand U6443 (N_6443,N_4781,N_5883);
and U6444 (N_6444,N_4741,N_4508);
xnor U6445 (N_6445,N_5987,N_4770);
nand U6446 (N_6446,N_5732,N_4768);
or U6447 (N_6447,N_5204,N_4569);
nand U6448 (N_6448,N_5715,N_5915);
or U6449 (N_6449,N_4965,N_4604);
nand U6450 (N_6450,N_5451,N_5826);
or U6451 (N_6451,N_5030,N_4599);
or U6452 (N_6452,N_5211,N_4577);
or U6453 (N_6453,N_4845,N_5130);
nor U6454 (N_6454,N_5023,N_4699);
and U6455 (N_6455,N_4774,N_4990);
nor U6456 (N_6456,N_5109,N_4895);
xor U6457 (N_6457,N_5818,N_5752);
nor U6458 (N_6458,N_4830,N_4961);
nor U6459 (N_6459,N_5850,N_5734);
nand U6460 (N_6460,N_5457,N_4808);
or U6461 (N_6461,N_5147,N_5117);
xnor U6462 (N_6462,N_5831,N_4877);
and U6463 (N_6463,N_4621,N_5104);
nand U6464 (N_6464,N_5766,N_4925);
or U6465 (N_6465,N_5201,N_4866);
nor U6466 (N_6466,N_5927,N_5520);
xor U6467 (N_6467,N_5882,N_4629);
or U6468 (N_6468,N_4623,N_4854);
xnor U6469 (N_6469,N_4502,N_5686);
and U6470 (N_6470,N_5040,N_4963);
and U6471 (N_6471,N_5144,N_4750);
nand U6472 (N_6472,N_5372,N_4846);
xnor U6473 (N_6473,N_5022,N_5765);
and U6474 (N_6474,N_5676,N_4716);
nor U6475 (N_6475,N_5760,N_5343);
nand U6476 (N_6476,N_5150,N_5039);
nand U6477 (N_6477,N_4821,N_4646);
and U6478 (N_6478,N_5194,N_4639);
xor U6479 (N_6479,N_5648,N_5311);
nor U6480 (N_6480,N_5470,N_4986);
nand U6481 (N_6481,N_5371,N_4597);
nand U6482 (N_6482,N_4520,N_4727);
xor U6483 (N_6483,N_4732,N_5878);
xnor U6484 (N_6484,N_5645,N_4687);
nor U6485 (N_6485,N_5907,N_4603);
xnor U6486 (N_6486,N_5089,N_4940);
nor U6487 (N_6487,N_5939,N_5056);
nand U6488 (N_6488,N_4957,N_4738);
nor U6489 (N_6489,N_5182,N_5720);
nand U6490 (N_6490,N_4833,N_5560);
xor U6491 (N_6491,N_5459,N_4778);
nor U6492 (N_6492,N_5623,N_4779);
and U6493 (N_6493,N_5020,N_5556);
nor U6494 (N_6494,N_5830,N_5586);
and U6495 (N_6495,N_4996,N_5888);
nand U6496 (N_6496,N_5403,N_5529);
nand U6497 (N_6497,N_5601,N_4737);
nor U6498 (N_6498,N_5674,N_5025);
or U6499 (N_6499,N_5928,N_5633);
and U6500 (N_6500,N_4936,N_5391);
and U6501 (N_6501,N_4857,N_4602);
nand U6502 (N_6502,N_5895,N_5387);
xor U6503 (N_6503,N_4524,N_5545);
nor U6504 (N_6504,N_5799,N_4703);
nor U6505 (N_6505,N_4684,N_4880);
xnor U6506 (N_6506,N_5133,N_5414);
nand U6507 (N_6507,N_4701,N_4941);
xnor U6508 (N_6508,N_4532,N_5898);
nand U6509 (N_6509,N_5282,N_5235);
nor U6510 (N_6510,N_5421,N_5161);
nand U6511 (N_6511,N_5894,N_5301);
nor U6512 (N_6512,N_5060,N_5087);
xnor U6513 (N_6513,N_4824,N_5716);
or U6514 (N_6514,N_5702,N_4760);
xnor U6515 (N_6515,N_4542,N_4867);
xnor U6516 (N_6516,N_5808,N_5384);
nand U6517 (N_6517,N_5358,N_4584);
xnor U6518 (N_6518,N_5472,N_5785);
or U6519 (N_6519,N_4545,N_5806);
and U6520 (N_6520,N_5246,N_5776);
xnor U6521 (N_6521,N_5169,N_4771);
nor U6522 (N_6522,N_5699,N_4890);
nor U6523 (N_6523,N_5995,N_4679);
or U6524 (N_6524,N_4888,N_5490);
and U6525 (N_6525,N_4968,N_4786);
nand U6526 (N_6526,N_5578,N_4964);
nand U6527 (N_6527,N_5615,N_5256);
nand U6528 (N_6528,N_4860,N_5317);
xnor U6529 (N_6529,N_5748,N_4874);
xnor U6530 (N_6530,N_4521,N_5691);
nand U6531 (N_6531,N_5307,N_5597);
and U6532 (N_6532,N_5424,N_5621);
or U6533 (N_6533,N_5149,N_5792);
xnor U6534 (N_6534,N_4906,N_5954);
nor U6535 (N_6535,N_5909,N_4580);
nor U6536 (N_6536,N_5325,N_5779);
and U6537 (N_6537,N_5746,N_5276);
nor U6538 (N_6538,N_4930,N_5382);
or U6539 (N_6539,N_5338,N_5406);
nand U6540 (N_6540,N_4767,N_5036);
nor U6541 (N_6541,N_4573,N_5364);
nand U6542 (N_6542,N_5008,N_5731);
xor U6543 (N_6543,N_4650,N_5705);
or U6544 (N_6544,N_4949,N_5658);
nand U6545 (N_6545,N_5738,N_5389);
nor U6546 (N_6546,N_4649,N_5337);
xor U6547 (N_6547,N_4656,N_4531);
xor U6548 (N_6548,N_5736,N_5363);
and U6549 (N_6549,N_5662,N_4826);
xnor U6550 (N_6550,N_5139,N_5829);
and U6551 (N_6551,N_5678,N_5385);
nand U6552 (N_6552,N_5790,N_5283);
or U6553 (N_6553,N_5254,N_5549);
and U6554 (N_6554,N_5990,N_5270);
or U6555 (N_6555,N_5963,N_5179);
nand U6556 (N_6556,N_4625,N_5571);
nor U6557 (N_6557,N_4820,N_5865);
or U6558 (N_6558,N_5667,N_5770);
xnor U6559 (N_6559,N_4548,N_5938);
xnor U6560 (N_6560,N_5595,N_5813);
and U6561 (N_6561,N_5259,N_5626);
nor U6562 (N_6562,N_4505,N_5351);
and U6563 (N_6563,N_5861,N_5069);
nand U6564 (N_6564,N_4789,N_5456);
nand U6565 (N_6565,N_5617,N_4632);
xor U6566 (N_6566,N_4712,N_4518);
nor U6567 (N_6567,N_4541,N_4717);
nor U6568 (N_6568,N_5007,N_5489);
nand U6569 (N_6569,N_5050,N_5606);
xor U6570 (N_6570,N_4515,N_5693);
xnor U6571 (N_6571,N_5955,N_5190);
and U6572 (N_6572,N_5010,N_5544);
nand U6573 (N_6573,N_5750,N_4715);
and U6574 (N_6574,N_5646,N_4657);
xnor U6575 (N_6575,N_5365,N_4519);
and U6576 (N_6576,N_5362,N_5300);
xnor U6577 (N_6577,N_5131,N_4764);
nor U6578 (N_6578,N_5082,N_5035);
and U6579 (N_6579,N_5920,N_5562);
or U6580 (N_6580,N_4722,N_5864);
or U6581 (N_6581,N_4816,N_4923);
and U6582 (N_6582,N_5120,N_5501);
or U6583 (N_6583,N_4979,N_5506);
nand U6584 (N_6584,N_4935,N_5949);
nand U6585 (N_6585,N_5643,N_5127);
nand U6586 (N_6586,N_5775,N_4624);
or U6587 (N_6587,N_5462,N_4708);
nor U6588 (N_6588,N_4900,N_5463);
or U6589 (N_6589,N_4743,N_4668);
nor U6590 (N_6590,N_5306,N_5058);
nor U6591 (N_6591,N_5113,N_5918);
nor U6592 (N_6592,N_4533,N_5444);
nand U6593 (N_6593,N_5482,N_4572);
xor U6594 (N_6594,N_4946,N_5948);
nor U6595 (N_6595,N_5493,N_5105);
and U6596 (N_6596,N_5262,N_5759);
nor U6597 (N_6597,N_4847,N_4710);
or U6598 (N_6598,N_4803,N_4587);
xnor U6599 (N_6599,N_4751,N_5142);
nand U6600 (N_6600,N_5914,N_5852);
xor U6601 (N_6601,N_4654,N_5122);
xnor U6602 (N_6602,N_5318,N_5735);
or U6603 (N_6603,N_5787,N_5244);
nor U6604 (N_6604,N_5796,N_5369);
and U6605 (N_6605,N_4666,N_5838);
xor U6606 (N_6606,N_5053,N_4561);
nand U6607 (N_6607,N_5090,N_4613);
and U6608 (N_6608,N_5887,N_4939);
or U6609 (N_6609,N_4564,N_5797);
xnor U6610 (N_6610,N_4534,N_4622);
or U6611 (N_6611,N_4731,N_5170);
xor U6612 (N_6612,N_5483,N_4901);
or U6613 (N_6613,N_4817,N_5359);
nor U6614 (N_6614,N_4686,N_5599);
xnor U6615 (N_6615,N_4705,N_5216);
xor U6616 (N_6616,N_5835,N_5102);
xnor U6617 (N_6617,N_5791,N_4787);
and U6618 (N_6618,N_5357,N_5400);
and U6619 (N_6619,N_5373,N_4905);
and U6620 (N_6620,N_4662,N_5017);
and U6621 (N_6621,N_5903,N_5308);
nor U6622 (N_6622,N_4746,N_5580);
nor U6623 (N_6623,N_4927,N_5772);
xnor U6624 (N_6624,N_5758,N_5590);
or U6625 (N_6625,N_4730,N_5764);
or U6626 (N_6626,N_5156,N_5531);
or U6627 (N_6627,N_5728,N_4513);
or U6628 (N_6628,N_5886,N_5614);
or U6629 (N_6629,N_5178,N_5782);
xor U6630 (N_6630,N_5233,N_5905);
and U6631 (N_6631,N_4594,N_5249);
and U6632 (N_6632,N_5229,N_5455);
or U6633 (N_6633,N_5730,N_4659);
and U6634 (N_6634,N_5454,N_5135);
or U6635 (N_6635,N_5253,N_4678);
nand U6636 (N_6636,N_4631,N_4563);
and U6637 (N_6637,N_5118,N_4842);
and U6638 (N_6638,N_4947,N_5727);
and U6639 (N_6639,N_4908,N_5071);
nand U6640 (N_6640,N_5188,N_5885);
nor U6641 (N_6641,N_4546,N_5471);
or U6642 (N_6642,N_5215,N_4616);
nor U6643 (N_6643,N_5862,N_5034);
nor U6644 (N_6644,N_5527,N_5950);
nand U6645 (N_6645,N_4537,N_5353);
and U6646 (N_6646,N_5027,N_5047);
nand U6647 (N_6647,N_4972,N_5164);
nor U6648 (N_6648,N_5509,N_5440);
or U6649 (N_6649,N_5795,N_5596);
and U6650 (N_6650,N_5587,N_4798);
or U6651 (N_6651,N_5491,N_4503);
nand U6652 (N_6652,N_5913,N_5004);
nand U6653 (N_6653,N_4638,N_5559);
nand U6654 (N_6654,N_5514,N_4897);
and U6655 (N_6655,N_5555,N_5355);
nand U6656 (N_6656,N_4500,N_4922);
nand U6657 (N_6657,N_5969,N_5352);
and U6658 (N_6658,N_4829,N_5026);
nand U6659 (N_6659,N_5329,N_4619);
xnor U6660 (N_6660,N_5466,N_4512);
nand U6661 (N_6661,N_5624,N_5289);
or U6662 (N_6662,N_5858,N_5874);
xor U6663 (N_6663,N_5998,N_5847);
nand U6664 (N_6664,N_4605,N_5214);
nor U6665 (N_6665,N_5789,N_5125);
or U6666 (N_6666,N_5048,N_4819);
nand U6667 (N_6667,N_5447,N_5095);
xor U6668 (N_6668,N_5425,N_4618);
nor U6669 (N_6669,N_5184,N_4862);
or U6670 (N_6670,N_5093,N_5524);
and U6671 (N_6671,N_5566,N_5967);
nand U6672 (N_6672,N_4693,N_5342);
and U6673 (N_6673,N_5106,N_5952);
or U6674 (N_6674,N_4839,N_5756);
xor U6675 (N_6675,N_5688,N_5742);
nand U6676 (N_6676,N_4529,N_5037);
nor U6677 (N_6677,N_5198,N_5245);
and U6678 (N_6678,N_4628,N_4910);
nand U6679 (N_6679,N_5726,N_5445);
nand U6680 (N_6680,N_5801,N_5160);
xor U6681 (N_6681,N_5930,N_5248);
xor U6682 (N_6682,N_4726,N_5112);
or U6683 (N_6683,N_5429,N_5094);
and U6684 (N_6684,N_5632,N_5884);
xnor U6685 (N_6685,N_4815,N_5846);
xor U6686 (N_6686,N_5901,N_5436);
nor U6687 (N_6687,N_5175,N_5879);
nor U6688 (N_6688,N_4993,N_5223);
and U6689 (N_6689,N_4581,N_5291);
xor U6690 (N_6690,N_5153,N_4589);
or U6691 (N_6691,N_5163,N_5368);
or U6692 (N_6692,N_5659,N_4796);
nand U6693 (N_6693,N_5018,N_5461);
nand U6694 (N_6694,N_5780,N_5441);
nor U6695 (N_6695,N_5747,N_4592);
and U6696 (N_6696,N_4971,N_5889);
nor U6697 (N_6697,N_4570,N_5822);
or U6698 (N_6698,N_4590,N_5550);
nand U6699 (N_6699,N_4514,N_5167);
xor U6700 (N_6700,N_4831,N_4920);
and U6701 (N_6701,N_5119,N_5935);
xnor U6702 (N_6702,N_5041,N_4642);
and U6703 (N_6703,N_4994,N_5537);
and U6704 (N_6704,N_5620,N_5855);
and U6705 (N_6705,N_5044,N_4747);
and U6706 (N_6706,N_4912,N_5554);
nor U6707 (N_6707,N_5622,N_5227);
and U6708 (N_6708,N_5478,N_4810);
and U6709 (N_6709,N_5181,N_5872);
nand U6710 (N_6710,N_5322,N_5793);
and U6711 (N_6711,N_4735,N_5652);
xor U6712 (N_6712,N_5475,N_5393);
or U6713 (N_6713,N_5114,N_5870);
and U6714 (N_6714,N_5148,N_5919);
and U6715 (N_6715,N_4835,N_5985);
xor U6716 (N_6716,N_5086,N_5528);
nor U6717 (N_6717,N_5339,N_5666);
and U6718 (N_6718,N_5024,N_4757);
nand U6719 (N_6719,N_4688,N_5180);
xor U6720 (N_6720,N_5769,N_4998);
nor U6721 (N_6721,N_5744,N_4933);
xor U6722 (N_6722,N_4921,N_5103);
xnor U6723 (N_6723,N_5054,N_4794);
and U6724 (N_6724,N_4611,N_5851);
xnor U6725 (N_6725,N_5827,N_5108);
nor U6726 (N_6726,N_5943,N_5251);
and U6727 (N_6727,N_5206,N_4579);
nor U6728 (N_6728,N_4942,N_5707);
or U6729 (N_6729,N_5460,N_5021);
nand U6730 (N_6730,N_4950,N_4670);
xnor U6731 (N_6731,N_4718,N_5946);
nor U6732 (N_6732,N_5390,N_5737);
nand U6733 (N_6733,N_4872,N_5800);
or U6734 (N_6734,N_5849,N_4755);
and U6735 (N_6735,N_5433,N_5218);
xnor U6736 (N_6736,N_5415,N_5132);
nor U6737 (N_6737,N_5798,N_5921);
nand U6738 (N_6738,N_5655,N_5684);
nor U6739 (N_6739,N_4932,N_5548);
and U6740 (N_6740,N_5423,N_4937);
or U6741 (N_6741,N_5293,N_5925);
or U6742 (N_6742,N_4506,N_5942);
or U6743 (N_6743,N_5346,N_4640);
or U6744 (N_6744,N_5768,N_5557);
nor U6745 (N_6745,N_4902,N_5812);
and U6746 (N_6746,N_5819,N_5379);
or U6747 (N_6747,N_5360,N_4882);
and U6748 (N_6748,N_5868,N_5073);
xnor U6749 (N_6749,N_5848,N_5959);
nor U6750 (N_6750,N_5884,N_5109);
nand U6751 (N_6751,N_4911,N_4524);
or U6752 (N_6752,N_4508,N_5435);
nand U6753 (N_6753,N_5560,N_5751);
nor U6754 (N_6754,N_5747,N_5794);
xor U6755 (N_6755,N_5512,N_4927);
nor U6756 (N_6756,N_5349,N_5675);
or U6757 (N_6757,N_5826,N_5590);
nand U6758 (N_6758,N_5231,N_4720);
or U6759 (N_6759,N_4891,N_5766);
nand U6760 (N_6760,N_5220,N_5052);
or U6761 (N_6761,N_4794,N_5752);
or U6762 (N_6762,N_5999,N_5755);
nand U6763 (N_6763,N_5852,N_5959);
xor U6764 (N_6764,N_4977,N_4779);
xnor U6765 (N_6765,N_5233,N_5012);
or U6766 (N_6766,N_5065,N_5369);
nor U6767 (N_6767,N_4506,N_4994);
and U6768 (N_6768,N_5957,N_5162);
nand U6769 (N_6769,N_5612,N_4614);
and U6770 (N_6770,N_5071,N_4553);
nand U6771 (N_6771,N_5318,N_4922);
and U6772 (N_6772,N_5590,N_5550);
nor U6773 (N_6773,N_4715,N_5197);
nand U6774 (N_6774,N_5336,N_5509);
nand U6775 (N_6775,N_5991,N_5110);
and U6776 (N_6776,N_5373,N_5832);
nand U6777 (N_6777,N_5687,N_5679);
nand U6778 (N_6778,N_4982,N_5819);
nand U6779 (N_6779,N_5349,N_4909);
nor U6780 (N_6780,N_5386,N_5481);
xnor U6781 (N_6781,N_5125,N_4648);
and U6782 (N_6782,N_5195,N_5180);
xnor U6783 (N_6783,N_5732,N_5020);
xor U6784 (N_6784,N_5014,N_5139);
nand U6785 (N_6785,N_5932,N_4792);
nand U6786 (N_6786,N_5016,N_5389);
nor U6787 (N_6787,N_5975,N_5586);
xnor U6788 (N_6788,N_5153,N_5519);
and U6789 (N_6789,N_4621,N_4960);
nor U6790 (N_6790,N_5219,N_4588);
or U6791 (N_6791,N_5228,N_5904);
or U6792 (N_6792,N_5242,N_5920);
or U6793 (N_6793,N_4662,N_5758);
nor U6794 (N_6794,N_5550,N_4578);
nor U6795 (N_6795,N_4607,N_5780);
nand U6796 (N_6796,N_4714,N_5572);
or U6797 (N_6797,N_5481,N_4877);
nor U6798 (N_6798,N_5485,N_4880);
nor U6799 (N_6799,N_5699,N_4566);
or U6800 (N_6800,N_4717,N_5963);
nor U6801 (N_6801,N_5296,N_5904);
nand U6802 (N_6802,N_4977,N_5589);
nand U6803 (N_6803,N_4677,N_5230);
xnor U6804 (N_6804,N_5671,N_5744);
or U6805 (N_6805,N_5129,N_4830);
nor U6806 (N_6806,N_5008,N_4749);
nor U6807 (N_6807,N_4828,N_5258);
nor U6808 (N_6808,N_4757,N_5893);
nand U6809 (N_6809,N_5268,N_4927);
xnor U6810 (N_6810,N_4790,N_4506);
xnor U6811 (N_6811,N_5193,N_4782);
and U6812 (N_6812,N_4910,N_4529);
nand U6813 (N_6813,N_4650,N_4627);
or U6814 (N_6814,N_5661,N_5734);
or U6815 (N_6815,N_5975,N_4556);
nor U6816 (N_6816,N_4605,N_5477);
or U6817 (N_6817,N_4805,N_5352);
or U6818 (N_6818,N_4936,N_5158);
nor U6819 (N_6819,N_5642,N_5880);
and U6820 (N_6820,N_4981,N_5488);
xnor U6821 (N_6821,N_5281,N_5975);
xnor U6822 (N_6822,N_5763,N_5235);
nor U6823 (N_6823,N_5290,N_5861);
nor U6824 (N_6824,N_4715,N_5211);
xor U6825 (N_6825,N_5466,N_5027);
xor U6826 (N_6826,N_4939,N_5570);
xor U6827 (N_6827,N_5291,N_5477);
xor U6828 (N_6828,N_5032,N_5747);
and U6829 (N_6829,N_4968,N_5762);
nand U6830 (N_6830,N_4829,N_4572);
or U6831 (N_6831,N_4983,N_5484);
nor U6832 (N_6832,N_5736,N_5575);
or U6833 (N_6833,N_5182,N_5253);
and U6834 (N_6834,N_5410,N_5263);
or U6835 (N_6835,N_5028,N_5079);
nor U6836 (N_6836,N_5624,N_5098);
nor U6837 (N_6837,N_5445,N_5759);
and U6838 (N_6838,N_5832,N_5238);
nor U6839 (N_6839,N_4676,N_5680);
nor U6840 (N_6840,N_4618,N_5365);
nor U6841 (N_6841,N_5721,N_4564);
or U6842 (N_6842,N_4615,N_5229);
xor U6843 (N_6843,N_5375,N_4579);
xor U6844 (N_6844,N_5002,N_4549);
or U6845 (N_6845,N_4915,N_5937);
xor U6846 (N_6846,N_5461,N_4889);
or U6847 (N_6847,N_5664,N_5530);
nand U6848 (N_6848,N_4576,N_5112);
and U6849 (N_6849,N_5878,N_5209);
and U6850 (N_6850,N_4852,N_5735);
or U6851 (N_6851,N_4538,N_4888);
nand U6852 (N_6852,N_4751,N_4806);
nor U6853 (N_6853,N_4530,N_5429);
xor U6854 (N_6854,N_5862,N_5040);
xor U6855 (N_6855,N_5449,N_5802);
nor U6856 (N_6856,N_5335,N_4981);
nor U6857 (N_6857,N_5057,N_5602);
nand U6858 (N_6858,N_4773,N_5180);
nor U6859 (N_6859,N_5526,N_4864);
or U6860 (N_6860,N_5305,N_5108);
or U6861 (N_6861,N_5340,N_4966);
or U6862 (N_6862,N_5500,N_5728);
or U6863 (N_6863,N_5875,N_4565);
nand U6864 (N_6864,N_5556,N_5960);
nor U6865 (N_6865,N_5424,N_4998);
xor U6866 (N_6866,N_4946,N_4681);
nand U6867 (N_6867,N_5485,N_4849);
nand U6868 (N_6868,N_5183,N_4886);
and U6869 (N_6869,N_5931,N_5763);
nand U6870 (N_6870,N_5858,N_5123);
and U6871 (N_6871,N_5325,N_5410);
or U6872 (N_6872,N_4584,N_4797);
and U6873 (N_6873,N_5155,N_5195);
nand U6874 (N_6874,N_5086,N_5278);
nand U6875 (N_6875,N_4893,N_5915);
nor U6876 (N_6876,N_5172,N_4818);
and U6877 (N_6877,N_4697,N_5670);
nor U6878 (N_6878,N_5947,N_5409);
xor U6879 (N_6879,N_5428,N_4831);
and U6880 (N_6880,N_5625,N_5951);
xnor U6881 (N_6881,N_5820,N_5662);
or U6882 (N_6882,N_4952,N_5183);
nand U6883 (N_6883,N_5222,N_4725);
nor U6884 (N_6884,N_5466,N_5594);
nand U6885 (N_6885,N_5143,N_4903);
xor U6886 (N_6886,N_4734,N_5965);
and U6887 (N_6887,N_5435,N_4797);
xnor U6888 (N_6888,N_5082,N_4742);
xnor U6889 (N_6889,N_4979,N_5869);
nand U6890 (N_6890,N_4646,N_5401);
or U6891 (N_6891,N_5961,N_4560);
and U6892 (N_6892,N_5789,N_5237);
xor U6893 (N_6893,N_5801,N_4834);
nand U6894 (N_6894,N_5779,N_4847);
nand U6895 (N_6895,N_5266,N_4955);
nand U6896 (N_6896,N_4627,N_4969);
nand U6897 (N_6897,N_5940,N_5247);
or U6898 (N_6898,N_5108,N_5360);
or U6899 (N_6899,N_5631,N_5350);
or U6900 (N_6900,N_5556,N_5964);
nand U6901 (N_6901,N_4614,N_5105);
and U6902 (N_6902,N_5247,N_4766);
nor U6903 (N_6903,N_5432,N_5880);
xor U6904 (N_6904,N_5098,N_5401);
nor U6905 (N_6905,N_5334,N_5084);
or U6906 (N_6906,N_5618,N_4759);
and U6907 (N_6907,N_5352,N_4501);
nor U6908 (N_6908,N_5291,N_5234);
and U6909 (N_6909,N_5607,N_5338);
xor U6910 (N_6910,N_5976,N_5310);
nand U6911 (N_6911,N_5812,N_5212);
nand U6912 (N_6912,N_5359,N_4930);
nor U6913 (N_6913,N_5245,N_5634);
nor U6914 (N_6914,N_5687,N_5916);
nand U6915 (N_6915,N_4906,N_4900);
or U6916 (N_6916,N_4705,N_4924);
and U6917 (N_6917,N_5696,N_5219);
and U6918 (N_6918,N_5982,N_4917);
nand U6919 (N_6919,N_5624,N_5018);
nor U6920 (N_6920,N_5272,N_5737);
or U6921 (N_6921,N_4742,N_4572);
or U6922 (N_6922,N_4898,N_5783);
and U6923 (N_6923,N_4652,N_5150);
nor U6924 (N_6924,N_5484,N_4840);
nor U6925 (N_6925,N_5232,N_5260);
nand U6926 (N_6926,N_4911,N_5073);
xor U6927 (N_6927,N_4731,N_4870);
and U6928 (N_6928,N_4771,N_5302);
or U6929 (N_6929,N_4749,N_4786);
nand U6930 (N_6930,N_5775,N_4573);
xnor U6931 (N_6931,N_5638,N_5536);
and U6932 (N_6932,N_5110,N_5061);
nand U6933 (N_6933,N_5067,N_5171);
xnor U6934 (N_6934,N_5108,N_4805);
nor U6935 (N_6935,N_5332,N_4917);
nand U6936 (N_6936,N_5989,N_5674);
xnor U6937 (N_6937,N_5591,N_4915);
and U6938 (N_6938,N_4654,N_5453);
xor U6939 (N_6939,N_4643,N_5289);
nor U6940 (N_6940,N_5620,N_5038);
nor U6941 (N_6941,N_5655,N_5208);
nand U6942 (N_6942,N_5531,N_5239);
nand U6943 (N_6943,N_4697,N_5807);
xnor U6944 (N_6944,N_4704,N_5708);
nor U6945 (N_6945,N_4815,N_5943);
nor U6946 (N_6946,N_5583,N_4873);
and U6947 (N_6947,N_5657,N_5684);
and U6948 (N_6948,N_5839,N_5069);
xnor U6949 (N_6949,N_4705,N_5929);
or U6950 (N_6950,N_4571,N_5865);
nand U6951 (N_6951,N_4805,N_4692);
xnor U6952 (N_6952,N_5232,N_4927);
xnor U6953 (N_6953,N_5385,N_4508);
xnor U6954 (N_6954,N_5438,N_5229);
xnor U6955 (N_6955,N_5891,N_5407);
and U6956 (N_6956,N_4555,N_4685);
nor U6957 (N_6957,N_5390,N_5336);
xnor U6958 (N_6958,N_5997,N_5832);
nand U6959 (N_6959,N_5582,N_5560);
or U6960 (N_6960,N_5544,N_5258);
nor U6961 (N_6961,N_5000,N_5266);
nor U6962 (N_6962,N_5439,N_5676);
nor U6963 (N_6963,N_5751,N_4969);
nand U6964 (N_6964,N_4879,N_5558);
or U6965 (N_6965,N_4729,N_5944);
xnor U6966 (N_6966,N_5620,N_5199);
or U6967 (N_6967,N_5593,N_5352);
or U6968 (N_6968,N_5027,N_4689);
nor U6969 (N_6969,N_4856,N_5505);
or U6970 (N_6970,N_5633,N_5939);
and U6971 (N_6971,N_5730,N_5020);
or U6972 (N_6972,N_5482,N_4853);
xnor U6973 (N_6973,N_5975,N_5998);
nor U6974 (N_6974,N_5408,N_4864);
and U6975 (N_6975,N_5239,N_5342);
xor U6976 (N_6976,N_4597,N_4956);
and U6977 (N_6977,N_4771,N_5410);
nor U6978 (N_6978,N_5075,N_5663);
and U6979 (N_6979,N_4756,N_5465);
or U6980 (N_6980,N_5146,N_5851);
nor U6981 (N_6981,N_5497,N_5592);
nand U6982 (N_6982,N_5532,N_5733);
xnor U6983 (N_6983,N_4840,N_4510);
nor U6984 (N_6984,N_4805,N_5549);
nand U6985 (N_6985,N_5735,N_5586);
or U6986 (N_6986,N_5570,N_5468);
and U6987 (N_6987,N_4580,N_5441);
nand U6988 (N_6988,N_5943,N_5176);
nor U6989 (N_6989,N_5647,N_5406);
xor U6990 (N_6990,N_5989,N_5285);
nand U6991 (N_6991,N_4780,N_4635);
nor U6992 (N_6992,N_5648,N_4694);
and U6993 (N_6993,N_5081,N_5367);
xor U6994 (N_6994,N_5892,N_4550);
xnor U6995 (N_6995,N_4958,N_4741);
and U6996 (N_6996,N_5160,N_4963);
or U6997 (N_6997,N_4588,N_5632);
or U6998 (N_6998,N_4620,N_5316);
nand U6999 (N_6999,N_4991,N_5158);
nor U7000 (N_7000,N_4863,N_5184);
and U7001 (N_7001,N_5652,N_5125);
xnor U7002 (N_7002,N_5096,N_5327);
and U7003 (N_7003,N_5110,N_4749);
xor U7004 (N_7004,N_4617,N_5014);
nand U7005 (N_7005,N_5879,N_5680);
or U7006 (N_7006,N_5016,N_4874);
nand U7007 (N_7007,N_4555,N_5428);
or U7008 (N_7008,N_4603,N_5526);
or U7009 (N_7009,N_5563,N_5899);
or U7010 (N_7010,N_5672,N_5742);
nand U7011 (N_7011,N_4544,N_4702);
nand U7012 (N_7012,N_5043,N_4849);
xor U7013 (N_7013,N_4983,N_5223);
xnor U7014 (N_7014,N_4550,N_4832);
nand U7015 (N_7015,N_5793,N_4634);
and U7016 (N_7016,N_5271,N_4666);
xor U7017 (N_7017,N_5844,N_5496);
and U7018 (N_7018,N_5549,N_4520);
xnor U7019 (N_7019,N_5123,N_5570);
nand U7020 (N_7020,N_5997,N_4778);
and U7021 (N_7021,N_4923,N_5442);
xor U7022 (N_7022,N_5602,N_4506);
or U7023 (N_7023,N_4662,N_4781);
or U7024 (N_7024,N_5909,N_5182);
nor U7025 (N_7025,N_4583,N_5617);
and U7026 (N_7026,N_5610,N_5473);
xnor U7027 (N_7027,N_5115,N_4835);
nor U7028 (N_7028,N_4624,N_5539);
or U7029 (N_7029,N_5412,N_5397);
and U7030 (N_7030,N_5214,N_5552);
and U7031 (N_7031,N_5041,N_5190);
or U7032 (N_7032,N_5241,N_4953);
and U7033 (N_7033,N_4752,N_5176);
nand U7034 (N_7034,N_5526,N_4940);
or U7035 (N_7035,N_5014,N_5082);
or U7036 (N_7036,N_5932,N_5317);
and U7037 (N_7037,N_5123,N_5697);
and U7038 (N_7038,N_5347,N_5539);
or U7039 (N_7039,N_5461,N_5161);
or U7040 (N_7040,N_5840,N_4930);
and U7041 (N_7041,N_5555,N_5654);
or U7042 (N_7042,N_5351,N_5525);
nand U7043 (N_7043,N_5400,N_4755);
nor U7044 (N_7044,N_5628,N_5153);
nand U7045 (N_7045,N_5757,N_5181);
nor U7046 (N_7046,N_5950,N_5326);
or U7047 (N_7047,N_5936,N_5144);
nand U7048 (N_7048,N_5922,N_5654);
nand U7049 (N_7049,N_4565,N_4608);
and U7050 (N_7050,N_5860,N_5941);
and U7051 (N_7051,N_4521,N_5226);
nand U7052 (N_7052,N_5246,N_4596);
and U7053 (N_7053,N_5064,N_5520);
and U7054 (N_7054,N_5021,N_4626);
nand U7055 (N_7055,N_4503,N_5879);
and U7056 (N_7056,N_4740,N_4811);
xnor U7057 (N_7057,N_5691,N_5013);
and U7058 (N_7058,N_5243,N_5648);
or U7059 (N_7059,N_5373,N_5740);
xor U7060 (N_7060,N_5498,N_4828);
xor U7061 (N_7061,N_5416,N_4943);
or U7062 (N_7062,N_5768,N_4997);
nand U7063 (N_7063,N_4739,N_5889);
or U7064 (N_7064,N_4502,N_5270);
nand U7065 (N_7065,N_5584,N_5407);
xor U7066 (N_7066,N_5269,N_5673);
nor U7067 (N_7067,N_4774,N_5985);
and U7068 (N_7068,N_5115,N_4913);
and U7069 (N_7069,N_5252,N_5265);
xnor U7070 (N_7070,N_5753,N_4537);
xnor U7071 (N_7071,N_5118,N_5514);
xor U7072 (N_7072,N_5364,N_5652);
xnor U7073 (N_7073,N_5657,N_4774);
and U7074 (N_7074,N_5675,N_5196);
and U7075 (N_7075,N_4873,N_4807);
nand U7076 (N_7076,N_4903,N_5876);
nand U7077 (N_7077,N_4904,N_4556);
or U7078 (N_7078,N_5239,N_5650);
or U7079 (N_7079,N_4871,N_4971);
and U7080 (N_7080,N_4743,N_5164);
nor U7081 (N_7081,N_5837,N_4647);
nand U7082 (N_7082,N_5489,N_5590);
or U7083 (N_7083,N_5569,N_5020);
nor U7084 (N_7084,N_5124,N_5680);
or U7085 (N_7085,N_4678,N_5341);
nand U7086 (N_7086,N_5674,N_4710);
nand U7087 (N_7087,N_5378,N_4606);
and U7088 (N_7088,N_4688,N_4842);
and U7089 (N_7089,N_5633,N_5934);
nor U7090 (N_7090,N_5714,N_5709);
or U7091 (N_7091,N_4532,N_5654);
xor U7092 (N_7092,N_5435,N_4968);
nand U7093 (N_7093,N_4764,N_5650);
xnor U7094 (N_7094,N_5973,N_5027);
xnor U7095 (N_7095,N_5009,N_5674);
nand U7096 (N_7096,N_4680,N_4584);
nor U7097 (N_7097,N_5546,N_5264);
and U7098 (N_7098,N_5120,N_5789);
nand U7099 (N_7099,N_5936,N_5331);
nor U7100 (N_7100,N_5274,N_5388);
xnor U7101 (N_7101,N_5134,N_5224);
or U7102 (N_7102,N_5439,N_5815);
nand U7103 (N_7103,N_5474,N_4500);
nand U7104 (N_7104,N_5640,N_5500);
or U7105 (N_7105,N_4886,N_4743);
xor U7106 (N_7106,N_5289,N_4602);
nor U7107 (N_7107,N_5842,N_5218);
and U7108 (N_7108,N_5249,N_5983);
and U7109 (N_7109,N_4910,N_5005);
nor U7110 (N_7110,N_5392,N_5141);
nor U7111 (N_7111,N_5740,N_5119);
or U7112 (N_7112,N_5592,N_4552);
xnor U7113 (N_7113,N_5085,N_5440);
nand U7114 (N_7114,N_4662,N_4674);
nand U7115 (N_7115,N_5320,N_5647);
and U7116 (N_7116,N_5578,N_5314);
and U7117 (N_7117,N_5293,N_4566);
or U7118 (N_7118,N_4599,N_4750);
xnor U7119 (N_7119,N_4775,N_4543);
xor U7120 (N_7120,N_5610,N_5160);
nor U7121 (N_7121,N_4691,N_5862);
nand U7122 (N_7122,N_5427,N_4819);
nor U7123 (N_7123,N_5322,N_4694);
xnor U7124 (N_7124,N_5009,N_5856);
and U7125 (N_7125,N_5987,N_5804);
nor U7126 (N_7126,N_4921,N_5241);
and U7127 (N_7127,N_5116,N_5415);
xor U7128 (N_7128,N_4611,N_4738);
nand U7129 (N_7129,N_5059,N_4911);
nor U7130 (N_7130,N_4872,N_5570);
nand U7131 (N_7131,N_4555,N_5989);
nor U7132 (N_7132,N_4693,N_5009);
or U7133 (N_7133,N_5804,N_5536);
nor U7134 (N_7134,N_5747,N_5290);
and U7135 (N_7135,N_4757,N_4905);
nor U7136 (N_7136,N_4637,N_4861);
nand U7137 (N_7137,N_5462,N_5558);
nand U7138 (N_7138,N_5280,N_5460);
xnor U7139 (N_7139,N_5616,N_5089);
nor U7140 (N_7140,N_5674,N_5498);
nor U7141 (N_7141,N_5437,N_5553);
and U7142 (N_7142,N_5928,N_4503);
nor U7143 (N_7143,N_5571,N_4952);
nor U7144 (N_7144,N_5253,N_5034);
xor U7145 (N_7145,N_4951,N_5493);
xor U7146 (N_7146,N_5299,N_4677);
and U7147 (N_7147,N_5755,N_4830);
xor U7148 (N_7148,N_5781,N_4861);
and U7149 (N_7149,N_5720,N_5427);
or U7150 (N_7150,N_5431,N_4897);
nand U7151 (N_7151,N_5983,N_5758);
or U7152 (N_7152,N_4698,N_5496);
or U7153 (N_7153,N_4917,N_5204);
and U7154 (N_7154,N_5804,N_5261);
nand U7155 (N_7155,N_5467,N_5864);
nor U7156 (N_7156,N_4887,N_5521);
nand U7157 (N_7157,N_5581,N_4600);
and U7158 (N_7158,N_5349,N_5465);
nand U7159 (N_7159,N_4872,N_5343);
and U7160 (N_7160,N_4989,N_5610);
and U7161 (N_7161,N_5959,N_5324);
nand U7162 (N_7162,N_5347,N_4983);
xnor U7163 (N_7163,N_4810,N_5515);
nand U7164 (N_7164,N_5752,N_5138);
and U7165 (N_7165,N_5097,N_5877);
nor U7166 (N_7166,N_5019,N_5671);
or U7167 (N_7167,N_5194,N_5784);
and U7168 (N_7168,N_5143,N_5118);
nand U7169 (N_7169,N_5771,N_4653);
nand U7170 (N_7170,N_4658,N_5276);
nor U7171 (N_7171,N_5525,N_5380);
or U7172 (N_7172,N_5067,N_5068);
nor U7173 (N_7173,N_5277,N_4696);
or U7174 (N_7174,N_4641,N_5256);
xnor U7175 (N_7175,N_4784,N_4665);
and U7176 (N_7176,N_5494,N_4539);
nand U7177 (N_7177,N_5570,N_4850);
or U7178 (N_7178,N_5598,N_5609);
nand U7179 (N_7179,N_4831,N_5483);
and U7180 (N_7180,N_4725,N_5081);
nor U7181 (N_7181,N_4955,N_5309);
and U7182 (N_7182,N_5769,N_5229);
nor U7183 (N_7183,N_4760,N_5627);
and U7184 (N_7184,N_4588,N_5655);
nor U7185 (N_7185,N_5397,N_5594);
nor U7186 (N_7186,N_5588,N_5822);
nand U7187 (N_7187,N_5096,N_4735);
xor U7188 (N_7188,N_4516,N_5425);
xnor U7189 (N_7189,N_5917,N_5539);
nor U7190 (N_7190,N_4656,N_5444);
and U7191 (N_7191,N_4557,N_4766);
nand U7192 (N_7192,N_4559,N_4587);
and U7193 (N_7193,N_4812,N_5387);
nor U7194 (N_7194,N_5924,N_5389);
xnor U7195 (N_7195,N_5325,N_4693);
xnor U7196 (N_7196,N_5468,N_5294);
xnor U7197 (N_7197,N_5607,N_5485);
and U7198 (N_7198,N_5994,N_5415);
or U7199 (N_7199,N_4804,N_4738);
or U7200 (N_7200,N_5269,N_4931);
nand U7201 (N_7201,N_4533,N_5908);
nor U7202 (N_7202,N_5664,N_5491);
nand U7203 (N_7203,N_5759,N_5087);
nand U7204 (N_7204,N_4629,N_5261);
and U7205 (N_7205,N_4907,N_4511);
xnor U7206 (N_7206,N_5919,N_5513);
nor U7207 (N_7207,N_4684,N_5762);
nand U7208 (N_7208,N_4912,N_5144);
or U7209 (N_7209,N_4582,N_5404);
and U7210 (N_7210,N_5586,N_5408);
and U7211 (N_7211,N_4599,N_4594);
nand U7212 (N_7212,N_4981,N_4611);
and U7213 (N_7213,N_5612,N_4710);
or U7214 (N_7214,N_4909,N_4789);
nor U7215 (N_7215,N_5190,N_5251);
and U7216 (N_7216,N_5901,N_5282);
or U7217 (N_7217,N_4902,N_5035);
and U7218 (N_7218,N_5182,N_5327);
and U7219 (N_7219,N_4979,N_5091);
nand U7220 (N_7220,N_4995,N_4684);
xor U7221 (N_7221,N_5646,N_5476);
xor U7222 (N_7222,N_5815,N_5656);
nand U7223 (N_7223,N_4766,N_5344);
xnor U7224 (N_7224,N_5429,N_5881);
or U7225 (N_7225,N_5452,N_5328);
nor U7226 (N_7226,N_5482,N_4540);
xnor U7227 (N_7227,N_4807,N_5922);
nand U7228 (N_7228,N_4619,N_5624);
or U7229 (N_7229,N_4759,N_5407);
or U7230 (N_7230,N_4534,N_5859);
and U7231 (N_7231,N_5789,N_5977);
nand U7232 (N_7232,N_5012,N_5516);
nor U7233 (N_7233,N_4840,N_4720);
nor U7234 (N_7234,N_5611,N_4635);
or U7235 (N_7235,N_4959,N_4664);
nand U7236 (N_7236,N_4987,N_5409);
xor U7237 (N_7237,N_4630,N_4619);
nand U7238 (N_7238,N_5787,N_5109);
nand U7239 (N_7239,N_4740,N_5735);
xor U7240 (N_7240,N_5026,N_4768);
nand U7241 (N_7241,N_5555,N_5023);
nor U7242 (N_7242,N_5166,N_5773);
nor U7243 (N_7243,N_5175,N_5012);
nor U7244 (N_7244,N_5098,N_4704);
xnor U7245 (N_7245,N_5633,N_5834);
nand U7246 (N_7246,N_4554,N_4646);
xor U7247 (N_7247,N_4810,N_4835);
xor U7248 (N_7248,N_5539,N_4596);
xor U7249 (N_7249,N_5651,N_5775);
nor U7250 (N_7250,N_5665,N_5058);
and U7251 (N_7251,N_5663,N_5335);
and U7252 (N_7252,N_4897,N_5583);
nor U7253 (N_7253,N_4655,N_5402);
and U7254 (N_7254,N_5611,N_5050);
and U7255 (N_7255,N_4980,N_5989);
nor U7256 (N_7256,N_5595,N_5033);
xnor U7257 (N_7257,N_5352,N_5768);
and U7258 (N_7258,N_5488,N_5896);
nor U7259 (N_7259,N_5400,N_5811);
xor U7260 (N_7260,N_5687,N_5910);
or U7261 (N_7261,N_4976,N_5388);
nand U7262 (N_7262,N_5387,N_4898);
nand U7263 (N_7263,N_4720,N_5440);
and U7264 (N_7264,N_4696,N_5441);
or U7265 (N_7265,N_5109,N_5210);
xor U7266 (N_7266,N_4586,N_5196);
nand U7267 (N_7267,N_5027,N_5292);
nand U7268 (N_7268,N_5689,N_5139);
nand U7269 (N_7269,N_5392,N_4775);
nor U7270 (N_7270,N_5948,N_4856);
nor U7271 (N_7271,N_5148,N_4621);
and U7272 (N_7272,N_5080,N_5345);
or U7273 (N_7273,N_4978,N_4652);
or U7274 (N_7274,N_4993,N_4678);
xnor U7275 (N_7275,N_4626,N_4543);
nand U7276 (N_7276,N_5523,N_5225);
nor U7277 (N_7277,N_4523,N_4977);
and U7278 (N_7278,N_5353,N_4877);
nand U7279 (N_7279,N_4753,N_5738);
xnor U7280 (N_7280,N_5435,N_5041);
nor U7281 (N_7281,N_5736,N_5770);
or U7282 (N_7282,N_5842,N_5572);
and U7283 (N_7283,N_5127,N_4611);
xnor U7284 (N_7284,N_5503,N_4987);
nand U7285 (N_7285,N_4617,N_5260);
nor U7286 (N_7286,N_5997,N_5214);
xnor U7287 (N_7287,N_4713,N_5782);
nand U7288 (N_7288,N_4942,N_5012);
xnor U7289 (N_7289,N_5455,N_5368);
nor U7290 (N_7290,N_5184,N_5762);
nor U7291 (N_7291,N_4969,N_5188);
or U7292 (N_7292,N_5813,N_5319);
or U7293 (N_7293,N_5890,N_4538);
nor U7294 (N_7294,N_5851,N_5936);
or U7295 (N_7295,N_4711,N_5006);
xor U7296 (N_7296,N_4614,N_4611);
nand U7297 (N_7297,N_5079,N_5243);
or U7298 (N_7298,N_5276,N_5656);
nand U7299 (N_7299,N_5858,N_4505);
nor U7300 (N_7300,N_5278,N_5390);
and U7301 (N_7301,N_5860,N_5638);
xnor U7302 (N_7302,N_5399,N_5663);
nor U7303 (N_7303,N_5387,N_4623);
or U7304 (N_7304,N_4710,N_5034);
nand U7305 (N_7305,N_5410,N_5460);
and U7306 (N_7306,N_5166,N_5024);
or U7307 (N_7307,N_5558,N_5304);
xor U7308 (N_7308,N_4962,N_5573);
or U7309 (N_7309,N_5176,N_5218);
nand U7310 (N_7310,N_4612,N_5945);
nand U7311 (N_7311,N_4702,N_5944);
and U7312 (N_7312,N_5745,N_4779);
nor U7313 (N_7313,N_4568,N_4587);
nor U7314 (N_7314,N_5420,N_4922);
nand U7315 (N_7315,N_4894,N_5407);
nand U7316 (N_7316,N_5148,N_5575);
nor U7317 (N_7317,N_5986,N_5537);
xor U7318 (N_7318,N_4896,N_4570);
or U7319 (N_7319,N_5456,N_4597);
and U7320 (N_7320,N_4895,N_5507);
or U7321 (N_7321,N_5559,N_5062);
nand U7322 (N_7322,N_5349,N_5065);
nand U7323 (N_7323,N_5991,N_5284);
or U7324 (N_7324,N_4861,N_5629);
or U7325 (N_7325,N_5366,N_4881);
and U7326 (N_7326,N_5561,N_5337);
and U7327 (N_7327,N_5594,N_4806);
xnor U7328 (N_7328,N_5711,N_5414);
nor U7329 (N_7329,N_5151,N_5906);
or U7330 (N_7330,N_5867,N_4681);
nor U7331 (N_7331,N_4774,N_5062);
nand U7332 (N_7332,N_5720,N_5924);
and U7333 (N_7333,N_4867,N_5683);
and U7334 (N_7334,N_5151,N_4698);
nor U7335 (N_7335,N_5630,N_5946);
nand U7336 (N_7336,N_5923,N_4518);
nor U7337 (N_7337,N_4719,N_4922);
or U7338 (N_7338,N_5851,N_4784);
nand U7339 (N_7339,N_4516,N_5976);
nand U7340 (N_7340,N_4637,N_4857);
and U7341 (N_7341,N_5892,N_4832);
nand U7342 (N_7342,N_4788,N_5814);
nand U7343 (N_7343,N_4959,N_5678);
nand U7344 (N_7344,N_5981,N_4979);
xor U7345 (N_7345,N_5999,N_5400);
nor U7346 (N_7346,N_4917,N_5598);
nor U7347 (N_7347,N_5158,N_5636);
nand U7348 (N_7348,N_5654,N_5958);
and U7349 (N_7349,N_5085,N_4769);
and U7350 (N_7350,N_5484,N_5268);
nor U7351 (N_7351,N_5485,N_4761);
or U7352 (N_7352,N_5245,N_5515);
nor U7353 (N_7353,N_4932,N_5563);
and U7354 (N_7354,N_5240,N_5197);
nor U7355 (N_7355,N_5880,N_5418);
nor U7356 (N_7356,N_4596,N_4788);
or U7357 (N_7357,N_5293,N_5084);
and U7358 (N_7358,N_5266,N_4701);
xnor U7359 (N_7359,N_5842,N_5959);
nor U7360 (N_7360,N_5658,N_5234);
and U7361 (N_7361,N_5000,N_5565);
nand U7362 (N_7362,N_5716,N_5841);
or U7363 (N_7363,N_5815,N_4589);
or U7364 (N_7364,N_4520,N_5798);
and U7365 (N_7365,N_5149,N_5269);
nand U7366 (N_7366,N_5091,N_5268);
nand U7367 (N_7367,N_5162,N_5408);
or U7368 (N_7368,N_4593,N_5917);
xor U7369 (N_7369,N_5650,N_4504);
or U7370 (N_7370,N_4845,N_5632);
or U7371 (N_7371,N_4785,N_5123);
nor U7372 (N_7372,N_5670,N_5603);
nand U7373 (N_7373,N_5088,N_5104);
nor U7374 (N_7374,N_5059,N_4988);
nand U7375 (N_7375,N_5475,N_5598);
nand U7376 (N_7376,N_5414,N_5366);
or U7377 (N_7377,N_5485,N_5424);
or U7378 (N_7378,N_5943,N_5133);
xnor U7379 (N_7379,N_5786,N_4943);
nand U7380 (N_7380,N_5415,N_4776);
or U7381 (N_7381,N_5903,N_4608);
xnor U7382 (N_7382,N_4957,N_5179);
nor U7383 (N_7383,N_4597,N_4989);
xor U7384 (N_7384,N_4924,N_5100);
xnor U7385 (N_7385,N_5013,N_5205);
nor U7386 (N_7386,N_5349,N_5304);
and U7387 (N_7387,N_5729,N_5313);
xor U7388 (N_7388,N_5474,N_5926);
and U7389 (N_7389,N_5026,N_5104);
or U7390 (N_7390,N_4777,N_4998);
xnor U7391 (N_7391,N_5315,N_5865);
or U7392 (N_7392,N_4622,N_4903);
nor U7393 (N_7393,N_5861,N_4976);
or U7394 (N_7394,N_5206,N_5328);
or U7395 (N_7395,N_5959,N_4795);
xnor U7396 (N_7396,N_5704,N_4823);
nand U7397 (N_7397,N_5588,N_4705);
and U7398 (N_7398,N_5260,N_5508);
xnor U7399 (N_7399,N_5990,N_5959);
nor U7400 (N_7400,N_4923,N_4702);
nand U7401 (N_7401,N_5077,N_5724);
nor U7402 (N_7402,N_5481,N_5988);
and U7403 (N_7403,N_4864,N_5381);
xnor U7404 (N_7404,N_5124,N_5695);
and U7405 (N_7405,N_5949,N_4665);
nor U7406 (N_7406,N_5804,N_5113);
xnor U7407 (N_7407,N_5901,N_5969);
nand U7408 (N_7408,N_5028,N_4753);
nand U7409 (N_7409,N_5638,N_5437);
or U7410 (N_7410,N_4593,N_5014);
xnor U7411 (N_7411,N_5845,N_5063);
and U7412 (N_7412,N_4995,N_4706);
nand U7413 (N_7413,N_4645,N_5888);
nand U7414 (N_7414,N_5224,N_5714);
or U7415 (N_7415,N_5569,N_4877);
nor U7416 (N_7416,N_5263,N_4560);
nor U7417 (N_7417,N_4829,N_5087);
and U7418 (N_7418,N_5382,N_4688);
nor U7419 (N_7419,N_4998,N_5242);
xnor U7420 (N_7420,N_4986,N_5792);
nor U7421 (N_7421,N_4551,N_5229);
xnor U7422 (N_7422,N_5413,N_5369);
nor U7423 (N_7423,N_5526,N_5118);
or U7424 (N_7424,N_5835,N_5446);
or U7425 (N_7425,N_5891,N_5465);
and U7426 (N_7426,N_5024,N_4933);
xor U7427 (N_7427,N_4896,N_5604);
and U7428 (N_7428,N_4936,N_4563);
xor U7429 (N_7429,N_4600,N_5925);
nor U7430 (N_7430,N_4676,N_4827);
nand U7431 (N_7431,N_5261,N_4977);
and U7432 (N_7432,N_5020,N_5995);
or U7433 (N_7433,N_5795,N_4967);
nand U7434 (N_7434,N_4507,N_5002);
xnor U7435 (N_7435,N_4693,N_4768);
nand U7436 (N_7436,N_5440,N_5441);
nand U7437 (N_7437,N_5126,N_5309);
nand U7438 (N_7438,N_4745,N_5220);
nor U7439 (N_7439,N_4883,N_4872);
and U7440 (N_7440,N_4833,N_4790);
or U7441 (N_7441,N_4842,N_5841);
or U7442 (N_7442,N_4804,N_5717);
nand U7443 (N_7443,N_4949,N_5245);
nand U7444 (N_7444,N_5343,N_5401);
and U7445 (N_7445,N_5574,N_4774);
or U7446 (N_7446,N_5279,N_5537);
nor U7447 (N_7447,N_4721,N_5947);
nand U7448 (N_7448,N_5162,N_4749);
xor U7449 (N_7449,N_5561,N_4920);
and U7450 (N_7450,N_5147,N_4841);
nand U7451 (N_7451,N_5981,N_5662);
and U7452 (N_7452,N_5145,N_5565);
or U7453 (N_7453,N_5747,N_5774);
nand U7454 (N_7454,N_4857,N_5185);
nand U7455 (N_7455,N_5250,N_5218);
nor U7456 (N_7456,N_5634,N_4623);
nand U7457 (N_7457,N_5296,N_4562);
or U7458 (N_7458,N_4682,N_5167);
nand U7459 (N_7459,N_5858,N_5729);
and U7460 (N_7460,N_5900,N_4949);
or U7461 (N_7461,N_5715,N_5460);
xor U7462 (N_7462,N_4601,N_5861);
xor U7463 (N_7463,N_5302,N_4979);
nor U7464 (N_7464,N_5428,N_5488);
xor U7465 (N_7465,N_5162,N_5006);
xnor U7466 (N_7466,N_5035,N_5490);
or U7467 (N_7467,N_5271,N_5798);
nand U7468 (N_7468,N_4615,N_4648);
nand U7469 (N_7469,N_4530,N_5924);
xnor U7470 (N_7470,N_5234,N_5002);
and U7471 (N_7471,N_5646,N_4712);
and U7472 (N_7472,N_5470,N_5898);
or U7473 (N_7473,N_4865,N_5659);
xnor U7474 (N_7474,N_4979,N_5189);
nand U7475 (N_7475,N_4707,N_5898);
or U7476 (N_7476,N_5843,N_5858);
xnor U7477 (N_7477,N_5685,N_5234);
nor U7478 (N_7478,N_5551,N_4994);
and U7479 (N_7479,N_5268,N_5938);
nor U7480 (N_7480,N_5480,N_4856);
and U7481 (N_7481,N_5971,N_5957);
nor U7482 (N_7482,N_5448,N_4964);
or U7483 (N_7483,N_5041,N_4802);
or U7484 (N_7484,N_4931,N_4664);
nand U7485 (N_7485,N_5832,N_5694);
nand U7486 (N_7486,N_5227,N_4615);
nor U7487 (N_7487,N_5436,N_4971);
and U7488 (N_7488,N_5568,N_4700);
xnor U7489 (N_7489,N_5192,N_5890);
xnor U7490 (N_7490,N_4938,N_5756);
or U7491 (N_7491,N_4691,N_5691);
and U7492 (N_7492,N_5197,N_4709);
nor U7493 (N_7493,N_4584,N_5453);
nand U7494 (N_7494,N_5034,N_5741);
or U7495 (N_7495,N_4550,N_5683);
and U7496 (N_7496,N_4930,N_4817);
xnor U7497 (N_7497,N_4828,N_5981);
nor U7498 (N_7498,N_5598,N_4560);
nor U7499 (N_7499,N_5053,N_4870);
nand U7500 (N_7500,N_6470,N_6518);
xor U7501 (N_7501,N_6073,N_7320);
nor U7502 (N_7502,N_7329,N_7478);
nand U7503 (N_7503,N_6219,N_6671);
xnor U7504 (N_7504,N_6315,N_6521);
nand U7505 (N_7505,N_7028,N_6304);
nand U7506 (N_7506,N_6772,N_7196);
nand U7507 (N_7507,N_6114,N_6798);
xnor U7508 (N_7508,N_7236,N_6620);
and U7509 (N_7509,N_7464,N_6306);
or U7510 (N_7510,N_7050,N_7430);
nor U7511 (N_7511,N_6871,N_7053);
xor U7512 (N_7512,N_7333,N_6686);
xor U7513 (N_7513,N_7176,N_7207);
nor U7514 (N_7514,N_7446,N_6055);
nand U7515 (N_7515,N_6478,N_7204);
nor U7516 (N_7516,N_6826,N_6978);
nand U7517 (N_7517,N_6591,N_6751);
nor U7518 (N_7518,N_7387,N_6577);
nor U7519 (N_7519,N_6157,N_7194);
xor U7520 (N_7520,N_6156,N_7095);
nor U7521 (N_7521,N_6496,N_7408);
and U7522 (N_7522,N_6380,N_6763);
xor U7523 (N_7523,N_6019,N_6746);
nor U7524 (N_7524,N_6024,N_6675);
nand U7525 (N_7525,N_6598,N_6350);
nand U7526 (N_7526,N_7096,N_6292);
and U7527 (N_7527,N_7315,N_6765);
nor U7528 (N_7528,N_6587,N_7070);
nand U7529 (N_7529,N_6660,N_7288);
or U7530 (N_7530,N_7227,N_6130);
xor U7531 (N_7531,N_7193,N_6464);
xor U7532 (N_7532,N_6678,N_7347);
xnor U7533 (N_7533,N_6316,N_6648);
nor U7534 (N_7534,N_6447,N_7382);
or U7535 (N_7535,N_6721,N_7367);
or U7536 (N_7536,N_6736,N_6050);
nand U7537 (N_7537,N_6031,N_6868);
or U7538 (N_7538,N_6855,N_6810);
xnor U7539 (N_7539,N_6749,N_6442);
nor U7540 (N_7540,N_7455,N_7286);
xor U7541 (N_7541,N_7266,N_7143);
nand U7542 (N_7542,N_7060,N_6597);
nand U7543 (N_7543,N_7006,N_6594);
nand U7544 (N_7544,N_6021,N_6621);
or U7545 (N_7545,N_6828,N_7044);
or U7546 (N_7546,N_6450,N_6667);
or U7547 (N_7547,N_6367,N_7308);
and U7548 (N_7548,N_7056,N_7327);
or U7549 (N_7549,N_6610,N_6806);
nor U7550 (N_7550,N_7232,N_7156);
or U7551 (N_7551,N_7088,N_7010);
nand U7552 (N_7552,N_6825,N_7147);
nand U7553 (N_7553,N_6102,N_7319);
and U7554 (N_7554,N_6153,N_7218);
nand U7555 (N_7555,N_6802,N_6561);
or U7556 (N_7556,N_6708,N_6116);
and U7557 (N_7557,N_6491,N_6891);
xor U7558 (N_7558,N_7324,N_6331);
xnor U7559 (N_7559,N_6724,N_6979);
nor U7560 (N_7560,N_6137,N_7090);
nor U7561 (N_7561,N_6115,N_6554);
and U7562 (N_7562,N_7228,N_6109);
and U7563 (N_7563,N_6712,N_7003);
or U7564 (N_7564,N_6862,N_6307);
or U7565 (N_7565,N_6344,N_7072);
and U7566 (N_7566,N_6499,N_6459);
xnor U7567 (N_7567,N_7079,N_6340);
nor U7568 (N_7568,N_6930,N_7303);
nor U7569 (N_7569,N_6112,N_6209);
xor U7570 (N_7570,N_6096,N_7233);
and U7571 (N_7571,N_6900,N_6537);
xor U7572 (N_7572,N_6040,N_7182);
or U7573 (N_7573,N_7191,N_6075);
nor U7574 (N_7574,N_7415,N_7486);
and U7575 (N_7575,N_6392,N_7113);
nor U7576 (N_7576,N_7073,N_6984);
nor U7577 (N_7577,N_7422,N_6070);
xnor U7578 (N_7578,N_6327,N_6127);
xor U7579 (N_7579,N_6542,N_6539);
or U7580 (N_7580,N_6989,N_6831);
and U7581 (N_7581,N_6707,N_7465);
xor U7582 (N_7582,N_6757,N_6025);
nand U7583 (N_7583,N_6808,N_6544);
nand U7584 (N_7584,N_7115,N_7302);
nand U7585 (N_7585,N_6579,N_6709);
nor U7586 (N_7586,N_6287,N_7471);
and U7587 (N_7587,N_6098,N_6702);
xor U7588 (N_7588,N_6433,N_6275);
and U7589 (N_7589,N_7104,N_6827);
nor U7590 (N_7590,N_7188,N_6844);
or U7591 (N_7591,N_6221,N_7238);
nand U7592 (N_7592,N_6782,N_6217);
nor U7593 (N_7593,N_6566,N_6687);
nand U7594 (N_7594,N_6502,N_7125);
xor U7595 (N_7595,N_6030,N_6389);
nand U7596 (N_7596,N_6458,N_6343);
nand U7597 (N_7597,N_7223,N_7005);
xor U7598 (N_7598,N_6557,N_6104);
or U7599 (N_7599,N_7151,N_6005);
and U7600 (N_7600,N_6929,N_7368);
nand U7601 (N_7601,N_6940,N_7277);
or U7602 (N_7602,N_6585,N_6800);
xnor U7603 (N_7603,N_6440,N_6311);
nand U7604 (N_7604,N_6171,N_6498);
or U7605 (N_7605,N_7311,N_6997);
nor U7606 (N_7606,N_7428,N_6135);
xor U7607 (N_7607,N_6391,N_6622);
nand U7608 (N_7608,N_7325,N_6305);
or U7609 (N_7609,N_7365,N_6425);
or U7610 (N_7610,N_6887,N_7015);
or U7611 (N_7611,N_7412,N_6322);
nand U7612 (N_7612,N_6903,N_6528);
or U7613 (N_7613,N_7374,N_7246);
nor U7614 (N_7614,N_7171,N_6013);
nand U7615 (N_7615,N_6875,N_6000);
nor U7616 (N_7616,N_6511,N_6501);
nand U7617 (N_7617,N_6923,N_6959);
xnor U7618 (N_7618,N_7034,N_6247);
and U7619 (N_7619,N_6371,N_7469);
nor U7620 (N_7620,N_7127,N_6890);
or U7621 (N_7621,N_7245,N_6342);
nand U7622 (N_7622,N_6638,N_6017);
and U7623 (N_7623,N_6069,N_7230);
and U7624 (N_7624,N_7298,N_6428);
xor U7625 (N_7625,N_7110,N_6260);
nand U7626 (N_7626,N_6796,N_7040);
xnor U7627 (N_7627,N_7112,N_6928);
nand U7628 (N_7628,N_6369,N_7419);
nor U7629 (N_7629,N_7370,N_7022);
and U7630 (N_7630,N_7305,N_7149);
and U7631 (N_7631,N_6485,N_7014);
nand U7632 (N_7632,N_7401,N_6099);
xnor U7633 (N_7633,N_6215,N_6444);
and U7634 (N_7634,N_6360,N_6599);
nand U7635 (N_7635,N_6227,N_7344);
nand U7636 (N_7636,N_6792,N_6908);
nand U7637 (N_7637,N_6644,N_7091);
nor U7638 (N_7638,N_6570,N_6457);
xor U7639 (N_7639,N_7362,N_6402);
xnor U7640 (N_7640,N_6089,N_6522);
or U7641 (N_7641,N_6397,N_6092);
nor U7642 (N_7642,N_7434,N_6011);
nand U7643 (N_7643,N_7123,N_7108);
or U7644 (N_7644,N_7267,N_7065);
and U7645 (N_7645,N_6507,N_6985);
nor U7646 (N_7646,N_6142,N_6455);
or U7647 (N_7647,N_7120,N_6347);
and U7648 (N_7648,N_7394,N_6144);
nor U7649 (N_7649,N_6590,N_6572);
xnor U7650 (N_7650,N_6230,N_6679);
and U7651 (N_7651,N_6362,N_6167);
or U7652 (N_7652,N_6718,N_6971);
or U7653 (N_7653,N_6880,N_7396);
nand U7654 (N_7654,N_7421,N_6879);
nor U7655 (N_7655,N_6035,N_6285);
or U7656 (N_7656,N_6974,N_6180);
and U7657 (N_7657,N_7285,N_6778);
and U7658 (N_7658,N_7290,N_7214);
nand U7659 (N_7659,N_6841,N_6582);
nor U7660 (N_7660,N_6226,N_6558);
xor U7661 (N_7661,N_6006,N_6152);
xnor U7662 (N_7662,N_6969,N_6436);
or U7663 (N_7663,N_7129,N_6711);
xor U7664 (N_7664,N_6149,N_6487);
or U7665 (N_7665,N_7106,N_6876);
nand U7666 (N_7666,N_6179,N_7045);
nand U7667 (N_7667,N_6308,N_6493);
nand U7668 (N_7668,N_6615,N_7435);
or U7669 (N_7669,N_6239,N_6432);
xnor U7670 (N_7670,N_6633,N_6435);
xnor U7671 (N_7671,N_6690,N_6155);
nor U7672 (N_7672,N_6376,N_7411);
nand U7673 (N_7673,N_6723,N_6071);
xor U7674 (N_7674,N_7358,N_6087);
or U7675 (N_7675,N_6947,N_6834);
nor U7676 (N_7676,N_6905,N_7429);
or U7677 (N_7677,N_6856,N_7025);
or U7678 (N_7678,N_6949,N_6366);
or U7679 (N_7679,N_6650,N_7485);
nor U7680 (N_7680,N_6699,N_6188);
and U7681 (N_7681,N_6510,N_7142);
nor U7682 (N_7682,N_7332,N_7121);
and U7683 (N_7683,N_7231,N_6895);
nand U7684 (N_7684,N_7269,N_6716);
and U7685 (N_7685,N_6294,N_6132);
or U7686 (N_7686,N_7016,N_7047);
nor U7687 (N_7687,N_7424,N_6913);
nor U7688 (N_7688,N_6338,N_7161);
and U7689 (N_7689,N_7036,N_6820);
nor U7690 (N_7690,N_6634,N_7076);
or U7691 (N_7691,N_6110,N_7128);
and U7692 (N_7692,N_7211,N_6753);
or U7693 (N_7693,N_7224,N_7386);
xor U7694 (N_7694,N_7484,N_7068);
or U7695 (N_7695,N_6661,N_6174);
nand U7696 (N_7696,N_6131,N_7206);
nand U7697 (N_7697,N_7283,N_6894);
nor U7698 (N_7698,N_6560,N_6613);
and U7699 (N_7699,N_6424,N_6355);
nand U7700 (N_7700,N_6664,N_7304);
nand U7701 (N_7701,N_7071,N_7312);
or U7702 (N_7702,N_6865,N_7440);
or U7703 (N_7703,N_6606,N_7062);
and U7704 (N_7704,N_7066,N_7219);
nor U7705 (N_7705,N_7268,N_7294);
xor U7706 (N_7706,N_7351,N_6245);
xor U7707 (N_7707,N_6377,N_6731);
nand U7708 (N_7708,N_6068,N_6257);
nand U7709 (N_7709,N_6846,N_6529);
and U7710 (N_7710,N_6359,N_7019);
nor U7711 (N_7711,N_6824,N_7355);
and U7712 (N_7712,N_6805,N_6818);
xor U7713 (N_7713,N_6264,N_6133);
nor U7714 (N_7714,N_6220,N_6405);
and U7715 (N_7715,N_7474,N_6672);
and U7716 (N_7716,N_6781,N_7322);
or U7717 (N_7717,N_6483,N_7461);
nor U7718 (N_7718,N_7102,N_6431);
and U7719 (N_7719,N_6028,N_6267);
nand U7720 (N_7720,N_7049,N_6462);
or U7721 (N_7721,N_6415,N_6655);
or U7722 (N_7722,N_6953,N_7221);
nor U7723 (N_7723,N_7496,N_7338);
nor U7724 (N_7724,N_7407,N_7378);
nor U7725 (N_7725,N_6237,N_7077);
or U7726 (N_7726,N_6559,N_6309);
xnor U7727 (N_7727,N_7089,N_6379);
nor U7728 (N_7728,N_7497,N_6669);
xnor U7729 (N_7729,N_6186,N_6922);
nor U7730 (N_7730,N_6172,N_6619);
or U7731 (N_7731,N_7078,N_7349);
nor U7732 (N_7732,N_6163,N_6787);
nand U7733 (N_7733,N_6255,N_7004);
xor U7734 (N_7734,N_6169,N_6385);
nor U7735 (N_7735,N_6991,N_6295);
xor U7736 (N_7736,N_6609,N_6277);
xnor U7737 (N_7737,N_6777,N_7155);
and U7738 (N_7738,N_6337,N_7406);
nand U7739 (N_7739,N_6999,N_6745);
xor U7740 (N_7740,N_6161,N_6289);
xnor U7741 (N_7741,N_7136,N_7114);
or U7742 (N_7742,N_7109,N_6748);
xnor U7743 (N_7743,N_6595,N_6696);
and U7744 (N_7744,N_6456,N_6565);
and U7745 (N_7745,N_7449,N_7400);
and U7746 (N_7746,N_7316,N_6231);
and U7747 (N_7747,N_6784,N_6983);
nand U7748 (N_7748,N_7197,N_6244);
or U7749 (N_7749,N_7243,N_7174);
nand U7750 (N_7750,N_7392,N_7080);
or U7751 (N_7751,N_6531,N_7041);
and U7752 (N_7752,N_6236,N_7187);
and U7753 (N_7753,N_6332,N_6370);
nand U7754 (N_7754,N_7132,N_6682);
and U7755 (N_7755,N_7289,N_7472);
and U7756 (N_7756,N_6363,N_6857);
and U7757 (N_7757,N_7052,N_6232);
xor U7758 (N_7758,N_7103,N_7234);
nand U7759 (N_7759,N_7397,N_6471);
nand U7760 (N_7760,N_6318,N_7458);
or U7761 (N_7761,N_6037,N_6437);
or U7762 (N_7762,N_6395,N_6048);
xor U7763 (N_7763,N_6326,N_6270);
or U7764 (N_7764,N_6119,N_6786);
nand U7765 (N_7765,N_6832,N_6600);
nor U7766 (N_7766,N_7463,N_6282);
or U7767 (N_7767,N_7439,N_7225);
nand U7768 (N_7768,N_6388,N_6045);
and U7769 (N_7769,N_6988,N_6383);
and U7770 (N_7770,N_6258,N_6698);
xor U7771 (N_7771,N_7248,N_6898);
nand U7772 (N_7772,N_7154,N_6489);
nand U7773 (N_7773,N_7490,N_6505);
and U7774 (N_7774,N_6183,N_7021);
nand U7775 (N_7775,N_6564,N_6365);
or U7776 (N_7776,N_6271,N_6012);
xnor U7777 (N_7777,N_7354,N_6516);
nor U7778 (N_7778,N_6512,N_6417);
nand U7779 (N_7779,N_7217,N_7100);
nand U7780 (N_7780,N_6358,N_7275);
xor U7781 (N_7781,N_7001,N_6297);
xor U7782 (N_7782,N_6795,N_6568);
or U7783 (N_7783,N_7420,N_6668);
nand U7784 (N_7784,N_7337,N_7342);
and U7785 (N_7785,N_6120,N_6335);
and U7786 (N_7786,N_6995,N_6198);
nor U7787 (N_7787,N_7146,N_7033);
or U7788 (N_7788,N_6914,N_6079);
xor U7789 (N_7789,N_6381,N_7292);
and U7790 (N_7790,N_6901,N_6536);
nor U7791 (N_7791,N_6044,N_6873);
nor U7792 (N_7792,N_7410,N_7479);
nand U7793 (N_7793,N_6977,N_6461);
xnor U7794 (N_7794,N_6532,N_6162);
nand U7795 (N_7795,N_7237,N_6486);
or U7796 (N_7796,N_7488,N_7160);
xnor U7797 (N_7797,N_6843,N_6761);
and U7798 (N_7798,N_6685,N_7069);
or U7799 (N_7799,N_6181,N_6176);
nand U7800 (N_7800,N_7220,N_7350);
xor U7801 (N_7801,N_7270,N_6627);
or U7802 (N_7802,N_6815,N_6029);
xor U7803 (N_7803,N_6280,N_6813);
or U7804 (N_7804,N_7326,N_6526);
or U7805 (N_7805,N_6733,N_6259);
and U7806 (N_7806,N_7423,N_6640);
and U7807 (N_7807,N_6147,N_6549);
or U7808 (N_7808,N_7007,N_6734);
xor U7809 (N_7809,N_6830,N_6009);
xor U7810 (N_7810,N_6225,N_6302);
nand U7811 (N_7811,N_6951,N_6943);
xor U7812 (N_7812,N_7371,N_7085);
xnor U7813 (N_7813,N_7139,N_6333);
xor U7814 (N_7814,N_6146,N_6208);
xnor U7815 (N_7815,N_6543,N_6414);
or U7816 (N_7816,N_7043,N_7175);
nor U7817 (N_7817,N_6883,N_7035);
or U7818 (N_7818,N_7063,N_7272);
nor U7819 (N_7819,N_6065,N_7157);
or U7820 (N_7820,N_7150,N_7475);
or U7821 (N_7821,N_6541,N_6224);
nor U7822 (N_7822,N_6603,N_6715);
nor U7823 (N_7823,N_6480,N_7301);
xor U7824 (N_7824,N_7170,N_7495);
nor U7825 (N_7825,N_6911,N_6907);
nand U7826 (N_7826,N_6047,N_7441);
or U7827 (N_7827,N_6918,N_7278);
or U7828 (N_7828,N_7013,N_6730);
or U7829 (N_7829,N_7306,N_7293);
and U7830 (N_7830,N_6845,N_6274);
nor U7831 (N_7831,N_7317,N_6090);
nor U7832 (N_7832,N_6159,N_6720);
and U7833 (N_7833,N_6842,N_7032);
or U7834 (N_7834,N_7087,N_6368);
and U7835 (N_7835,N_6975,N_6122);
nand U7836 (N_7836,N_6004,N_6580);
xor U7837 (N_7837,N_6330,N_7168);
nor U7838 (N_7838,N_7247,N_6240);
and U7839 (N_7839,N_7281,N_6527);
and U7840 (N_7840,N_6656,N_6662);
nor U7841 (N_7841,N_6623,N_6888);
nor U7842 (N_7842,N_6631,N_7433);
nand U7843 (N_7843,N_6027,N_7482);
nor U7844 (N_7844,N_7276,N_6472);
or U7845 (N_7845,N_6921,N_6348);
nand U7846 (N_7846,N_7083,N_6321);
or U7847 (N_7847,N_7369,N_6967);
nor U7848 (N_7848,N_6628,N_7082);
and U7849 (N_7849,N_7352,N_6896);
and U7850 (N_7850,N_7249,N_7235);
or U7851 (N_7851,N_7165,N_6552);
and U7852 (N_7852,N_6372,N_6482);
nor U7853 (N_7853,N_7166,N_6034);
xor U7854 (N_7854,N_6519,N_7336);
nor U7855 (N_7855,N_7456,N_6589);
or U7856 (N_7856,N_6445,N_6704);
nor U7857 (N_7857,N_7379,N_6517);
and U7858 (N_7858,N_7173,N_7002);
nand U7859 (N_7859,N_7124,N_7335);
xor U7860 (N_7860,N_7383,N_6881);
nor U7861 (N_7861,N_7381,N_6454);
nand U7862 (N_7862,N_6942,N_6927);
and U7863 (N_7863,N_6443,N_6755);
xnor U7864 (N_7864,N_6850,N_7388);
nand U7865 (N_7865,N_6413,N_7460);
nor U7866 (N_7866,N_6869,N_7118);
nor U7867 (N_7867,N_6955,N_6571);
and U7868 (N_7868,N_6262,N_6766);
nor U7869 (N_7869,N_6931,N_7395);
nor U7870 (N_7870,N_6423,N_6121);
nand U7871 (N_7871,N_7239,N_7481);
and U7872 (N_7872,N_6242,N_6067);
nor U7873 (N_7873,N_6173,N_6243);
nand U7874 (N_7874,N_6420,N_6750);
or U7875 (N_7875,N_6351,N_6148);
nor U7876 (N_7876,N_6015,N_7205);
or U7877 (N_7877,N_6460,N_6108);
nand U7878 (N_7878,N_6601,N_7020);
and U7879 (N_7879,N_6791,N_6713);
nor U7880 (N_7880,N_6972,N_6291);
nor U7881 (N_7881,N_6064,N_6094);
and U7882 (N_7882,N_7178,N_6465);
nand U7883 (N_7883,N_7180,N_6893);
xnor U7884 (N_7884,N_7222,N_7494);
nand U7885 (N_7885,N_6674,N_7164);
or U7886 (N_7886,N_7284,N_7017);
nand U7887 (N_7887,N_6575,N_6867);
and U7888 (N_7888,N_7012,N_6202);
nor U7889 (N_7889,N_7409,N_6143);
nand U7890 (N_7890,N_6848,N_6897);
nand U7891 (N_7891,N_7454,N_7448);
nand U7892 (N_7892,N_6775,N_6645);
xor U7893 (N_7893,N_6945,N_6919);
or U7894 (N_7894,N_6474,N_7075);
nand U7895 (N_7895,N_7307,N_7210);
nor U7896 (N_7896,N_7008,N_7055);
and U7897 (N_7897,N_6695,N_6807);
or U7898 (N_7898,N_6353,N_6548);
xor U7899 (N_7899,N_6593,N_6793);
nand U7900 (N_7900,N_6637,N_6550);
nor U7901 (N_7901,N_6126,N_6039);
xnor U7902 (N_7902,N_6384,N_6990);
xnor U7903 (N_7903,N_6288,N_6697);
and U7904 (N_7904,N_6688,N_6394);
xnor U7905 (N_7905,N_7009,N_7416);
and U7906 (N_7906,N_7300,N_6569);
and U7907 (N_7907,N_6700,N_6863);
and U7908 (N_7908,N_6049,N_6497);
or U7909 (N_7909,N_7190,N_6268);
xor U7910 (N_7910,N_6200,N_6197);
xnor U7911 (N_7911,N_7184,N_6182);
and U7912 (N_7912,N_6339,N_6816);
xor U7913 (N_7913,N_6319,N_6966);
or U7914 (N_7914,N_7030,N_7051);
or U7915 (N_7915,N_7264,N_6821);
xor U7916 (N_7916,N_6301,N_6253);
and U7917 (N_7917,N_6452,N_6626);
or U7918 (N_7918,N_6154,N_6754);
and U7919 (N_7919,N_6195,N_6705);
nor U7920 (N_7920,N_6658,N_6889);
nor U7921 (N_7921,N_6616,N_6107);
nand U7922 (N_7922,N_7404,N_6732);
or U7923 (N_7923,N_6278,N_6780);
xnor U7924 (N_7924,N_6213,N_7172);
xnor U7925 (N_7925,N_6833,N_7296);
or U7926 (N_7926,N_7084,N_6612);
and U7927 (N_7927,N_6973,N_7126);
nand U7928 (N_7928,N_6924,N_7054);
and U7929 (N_7929,N_7024,N_6082);
xor U7930 (N_7930,N_6588,N_6246);
nor U7931 (N_7931,N_6728,N_6910);
nor U7932 (N_7932,N_7287,N_6680);
nand U7933 (N_7933,N_6706,N_6506);
nor U7934 (N_7934,N_6007,N_6046);
and U7935 (N_7935,N_7466,N_7122);
xor U7936 (N_7936,N_7451,N_6393);
xor U7937 (N_7937,N_6520,N_6996);
nor U7938 (N_7938,N_6968,N_7133);
nor U7939 (N_7939,N_7313,N_7209);
and U7940 (N_7940,N_6904,N_6618);
nor U7941 (N_7941,N_6719,N_6141);
or U7942 (N_7942,N_7259,N_6357);
nand U7943 (N_7943,N_6515,N_6636);
nand U7944 (N_7944,N_6207,N_6553);
or U7945 (N_7945,N_6158,N_6939);
nor U7946 (N_7946,N_6817,N_6022);
nand U7947 (N_7947,N_6421,N_7037);
nand U7948 (N_7948,N_6053,N_6074);
or U7949 (N_7949,N_6016,N_6877);
and U7950 (N_7950,N_6438,N_6191);
nor U7951 (N_7951,N_7163,N_6160);
nand U7952 (N_7952,N_6653,N_6139);
or U7953 (N_7953,N_6422,N_6814);
nand U7954 (N_7954,N_7380,N_7310);
nand U7955 (N_7955,N_7413,N_6241);
xnor U7956 (N_7956,N_7200,N_6124);
xor U7957 (N_7957,N_7452,N_7208);
nor U7958 (N_7958,N_6426,N_7339);
and U7959 (N_7959,N_7116,N_6938);
xor U7960 (N_7960,N_6629,N_6965);
and U7961 (N_7961,N_7099,N_6899);
or U7962 (N_7962,N_6915,N_6555);
nor U7963 (N_7963,N_7244,N_6596);
nor U7964 (N_7964,N_7203,N_7373);
and U7965 (N_7965,N_7081,N_6453);
and U7966 (N_7966,N_6170,N_6375);
xor U7967 (N_7967,N_6468,N_7098);
or U7968 (N_7968,N_6313,N_7000);
nand U7969 (N_7969,N_6352,N_6934);
or U7970 (N_7970,N_7468,N_7363);
nand U7971 (N_7971,N_6773,N_6926);
or U7972 (N_7972,N_6625,N_6329);
nand U7973 (N_7973,N_6964,N_6088);
xor U7974 (N_7974,N_6574,N_6982);
nand U7975 (N_7975,N_6860,N_6774);
nor U7976 (N_7976,N_6884,N_6466);
nor U7977 (N_7977,N_6051,N_7107);
xnor U7978 (N_7978,N_6925,N_6611);
nor U7979 (N_7979,N_6513,N_6100);
xor U7980 (N_7980,N_6314,N_6906);
nor U7981 (N_7981,N_7274,N_6562);
xor U7982 (N_7982,N_6535,N_6398);
nand U7983 (N_7983,N_6592,N_6932);
nor U7984 (N_7984,N_6494,N_7476);
and U7985 (N_7985,N_6654,N_7436);
nor U7986 (N_7986,N_6150,N_6673);
nand U7987 (N_7987,N_6411,N_6193);
or U7988 (N_7988,N_7158,N_6429);
or U7989 (N_7989,N_6663,N_7295);
nor U7990 (N_7990,N_6178,N_7331);
nor U7991 (N_7991,N_6917,N_6020);
nor U7992 (N_7992,N_6036,N_6003);
xnor U7993 (N_7993,N_7042,N_6477);
or U7994 (N_7994,N_7291,N_7442);
or U7995 (N_7995,N_6364,N_6801);
nand U7996 (N_7996,N_6324,N_7195);
or U7997 (N_7997,N_6771,N_6134);
or U7998 (N_7998,N_6849,N_6681);
xor U7999 (N_7999,N_6401,N_6449);
nand U8000 (N_8000,N_6776,N_6113);
or U8001 (N_8001,N_6076,N_6737);
nand U8002 (N_8002,N_6269,N_7064);
or U8003 (N_8003,N_6783,N_6851);
or U8004 (N_8004,N_6266,N_6649);
nor U8005 (N_8005,N_6912,N_6410);
xnor U8006 (N_8006,N_6799,N_6878);
or U8007 (N_8007,N_7366,N_6083);
nor U8008 (N_8008,N_6117,N_7240);
or U8009 (N_8009,N_6403,N_6281);
nor U8010 (N_8010,N_6635,N_6525);
nand U8011 (N_8011,N_6233,N_7273);
and U8012 (N_8012,N_7153,N_6320);
and U8013 (N_8013,N_6323,N_6328);
or U8014 (N_8014,N_6263,N_6794);
or U8015 (N_8015,N_6008,N_6717);
nor U8016 (N_8016,N_7145,N_6312);
and U8017 (N_8017,N_6060,N_6105);
or U8018 (N_8018,N_6206,N_7131);
nand U8019 (N_8019,N_6578,N_6847);
nand U8020 (N_8020,N_6659,N_6145);
xor U8021 (N_8021,N_7345,N_6481);
nor U8022 (N_8022,N_6981,N_6138);
and U8023 (N_8023,N_7250,N_6740);
nor U8024 (N_8024,N_6933,N_7257);
nor U8025 (N_8025,N_6683,N_7138);
nor U8026 (N_8026,N_7202,N_7390);
and U8027 (N_8027,N_6451,N_6234);
nand U8028 (N_8028,N_7393,N_6838);
nand U8029 (N_8029,N_6164,N_6373);
or U8030 (N_8030,N_6962,N_6882);
nor U8031 (N_8031,N_7260,N_6509);
nor U8032 (N_8032,N_7389,N_6467);
and U8033 (N_8033,N_7437,N_6937);
nor U8034 (N_8034,N_7144,N_7470);
nand U8035 (N_8035,N_7130,N_7361);
and U8036 (N_8036,N_7212,N_6283);
nor U8037 (N_8037,N_6054,N_6205);
and U8038 (N_8038,N_6747,N_7152);
nand U8039 (N_8039,N_6811,N_7357);
or U8040 (N_8040,N_6874,N_6187);
nor U8041 (N_8041,N_6759,N_7216);
nand U8042 (N_8042,N_6872,N_6722);
nor U8043 (N_8043,N_7263,N_6909);
nor U8044 (N_8044,N_7167,N_7261);
nand U8045 (N_8045,N_6129,N_6630);
xor U8046 (N_8046,N_6743,N_6059);
or U8047 (N_8047,N_6341,N_6556);
and U8048 (N_8048,N_6014,N_6551);
nand U8049 (N_8049,N_6299,N_6387);
and U8050 (N_8050,N_7058,N_6986);
xnor U8051 (N_8051,N_6408,N_7258);
nand U8052 (N_8052,N_6211,N_6463);
or U8053 (N_8053,N_6298,N_6086);
or U8054 (N_8054,N_7499,N_7444);
nor U8055 (N_8055,N_6093,N_7391);
and U8056 (N_8056,N_6473,N_6785);
xnor U8057 (N_8057,N_6670,N_7321);
nor U8058 (N_8058,N_7417,N_6390);
xnor U8059 (N_8059,N_6866,N_6767);
xnor U8060 (N_8060,N_6041,N_7453);
nand U8061 (N_8061,N_6165,N_6249);
and U8062 (N_8062,N_6738,N_6400);
nand U8063 (N_8063,N_6168,N_7057);
nor U8064 (N_8064,N_6958,N_7348);
nor U8065 (N_8065,N_6261,N_7135);
nand U8066 (N_8066,N_7399,N_7226);
nor U8067 (N_8067,N_7169,N_6430);
or U8068 (N_8068,N_7473,N_6484);
xnor U8069 (N_8069,N_7402,N_6272);
nand U8070 (N_8070,N_6427,N_6488);
xnor U8071 (N_8071,N_7097,N_6797);
nand U8072 (N_8072,N_7046,N_6665);
or U8073 (N_8073,N_6111,N_6023);
or U8074 (N_8074,N_6533,N_6547);
xor U8075 (N_8075,N_6214,N_6508);
or U8076 (N_8076,N_6835,N_6177);
xor U8077 (N_8077,N_6080,N_6534);
and U8078 (N_8078,N_6396,N_6290);
or U8079 (N_8079,N_7346,N_7198);
or U8080 (N_8080,N_6439,N_6346);
xnor U8081 (N_8081,N_6057,N_6992);
nand U8082 (N_8082,N_6605,N_6500);
or U8083 (N_8083,N_6652,N_6651);
xnor U8084 (N_8084,N_6729,N_6530);
and U8085 (N_8085,N_6334,N_7186);
nor U8086 (N_8086,N_7059,N_6196);
and U8087 (N_8087,N_6406,N_6033);
nand U8088 (N_8088,N_6762,N_6916);
xor U8089 (N_8089,N_7179,N_7134);
or U8090 (N_8090,N_7023,N_6216);
nor U8091 (N_8091,N_6952,N_7256);
nor U8092 (N_8092,N_6078,N_7092);
xor U8093 (N_8093,N_7141,N_6018);
or U8094 (N_8094,N_6123,N_6804);
or U8095 (N_8095,N_6286,N_6125);
nand U8096 (N_8096,N_6032,N_6701);
xor U8097 (N_8097,N_6254,N_6584);
and U8098 (N_8098,N_7483,N_6920);
nand U8099 (N_8099,N_6676,N_6476);
and U8100 (N_8100,N_7341,N_6886);
nor U8101 (N_8101,N_6223,N_6345);
nand U8102 (N_8102,N_6563,N_7265);
nand U8103 (N_8103,N_6118,N_6140);
xor U8104 (N_8104,N_7199,N_6336);
nor U8105 (N_8105,N_6354,N_6987);
or U8106 (N_8106,N_6190,N_6864);
nor U8107 (N_8107,N_6752,N_6256);
nor U8108 (N_8108,N_6727,N_6950);
nand U8109 (N_8109,N_6043,N_7375);
xor U8110 (N_8110,N_7011,N_7101);
nor U8111 (N_8111,N_7330,N_6694);
nand U8112 (N_8112,N_6418,N_6052);
xor U8113 (N_8113,N_6789,N_6434);
or U8114 (N_8114,N_6416,N_6106);
or U8115 (N_8115,N_6409,N_6222);
and U8116 (N_8116,N_6545,N_6540);
nor U8117 (N_8117,N_6399,N_6935);
or U8118 (N_8118,N_6604,N_7405);
and U8119 (N_8119,N_6523,N_6858);
xor U8120 (N_8120,N_6235,N_7271);
nand U8121 (N_8121,N_6735,N_7299);
nand U8122 (N_8122,N_6859,N_7111);
nor U8123 (N_8123,N_7038,N_6210);
and U8124 (N_8124,N_7398,N_7061);
and U8125 (N_8125,N_6103,N_7353);
or U8126 (N_8126,N_6300,N_7215);
nand U8127 (N_8127,N_6642,N_6097);
or U8128 (N_8128,N_6166,N_6446);
nand U8129 (N_8129,N_6726,N_6836);
and U8130 (N_8130,N_6870,N_7489);
nand U8131 (N_8131,N_6853,N_7177);
nand U8132 (N_8132,N_7450,N_6583);
xor U8133 (N_8133,N_6936,N_6475);
or U8134 (N_8134,N_7438,N_6469);
or U8135 (N_8135,N_7372,N_6349);
or U8136 (N_8136,N_6837,N_6095);
nand U8137 (N_8137,N_6063,N_7477);
and U8138 (N_8138,N_7253,N_7162);
or U8139 (N_8139,N_7039,N_7026);
or U8140 (N_8140,N_6742,N_7364);
or U8141 (N_8141,N_7282,N_6279);
nor U8142 (N_8142,N_6229,N_7094);
or U8143 (N_8143,N_6382,N_6407);
xnor U8144 (N_8144,N_6010,N_6960);
and U8145 (N_8145,N_6492,N_6151);
nor U8146 (N_8146,N_6567,N_6317);
nand U8147 (N_8147,N_7117,N_6963);
xor U8148 (N_8148,N_6081,N_6994);
and U8149 (N_8149,N_6647,N_6303);
and U8150 (N_8150,N_6714,N_6546);
or U8151 (N_8151,N_6001,N_7262);
xnor U8152 (N_8152,N_7279,N_6265);
or U8153 (N_8153,N_7385,N_7487);
nand U8154 (N_8154,N_6252,N_6404);
xnor U8155 (N_8155,N_6293,N_7309);
xnor U8156 (N_8156,N_7189,N_6809);
xor U8157 (N_8157,N_6228,N_7027);
xnor U8158 (N_8158,N_7377,N_7086);
or U8159 (N_8159,N_7297,N_6948);
nor U8160 (N_8160,N_7241,N_7459);
nor U8161 (N_8161,N_7492,N_6725);
and U8162 (N_8162,N_6944,N_7252);
or U8163 (N_8163,N_6284,N_6614);
nand U8164 (N_8164,N_6976,N_7328);
and U8165 (N_8165,N_7185,N_6378);
or U8166 (N_8166,N_6980,N_7414);
and U8167 (N_8167,N_6084,N_7140);
nand U8168 (N_8168,N_7251,N_7093);
and U8169 (N_8169,N_6204,N_7493);
nand U8170 (N_8170,N_7447,N_7074);
xnor U8171 (N_8171,N_7192,N_6026);
nor U8172 (N_8172,N_7323,N_7418);
nand U8173 (N_8173,N_7480,N_6441);
nor U8174 (N_8174,N_6361,N_7183);
nand U8175 (N_8175,N_6276,N_6576);
nand U8176 (N_8176,N_7213,N_7334);
xor U8177 (N_8177,N_6892,N_7360);
and U8178 (N_8178,N_6128,N_6412);
xor U8179 (N_8179,N_6758,N_6514);
nand U8180 (N_8180,N_6251,N_6956);
and U8181 (N_8181,N_7181,N_6941);
xor U8182 (N_8182,N_6201,N_6998);
xor U8183 (N_8183,N_6524,N_6861);
xnor U8184 (N_8184,N_7425,N_6770);
nand U8185 (N_8185,N_6768,N_6839);
or U8186 (N_8186,N_7255,N_6885);
nand U8187 (N_8187,N_6756,N_6538);
xor U8188 (N_8188,N_6199,N_6829);
and U8189 (N_8189,N_6218,N_7431);
xnor U8190 (N_8190,N_7018,N_6760);
nor U8191 (N_8191,N_6448,N_7137);
and U8192 (N_8192,N_6769,N_6788);
nand U8193 (N_8193,N_7314,N_6504);
or U8194 (N_8194,N_7048,N_6101);
or U8195 (N_8195,N_6703,N_6607);
xnor U8196 (N_8196,N_6691,N_7491);
or U8197 (N_8197,N_6689,N_6175);
or U8198 (N_8198,N_6077,N_6823);
and U8199 (N_8199,N_6503,N_6038);
nand U8200 (N_8200,N_6602,N_6586);
or U8201 (N_8201,N_6194,N_6946);
nand U8202 (N_8202,N_6744,N_6993);
and U8203 (N_8203,N_6273,N_6184);
and U8204 (N_8204,N_6356,N_6779);
or U8205 (N_8205,N_7242,N_6189);
and U8206 (N_8206,N_7148,N_6639);
nand U8207 (N_8207,N_6581,N_6066);
nand U8208 (N_8208,N_6310,N_6822);
nand U8209 (N_8209,N_6819,N_6852);
and U8210 (N_8210,N_6854,N_6840);
or U8211 (N_8211,N_6617,N_7201);
and U8212 (N_8212,N_6790,N_6325);
xor U8213 (N_8213,N_7340,N_6970);
and U8214 (N_8214,N_6693,N_7376);
nand U8215 (N_8215,N_6479,N_6666);
nor U8216 (N_8216,N_6248,N_6062);
xor U8217 (N_8217,N_6203,N_6657);
nand U8218 (N_8218,N_6212,N_6072);
and U8219 (N_8219,N_6624,N_7403);
nor U8220 (N_8220,N_6042,N_6136);
nor U8221 (N_8221,N_7029,N_6608);
or U8222 (N_8222,N_7443,N_6185);
and U8223 (N_8223,N_7254,N_7427);
nor U8224 (N_8224,N_6296,N_7356);
or U8225 (N_8225,N_7343,N_7467);
xor U8226 (N_8226,N_6091,N_6250);
nor U8227 (N_8227,N_6056,N_7359);
and U8228 (N_8228,N_6710,N_6061);
xnor U8229 (N_8229,N_6957,N_6192);
nor U8230 (N_8230,N_7159,N_6812);
nand U8231 (N_8231,N_6085,N_6646);
or U8232 (N_8232,N_6419,N_7498);
or U8233 (N_8233,N_6495,N_6386);
nand U8234 (N_8234,N_7105,N_6490);
nand U8235 (N_8235,N_6739,N_6632);
and U8236 (N_8236,N_7462,N_7457);
nand U8237 (N_8237,N_7067,N_6741);
nand U8238 (N_8238,N_7031,N_6803);
nor U8239 (N_8239,N_6573,N_6961);
or U8240 (N_8240,N_7432,N_6954);
xnor U8241 (N_8241,N_6374,N_6764);
nand U8242 (N_8242,N_6692,N_6058);
nor U8243 (N_8243,N_6641,N_7384);
xor U8244 (N_8244,N_7119,N_6238);
and U8245 (N_8245,N_7280,N_6902);
and U8246 (N_8246,N_6684,N_6002);
and U8247 (N_8247,N_6677,N_7318);
or U8248 (N_8248,N_7229,N_6643);
and U8249 (N_8249,N_7445,N_7426);
and U8250 (N_8250,N_7075,N_6711);
nand U8251 (N_8251,N_6159,N_6816);
xnor U8252 (N_8252,N_6285,N_6335);
or U8253 (N_8253,N_6491,N_7334);
nor U8254 (N_8254,N_6479,N_6378);
nor U8255 (N_8255,N_6675,N_6256);
and U8256 (N_8256,N_6674,N_6443);
or U8257 (N_8257,N_6961,N_7289);
xnor U8258 (N_8258,N_6446,N_6619);
or U8259 (N_8259,N_7422,N_6757);
xnor U8260 (N_8260,N_7235,N_6466);
nand U8261 (N_8261,N_6328,N_6600);
and U8262 (N_8262,N_6977,N_6148);
nand U8263 (N_8263,N_6806,N_6751);
xnor U8264 (N_8264,N_6308,N_7386);
xnor U8265 (N_8265,N_6213,N_6003);
and U8266 (N_8266,N_7407,N_6632);
or U8267 (N_8267,N_6855,N_7228);
xor U8268 (N_8268,N_6770,N_6919);
nor U8269 (N_8269,N_7142,N_6050);
or U8270 (N_8270,N_6864,N_7328);
and U8271 (N_8271,N_7440,N_7164);
nand U8272 (N_8272,N_7272,N_7340);
or U8273 (N_8273,N_7400,N_6796);
and U8274 (N_8274,N_6413,N_7214);
or U8275 (N_8275,N_7052,N_6945);
or U8276 (N_8276,N_6702,N_6865);
or U8277 (N_8277,N_6696,N_6549);
nor U8278 (N_8278,N_6122,N_6690);
xnor U8279 (N_8279,N_7226,N_6525);
xnor U8280 (N_8280,N_6013,N_6106);
nand U8281 (N_8281,N_6532,N_7249);
and U8282 (N_8282,N_6310,N_7134);
nor U8283 (N_8283,N_6127,N_6967);
nand U8284 (N_8284,N_7259,N_6018);
nor U8285 (N_8285,N_6666,N_6476);
and U8286 (N_8286,N_6085,N_6975);
nand U8287 (N_8287,N_6648,N_7453);
nand U8288 (N_8288,N_6187,N_6362);
or U8289 (N_8289,N_6359,N_7011);
or U8290 (N_8290,N_7428,N_6646);
and U8291 (N_8291,N_7219,N_6496);
nor U8292 (N_8292,N_6797,N_6073);
nor U8293 (N_8293,N_6028,N_6003);
or U8294 (N_8294,N_7430,N_6917);
nand U8295 (N_8295,N_6711,N_6859);
and U8296 (N_8296,N_7469,N_7152);
nand U8297 (N_8297,N_6709,N_7019);
nor U8298 (N_8298,N_6838,N_6930);
and U8299 (N_8299,N_7000,N_6491);
nand U8300 (N_8300,N_7296,N_6717);
and U8301 (N_8301,N_6695,N_6487);
nor U8302 (N_8302,N_6805,N_7050);
nor U8303 (N_8303,N_7028,N_7333);
nand U8304 (N_8304,N_6818,N_7130);
or U8305 (N_8305,N_6815,N_7205);
and U8306 (N_8306,N_6189,N_6182);
nor U8307 (N_8307,N_6310,N_7142);
and U8308 (N_8308,N_7089,N_6269);
nor U8309 (N_8309,N_6230,N_6516);
or U8310 (N_8310,N_6304,N_6076);
and U8311 (N_8311,N_6988,N_6908);
or U8312 (N_8312,N_6609,N_7083);
or U8313 (N_8313,N_6556,N_7076);
nor U8314 (N_8314,N_6055,N_6467);
or U8315 (N_8315,N_7338,N_7467);
or U8316 (N_8316,N_6756,N_7410);
and U8317 (N_8317,N_6080,N_6930);
xnor U8318 (N_8318,N_7232,N_6182);
or U8319 (N_8319,N_7153,N_7043);
xnor U8320 (N_8320,N_6241,N_6646);
nor U8321 (N_8321,N_7099,N_6101);
nand U8322 (N_8322,N_7416,N_7326);
xnor U8323 (N_8323,N_7013,N_6154);
xnor U8324 (N_8324,N_6733,N_6666);
and U8325 (N_8325,N_6074,N_6761);
nand U8326 (N_8326,N_7010,N_6269);
xor U8327 (N_8327,N_7462,N_7368);
xor U8328 (N_8328,N_7401,N_6219);
and U8329 (N_8329,N_6988,N_6113);
or U8330 (N_8330,N_7359,N_6734);
nand U8331 (N_8331,N_7073,N_6929);
nand U8332 (N_8332,N_7334,N_6202);
xnor U8333 (N_8333,N_6161,N_7292);
and U8334 (N_8334,N_6291,N_7223);
or U8335 (N_8335,N_6206,N_7370);
nand U8336 (N_8336,N_6432,N_6063);
or U8337 (N_8337,N_6232,N_6112);
nor U8338 (N_8338,N_6792,N_6658);
xor U8339 (N_8339,N_6318,N_6927);
xnor U8340 (N_8340,N_6170,N_7456);
nor U8341 (N_8341,N_7482,N_6464);
xor U8342 (N_8342,N_6594,N_6123);
nor U8343 (N_8343,N_7452,N_7223);
nand U8344 (N_8344,N_6981,N_6747);
nor U8345 (N_8345,N_6682,N_6114);
or U8346 (N_8346,N_7383,N_6312);
or U8347 (N_8347,N_7067,N_7199);
xnor U8348 (N_8348,N_6927,N_7448);
nand U8349 (N_8349,N_6109,N_6217);
xnor U8350 (N_8350,N_7274,N_6083);
nor U8351 (N_8351,N_6146,N_6862);
nand U8352 (N_8352,N_6785,N_6368);
or U8353 (N_8353,N_6505,N_6292);
xnor U8354 (N_8354,N_7145,N_6591);
nand U8355 (N_8355,N_6770,N_7383);
nand U8356 (N_8356,N_6957,N_6235);
xnor U8357 (N_8357,N_7456,N_6981);
nand U8358 (N_8358,N_6161,N_7268);
xnor U8359 (N_8359,N_6870,N_7424);
nor U8360 (N_8360,N_7162,N_7051);
or U8361 (N_8361,N_6605,N_7229);
xnor U8362 (N_8362,N_6369,N_7310);
nand U8363 (N_8363,N_7376,N_6476);
or U8364 (N_8364,N_6959,N_6587);
nor U8365 (N_8365,N_7101,N_6611);
xnor U8366 (N_8366,N_7421,N_6840);
or U8367 (N_8367,N_7129,N_6665);
nand U8368 (N_8368,N_6550,N_6954);
nand U8369 (N_8369,N_6531,N_7084);
xor U8370 (N_8370,N_6026,N_7441);
xor U8371 (N_8371,N_6254,N_7163);
nor U8372 (N_8372,N_7329,N_6744);
or U8373 (N_8373,N_6015,N_6703);
xor U8374 (N_8374,N_6241,N_6572);
nor U8375 (N_8375,N_7180,N_6325);
or U8376 (N_8376,N_7153,N_6338);
or U8377 (N_8377,N_7103,N_6310);
or U8378 (N_8378,N_7386,N_6795);
and U8379 (N_8379,N_6985,N_6524);
nor U8380 (N_8380,N_7337,N_6404);
nor U8381 (N_8381,N_6756,N_7473);
nand U8382 (N_8382,N_6818,N_7139);
and U8383 (N_8383,N_6246,N_6574);
xnor U8384 (N_8384,N_7448,N_6215);
and U8385 (N_8385,N_6862,N_7131);
and U8386 (N_8386,N_6984,N_6628);
or U8387 (N_8387,N_6382,N_6589);
or U8388 (N_8388,N_6089,N_7405);
and U8389 (N_8389,N_7024,N_7326);
or U8390 (N_8390,N_7311,N_6660);
xnor U8391 (N_8391,N_6835,N_6526);
xor U8392 (N_8392,N_6206,N_6447);
and U8393 (N_8393,N_6660,N_7153);
nor U8394 (N_8394,N_6801,N_6681);
nand U8395 (N_8395,N_6348,N_6589);
or U8396 (N_8396,N_6006,N_7046);
nand U8397 (N_8397,N_6212,N_7088);
nor U8398 (N_8398,N_7156,N_7143);
nor U8399 (N_8399,N_6144,N_7492);
nand U8400 (N_8400,N_6605,N_6321);
xor U8401 (N_8401,N_6993,N_7037);
nor U8402 (N_8402,N_7004,N_6607);
nand U8403 (N_8403,N_7253,N_7421);
xnor U8404 (N_8404,N_6802,N_6592);
nor U8405 (N_8405,N_6841,N_6324);
nor U8406 (N_8406,N_6009,N_6915);
or U8407 (N_8407,N_6873,N_6618);
nand U8408 (N_8408,N_6548,N_6959);
and U8409 (N_8409,N_7167,N_6549);
nor U8410 (N_8410,N_6101,N_7215);
nand U8411 (N_8411,N_6455,N_7386);
and U8412 (N_8412,N_7111,N_7029);
nand U8413 (N_8413,N_6202,N_7009);
or U8414 (N_8414,N_6051,N_6124);
and U8415 (N_8415,N_6289,N_6153);
xnor U8416 (N_8416,N_6015,N_7489);
nand U8417 (N_8417,N_7446,N_6215);
or U8418 (N_8418,N_7009,N_6519);
or U8419 (N_8419,N_6056,N_6094);
and U8420 (N_8420,N_6568,N_6435);
nand U8421 (N_8421,N_6324,N_6954);
or U8422 (N_8422,N_7299,N_6834);
nand U8423 (N_8423,N_6585,N_7307);
or U8424 (N_8424,N_6406,N_6594);
nand U8425 (N_8425,N_6952,N_6639);
and U8426 (N_8426,N_6732,N_7051);
xor U8427 (N_8427,N_7222,N_6198);
nor U8428 (N_8428,N_6976,N_6149);
nand U8429 (N_8429,N_6794,N_7308);
nand U8430 (N_8430,N_6410,N_7161);
or U8431 (N_8431,N_6150,N_6313);
or U8432 (N_8432,N_7161,N_6876);
and U8433 (N_8433,N_6790,N_7064);
nand U8434 (N_8434,N_6273,N_6754);
nor U8435 (N_8435,N_7320,N_6965);
nor U8436 (N_8436,N_6799,N_6122);
nor U8437 (N_8437,N_6147,N_6379);
nor U8438 (N_8438,N_6542,N_7198);
nand U8439 (N_8439,N_7300,N_7121);
nand U8440 (N_8440,N_7227,N_6945);
xor U8441 (N_8441,N_6997,N_6831);
nor U8442 (N_8442,N_6449,N_6611);
nor U8443 (N_8443,N_6323,N_6635);
xor U8444 (N_8444,N_6839,N_6431);
xor U8445 (N_8445,N_6024,N_6343);
xor U8446 (N_8446,N_6468,N_6414);
nand U8447 (N_8447,N_6664,N_7349);
nor U8448 (N_8448,N_7215,N_6105);
nand U8449 (N_8449,N_6439,N_7352);
nand U8450 (N_8450,N_6762,N_7296);
xor U8451 (N_8451,N_6215,N_6568);
nand U8452 (N_8452,N_6116,N_6770);
xnor U8453 (N_8453,N_6336,N_6879);
or U8454 (N_8454,N_7310,N_7172);
or U8455 (N_8455,N_7297,N_6022);
or U8456 (N_8456,N_7477,N_6935);
and U8457 (N_8457,N_7497,N_6676);
and U8458 (N_8458,N_6783,N_6662);
and U8459 (N_8459,N_7432,N_6690);
or U8460 (N_8460,N_7041,N_6664);
xnor U8461 (N_8461,N_7442,N_6471);
xnor U8462 (N_8462,N_6444,N_6642);
and U8463 (N_8463,N_6357,N_7205);
xor U8464 (N_8464,N_6942,N_6042);
or U8465 (N_8465,N_6859,N_6690);
nor U8466 (N_8466,N_6821,N_6492);
and U8467 (N_8467,N_7038,N_6571);
and U8468 (N_8468,N_6997,N_6948);
nor U8469 (N_8469,N_6177,N_6925);
nand U8470 (N_8470,N_7245,N_6304);
xnor U8471 (N_8471,N_6012,N_7199);
and U8472 (N_8472,N_6888,N_6498);
and U8473 (N_8473,N_6719,N_6178);
or U8474 (N_8474,N_7411,N_7440);
nand U8475 (N_8475,N_6886,N_6188);
xor U8476 (N_8476,N_7294,N_6325);
and U8477 (N_8477,N_6700,N_6014);
nor U8478 (N_8478,N_7376,N_6828);
and U8479 (N_8479,N_6148,N_7343);
nand U8480 (N_8480,N_7371,N_6226);
and U8481 (N_8481,N_6941,N_6785);
nand U8482 (N_8482,N_6770,N_7243);
xnor U8483 (N_8483,N_6945,N_6025);
nor U8484 (N_8484,N_6795,N_7208);
and U8485 (N_8485,N_6716,N_6206);
and U8486 (N_8486,N_6138,N_7246);
and U8487 (N_8487,N_7357,N_7135);
nand U8488 (N_8488,N_7364,N_6346);
nor U8489 (N_8489,N_6855,N_6417);
xor U8490 (N_8490,N_7090,N_6235);
nor U8491 (N_8491,N_7046,N_7453);
and U8492 (N_8492,N_6535,N_6639);
xnor U8493 (N_8493,N_7255,N_6006);
or U8494 (N_8494,N_6534,N_6962);
and U8495 (N_8495,N_6648,N_6617);
or U8496 (N_8496,N_7074,N_6554);
and U8497 (N_8497,N_6605,N_6995);
or U8498 (N_8498,N_6981,N_6028);
nand U8499 (N_8499,N_6189,N_6485);
or U8500 (N_8500,N_6958,N_7490);
nor U8501 (N_8501,N_7433,N_6693);
and U8502 (N_8502,N_6390,N_6618);
or U8503 (N_8503,N_6888,N_6319);
nand U8504 (N_8504,N_6988,N_6213);
or U8505 (N_8505,N_6880,N_7425);
nand U8506 (N_8506,N_6828,N_6014);
xnor U8507 (N_8507,N_7087,N_6641);
or U8508 (N_8508,N_6978,N_6799);
nand U8509 (N_8509,N_7072,N_6881);
or U8510 (N_8510,N_6553,N_6165);
xnor U8511 (N_8511,N_6830,N_6475);
and U8512 (N_8512,N_6610,N_6893);
or U8513 (N_8513,N_6868,N_6163);
or U8514 (N_8514,N_6375,N_6528);
nand U8515 (N_8515,N_6204,N_6447);
or U8516 (N_8516,N_6532,N_6812);
and U8517 (N_8517,N_7268,N_6017);
nand U8518 (N_8518,N_7279,N_7024);
or U8519 (N_8519,N_7137,N_7034);
or U8520 (N_8520,N_7399,N_6686);
or U8521 (N_8521,N_6448,N_6978);
nand U8522 (N_8522,N_6341,N_7154);
nor U8523 (N_8523,N_6049,N_6474);
nand U8524 (N_8524,N_6499,N_6687);
xor U8525 (N_8525,N_7225,N_7155);
or U8526 (N_8526,N_6287,N_6506);
xnor U8527 (N_8527,N_7305,N_6463);
nand U8528 (N_8528,N_6288,N_6342);
nand U8529 (N_8529,N_6193,N_6802);
or U8530 (N_8530,N_6808,N_7056);
and U8531 (N_8531,N_6050,N_6605);
nand U8532 (N_8532,N_6957,N_6229);
or U8533 (N_8533,N_6814,N_7241);
nor U8534 (N_8534,N_6909,N_6315);
nor U8535 (N_8535,N_6321,N_6390);
nor U8536 (N_8536,N_7327,N_7384);
nor U8537 (N_8537,N_6206,N_7441);
nor U8538 (N_8538,N_6095,N_7138);
or U8539 (N_8539,N_7146,N_6216);
or U8540 (N_8540,N_6199,N_7150);
or U8541 (N_8541,N_7239,N_7034);
nor U8542 (N_8542,N_6998,N_6665);
and U8543 (N_8543,N_6311,N_7248);
nand U8544 (N_8544,N_6444,N_6729);
nor U8545 (N_8545,N_7245,N_6505);
nor U8546 (N_8546,N_6728,N_6138);
nand U8547 (N_8547,N_7057,N_6036);
nor U8548 (N_8548,N_7397,N_6144);
or U8549 (N_8549,N_6085,N_6665);
or U8550 (N_8550,N_6375,N_6983);
or U8551 (N_8551,N_6330,N_6996);
nand U8552 (N_8552,N_7249,N_6203);
nor U8553 (N_8553,N_7105,N_6510);
nand U8554 (N_8554,N_7082,N_7496);
nor U8555 (N_8555,N_6020,N_7282);
nor U8556 (N_8556,N_6539,N_6797);
xor U8557 (N_8557,N_6587,N_6949);
or U8558 (N_8558,N_6689,N_6013);
and U8559 (N_8559,N_6416,N_6417);
or U8560 (N_8560,N_7044,N_6876);
or U8561 (N_8561,N_6284,N_6654);
xnor U8562 (N_8562,N_7299,N_6271);
and U8563 (N_8563,N_6310,N_6594);
nor U8564 (N_8564,N_6754,N_7419);
or U8565 (N_8565,N_6394,N_6959);
and U8566 (N_8566,N_6074,N_6927);
nor U8567 (N_8567,N_6070,N_7077);
and U8568 (N_8568,N_7268,N_6451);
nand U8569 (N_8569,N_6657,N_6434);
or U8570 (N_8570,N_6548,N_6628);
nor U8571 (N_8571,N_6921,N_6826);
and U8572 (N_8572,N_7212,N_7163);
xnor U8573 (N_8573,N_7339,N_7178);
xor U8574 (N_8574,N_6524,N_6028);
nor U8575 (N_8575,N_6006,N_6937);
xnor U8576 (N_8576,N_6735,N_6716);
nor U8577 (N_8577,N_6347,N_6201);
nor U8578 (N_8578,N_6115,N_6366);
xnor U8579 (N_8579,N_7428,N_6075);
nor U8580 (N_8580,N_6556,N_6055);
and U8581 (N_8581,N_6751,N_7127);
and U8582 (N_8582,N_6310,N_6785);
nand U8583 (N_8583,N_7252,N_6056);
nor U8584 (N_8584,N_6714,N_7123);
or U8585 (N_8585,N_6949,N_7352);
nand U8586 (N_8586,N_7240,N_6461);
or U8587 (N_8587,N_6978,N_7242);
xnor U8588 (N_8588,N_6703,N_7009);
nand U8589 (N_8589,N_6311,N_6891);
and U8590 (N_8590,N_7107,N_7452);
xor U8591 (N_8591,N_6854,N_6773);
and U8592 (N_8592,N_6567,N_6295);
or U8593 (N_8593,N_6371,N_7363);
and U8594 (N_8594,N_6975,N_7060);
and U8595 (N_8595,N_7117,N_7021);
nor U8596 (N_8596,N_6336,N_6021);
xnor U8597 (N_8597,N_6547,N_6490);
nor U8598 (N_8598,N_7300,N_6379);
xnor U8599 (N_8599,N_6709,N_6723);
nor U8600 (N_8600,N_6122,N_6232);
or U8601 (N_8601,N_7146,N_7168);
and U8602 (N_8602,N_7099,N_6239);
xnor U8603 (N_8603,N_7013,N_6948);
nand U8604 (N_8604,N_7409,N_6799);
xnor U8605 (N_8605,N_6548,N_6236);
xnor U8606 (N_8606,N_6481,N_7490);
nand U8607 (N_8607,N_6737,N_6383);
nand U8608 (N_8608,N_6702,N_6672);
xnor U8609 (N_8609,N_6582,N_6565);
and U8610 (N_8610,N_6386,N_6325);
xnor U8611 (N_8611,N_7472,N_6165);
xnor U8612 (N_8612,N_6221,N_6751);
nand U8613 (N_8613,N_6930,N_7299);
xnor U8614 (N_8614,N_6677,N_6707);
and U8615 (N_8615,N_6124,N_7349);
nor U8616 (N_8616,N_6166,N_6477);
nor U8617 (N_8617,N_6173,N_6579);
xnor U8618 (N_8618,N_6554,N_6241);
nand U8619 (N_8619,N_7088,N_6221);
nand U8620 (N_8620,N_6970,N_6633);
nand U8621 (N_8621,N_6308,N_7494);
nor U8622 (N_8622,N_6365,N_6373);
nor U8623 (N_8623,N_6402,N_6569);
and U8624 (N_8624,N_6281,N_6873);
nand U8625 (N_8625,N_6577,N_7356);
xor U8626 (N_8626,N_6968,N_6100);
nor U8627 (N_8627,N_7111,N_7131);
xor U8628 (N_8628,N_6436,N_7016);
xnor U8629 (N_8629,N_6877,N_7282);
xor U8630 (N_8630,N_6896,N_7193);
and U8631 (N_8631,N_6245,N_6490);
xnor U8632 (N_8632,N_7005,N_6082);
or U8633 (N_8633,N_6851,N_7239);
nor U8634 (N_8634,N_6518,N_7086);
xor U8635 (N_8635,N_6879,N_6506);
nor U8636 (N_8636,N_6234,N_6962);
nor U8637 (N_8637,N_6486,N_7009);
xnor U8638 (N_8638,N_6934,N_7403);
nand U8639 (N_8639,N_6104,N_7445);
nor U8640 (N_8640,N_6884,N_6623);
or U8641 (N_8641,N_6124,N_6306);
xor U8642 (N_8642,N_7132,N_6332);
xor U8643 (N_8643,N_6288,N_6637);
nor U8644 (N_8644,N_6136,N_7211);
xor U8645 (N_8645,N_7279,N_6793);
nor U8646 (N_8646,N_7259,N_6432);
or U8647 (N_8647,N_6869,N_7398);
or U8648 (N_8648,N_6761,N_6797);
and U8649 (N_8649,N_6493,N_6143);
nor U8650 (N_8650,N_7293,N_7158);
nand U8651 (N_8651,N_6285,N_6855);
xnor U8652 (N_8652,N_6316,N_7208);
nand U8653 (N_8653,N_7094,N_6606);
nor U8654 (N_8654,N_6102,N_7375);
xnor U8655 (N_8655,N_7449,N_6307);
and U8656 (N_8656,N_6620,N_6797);
or U8657 (N_8657,N_6910,N_6347);
xor U8658 (N_8658,N_6021,N_7004);
xor U8659 (N_8659,N_6254,N_6467);
xnor U8660 (N_8660,N_7318,N_6834);
nor U8661 (N_8661,N_7198,N_7044);
xor U8662 (N_8662,N_6244,N_6313);
nor U8663 (N_8663,N_7003,N_6161);
nor U8664 (N_8664,N_6806,N_7379);
and U8665 (N_8665,N_6126,N_6601);
and U8666 (N_8666,N_6033,N_7039);
nand U8667 (N_8667,N_6519,N_6742);
and U8668 (N_8668,N_6473,N_7159);
xnor U8669 (N_8669,N_7153,N_6750);
and U8670 (N_8670,N_6781,N_6191);
or U8671 (N_8671,N_6276,N_6903);
xor U8672 (N_8672,N_7325,N_7486);
nand U8673 (N_8673,N_6923,N_7177);
and U8674 (N_8674,N_6696,N_7257);
nand U8675 (N_8675,N_6874,N_7487);
or U8676 (N_8676,N_7386,N_6638);
xnor U8677 (N_8677,N_7016,N_7254);
and U8678 (N_8678,N_7162,N_6493);
and U8679 (N_8679,N_6397,N_6608);
nand U8680 (N_8680,N_6181,N_6546);
nor U8681 (N_8681,N_7397,N_6570);
nor U8682 (N_8682,N_7482,N_6485);
nor U8683 (N_8683,N_7426,N_6047);
nand U8684 (N_8684,N_7478,N_6643);
xor U8685 (N_8685,N_7453,N_6710);
and U8686 (N_8686,N_7064,N_7397);
or U8687 (N_8687,N_7177,N_6580);
xnor U8688 (N_8688,N_6494,N_6275);
or U8689 (N_8689,N_6113,N_6775);
nand U8690 (N_8690,N_7040,N_6753);
or U8691 (N_8691,N_7369,N_7201);
nor U8692 (N_8692,N_6366,N_6519);
nor U8693 (N_8693,N_7302,N_6465);
xnor U8694 (N_8694,N_7132,N_7010);
nor U8695 (N_8695,N_7196,N_7430);
nand U8696 (N_8696,N_6100,N_7438);
xor U8697 (N_8697,N_7344,N_6529);
nand U8698 (N_8698,N_6134,N_6923);
nand U8699 (N_8699,N_7461,N_7356);
nand U8700 (N_8700,N_7151,N_6073);
or U8701 (N_8701,N_7378,N_7057);
nand U8702 (N_8702,N_7022,N_6295);
xor U8703 (N_8703,N_6109,N_6711);
xnor U8704 (N_8704,N_6815,N_6274);
and U8705 (N_8705,N_6098,N_6262);
and U8706 (N_8706,N_7147,N_6787);
or U8707 (N_8707,N_6726,N_7280);
nor U8708 (N_8708,N_6703,N_6042);
and U8709 (N_8709,N_6545,N_6323);
nand U8710 (N_8710,N_6215,N_7424);
xor U8711 (N_8711,N_6556,N_7277);
or U8712 (N_8712,N_6882,N_6362);
and U8713 (N_8713,N_6745,N_6554);
and U8714 (N_8714,N_7023,N_6007);
and U8715 (N_8715,N_6924,N_7108);
xnor U8716 (N_8716,N_6047,N_6964);
xnor U8717 (N_8717,N_7483,N_6870);
and U8718 (N_8718,N_7483,N_6008);
nor U8719 (N_8719,N_7302,N_6071);
nand U8720 (N_8720,N_6628,N_6058);
nor U8721 (N_8721,N_6334,N_7430);
nand U8722 (N_8722,N_7364,N_7415);
or U8723 (N_8723,N_6657,N_6879);
and U8724 (N_8724,N_7491,N_7376);
nand U8725 (N_8725,N_6020,N_6231);
nor U8726 (N_8726,N_6920,N_6418);
and U8727 (N_8727,N_6104,N_6459);
or U8728 (N_8728,N_7063,N_6346);
nand U8729 (N_8729,N_6658,N_7396);
xnor U8730 (N_8730,N_7171,N_6412);
and U8731 (N_8731,N_7195,N_6624);
xor U8732 (N_8732,N_6002,N_6444);
nor U8733 (N_8733,N_7337,N_7444);
or U8734 (N_8734,N_6323,N_6067);
xor U8735 (N_8735,N_6475,N_6603);
or U8736 (N_8736,N_6175,N_6736);
xor U8737 (N_8737,N_6133,N_6332);
and U8738 (N_8738,N_6096,N_7339);
nor U8739 (N_8739,N_6065,N_6818);
nor U8740 (N_8740,N_7425,N_6849);
or U8741 (N_8741,N_6168,N_6644);
or U8742 (N_8742,N_6512,N_7444);
nor U8743 (N_8743,N_6722,N_7163);
nor U8744 (N_8744,N_7086,N_6935);
xor U8745 (N_8745,N_6668,N_6546);
nor U8746 (N_8746,N_6000,N_6992);
xor U8747 (N_8747,N_6566,N_6070);
xnor U8748 (N_8748,N_6346,N_6986);
nor U8749 (N_8749,N_6301,N_6636);
and U8750 (N_8750,N_6779,N_6589);
or U8751 (N_8751,N_6371,N_7002);
xnor U8752 (N_8752,N_7124,N_6571);
xnor U8753 (N_8753,N_7019,N_6804);
xor U8754 (N_8754,N_6762,N_7226);
and U8755 (N_8755,N_7214,N_6627);
and U8756 (N_8756,N_7059,N_6295);
nor U8757 (N_8757,N_6549,N_6094);
xor U8758 (N_8758,N_7392,N_6987);
xnor U8759 (N_8759,N_6115,N_7048);
nor U8760 (N_8760,N_6547,N_6756);
and U8761 (N_8761,N_7312,N_6521);
or U8762 (N_8762,N_6515,N_6250);
nor U8763 (N_8763,N_6564,N_7199);
and U8764 (N_8764,N_6434,N_6871);
nor U8765 (N_8765,N_6515,N_7014);
nor U8766 (N_8766,N_6617,N_7190);
xnor U8767 (N_8767,N_6891,N_6317);
nor U8768 (N_8768,N_7019,N_7039);
xnor U8769 (N_8769,N_7306,N_6952);
nand U8770 (N_8770,N_6215,N_7087);
nor U8771 (N_8771,N_6897,N_7038);
and U8772 (N_8772,N_6619,N_6527);
or U8773 (N_8773,N_6600,N_6921);
xor U8774 (N_8774,N_6723,N_7162);
nor U8775 (N_8775,N_6432,N_6007);
xnor U8776 (N_8776,N_6702,N_7131);
nand U8777 (N_8777,N_7244,N_6309);
nand U8778 (N_8778,N_7052,N_6782);
nand U8779 (N_8779,N_6565,N_6025);
nand U8780 (N_8780,N_6794,N_7084);
or U8781 (N_8781,N_7332,N_6765);
nand U8782 (N_8782,N_6690,N_6284);
nor U8783 (N_8783,N_7001,N_7406);
nor U8784 (N_8784,N_7021,N_6875);
and U8785 (N_8785,N_7422,N_6269);
and U8786 (N_8786,N_6685,N_7028);
nor U8787 (N_8787,N_6667,N_6295);
nor U8788 (N_8788,N_7435,N_7075);
nand U8789 (N_8789,N_6834,N_6582);
or U8790 (N_8790,N_6356,N_6104);
xnor U8791 (N_8791,N_6587,N_6586);
nand U8792 (N_8792,N_6115,N_6385);
and U8793 (N_8793,N_6028,N_6124);
nor U8794 (N_8794,N_6683,N_6184);
xor U8795 (N_8795,N_6227,N_6755);
nand U8796 (N_8796,N_6910,N_7091);
and U8797 (N_8797,N_6516,N_6214);
or U8798 (N_8798,N_7122,N_6545);
xnor U8799 (N_8799,N_6625,N_6442);
and U8800 (N_8800,N_6353,N_6588);
and U8801 (N_8801,N_6469,N_6938);
or U8802 (N_8802,N_6825,N_6813);
nand U8803 (N_8803,N_6956,N_6742);
nand U8804 (N_8804,N_7422,N_6556);
nand U8805 (N_8805,N_6683,N_7263);
or U8806 (N_8806,N_6981,N_6547);
nand U8807 (N_8807,N_6171,N_7408);
nand U8808 (N_8808,N_7481,N_7202);
nor U8809 (N_8809,N_6910,N_6352);
or U8810 (N_8810,N_7467,N_6661);
xor U8811 (N_8811,N_7123,N_6509);
or U8812 (N_8812,N_7029,N_6109);
or U8813 (N_8813,N_7297,N_6926);
xnor U8814 (N_8814,N_6659,N_7429);
or U8815 (N_8815,N_7169,N_7262);
xnor U8816 (N_8816,N_7220,N_6525);
xnor U8817 (N_8817,N_7165,N_7008);
nand U8818 (N_8818,N_7065,N_7245);
and U8819 (N_8819,N_7491,N_6283);
nor U8820 (N_8820,N_7213,N_6268);
nand U8821 (N_8821,N_6243,N_7266);
xnor U8822 (N_8822,N_6629,N_7349);
xor U8823 (N_8823,N_6402,N_6278);
nor U8824 (N_8824,N_7312,N_7451);
nand U8825 (N_8825,N_6484,N_6126);
nand U8826 (N_8826,N_6457,N_7014);
or U8827 (N_8827,N_7271,N_7363);
and U8828 (N_8828,N_6830,N_7258);
xor U8829 (N_8829,N_7218,N_6383);
nand U8830 (N_8830,N_7254,N_6570);
nand U8831 (N_8831,N_6283,N_6909);
and U8832 (N_8832,N_6926,N_6493);
xnor U8833 (N_8833,N_6498,N_6485);
nor U8834 (N_8834,N_6552,N_6996);
or U8835 (N_8835,N_7390,N_7331);
xnor U8836 (N_8836,N_6389,N_6996);
or U8837 (N_8837,N_6827,N_6020);
or U8838 (N_8838,N_7254,N_6810);
nor U8839 (N_8839,N_7047,N_7427);
nor U8840 (N_8840,N_6106,N_6520);
or U8841 (N_8841,N_6365,N_7164);
nor U8842 (N_8842,N_6241,N_7297);
and U8843 (N_8843,N_6939,N_7044);
xnor U8844 (N_8844,N_6290,N_7055);
nor U8845 (N_8845,N_6582,N_6238);
xor U8846 (N_8846,N_6203,N_7398);
or U8847 (N_8847,N_6802,N_7324);
nand U8848 (N_8848,N_6397,N_7081);
and U8849 (N_8849,N_6493,N_6272);
nor U8850 (N_8850,N_6179,N_7454);
and U8851 (N_8851,N_7073,N_6876);
xnor U8852 (N_8852,N_7451,N_6076);
or U8853 (N_8853,N_7149,N_7248);
nor U8854 (N_8854,N_7254,N_7251);
nor U8855 (N_8855,N_6200,N_6274);
or U8856 (N_8856,N_6920,N_7423);
nand U8857 (N_8857,N_6757,N_6962);
nand U8858 (N_8858,N_6066,N_7254);
nor U8859 (N_8859,N_6719,N_6680);
nand U8860 (N_8860,N_6284,N_6785);
nand U8861 (N_8861,N_6576,N_6599);
nand U8862 (N_8862,N_6315,N_6245);
nor U8863 (N_8863,N_7056,N_6364);
or U8864 (N_8864,N_6633,N_6015);
and U8865 (N_8865,N_6762,N_6655);
or U8866 (N_8866,N_7174,N_6934);
xor U8867 (N_8867,N_6251,N_6086);
nor U8868 (N_8868,N_7090,N_7442);
nor U8869 (N_8869,N_6772,N_7479);
xnor U8870 (N_8870,N_6594,N_6399);
xor U8871 (N_8871,N_6999,N_7301);
and U8872 (N_8872,N_7098,N_7249);
nand U8873 (N_8873,N_6387,N_7438);
nand U8874 (N_8874,N_6039,N_6266);
or U8875 (N_8875,N_6779,N_6437);
nand U8876 (N_8876,N_6898,N_6578);
or U8877 (N_8877,N_7052,N_6570);
nand U8878 (N_8878,N_7230,N_7381);
xor U8879 (N_8879,N_6838,N_6049);
or U8880 (N_8880,N_7375,N_6591);
and U8881 (N_8881,N_6820,N_7240);
and U8882 (N_8882,N_6164,N_7367);
nor U8883 (N_8883,N_7498,N_6290);
xnor U8884 (N_8884,N_7440,N_7184);
or U8885 (N_8885,N_6344,N_6037);
or U8886 (N_8886,N_6844,N_7214);
nor U8887 (N_8887,N_6908,N_6017);
and U8888 (N_8888,N_6541,N_6891);
or U8889 (N_8889,N_6544,N_6067);
nor U8890 (N_8890,N_6022,N_7195);
nor U8891 (N_8891,N_7462,N_7327);
xor U8892 (N_8892,N_6815,N_6220);
and U8893 (N_8893,N_6956,N_6655);
nand U8894 (N_8894,N_6882,N_7259);
nand U8895 (N_8895,N_6854,N_6762);
nand U8896 (N_8896,N_6768,N_6615);
and U8897 (N_8897,N_6332,N_7314);
xor U8898 (N_8898,N_7418,N_6594);
nand U8899 (N_8899,N_7098,N_6601);
or U8900 (N_8900,N_6551,N_6598);
and U8901 (N_8901,N_7054,N_6651);
nand U8902 (N_8902,N_6422,N_6115);
nor U8903 (N_8903,N_7045,N_7085);
xnor U8904 (N_8904,N_6700,N_6028);
nor U8905 (N_8905,N_6352,N_6141);
or U8906 (N_8906,N_7296,N_6552);
xor U8907 (N_8907,N_6720,N_7437);
or U8908 (N_8908,N_7413,N_6302);
nor U8909 (N_8909,N_6689,N_6305);
nand U8910 (N_8910,N_7483,N_7260);
xnor U8911 (N_8911,N_7249,N_7494);
and U8912 (N_8912,N_6142,N_6119);
nand U8913 (N_8913,N_6933,N_6008);
or U8914 (N_8914,N_6067,N_6248);
xor U8915 (N_8915,N_7120,N_6073);
xor U8916 (N_8916,N_6902,N_7445);
or U8917 (N_8917,N_6109,N_7491);
nand U8918 (N_8918,N_7007,N_7172);
nor U8919 (N_8919,N_7130,N_6194);
nor U8920 (N_8920,N_7376,N_6986);
nor U8921 (N_8921,N_6509,N_6445);
and U8922 (N_8922,N_7220,N_7459);
and U8923 (N_8923,N_7482,N_6549);
nor U8924 (N_8924,N_7155,N_7062);
nor U8925 (N_8925,N_6633,N_6722);
xor U8926 (N_8926,N_6651,N_6305);
nand U8927 (N_8927,N_7189,N_6210);
or U8928 (N_8928,N_6090,N_7023);
and U8929 (N_8929,N_6284,N_6475);
and U8930 (N_8930,N_6236,N_6349);
and U8931 (N_8931,N_7498,N_6008);
and U8932 (N_8932,N_6701,N_6679);
or U8933 (N_8933,N_6612,N_7411);
or U8934 (N_8934,N_6470,N_6673);
or U8935 (N_8935,N_6898,N_7056);
nand U8936 (N_8936,N_6944,N_6429);
nand U8937 (N_8937,N_6063,N_7134);
xor U8938 (N_8938,N_7064,N_6560);
and U8939 (N_8939,N_6044,N_6303);
nor U8940 (N_8940,N_6019,N_7357);
xor U8941 (N_8941,N_6713,N_6313);
or U8942 (N_8942,N_7130,N_6491);
xor U8943 (N_8943,N_6071,N_7246);
or U8944 (N_8944,N_6328,N_6586);
or U8945 (N_8945,N_6805,N_6012);
nand U8946 (N_8946,N_6672,N_7396);
xor U8947 (N_8947,N_6745,N_6074);
or U8948 (N_8948,N_7042,N_7251);
xor U8949 (N_8949,N_6951,N_7330);
nand U8950 (N_8950,N_6919,N_6982);
or U8951 (N_8951,N_7480,N_6583);
xnor U8952 (N_8952,N_7397,N_6708);
and U8953 (N_8953,N_6025,N_6108);
nand U8954 (N_8954,N_6314,N_7041);
nor U8955 (N_8955,N_6317,N_7123);
or U8956 (N_8956,N_7404,N_6193);
and U8957 (N_8957,N_6820,N_6900);
nor U8958 (N_8958,N_7027,N_7335);
nor U8959 (N_8959,N_6500,N_6766);
or U8960 (N_8960,N_6945,N_6819);
nand U8961 (N_8961,N_7273,N_7370);
or U8962 (N_8962,N_7425,N_6532);
and U8963 (N_8963,N_7304,N_6766);
and U8964 (N_8964,N_7466,N_6305);
or U8965 (N_8965,N_6672,N_7128);
or U8966 (N_8966,N_6663,N_7321);
or U8967 (N_8967,N_6154,N_6803);
nand U8968 (N_8968,N_6852,N_7104);
and U8969 (N_8969,N_7336,N_6423);
xor U8970 (N_8970,N_6551,N_6851);
nand U8971 (N_8971,N_6423,N_7037);
nand U8972 (N_8972,N_6734,N_6039);
nand U8973 (N_8973,N_6143,N_6477);
nor U8974 (N_8974,N_6949,N_7128);
or U8975 (N_8975,N_7032,N_6130);
nor U8976 (N_8976,N_6327,N_6884);
and U8977 (N_8977,N_6467,N_6249);
and U8978 (N_8978,N_7378,N_7100);
and U8979 (N_8979,N_6455,N_6219);
and U8980 (N_8980,N_6591,N_6142);
xnor U8981 (N_8981,N_6415,N_6869);
and U8982 (N_8982,N_6087,N_6798);
nor U8983 (N_8983,N_6181,N_6708);
nand U8984 (N_8984,N_6913,N_7482);
or U8985 (N_8985,N_6001,N_6399);
nor U8986 (N_8986,N_6382,N_7165);
nor U8987 (N_8987,N_6005,N_6227);
nand U8988 (N_8988,N_7234,N_7493);
or U8989 (N_8989,N_6862,N_6246);
and U8990 (N_8990,N_6793,N_6193);
nand U8991 (N_8991,N_7010,N_7075);
nand U8992 (N_8992,N_6911,N_6060);
nor U8993 (N_8993,N_6956,N_7129);
xnor U8994 (N_8994,N_6897,N_6328);
xnor U8995 (N_8995,N_7170,N_6932);
nand U8996 (N_8996,N_6450,N_6444);
and U8997 (N_8997,N_6390,N_6751);
nor U8998 (N_8998,N_7248,N_7378);
nand U8999 (N_8999,N_6180,N_7496);
or U9000 (N_9000,N_7680,N_8220);
nor U9001 (N_9001,N_8621,N_8329);
or U9002 (N_9002,N_8385,N_8663);
nand U9003 (N_9003,N_7873,N_7523);
nand U9004 (N_9004,N_8275,N_8611);
nand U9005 (N_9005,N_7593,N_8752);
or U9006 (N_9006,N_8513,N_8521);
and U9007 (N_9007,N_8880,N_7627);
and U9008 (N_9008,N_7844,N_7674);
xor U9009 (N_9009,N_8046,N_8398);
nor U9010 (N_9010,N_8977,N_8133);
and U9011 (N_9011,N_7571,N_8170);
and U9012 (N_9012,N_8440,N_7561);
and U9013 (N_9013,N_7541,N_8273);
xnor U9014 (N_9014,N_8647,N_7800);
xor U9015 (N_9015,N_8569,N_8475);
or U9016 (N_9016,N_8294,N_8684);
xor U9017 (N_9017,N_8915,N_8137);
nor U9018 (N_9018,N_8856,N_7679);
nor U9019 (N_9019,N_8733,N_8819);
or U9020 (N_9020,N_7897,N_7756);
and U9021 (N_9021,N_8750,N_7748);
and U9022 (N_9022,N_7849,N_8797);
or U9023 (N_9023,N_7799,N_8091);
xnor U9024 (N_9024,N_7514,N_7696);
nor U9025 (N_9025,N_8051,N_8575);
nor U9026 (N_9026,N_8512,N_8337);
or U9027 (N_9027,N_8914,N_8140);
nor U9028 (N_9028,N_8911,N_8672);
and U9029 (N_9029,N_8480,N_8762);
or U9030 (N_9030,N_7763,N_8279);
or U9031 (N_9031,N_7681,N_8526);
xor U9032 (N_9032,N_7770,N_8773);
xor U9033 (N_9033,N_8820,N_7911);
and U9034 (N_9034,N_8686,N_8678);
and U9035 (N_9035,N_8290,N_8844);
and U9036 (N_9036,N_7961,N_8543);
or U9037 (N_9037,N_7948,N_8607);
nor U9038 (N_9038,N_8461,N_7537);
xnor U9039 (N_9039,N_8782,N_7666);
and U9040 (N_9040,N_8740,N_8642);
and U9041 (N_9041,N_7869,N_8434);
nand U9042 (N_9042,N_8587,N_8809);
nor U9043 (N_9043,N_8816,N_8921);
and U9044 (N_9044,N_8136,N_8522);
or U9045 (N_9045,N_8549,N_8961);
nor U9046 (N_9046,N_7927,N_8084);
or U9047 (N_9047,N_8511,N_8793);
nand U9048 (N_9048,N_7675,N_7944);
nand U9049 (N_9049,N_8690,N_8808);
nand U9050 (N_9050,N_8324,N_8747);
and U9051 (N_9051,N_8426,N_7735);
and U9052 (N_9052,N_7881,N_7736);
xnor U9053 (N_9053,N_8547,N_8601);
and U9054 (N_9054,N_7823,N_7802);
nand U9055 (N_9055,N_8149,N_8244);
nor U9056 (N_9056,N_7574,N_8253);
xor U9057 (N_9057,N_7996,N_8383);
nor U9058 (N_9058,N_8008,N_7812);
or U9059 (N_9059,N_7724,N_8414);
nor U9060 (N_9060,N_8577,N_8363);
nand U9061 (N_9061,N_8075,N_8318);
nand U9062 (N_9062,N_8882,N_7580);
nand U9063 (N_9063,N_8377,N_8720);
or U9064 (N_9064,N_7762,N_8757);
or U9065 (N_9065,N_7884,N_7865);
and U9066 (N_9066,N_8218,N_8934);
nand U9067 (N_9067,N_7538,N_7781);
nor U9068 (N_9068,N_8506,N_8903);
or U9069 (N_9069,N_7941,N_7749);
and U9070 (N_9070,N_8216,N_7525);
nand U9071 (N_9071,N_8109,N_8291);
xor U9072 (N_9072,N_8852,N_7755);
and U9073 (N_9073,N_7728,N_8286);
and U9074 (N_9074,N_7693,N_7792);
nand U9075 (N_9075,N_8834,N_7654);
xor U9076 (N_9076,N_7786,N_7940);
or U9077 (N_9077,N_8950,N_8194);
xor U9078 (N_9078,N_8765,N_8894);
or U9079 (N_9079,N_8272,N_8325);
nand U9080 (N_9080,N_7533,N_8764);
xor U9081 (N_9081,N_7874,N_7650);
nor U9082 (N_9082,N_7697,N_8251);
nor U9083 (N_9083,N_8261,N_8004);
or U9084 (N_9084,N_8925,N_8312);
nor U9085 (N_9085,N_8789,N_7958);
nand U9086 (N_9086,N_8567,N_8270);
xor U9087 (N_9087,N_8357,N_8323);
and U9088 (N_9088,N_8725,N_8947);
or U9089 (N_9089,N_7831,N_8722);
and U9090 (N_9090,N_7867,N_8496);
or U9091 (N_9091,N_8717,N_8959);
xor U9092 (N_9092,N_7935,N_7767);
xnor U9093 (N_9093,N_7742,N_8365);
xnor U9094 (N_9094,N_8088,N_8835);
nor U9095 (N_9095,N_8016,N_8281);
nor U9096 (N_9096,N_8192,N_8166);
or U9097 (N_9097,N_8104,N_8516);
and U9098 (N_9098,N_8813,N_8002);
nor U9099 (N_9099,N_7965,N_8085);
or U9100 (N_9100,N_8862,N_8198);
nor U9101 (N_9101,N_8157,N_8126);
xor U9102 (N_9102,N_8560,N_8850);
xor U9103 (N_9103,N_8268,N_8451);
and U9104 (N_9104,N_8050,N_7818);
and U9105 (N_9105,N_8580,N_7511);
or U9106 (N_9106,N_7592,N_8349);
nor U9107 (N_9107,N_7885,N_7597);
nor U9108 (N_9108,N_7853,N_8040);
nor U9109 (N_9109,N_8299,N_8769);
xnor U9110 (N_9110,N_7698,N_8129);
nor U9111 (N_9111,N_8909,N_8645);
nand U9112 (N_9112,N_8651,N_8558);
xor U9113 (N_9113,N_7840,N_8112);
or U9114 (N_9114,N_8207,N_7783);
xor U9115 (N_9115,N_8732,N_8228);
or U9116 (N_9116,N_8848,N_8308);
nor U9117 (N_9117,N_7512,N_8276);
nand U9118 (N_9118,N_8726,N_8083);
nand U9119 (N_9119,N_8252,N_7531);
nor U9120 (N_9120,N_8231,N_8529);
and U9121 (N_9121,N_8095,N_7667);
xor U9122 (N_9122,N_8055,N_8379);
and U9123 (N_9123,N_8156,N_8185);
xor U9124 (N_9124,N_8641,N_7707);
xor U9125 (N_9125,N_8518,N_8763);
or U9126 (N_9126,N_8135,N_8067);
xor U9127 (N_9127,N_8904,N_8869);
nand U9128 (N_9128,N_8910,N_8173);
xor U9129 (N_9129,N_8593,N_7968);
nand U9130 (N_9130,N_8791,N_8130);
and U9131 (N_9131,N_8954,N_8553);
xnor U9132 (N_9132,N_7590,N_8982);
nand U9133 (N_9133,N_8563,N_8366);
nor U9134 (N_9134,N_8145,N_8396);
xor U9135 (N_9135,N_7662,N_7625);
xnor U9136 (N_9136,N_8650,N_7851);
xor U9137 (N_9137,N_8627,N_7551);
nand U9138 (N_9138,N_8502,N_8939);
nor U9139 (N_9139,N_8892,N_8917);
xnor U9140 (N_9140,N_8952,N_8468);
or U9141 (N_9141,N_8515,N_7753);
xnor U9142 (N_9142,N_8096,N_7855);
xor U9143 (N_9143,N_8680,N_7955);
or U9144 (N_9144,N_7578,N_8825);
xnor U9145 (N_9145,N_7614,N_8221);
and U9146 (N_9146,N_7774,N_8519);
or U9147 (N_9147,N_7655,N_7761);
and U9148 (N_9148,N_8940,N_8382);
xor U9149 (N_9149,N_7923,N_8989);
and U9150 (N_9150,N_8744,N_7782);
or U9151 (N_9151,N_8566,N_7673);
or U9152 (N_9152,N_7685,N_8146);
or U9153 (N_9153,N_8527,N_7563);
xor U9154 (N_9154,N_7721,N_8184);
nor U9155 (N_9155,N_8668,N_7622);
nor U9156 (N_9156,N_8018,N_8230);
and U9157 (N_9157,N_7604,N_7631);
xor U9158 (N_9158,N_8817,N_8235);
nand U9159 (N_9159,N_7913,N_8304);
or U9160 (N_9160,N_8333,N_8514);
nor U9161 (N_9161,N_8435,N_8520);
or U9162 (N_9162,N_7956,N_8760);
nand U9163 (N_9163,N_8009,N_8854);
nor U9164 (N_9164,N_8634,N_7539);
nand U9165 (N_9165,N_7505,N_8043);
or U9166 (N_9166,N_7513,N_7569);
nor U9167 (N_9167,N_7630,N_8079);
and U9168 (N_9168,N_8024,N_7718);
or U9169 (N_9169,N_7854,N_8759);
and U9170 (N_9170,N_8080,N_7725);
and U9171 (N_9171,N_8188,N_8618);
nand U9172 (N_9172,N_8070,N_8661);
xor U9173 (N_9173,N_7745,N_8362);
nand U9174 (N_9174,N_8846,N_8479);
xnor U9175 (N_9175,N_8073,N_8005);
and U9176 (N_9176,N_8400,N_8222);
nor U9177 (N_9177,N_8197,N_8913);
or U9178 (N_9178,N_8795,N_8658);
and U9179 (N_9179,N_8017,N_8905);
or U9180 (N_9180,N_8169,N_8983);
xor U9181 (N_9181,N_7572,N_8422);
and U9182 (N_9182,N_8738,N_8855);
nand U9183 (N_9183,N_8219,N_8403);
nand U9184 (N_9184,N_7902,N_8102);
xnor U9185 (N_9185,N_7652,N_8978);
and U9186 (N_9186,N_8237,N_7757);
nor U9187 (N_9187,N_8401,N_7723);
xor U9188 (N_9188,N_7967,N_8491);
or U9189 (N_9189,N_8701,N_7957);
and U9190 (N_9190,N_8597,N_8500);
or U9191 (N_9191,N_8867,N_7586);
xnor U9192 (N_9192,N_8388,N_8614);
or U9193 (N_9193,N_8837,N_7752);
nand U9194 (N_9194,N_8545,N_8444);
nand U9195 (N_9195,N_8162,N_7637);
nand U9196 (N_9196,N_7613,N_7676);
nand U9197 (N_9197,N_8920,N_8001);
nor U9198 (N_9198,N_8035,N_7889);
and U9199 (N_9199,N_8739,N_8250);
nand U9200 (N_9200,N_7678,N_8014);
nor U9201 (N_9201,N_8257,N_8041);
nor U9202 (N_9202,N_8537,N_8639);
nor U9203 (N_9203,N_8822,N_8469);
xnor U9204 (N_9204,N_7908,N_8420);
nand U9205 (N_9205,N_8624,N_8840);
or U9206 (N_9206,N_8929,N_8196);
and U9207 (N_9207,N_7542,N_8699);
xor U9208 (N_9208,N_7960,N_7909);
and U9209 (N_9209,N_7722,N_8153);
and U9210 (N_9210,N_7704,N_7937);
nor U9211 (N_9211,N_8212,N_8175);
and U9212 (N_9212,N_7875,N_7779);
or U9213 (N_9213,N_7611,N_7553);
nand U9214 (N_9214,N_8182,N_8234);
xnor U9215 (N_9215,N_7915,N_8359);
or U9216 (N_9216,N_7953,N_8742);
or U9217 (N_9217,N_7835,N_7547);
or U9218 (N_9218,N_8829,N_8360);
nand U9219 (N_9219,N_7747,N_7608);
nor U9220 (N_9220,N_7978,N_7946);
nor U9221 (N_9221,N_7609,N_8478);
and U9222 (N_9222,N_8408,N_8441);
and U9223 (N_9223,N_8761,N_7558);
nand U9224 (N_9224,N_8926,N_8991);
xor U9225 (N_9225,N_8698,N_8554);
xnor U9226 (N_9226,N_7519,N_7585);
or U9227 (N_9227,N_7933,N_8011);
and U9228 (N_9228,N_7975,N_8147);
nand U9229 (N_9229,N_8199,N_8373);
nand U9230 (N_9230,N_7936,N_7841);
or U9231 (N_9231,N_8657,N_8729);
nor U9232 (N_9232,N_8395,N_8372);
or U9233 (N_9233,N_8332,N_8280);
or U9234 (N_9234,N_7938,N_8524);
nor U9235 (N_9235,N_8038,N_7529);
nand U9236 (N_9236,N_8633,N_8893);
and U9237 (N_9237,N_8881,N_8833);
xnor U9238 (N_9238,N_8301,N_7887);
nand U9239 (N_9239,N_7890,N_7963);
or U9240 (N_9240,N_7738,N_8531);
nand U9241 (N_9241,N_8066,N_7924);
xor U9242 (N_9242,N_8223,N_8314);
nand U9243 (N_9243,N_8159,N_7508);
nor U9244 (N_9244,N_8510,N_8667);
and U9245 (N_9245,N_8836,N_7517);
or U9246 (N_9246,N_8802,N_8858);
nand U9247 (N_9247,N_8239,N_8433);
or U9248 (N_9248,N_7570,N_8417);
and U9249 (N_9249,N_8081,N_7751);
xor U9250 (N_9250,N_8955,N_8517);
and U9251 (N_9251,N_8736,N_8564);
nor U9252 (N_9252,N_8203,N_7651);
xor U9253 (N_9253,N_8671,N_7832);
nand U9254 (N_9254,N_8805,N_8151);
or U9255 (N_9255,N_8709,N_7863);
xnor U9256 (N_9256,N_8509,N_8631);
or U9257 (N_9257,N_8148,N_8064);
nor U9258 (N_9258,N_8540,N_7646);
nor U9259 (N_9259,N_8338,N_8505);
nand U9260 (N_9260,N_7601,N_8924);
or U9261 (N_9261,N_7600,N_8985);
nand U9262 (N_9262,N_7907,N_7997);
and U9263 (N_9263,N_7794,N_8056);
or U9264 (N_9264,N_8503,N_7943);
nor U9265 (N_9265,N_7916,N_7573);
nor U9266 (N_9266,N_8020,N_7871);
or U9267 (N_9267,N_7862,N_8226);
and U9268 (N_9268,N_8656,N_7746);
or U9269 (N_9269,N_7606,N_8895);
and U9270 (N_9270,N_7828,N_8603);
xnor U9271 (N_9271,N_8027,N_7929);
and U9272 (N_9272,N_8107,N_8225);
or U9273 (N_9273,N_8958,N_7983);
and U9274 (N_9274,N_8785,N_7920);
and U9275 (N_9275,N_7554,N_8437);
xnor U9276 (N_9276,N_8679,N_7641);
nor U9277 (N_9277,N_7521,N_7820);
or U9278 (N_9278,N_8625,N_7649);
nand U9279 (N_9279,N_7977,N_8240);
nor U9280 (N_9280,N_8715,N_8103);
nor U9281 (N_9281,N_7535,N_8800);
and U9282 (N_9282,N_8346,N_7526);
nor U9283 (N_9283,N_8048,N_8779);
or U9284 (N_9284,N_8898,N_8692);
or U9285 (N_9285,N_7833,N_8158);
xnor U9286 (N_9286,N_7550,N_8556);
nor U9287 (N_9287,N_8853,N_8421);
xnor U9288 (N_9288,N_7502,N_7717);
xor U9289 (N_9289,N_7804,N_7733);
or U9290 (N_9290,N_8777,N_7981);
nand U9291 (N_9291,N_8908,N_8849);
or U9292 (N_9292,N_8968,N_8187);
or U9293 (N_9293,N_8755,N_8675);
or U9294 (N_9294,N_8052,N_8155);
nor U9295 (N_9295,N_8964,N_8447);
nand U9296 (N_9296,N_8248,N_7633);
nor U9297 (N_9297,N_8013,N_8271);
xor U9298 (N_9298,N_8878,N_8034);
nor U9299 (N_9299,N_8786,N_8695);
or U9300 (N_9300,N_7877,N_8758);
or U9301 (N_9301,N_7599,N_7626);
or U9302 (N_9302,N_8003,N_7653);
and U9303 (N_9303,N_7805,N_8328);
nor U9304 (N_9304,N_7524,N_8264);
xor U9305 (N_9305,N_8037,N_8347);
nor U9306 (N_9306,N_8063,N_8242);
and U9307 (N_9307,N_7669,N_8093);
nand U9308 (N_9308,N_8811,N_8458);
nand U9309 (N_9309,N_8443,N_8967);
nor U9310 (N_9310,N_7703,N_8453);
or U9311 (N_9311,N_8442,N_8106);
and U9312 (N_9312,N_7509,N_8766);
nand U9313 (N_9313,N_8306,N_8774);
nand U9314 (N_9314,N_7711,N_7584);
nand U9315 (N_9315,N_8288,N_8718);
and U9316 (N_9316,N_7565,N_8439);
or U9317 (N_9317,N_8044,N_7719);
nor U9318 (N_9318,N_7971,N_8352);
and U9319 (N_9319,N_8380,N_8945);
xor U9320 (N_9320,N_8525,N_7917);
and U9321 (N_9321,N_8142,N_8803);
or U9322 (N_9322,N_8781,N_8019);
and U9323 (N_9323,N_8429,N_7817);
xnor U9324 (N_9324,N_7684,N_7620);
and U9325 (N_9325,N_8128,N_8857);
nor U9326 (N_9326,N_8392,N_7951);
nor U9327 (N_9327,N_7821,N_8074);
nor U9328 (N_9328,N_7836,N_8931);
xor U9329 (N_9329,N_8445,N_8605);
nand U9330 (N_9330,N_8416,N_8042);
xor U9331 (N_9331,N_7990,N_8704);
xor U9332 (N_9332,N_8410,N_8277);
or U9333 (N_9333,N_8399,N_8804);
xnor U9334 (N_9334,N_8204,N_7589);
xor U9335 (N_9335,N_8665,N_7824);
or U9336 (N_9336,N_7772,N_8600);
nand U9337 (N_9337,N_8381,N_8694);
nor U9338 (N_9338,N_8935,N_8007);
nor U9339 (N_9339,N_8201,N_8211);
or U9340 (N_9340,N_8648,N_7921);
nand U9341 (N_9341,N_8462,N_8713);
nor U9342 (N_9342,N_8430,N_8446);
xnor U9343 (N_9343,N_7618,N_8523);
nor U9344 (N_9344,N_7577,N_8161);
xor U9345 (N_9345,N_8636,N_8590);
or U9346 (N_9346,N_7617,N_7901);
xnor U9347 (N_9347,N_8812,N_8472);
nand U9348 (N_9348,N_8144,N_8743);
and U9349 (N_9349,N_7857,N_7516);
nor U9350 (N_9350,N_7788,N_8942);
xnor U9351 (N_9351,N_7560,N_8615);
nand U9352 (N_9352,N_8351,N_8229);
and U9353 (N_9353,N_7880,N_7744);
nand U9354 (N_9354,N_8899,N_8452);
nor U9355 (N_9355,N_8374,N_8859);
xnor U9356 (N_9356,N_7769,N_8266);
nor U9357 (N_9357,N_8449,N_7904);
xnor U9358 (N_9358,N_7632,N_8981);
xor U9359 (N_9359,N_8190,N_7985);
nand U9360 (N_9360,N_7891,N_8330);
xor U9361 (N_9361,N_8975,N_8623);
and U9362 (N_9362,N_7966,N_8206);
nand U9363 (N_9363,N_8721,N_7979);
xnor U9364 (N_9364,N_7730,N_8616);
xnor U9365 (N_9365,N_8045,N_8053);
nand U9366 (N_9366,N_8866,N_8404);
nand U9367 (N_9367,N_8233,N_8711);
and U9368 (N_9368,N_7830,N_8501);
nand U9369 (N_9369,N_7939,N_7850);
and U9370 (N_9370,N_8393,N_7647);
xnor U9371 (N_9371,N_7713,N_7665);
nand U9372 (N_9372,N_8387,N_7528);
nand U9373 (N_9373,N_8585,N_8719);
nand U9374 (N_9374,N_7648,N_8303);
xnor U9375 (N_9375,N_7540,N_8415);
or U9376 (N_9376,N_8326,N_7795);
nand U9377 (N_9377,N_7995,N_8630);
nor U9378 (N_9378,N_7546,N_7635);
nand U9379 (N_9379,N_8541,N_8431);
nor U9380 (N_9380,N_7670,N_8652);
xnor U9381 (N_9381,N_8928,N_8728);
or U9382 (N_9382,N_8824,N_7822);
and U9383 (N_9383,N_7544,N_8171);
xor U9384 (N_9384,N_7692,N_8214);
nand U9385 (N_9385,N_8141,N_8573);
and U9386 (N_9386,N_8730,N_7700);
and U9387 (N_9387,N_7623,N_8487);
and U9388 (N_9388,N_7741,N_8492);
and U9389 (N_9389,N_8953,N_7798);
xor U9390 (N_9390,N_7643,N_8973);
nand U9391 (N_9391,N_8464,N_8823);
and U9392 (N_9392,N_7624,N_7559);
xnor U9393 (N_9393,N_7825,N_8300);
or U9394 (N_9394,N_8448,N_8960);
nor U9395 (N_9395,N_8342,N_8310);
xnor U9396 (N_9396,N_7743,N_8267);
nand U9397 (N_9397,N_8714,N_8845);
nor U9398 (N_9398,N_7500,N_8406);
or U9399 (N_9399,N_8653,N_8937);
xor U9400 (N_9400,N_7843,N_8168);
or U9401 (N_9401,N_8613,N_8912);
or U9402 (N_9402,N_8193,N_8598);
xor U9403 (N_9403,N_8473,N_8205);
nand U9404 (N_9404,N_8897,N_7846);
nor U9405 (N_9405,N_8274,N_8154);
nor U9406 (N_9406,N_8317,N_8655);
nand U9407 (N_9407,N_7898,N_7686);
xor U9408 (N_9408,N_8122,N_8643);
and U9409 (N_9409,N_8990,N_8980);
and U9410 (N_9410,N_7878,N_8476);
nor U9411 (N_9411,N_8322,N_8389);
xor U9412 (N_9412,N_8532,N_8535);
nand U9413 (N_9413,N_7612,N_8423);
xor U9414 (N_9414,N_8710,N_8504);
nor U9415 (N_9415,N_8456,N_7702);
nand U9416 (N_9416,N_8936,N_8427);
and U9417 (N_9417,N_7720,N_7950);
nor U9418 (N_9418,N_7709,N_7972);
and U9419 (N_9419,N_8681,N_7914);
nand U9420 (N_9420,N_7727,N_7510);
nand U9421 (N_9421,N_8565,N_7656);
or U9422 (N_9422,N_7912,N_8798);
nand U9423 (N_9423,N_8467,N_8930);
xor U9424 (N_9424,N_8818,N_8588);
nor U9425 (N_9425,N_7789,N_8375);
nand U9426 (N_9426,N_7954,N_7664);
xor U9427 (N_9427,N_7785,N_8831);
or U9428 (N_9428,N_8873,N_8622);
or U9429 (N_9429,N_8489,N_8999);
xor U9430 (N_9430,N_7715,N_8599);
nor U9431 (N_9431,N_8200,N_8341);
nand U9432 (N_9432,N_8006,N_7731);
nand U9433 (N_9433,N_7910,N_8794);
or U9434 (N_9434,N_8485,N_8238);
or U9435 (N_9435,N_7861,N_8246);
nor U9436 (N_9436,N_8963,N_8249);
and U9437 (N_9437,N_7811,N_8883);
xnor U9438 (N_9438,N_8696,N_7903);
and U9439 (N_9439,N_7932,N_8413);
nor U9440 (N_9440,N_7587,N_8863);
xor U9441 (N_9441,N_7919,N_8499);
nor U9442 (N_9442,N_8886,N_8176);
xnor U9443 (N_9443,N_7900,N_8775);
xor U9444 (N_9444,N_7708,N_8570);
or U9445 (N_9445,N_8646,N_7754);
or U9446 (N_9446,N_7661,N_8108);
xor U9447 (N_9447,N_8402,N_8315);
nand U9448 (N_9448,N_7668,N_8123);
and U9449 (N_9449,N_8425,N_8748);
nor U9450 (N_9450,N_8832,N_8640);
nor U9451 (N_9451,N_8896,N_7806);
or U9452 (N_9452,N_8689,N_8183);
nand U9453 (N_9453,N_7712,N_8311);
nand U9454 (N_9454,N_8023,N_8944);
xor U9455 (N_9455,N_8345,N_8984);
nor U9456 (N_9456,N_7596,N_8029);
nand U9457 (N_9457,N_8305,N_8932);
nor U9458 (N_9458,N_8971,N_8826);
xor U9459 (N_9459,N_8807,N_8993);
nor U9460 (N_9460,N_7575,N_7866);
nand U9461 (N_9461,N_8484,N_8436);
nand U9462 (N_9462,N_8581,N_8787);
or U9463 (N_9463,N_8576,N_7530);
nand U9464 (N_9464,N_7964,N_8716);
or U9465 (N_9465,N_8282,N_7706);
nor U9466 (N_9466,N_7607,N_8179);
nor U9467 (N_9467,N_8355,N_7998);
xnor U9468 (N_9468,N_8210,N_8877);
nor U9469 (N_9469,N_8327,N_8181);
or U9470 (N_9470,N_8788,N_8965);
or U9471 (N_9471,N_7628,N_8058);
xnor U9472 (N_9472,N_8778,N_8997);
and U9473 (N_9473,N_8087,N_7549);
or U9474 (N_9474,N_8927,N_8839);
xor U9475 (N_9475,N_8700,N_7520);
nor U9476 (N_9476,N_7899,N_8608);
nand U9477 (N_9477,N_7598,N_7845);
and U9478 (N_9478,N_8674,N_8702);
and U9479 (N_9479,N_8049,N_8933);
nor U9480 (N_9480,N_8298,N_8247);
nand U9481 (N_9481,N_8293,N_8466);
or U9482 (N_9482,N_8806,N_7922);
nand U9483 (N_9483,N_7882,N_7839);
or U9484 (N_9484,N_7615,N_8586);
or U9485 (N_9485,N_8285,N_8028);
or U9486 (N_9486,N_8054,N_8707);
nor U9487 (N_9487,N_8497,N_8113);
xnor U9488 (N_9488,N_7816,N_7532);
nand U9489 (N_9489,N_8255,N_8772);
xor U9490 (N_9490,N_7994,N_7988);
nor U9491 (N_9491,N_8068,N_8870);
and U9492 (N_9492,N_8364,N_8987);
nor U9493 (N_9493,N_7543,N_8691);
and U9494 (N_9494,N_8477,N_7888);
nand U9495 (N_9495,N_8098,N_8801);
xor U9496 (N_9496,N_8884,N_7689);
nand U9497 (N_9497,N_7945,N_8574);
xnor U9498 (N_9498,N_7659,N_8589);
nor U9499 (N_9499,N_7567,N_7758);
or U9500 (N_9500,N_7619,N_7581);
nor U9501 (N_9501,N_8089,N_8891);
xor U9502 (N_9502,N_8284,N_7644);
and U9503 (N_9503,N_8872,N_7974);
or U9504 (N_9504,N_7829,N_8262);
nand U9505 (N_9505,N_8010,N_8637);
nor U9506 (N_9506,N_7773,N_8026);
xor U9507 (N_9507,N_7694,N_8705);
and U9508 (N_9508,N_8974,N_8557);
nor U9509 (N_9509,N_8507,N_8213);
xor U9510 (N_9510,N_7959,N_8916);
or U9511 (N_9511,N_7942,N_8751);
nor U9512 (N_9512,N_8482,N_8919);
and U9513 (N_9513,N_8114,N_8568);
nor U9514 (N_9514,N_8097,N_8457);
xnor U9515 (N_9515,N_8343,N_8941);
nand U9516 (N_9516,N_7507,N_8998);
nor U9517 (N_9517,N_8796,N_7864);
xor U9518 (N_9518,N_8612,N_8923);
xor U9519 (N_9519,N_8687,N_8992);
xnor U9520 (N_9520,N_8731,N_8583);
and U9521 (N_9521,N_8508,N_8358);
or U9522 (N_9522,N_7928,N_8888);
nor U9523 (N_9523,N_8956,N_8948);
nor U9524 (N_9524,N_8160,N_7699);
or U9525 (N_9525,N_8619,N_8178);
nand U9526 (N_9526,N_8768,N_8712);
nor U9527 (N_9527,N_7847,N_8092);
xor U9528 (N_9528,N_8208,N_8459);
and U9529 (N_9529,N_7583,N_8970);
and U9530 (N_9530,N_7695,N_7992);
and U9531 (N_9531,N_7886,N_7645);
nor U9532 (N_9532,N_8030,N_7701);
or U9533 (N_9533,N_7791,N_7732);
nor U9534 (N_9534,N_8180,N_8031);
nor U9535 (N_9535,N_7796,N_7784);
nand U9536 (N_9536,N_8295,N_8076);
or U9537 (N_9537,N_7595,N_8313);
and U9538 (N_9538,N_8594,N_7568);
nand U9539 (N_9539,N_8683,N_8943);
and U9540 (N_9540,N_8629,N_7895);
xnor U9541 (N_9541,N_8538,N_7737);
or U9542 (N_9542,N_8724,N_8125);
xnor U9543 (N_9543,N_7765,N_8438);
or U9544 (N_9544,N_7970,N_8174);
xor U9545 (N_9545,N_8059,N_8376);
xnor U9546 (N_9546,N_8450,N_8117);
or U9547 (N_9547,N_8561,N_7582);
nand U9548 (N_9548,N_7973,N_8138);
and U9549 (N_9549,N_8749,N_8348);
nand U9550 (N_9550,N_8039,N_8077);
or U9551 (N_9551,N_8617,N_7787);
and U9552 (N_9552,N_8810,N_7671);
nor U9553 (N_9553,N_8127,N_8022);
or U9554 (N_9554,N_8843,N_8688);
nand U9555 (N_9555,N_8105,N_7603);
nand U9556 (N_9556,N_7848,N_8021);
xor U9557 (N_9557,N_8409,N_7677);
nor U9558 (N_9558,N_8771,N_8697);
nor U9559 (N_9559,N_7726,N_8132);
and U9560 (N_9560,N_8792,N_8596);
and U9561 (N_9561,N_8745,N_8195);
or U9562 (N_9562,N_8134,N_8163);
and U9563 (N_9563,N_8094,N_8165);
or U9564 (N_9564,N_8670,N_7790);
nand U9565 (N_9565,N_8783,N_8120);
nand U9566 (N_9566,N_7518,N_8790);
nor U9567 (N_9567,N_7993,N_8685);
or U9568 (N_9568,N_8033,N_7989);
and U9569 (N_9569,N_7777,N_8302);
nor U9570 (N_9570,N_8000,N_8591);
nand U9571 (N_9571,N_8498,N_7638);
and U9572 (N_9572,N_8386,N_8407);
nor U9573 (N_9573,N_8620,N_8542);
nand U9574 (N_9574,N_8258,N_8259);
xnor U9575 (N_9575,N_8065,N_7949);
nand U9576 (N_9576,N_7610,N_8962);
nand U9577 (N_9577,N_8546,N_8994);
and U9578 (N_9578,N_8842,N_8536);
or U9579 (N_9579,N_7771,N_8951);
nor U9580 (N_9580,N_7984,N_8036);
nand U9581 (N_9581,N_8465,N_8815);
and U9582 (N_9582,N_7602,N_7760);
nor U9583 (N_9583,N_7534,N_8283);
or U9584 (N_9584,N_8032,N_8224);
and U9585 (N_9585,N_8390,N_8186);
nor U9586 (N_9586,N_8101,N_8753);
nand U9587 (N_9587,N_7976,N_7527);
and U9588 (N_9588,N_7892,N_8493);
xor U9589 (N_9589,N_7872,N_7688);
nand U9590 (N_9590,N_8544,N_8432);
nor U9591 (N_9591,N_8394,N_8734);
or U9592 (N_9592,N_8256,N_7594);
xnor U9593 (N_9593,N_7780,N_7766);
or U9594 (N_9594,N_7672,N_8918);
nor U9595 (N_9595,N_8397,N_7893);
xnor U9596 (N_9596,N_8676,N_8938);
or U9597 (N_9597,N_8307,N_7687);
nor U9598 (N_9598,N_7819,N_8061);
nand U9599 (N_9599,N_8189,N_7750);
nor U9600 (N_9600,N_8118,N_7883);
nand U9601 (N_9601,N_8900,N_8865);
nand U9602 (N_9602,N_8350,N_8828);
or U9603 (N_9603,N_7579,N_8289);
or U9604 (N_9604,N_8976,N_7710);
nor U9605 (N_9605,N_8770,N_7815);
and U9606 (N_9606,N_8405,N_7634);
xnor U9607 (N_9607,N_8334,N_7962);
nand U9608 (N_9608,N_7803,N_7555);
nor U9609 (N_9609,N_8682,N_8419);
nand U9610 (N_9610,N_8551,N_7856);
or U9611 (N_9611,N_7860,N_7797);
and U9612 (N_9612,N_8703,N_8610);
or U9613 (N_9613,N_7729,N_8669);
xnor U9614 (N_9614,N_8602,N_8552);
nor U9615 (N_9615,N_8604,N_8340);
and U9616 (N_9616,N_8490,N_8767);
nor U9617 (N_9617,N_8821,N_8628);
nand U9618 (N_9618,N_7764,N_7657);
and U9619 (N_9619,N_8784,N_8548);
nor U9620 (N_9620,N_7683,N_8539);
nand U9621 (N_9621,N_8638,N_8331);
and U9622 (N_9622,N_8470,N_8411);
xnor U9623 (N_9623,N_8606,N_8996);
nand U9624 (N_9624,N_8245,N_8582);
or U9625 (N_9625,N_8874,N_8115);
and U9626 (N_9626,N_8335,N_8609);
nor U9627 (N_9627,N_7931,N_7776);
nand U9628 (N_9628,N_7768,N_8143);
and U9629 (N_9629,N_7640,N_8116);
or U9630 (N_9630,N_8412,N_8172);
or U9631 (N_9631,N_7739,N_8460);
nand U9632 (N_9632,N_8799,N_8885);
nand U9633 (N_9633,N_8015,N_8868);
nand U9634 (N_9634,N_7576,N_8995);
or U9635 (N_9635,N_8025,N_7982);
or U9636 (N_9636,N_8654,N_8579);
or U9637 (N_9637,N_8889,N_8369);
or U9638 (N_9638,N_8693,N_7552);
nand U9639 (N_9639,N_8191,N_8746);
nand U9640 (N_9640,N_7999,N_8111);
or U9641 (N_9641,N_8428,N_8265);
and U9642 (N_9642,N_8528,N_8887);
nand U9643 (N_9643,N_7807,N_7591);
xor U9644 (N_9644,N_7536,N_7837);
and U9645 (N_9645,N_8861,N_7548);
and U9646 (N_9646,N_8534,N_7894);
and U9647 (N_9647,N_8319,N_7663);
xor U9648 (N_9648,N_8741,N_7588);
nand U9649 (N_9649,N_7896,N_8481);
xor U9650 (N_9650,N_7564,N_7980);
xnor U9651 (N_9651,N_8901,N_8167);
nor U9652 (N_9652,N_8012,N_8152);
nand U9653 (N_9653,N_8321,N_8047);
nand U9654 (N_9654,N_8562,N_8227);
nand U9655 (N_9655,N_8278,N_8424);
nor U9656 (N_9656,N_7879,N_7801);
xor U9657 (N_9657,N_8780,N_8361);
or U9658 (N_9658,N_7952,N_8592);
xnor U9659 (N_9659,N_8875,N_7682);
and U9660 (N_9660,N_7557,N_8296);
and U9661 (N_9661,N_8418,N_8370);
nor U9662 (N_9662,N_7504,N_8217);
and U9663 (N_9663,N_7566,N_8486);
nor U9664 (N_9664,N_8907,N_7876);
or U9665 (N_9665,N_8241,N_7969);
xor U9666 (N_9666,N_8356,N_7947);
and U9667 (N_9667,N_8287,N_8090);
or U9668 (N_9668,N_8336,N_8595);
nor U9669 (N_9669,N_7501,N_8215);
or U9670 (N_9670,N_8354,N_8814);
and U9671 (N_9671,N_8071,N_8673);
nand U9672 (N_9672,N_8644,N_8635);
xnor U9673 (N_9673,N_8320,N_7842);
nor U9674 (N_9674,N_8578,N_8474);
or U9675 (N_9675,N_7926,N_8062);
nand U9676 (N_9676,N_7515,N_7714);
xor U9677 (N_9677,N_7834,N_7905);
nand U9678 (N_9678,N_7859,N_7868);
nand U9679 (N_9679,N_8384,N_7987);
xnor U9680 (N_9680,N_8371,N_7852);
and U9681 (N_9681,N_7793,N_8078);
nor U9682 (N_9682,N_8946,N_8344);
nor U9683 (N_9683,N_7813,N_7906);
nor U9684 (N_9684,N_8463,N_8150);
xnor U9685 (N_9685,N_7986,N_8530);
nor U9686 (N_9686,N_7826,N_8254);
nor U9687 (N_9687,N_8269,N_8966);
nor U9688 (N_9688,N_8876,N_8584);
xnor U9689 (N_9689,N_7605,N_7870);
or U9690 (N_9690,N_8209,N_8659);
nor U9691 (N_9691,N_7810,N_8626);
nand U9692 (N_9692,N_7658,N_8494);
or U9693 (N_9693,N_8177,N_8851);
nor U9694 (N_9694,N_7636,N_7691);
nor U9695 (N_9695,N_8297,N_8969);
xor U9696 (N_9696,N_8664,N_8708);
or U9697 (N_9697,N_8368,N_8121);
nor U9698 (N_9698,N_8455,N_8100);
and U9699 (N_9699,N_7629,N_8260);
nand U9700 (N_9700,N_8057,N_8571);
nor U9701 (N_9701,N_7858,N_8082);
and U9702 (N_9702,N_8533,N_8838);
or U9703 (N_9703,N_8139,N_7639);
nand U9704 (N_9704,N_8110,N_8660);
xor U9705 (N_9705,N_7991,N_8864);
nand U9706 (N_9706,N_8495,N_7838);
nor U9707 (N_9707,N_8072,N_8949);
and U9708 (N_9708,N_8488,N_7522);
xor U9709 (N_9709,N_8483,N_8339);
nand U9710 (N_9710,N_8202,N_7690);
and U9711 (N_9711,N_8756,N_8131);
xnor U9712 (N_9712,N_8555,N_8737);
nand U9713 (N_9713,N_8316,N_7734);
xnor U9714 (N_9714,N_8119,N_8086);
or U9715 (N_9715,N_8879,N_8471);
nor U9716 (N_9716,N_7660,N_8367);
and U9717 (N_9717,N_7827,N_8124);
nand U9718 (N_9718,N_7506,N_8972);
and U9719 (N_9719,N_8550,N_7808);
nand U9720 (N_9720,N_8666,N_7556);
nor U9721 (N_9721,N_7642,N_8232);
or U9722 (N_9722,N_8890,N_8164);
and U9723 (N_9723,N_8860,N_8988);
nand U9724 (N_9724,N_8632,N_8871);
or U9725 (N_9725,N_7925,N_7545);
nor U9726 (N_9726,N_8263,N_8847);
nand U9727 (N_9727,N_7740,N_8677);
or U9728 (N_9728,N_7562,N_7918);
nor U9729 (N_9729,N_8827,N_7616);
and U9730 (N_9730,N_8572,N_8662);
and U9731 (N_9731,N_8986,N_7930);
nand U9732 (N_9732,N_8378,N_7814);
nor U9733 (N_9733,N_7716,N_8754);
or U9734 (N_9734,N_8776,N_7809);
nor U9735 (N_9735,N_8979,N_7934);
nand U9736 (N_9736,N_8906,N_7503);
nor U9737 (N_9737,N_8735,N_8957);
or U9738 (N_9738,N_8060,N_8706);
xnor U9739 (N_9739,N_8309,N_8922);
nand U9740 (N_9740,N_8830,N_7778);
nand U9741 (N_9741,N_8727,N_8391);
nor U9742 (N_9742,N_8559,N_8841);
xnor U9743 (N_9743,N_8099,N_8649);
nor U9744 (N_9744,N_8353,N_8723);
or U9745 (N_9745,N_8292,N_8243);
xor U9746 (N_9746,N_8454,N_7621);
or U9747 (N_9747,N_8069,N_7759);
xor U9748 (N_9748,N_8902,N_8236);
and U9749 (N_9749,N_7775,N_7705);
or U9750 (N_9750,N_8534,N_8785);
nand U9751 (N_9751,N_8577,N_8499);
and U9752 (N_9752,N_7967,N_8257);
nand U9753 (N_9753,N_7718,N_8052);
xnor U9754 (N_9754,N_7917,N_8581);
xor U9755 (N_9755,N_8924,N_8199);
or U9756 (N_9756,N_7998,N_7610);
xnor U9757 (N_9757,N_7587,N_8755);
or U9758 (N_9758,N_8176,N_8548);
nor U9759 (N_9759,N_7806,N_8606);
nor U9760 (N_9760,N_8987,N_8030);
and U9761 (N_9761,N_7795,N_8668);
or U9762 (N_9762,N_8700,N_8194);
and U9763 (N_9763,N_8998,N_8461);
xor U9764 (N_9764,N_8286,N_7828);
xnor U9765 (N_9765,N_7860,N_8578);
or U9766 (N_9766,N_8732,N_8838);
xnor U9767 (N_9767,N_8456,N_8394);
nand U9768 (N_9768,N_8845,N_7562);
and U9769 (N_9769,N_8817,N_7614);
nor U9770 (N_9770,N_8736,N_7622);
nor U9771 (N_9771,N_7549,N_8578);
or U9772 (N_9772,N_7933,N_7731);
nor U9773 (N_9773,N_7699,N_7725);
or U9774 (N_9774,N_7582,N_8822);
and U9775 (N_9775,N_7501,N_7883);
xor U9776 (N_9776,N_8027,N_8014);
nor U9777 (N_9777,N_8829,N_7953);
nand U9778 (N_9778,N_7829,N_8410);
nor U9779 (N_9779,N_8650,N_7719);
nor U9780 (N_9780,N_8310,N_7781);
or U9781 (N_9781,N_7574,N_8411);
and U9782 (N_9782,N_7685,N_8882);
and U9783 (N_9783,N_8380,N_8980);
and U9784 (N_9784,N_8703,N_7650);
and U9785 (N_9785,N_8033,N_8799);
nor U9786 (N_9786,N_8379,N_8361);
nor U9787 (N_9787,N_8052,N_7994);
nor U9788 (N_9788,N_8177,N_7812);
nand U9789 (N_9789,N_8569,N_8633);
nand U9790 (N_9790,N_7580,N_8121);
or U9791 (N_9791,N_7928,N_8974);
nand U9792 (N_9792,N_8625,N_8670);
nand U9793 (N_9793,N_8146,N_8560);
nor U9794 (N_9794,N_8592,N_8365);
nand U9795 (N_9795,N_8513,N_8922);
or U9796 (N_9796,N_8462,N_8475);
nor U9797 (N_9797,N_8419,N_8561);
xor U9798 (N_9798,N_8909,N_8847);
and U9799 (N_9799,N_8091,N_8620);
and U9800 (N_9800,N_7874,N_7710);
or U9801 (N_9801,N_8870,N_8254);
xnor U9802 (N_9802,N_7613,N_7549);
and U9803 (N_9803,N_7926,N_7995);
nand U9804 (N_9804,N_8305,N_7975);
xor U9805 (N_9805,N_7648,N_8995);
nor U9806 (N_9806,N_8800,N_8789);
xnor U9807 (N_9807,N_8603,N_8341);
xor U9808 (N_9808,N_7886,N_8468);
xor U9809 (N_9809,N_7811,N_7794);
and U9810 (N_9810,N_7675,N_8506);
nor U9811 (N_9811,N_8115,N_8283);
or U9812 (N_9812,N_7637,N_7739);
xor U9813 (N_9813,N_8097,N_8257);
or U9814 (N_9814,N_8848,N_8935);
and U9815 (N_9815,N_7826,N_8403);
nor U9816 (N_9816,N_8703,N_8201);
or U9817 (N_9817,N_7559,N_8026);
or U9818 (N_9818,N_8811,N_8053);
nand U9819 (N_9819,N_8852,N_7594);
or U9820 (N_9820,N_8372,N_7838);
nand U9821 (N_9821,N_8320,N_8351);
nand U9822 (N_9822,N_7539,N_8976);
xnor U9823 (N_9823,N_8492,N_7682);
nand U9824 (N_9824,N_7994,N_8735);
and U9825 (N_9825,N_8275,N_7833);
or U9826 (N_9826,N_7668,N_8547);
nand U9827 (N_9827,N_7965,N_8237);
nand U9828 (N_9828,N_8685,N_8333);
nor U9829 (N_9829,N_8896,N_7906);
nor U9830 (N_9830,N_7766,N_8109);
xnor U9831 (N_9831,N_8402,N_8519);
nor U9832 (N_9832,N_8337,N_8862);
and U9833 (N_9833,N_8260,N_7735);
nor U9834 (N_9834,N_8710,N_8299);
or U9835 (N_9835,N_7658,N_7968);
xnor U9836 (N_9836,N_8831,N_8794);
and U9837 (N_9837,N_8644,N_7951);
or U9838 (N_9838,N_7805,N_8077);
nand U9839 (N_9839,N_7653,N_8687);
nor U9840 (N_9840,N_8424,N_8829);
xor U9841 (N_9841,N_8274,N_8412);
xor U9842 (N_9842,N_8085,N_8585);
xor U9843 (N_9843,N_8545,N_7580);
nor U9844 (N_9844,N_7783,N_8796);
nand U9845 (N_9845,N_8588,N_7958);
and U9846 (N_9846,N_8851,N_7500);
or U9847 (N_9847,N_7655,N_8506);
nor U9848 (N_9848,N_8160,N_8382);
and U9849 (N_9849,N_7621,N_7936);
xnor U9850 (N_9850,N_7811,N_8371);
or U9851 (N_9851,N_8686,N_8416);
and U9852 (N_9852,N_7996,N_8579);
nand U9853 (N_9853,N_7898,N_8079);
nor U9854 (N_9854,N_7938,N_7950);
nand U9855 (N_9855,N_7703,N_8883);
and U9856 (N_9856,N_7965,N_8460);
nor U9857 (N_9857,N_7701,N_8924);
or U9858 (N_9858,N_8973,N_7911);
xnor U9859 (N_9859,N_7558,N_8289);
xnor U9860 (N_9860,N_7676,N_8341);
nand U9861 (N_9861,N_8317,N_8793);
nor U9862 (N_9862,N_8415,N_8203);
nor U9863 (N_9863,N_8763,N_8277);
nand U9864 (N_9864,N_8276,N_8643);
nand U9865 (N_9865,N_8083,N_7780);
or U9866 (N_9866,N_7544,N_8209);
nand U9867 (N_9867,N_8210,N_7856);
or U9868 (N_9868,N_8750,N_8446);
xnor U9869 (N_9869,N_7722,N_8220);
xor U9870 (N_9870,N_7854,N_8429);
nor U9871 (N_9871,N_7540,N_8401);
nand U9872 (N_9872,N_8550,N_7832);
and U9873 (N_9873,N_8220,N_8688);
or U9874 (N_9874,N_8080,N_8865);
nand U9875 (N_9875,N_8707,N_8647);
nand U9876 (N_9876,N_8231,N_7664);
nand U9877 (N_9877,N_8583,N_8861);
and U9878 (N_9878,N_8407,N_8648);
or U9879 (N_9879,N_8297,N_8674);
xor U9880 (N_9880,N_8395,N_8568);
nand U9881 (N_9881,N_8310,N_8106);
nand U9882 (N_9882,N_8681,N_8701);
and U9883 (N_9883,N_7685,N_8476);
nand U9884 (N_9884,N_8466,N_7984);
and U9885 (N_9885,N_8137,N_8612);
and U9886 (N_9886,N_8547,N_8997);
nand U9887 (N_9887,N_8411,N_8607);
nand U9888 (N_9888,N_8936,N_7944);
and U9889 (N_9889,N_8924,N_7905);
nand U9890 (N_9890,N_8741,N_8533);
nand U9891 (N_9891,N_8421,N_7530);
and U9892 (N_9892,N_7661,N_8964);
nand U9893 (N_9893,N_7869,N_8322);
or U9894 (N_9894,N_8504,N_7984);
xor U9895 (N_9895,N_8543,N_8822);
nand U9896 (N_9896,N_7546,N_7513);
nand U9897 (N_9897,N_7708,N_8847);
xor U9898 (N_9898,N_8482,N_8738);
nor U9899 (N_9899,N_7510,N_7608);
xor U9900 (N_9900,N_8582,N_8816);
nor U9901 (N_9901,N_7668,N_8194);
nand U9902 (N_9902,N_7639,N_8565);
nand U9903 (N_9903,N_7931,N_8056);
xnor U9904 (N_9904,N_8373,N_8323);
nor U9905 (N_9905,N_7755,N_8318);
nand U9906 (N_9906,N_7651,N_7567);
and U9907 (N_9907,N_8639,N_8536);
nand U9908 (N_9908,N_7940,N_8210);
xnor U9909 (N_9909,N_8040,N_8150);
or U9910 (N_9910,N_7967,N_8062);
nor U9911 (N_9911,N_8082,N_8737);
nand U9912 (N_9912,N_8088,N_8248);
or U9913 (N_9913,N_7858,N_8941);
nor U9914 (N_9914,N_8425,N_7607);
nor U9915 (N_9915,N_7909,N_8102);
xor U9916 (N_9916,N_7639,N_8997);
or U9917 (N_9917,N_8578,N_8714);
nand U9918 (N_9918,N_8772,N_8089);
and U9919 (N_9919,N_8254,N_8203);
xor U9920 (N_9920,N_7942,N_8774);
nor U9921 (N_9921,N_7836,N_8693);
nand U9922 (N_9922,N_7595,N_8764);
nand U9923 (N_9923,N_8534,N_7975);
and U9924 (N_9924,N_7867,N_8221);
nand U9925 (N_9925,N_8924,N_8064);
or U9926 (N_9926,N_8493,N_7523);
xnor U9927 (N_9927,N_7685,N_8544);
and U9928 (N_9928,N_8216,N_8475);
nor U9929 (N_9929,N_7900,N_8706);
nand U9930 (N_9930,N_8171,N_7883);
nor U9931 (N_9931,N_8425,N_7553);
nor U9932 (N_9932,N_8224,N_8574);
xor U9933 (N_9933,N_8857,N_8880);
nand U9934 (N_9934,N_8139,N_8199);
or U9935 (N_9935,N_7608,N_7905);
xnor U9936 (N_9936,N_7806,N_8310);
nand U9937 (N_9937,N_8218,N_8830);
or U9938 (N_9938,N_8734,N_8155);
and U9939 (N_9939,N_8773,N_8809);
or U9940 (N_9940,N_8941,N_8258);
or U9941 (N_9941,N_7704,N_7552);
and U9942 (N_9942,N_8632,N_8115);
or U9943 (N_9943,N_8063,N_8177);
nand U9944 (N_9944,N_7822,N_8087);
nand U9945 (N_9945,N_8849,N_8037);
nand U9946 (N_9946,N_8324,N_7638);
or U9947 (N_9947,N_8464,N_8387);
and U9948 (N_9948,N_8858,N_7667);
or U9949 (N_9949,N_7621,N_8673);
nor U9950 (N_9950,N_7759,N_8991);
xor U9951 (N_9951,N_8832,N_8127);
nand U9952 (N_9952,N_8109,N_8305);
xnor U9953 (N_9953,N_8392,N_8191);
nand U9954 (N_9954,N_8759,N_8775);
nor U9955 (N_9955,N_7888,N_8188);
nand U9956 (N_9956,N_8570,N_7522);
nor U9957 (N_9957,N_8929,N_8230);
nand U9958 (N_9958,N_8499,N_8185);
nand U9959 (N_9959,N_8368,N_8940);
nand U9960 (N_9960,N_7696,N_8771);
xor U9961 (N_9961,N_8379,N_8511);
or U9962 (N_9962,N_8657,N_8032);
or U9963 (N_9963,N_8043,N_7837);
nand U9964 (N_9964,N_8296,N_7738);
nand U9965 (N_9965,N_8002,N_8216);
nand U9966 (N_9966,N_7920,N_7681);
xor U9967 (N_9967,N_8946,N_7942);
or U9968 (N_9968,N_7736,N_8346);
and U9969 (N_9969,N_8992,N_8229);
xor U9970 (N_9970,N_8152,N_8534);
and U9971 (N_9971,N_8077,N_7579);
or U9972 (N_9972,N_7634,N_8796);
and U9973 (N_9973,N_8651,N_8215);
xnor U9974 (N_9974,N_8559,N_8515);
or U9975 (N_9975,N_7781,N_8412);
or U9976 (N_9976,N_8999,N_8152);
nand U9977 (N_9977,N_8952,N_8985);
and U9978 (N_9978,N_8184,N_8859);
xnor U9979 (N_9979,N_7923,N_7547);
or U9980 (N_9980,N_8300,N_8964);
nand U9981 (N_9981,N_8244,N_8206);
or U9982 (N_9982,N_8821,N_8880);
and U9983 (N_9983,N_8713,N_8243);
and U9984 (N_9984,N_8981,N_8475);
nand U9985 (N_9985,N_8652,N_7619);
nor U9986 (N_9986,N_8886,N_8669);
and U9987 (N_9987,N_8977,N_7746);
nand U9988 (N_9988,N_7958,N_7587);
and U9989 (N_9989,N_8757,N_8441);
and U9990 (N_9990,N_8935,N_7733);
and U9991 (N_9991,N_8970,N_7803);
or U9992 (N_9992,N_8331,N_8420);
xor U9993 (N_9993,N_7984,N_8794);
and U9994 (N_9994,N_8493,N_7646);
or U9995 (N_9995,N_8969,N_8818);
or U9996 (N_9996,N_7634,N_8880);
nor U9997 (N_9997,N_8809,N_7770);
or U9998 (N_9998,N_7897,N_8138);
and U9999 (N_9999,N_8804,N_7927);
xnor U10000 (N_10000,N_8752,N_8323);
and U10001 (N_10001,N_7899,N_8539);
xor U10002 (N_10002,N_8497,N_8183);
nor U10003 (N_10003,N_8736,N_8914);
nor U10004 (N_10004,N_8071,N_8840);
or U10005 (N_10005,N_7567,N_8494);
nand U10006 (N_10006,N_8893,N_7870);
nor U10007 (N_10007,N_7572,N_8957);
nor U10008 (N_10008,N_7761,N_8124);
or U10009 (N_10009,N_8292,N_8198);
or U10010 (N_10010,N_7689,N_8533);
and U10011 (N_10011,N_7570,N_7592);
and U10012 (N_10012,N_8366,N_7878);
xor U10013 (N_10013,N_8336,N_8051);
or U10014 (N_10014,N_8517,N_8542);
nand U10015 (N_10015,N_7935,N_7547);
or U10016 (N_10016,N_8784,N_8326);
and U10017 (N_10017,N_8769,N_8226);
xnor U10018 (N_10018,N_8111,N_8280);
nand U10019 (N_10019,N_8961,N_8128);
nor U10020 (N_10020,N_7859,N_7995);
nor U10021 (N_10021,N_7914,N_8348);
xor U10022 (N_10022,N_7602,N_8029);
nand U10023 (N_10023,N_7533,N_8329);
nand U10024 (N_10024,N_7758,N_7717);
or U10025 (N_10025,N_7969,N_8895);
or U10026 (N_10026,N_8499,N_7758);
and U10027 (N_10027,N_8852,N_8115);
nor U10028 (N_10028,N_7861,N_8603);
nand U10029 (N_10029,N_8737,N_8203);
nand U10030 (N_10030,N_8242,N_8462);
and U10031 (N_10031,N_8804,N_7640);
nand U10032 (N_10032,N_8925,N_7691);
nand U10033 (N_10033,N_8890,N_8647);
nand U10034 (N_10034,N_8844,N_7735);
nand U10035 (N_10035,N_8441,N_7918);
nand U10036 (N_10036,N_8906,N_7698);
xnor U10037 (N_10037,N_8980,N_8417);
xnor U10038 (N_10038,N_8764,N_8342);
nor U10039 (N_10039,N_8295,N_7668);
or U10040 (N_10040,N_8374,N_7784);
and U10041 (N_10041,N_8182,N_8325);
or U10042 (N_10042,N_8581,N_7839);
nand U10043 (N_10043,N_8791,N_7825);
or U10044 (N_10044,N_8845,N_7535);
or U10045 (N_10045,N_7507,N_7981);
nor U10046 (N_10046,N_8031,N_8344);
nor U10047 (N_10047,N_7560,N_8806);
nor U10048 (N_10048,N_8115,N_8137);
nor U10049 (N_10049,N_7717,N_7622);
xnor U10050 (N_10050,N_7757,N_8474);
nand U10051 (N_10051,N_8008,N_8957);
and U10052 (N_10052,N_8955,N_8888);
and U10053 (N_10053,N_7711,N_7814);
xor U10054 (N_10054,N_8527,N_8981);
nor U10055 (N_10055,N_7733,N_8359);
and U10056 (N_10056,N_7972,N_8909);
xnor U10057 (N_10057,N_8685,N_7861);
nor U10058 (N_10058,N_8588,N_8374);
xor U10059 (N_10059,N_8631,N_7854);
or U10060 (N_10060,N_8491,N_7915);
and U10061 (N_10061,N_7726,N_7856);
nor U10062 (N_10062,N_8182,N_7907);
nand U10063 (N_10063,N_8550,N_7798);
nor U10064 (N_10064,N_7852,N_7637);
nor U10065 (N_10065,N_8335,N_8554);
xor U10066 (N_10066,N_7997,N_8928);
xor U10067 (N_10067,N_8991,N_8538);
and U10068 (N_10068,N_8911,N_8889);
nand U10069 (N_10069,N_8031,N_8643);
nor U10070 (N_10070,N_7890,N_8948);
or U10071 (N_10071,N_8735,N_8916);
nor U10072 (N_10072,N_8442,N_8685);
nand U10073 (N_10073,N_8289,N_8604);
and U10074 (N_10074,N_8057,N_7957);
xor U10075 (N_10075,N_8256,N_8953);
nor U10076 (N_10076,N_7680,N_7846);
or U10077 (N_10077,N_7581,N_8252);
nand U10078 (N_10078,N_8332,N_7675);
nand U10079 (N_10079,N_8701,N_8355);
and U10080 (N_10080,N_7765,N_8912);
nand U10081 (N_10081,N_8409,N_7930);
nand U10082 (N_10082,N_8778,N_7573);
and U10083 (N_10083,N_8990,N_8988);
and U10084 (N_10084,N_8054,N_8340);
and U10085 (N_10085,N_8611,N_8116);
nor U10086 (N_10086,N_7987,N_7562);
nor U10087 (N_10087,N_7904,N_7655);
nand U10088 (N_10088,N_8781,N_8977);
and U10089 (N_10089,N_8226,N_8664);
nand U10090 (N_10090,N_8208,N_7713);
and U10091 (N_10091,N_7865,N_8543);
nand U10092 (N_10092,N_8485,N_8793);
or U10093 (N_10093,N_7659,N_8671);
xnor U10094 (N_10094,N_8157,N_7741);
nand U10095 (N_10095,N_7868,N_8514);
and U10096 (N_10096,N_8698,N_8649);
nand U10097 (N_10097,N_8156,N_7714);
or U10098 (N_10098,N_8487,N_8398);
nand U10099 (N_10099,N_8532,N_8755);
and U10100 (N_10100,N_7635,N_7855);
or U10101 (N_10101,N_8297,N_7630);
or U10102 (N_10102,N_8999,N_8764);
or U10103 (N_10103,N_7980,N_8329);
xor U10104 (N_10104,N_7579,N_7525);
or U10105 (N_10105,N_7870,N_8366);
and U10106 (N_10106,N_7793,N_8094);
nor U10107 (N_10107,N_8776,N_7704);
nor U10108 (N_10108,N_8698,N_8283);
xor U10109 (N_10109,N_7629,N_7784);
xnor U10110 (N_10110,N_8096,N_8987);
nor U10111 (N_10111,N_8174,N_8937);
or U10112 (N_10112,N_8223,N_8769);
xnor U10113 (N_10113,N_7964,N_8895);
nand U10114 (N_10114,N_8302,N_8089);
or U10115 (N_10115,N_7621,N_8797);
nor U10116 (N_10116,N_8981,N_8234);
nand U10117 (N_10117,N_8882,N_8524);
xnor U10118 (N_10118,N_8904,N_8582);
xnor U10119 (N_10119,N_8591,N_7501);
xor U10120 (N_10120,N_7914,N_8264);
or U10121 (N_10121,N_7996,N_8574);
nand U10122 (N_10122,N_8419,N_8536);
and U10123 (N_10123,N_7711,N_7514);
and U10124 (N_10124,N_8819,N_7860);
or U10125 (N_10125,N_7725,N_7509);
nand U10126 (N_10126,N_8631,N_8427);
nor U10127 (N_10127,N_8415,N_8284);
nand U10128 (N_10128,N_8537,N_8306);
nand U10129 (N_10129,N_8687,N_7814);
nand U10130 (N_10130,N_8013,N_8990);
nor U10131 (N_10131,N_8596,N_8163);
xor U10132 (N_10132,N_8062,N_7513);
nand U10133 (N_10133,N_7535,N_8592);
and U10134 (N_10134,N_7743,N_8549);
nand U10135 (N_10135,N_7687,N_8558);
nor U10136 (N_10136,N_8237,N_8985);
and U10137 (N_10137,N_8367,N_7895);
and U10138 (N_10138,N_7638,N_7724);
or U10139 (N_10139,N_7803,N_8335);
nor U10140 (N_10140,N_8774,N_7575);
and U10141 (N_10141,N_8300,N_7980);
and U10142 (N_10142,N_7593,N_7699);
xor U10143 (N_10143,N_8370,N_8627);
or U10144 (N_10144,N_8101,N_8870);
or U10145 (N_10145,N_7992,N_7940);
nand U10146 (N_10146,N_8443,N_7815);
nand U10147 (N_10147,N_8152,N_8673);
and U10148 (N_10148,N_7793,N_8884);
and U10149 (N_10149,N_8539,N_7632);
and U10150 (N_10150,N_8214,N_7603);
or U10151 (N_10151,N_8850,N_8624);
or U10152 (N_10152,N_8310,N_7990);
nor U10153 (N_10153,N_8866,N_8856);
and U10154 (N_10154,N_8589,N_8152);
xnor U10155 (N_10155,N_7919,N_7638);
and U10156 (N_10156,N_7986,N_8633);
nand U10157 (N_10157,N_8934,N_8442);
xor U10158 (N_10158,N_7748,N_8853);
nor U10159 (N_10159,N_8164,N_8938);
or U10160 (N_10160,N_8041,N_7654);
xor U10161 (N_10161,N_7962,N_8134);
nand U10162 (N_10162,N_7995,N_7791);
nand U10163 (N_10163,N_8986,N_7743);
nand U10164 (N_10164,N_8959,N_8474);
nor U10165 (N_10165,N_8432,N_8898);
and U10166 (N_10166,N_8264,N_8340);
nor U10167 (N_10167,N_8230,N_8623);
xor U10168 (N_10168,N_8946,N_7755);
nand U10169 (N_10169,N_8521,N_7754);
nor U10170 (N_10170,N_7962,N_8109);
nand U10171 (N_10171,N_7890,N_7779);
nor U10172 (N_10172,N_8310,N_8986);
xor U10173 (N_10173,N_8678,N_8270);
xnor U10174 (N_10174,N_8008,N_8177);
nand U10175 (N_10175,N_7779,N_7515);
and U10176 (N_10176,N_8933,N_7732);
or U10177 (N_10177,N_8199,N_7789);
or U10178 (N_10178,N_8187,N_8895);
xnor U10179 (N_10179,N_7669,N_7989);
xnor U10180 (N_10180,N_7908,N_7618);
or U10181 (N_10181,N_7699,N_7552);
xnor U10182 (N_10182,N_8053,N_8731);
xnor U10183 (N_10183,N_7814,N_8387);
nor U10184 (N_10184,N_8893,N_8554);
xnor U10185 (N_10185,N_8748,N_8873);
or U10186 (N_10186,N_8174,N_8245);
xnor U10187 (N_10187,N_8220,N_8079);
and U10188 (N_10188,N_8489,N_7580);
xor U10189 (N_10189,N_8688,N_8264);
xnor U10190 (N_10190,N_7662,N_8312);
and U10191 (N_10191,N_8267,N_8981);
nor U10192 (N_10192,N_8813,N_8411);
or U10193 (N_10193,N_7872,N_8521);
xnor U10194 (N_10194,N_8629,N_7654);
nand U10195 (N_10195,N_8054,N_8678);
nand U10196 (N_10196,N_7642,N_8031);
and U10197 (N_10197,N_7670,N_8538);
nand U10198 (N_10198,N_8110,N_8196);
and U10199 (N_10199,N_8926,N_8214);
nand U10200 (N_10200,N_8125,N_8442);
xor U10201 (N_10201,N_8589,N_8790);
nor U10202 (N_10202,N_8525,N_7912);
nor U10203 (N_10203,N_8551,N_8678);
or U10204 (N_10204,N_7501,N_7600);
and U10205 (N_10205,N_8176,N_7754);
nor U10206 (N_10206,N_8407,N_7545);
nor U10207 (N_10207,N_8079,N_8339);
or U10208 (N_10208,N_7919,N_7643);
nor U10209 (N_10209,N_8127,N_7832);
nand U10210 (N_10210,N_7976,N_7759);
nor U10211 (N_10211,N_8963,N_8880);
or U10212 (N_10212,N_8665,N_8060);
nand U10213 (N_10213,N_8854,N_7574);
or U10214 (N_10214,N_7552,N_8672);
xnor U10215 (N_10215,N_8264,N_8161);
xnor U10216 (N_10216,N_8848,N_8707);
and U10217 (N_10217,N_8366,N_7942);
and U10218 (N_10218,N_8988,N_8032);
nand U10219 (N_10219,N_7939,N_8401);
nand U10220 (N_10220,N_8272,N_8980);
nand U10221 (N_10221,N_7628,N_7686);
and U10222 (N_10222,N_8532,N_8304);
and U10223 (N_10223,N_8935,N_8494);
or U10224 (N_10224,N_8471,N_8156);
and U10225 (N_10225,N_8025,N_8077);
or U10226 (N_10226,N_7960,N_8663);
nand U10227 (N_10227,N_8718,N_7860);
nor U10228 (N_10228,N_8582,N_8286);
nand U10229 (N_10229,N_7641,N_8064);
or U10230 (N_10230,N_8788,N_8338);
nand U10231 (N_10231,N_8533,N_8103);
xnor U10232 (N_10232,N_7773,N_8375);
xnor U10233 (N_10233,N_8145,N_8136);
xnor U10234 (N_10234,N_8931,N_8896);
and U10235 (N_10235,N_8408,N_8241);
and U10236 (N_10236,N_7874,N_8260);
nand U10237 (N_10237,N_8548,N_7977);
nand U10238 (N_10238,N_8439,N_8411);
or U10239 (N_10239,N_7666,N_8555);
xnor U10240 (N_10240,N_7598,N_8866);
xnor U10241 (N_10241,N_8352,N_8302);
and U10242 (N_10242,N_8205,N_7541);
or U10243 (N_10243,N_8183,N_8586);
nor U10244 (N_10244,N_7902,N_8553);
nand U10245 (N_10245,N_8634,N_7775);
nand U10246 (N_10246,N_8701,N_8474);
nand U10247 (N_10247,N_7819,N_8464);
nor U10248 (N_10248,N_8857,N_8919);
nand U10249 (N_10249,N_7514,N_8074);
nand U10250 (N_10250,N_8120,N_8708);
nor U10251 (N_10251,N_7906,N_8191);
nand U10252 (N_10252,N_8828,N_7801);
and U10253 (N_10253,N_7524,N_7760);
or U10254 (N_10254,N_8816,N_7656);
nor U10255 (N_10255,N_7760,N_8845);
nor U10256 (N_10256,N_7765,N_7908);
nand U10257 (N_10257,N_8124,N_8286);
and U10258 (N_10258,N_7809,N_7787);
xor U10259 (N_10259,N_7706,N_8635);
xnor U10260 (N_10260,N_8453,N_7884);
and U10261 (N_10261,N_7777,N_8134);
xor U10262 (N_10262,N_8777,N_8724);
nor U10263 (N_10263,N_8016,N_8563);
nand U10264 (N_10264,N_8132,N_8131);
nand U10265 (N_10265,N_8237,N_7924);
or U10266 (N_10266,N_7631,N_7518);
xnor U10267 (N_10267,N_8237,N_8686);
xnor U10268 (N_10268,N_8210,N_7583);
xor U10269 (N_10269,N_8359,N_8195);
nand U10270 (N_10270,N_8697,N_7804);
xor U10271 (N_10271,N_8495,N_8988);
xor U10272 (N_10272,N_8937,N_8137);
nand U10273 (N_10273,N_8740,N_8694);
nor U10274 (N_10274,N_8629,N_8845);
nand U10275 (N_10275,N_7839,N_7887);
xnor U10276 (N_10276,N_8278,N_8123);
xor U10277 (N_10277,N_7585,N_8117);
nor U10278 (N_10278,N_8082,N_8460);
xnor U10279 (N_10279,N_8064,N_8947);
nor U10280 (N_10280,N_7834,N_8341);
or U10281 (N_10281,N_7990,N_8525);
xnor U10282 (N_10282,N_8455,N_8451);
and U10283 (N_10283,N_8431,N_8181);
nor U10284 (N_10284,N_8760,N_8718);
nor U10285 (N_10285,N_8728,N_7845);
nand U10286 (N_10286,N_8543,N_7592);
nor U10287 (N_10287,N_8506,N_7774);
or U10288 (N_10288,N_7814,N_8226);
nor U10289 (N_10289,N_8593,N_7828);
xor U10290 (N_10290,N_7882,N_8325);
nor U10291 (N_10291,N_8221,N_8902);
nor U10292 (N_10292,N_7814,N_8863);
nand U10293 (N_10293,N_8709,N_7573);
xor U10294 (N_10294,N_8086,N_8915);
or U10295 (N_10295,N_8515,N_8130);
xnor U10296 (N_10296,N_8636,N_8807);
or U10297 (N_10297,N_8261,N_8543);
and U10298 (N_10298,N_7924,N_8789);
nand U10299 (N_10299,N_8314,N_7961);
nand U10300 (N_10300,N_7997,N_7613);
xor U10301 (N_10301,N_7906,N_8073);
xor U10302 (N_10302,N_7992,N_7813);
xnor U10303 (N_10303,N_7930,N_8365);
xor U10304 (N_10304,N_8667,N_8392);
or U10305 (N_10305,N_8006,N_8712);
nor U10306 (N_10306,N_8122,N_8166);
xor U10307 (N_10307,N_8739,N_8407);
and U10308 (N_10308,N_8089,N_8665);
or U10309 (N_10309,N_7690,N_8332);
and U10310 (N_10310,N_8648,N_8668);
or U10311 (N_10311,N_8963,N_8428);
nor U10312 (N_10312,N_8865,N_8370);
nand U10313 (N_10313,N_8183,N_7842);
nor U10314 (N_10314,N_7925,N_7884);
nor U10315 (N_10315,N_8778,N_8565);
nand U10316 (N_10316,N_7647,N_8401);
nand U10317 (N_10317,N_8014,N_8855);
nor U10318 (N_10318,N_8658,N_8784);
xnor U10319 (N_10319,N_8049,N_8266);
or U10320 (N_10320,N_8184,N_8917);
xnor U10321 (N_10321,N_8796,N_8939);
or U10322 (N_10322,N_7853,N_8819);
nor U10323 (N_10323,N_8107,N_8477);
nor U10324 (N_10324,N_8148,N_8189);
or U10325 (N_10325,N_8021,N_8444);
or U10326 (N_10326,N_7937,N_7814);
and U10327 (N_10327,N_7981,N_8007);
nor U10328 (N_10328,N_8537,N_8338);
or U10329 (N_10329,N_8498,N_7634);
xnor U10330 (N_10330,N_8000,N_8610);
nor U10331 (N_10331,N_8397,N_8591);
and U10332 (N_10332,N_8728,N_7707);
nor U10333 (N_10333,N_8374,N_7733);
or U10334 (N_10334,N_8025,N_8782);
xnor U10335 (N_10335,N_8310,N_8455);
nand U10336 (N_10336,N_7960,N_7518);
or U10337 (N_10337,N_7679,N_7762);
and U10338 (N_10338,N_8219,N_8767);
and U10339 (N_10339,N_7636,N_7630);
or U10340 (N_10340,N_8286,N_7620);
or U10341 (N_10341,N_7738,N_8388);
nor U10342 (N_10342,N_7986,N_8598);
xor U10343 (N_10343,N_7740,N_7612);
or U10344 (N_10344,N_7804,N_7822);
or U10345 (N_10345,N_8856,N_8545);
nor U10346 (N_10346,N_8041,N_7873);
xnor U10347 (N_10347,N_7647,N_8196);
nand U10348 (N_10348,N_8114,N_7953);
or U10349 (N_10349,N_8313,N_8834);
nand U10350 (N_10350,N_7579,N_7530);
nor U10351 (N_10351,N_8749,N_8116);
xor U10352 (N_10352,N_8593,N_8944);
or U10353 (N_10353,N_8739,N_7711);
xor U10354 (N_10354,N_8767,N_8038);
or U10355 (N_10355,N_7825,N_8910);
nand U10356 (N_10356,N_8103,N_8004);
and U10357 (N_10357,N_8651,N_8166);
xnor U10358 (N_10358,N_7862,N_8980);
or U10359 (N_10359,N_8236,N_8931);
and U10360 (N_10360,N_8988,N_8430);
xor U10361 (N_10361,N_8477,N_8295);
nor U10362 (N_10362,N_8409,N_8481);
and U10363 (N_10363,N_7887,N_8342);
or U10364 (N_10364,N_8575,N_8935);
or U10365 (N_10365,N_8310,N_7955);
xor U10366 (N_10366,N_7886,N_8677);
or U10367 (N_10367,N_7722,N_7597);
and U10368 (N_10368,N_7546,N_7828);
nor U10369 (N_10369,N_7661,N_7775);
xor U10370 (N_10370,N_7806,N_7553);
and U10371 (N_10371,N_8734,N_8629);
nand U10372 (N_10372,N_8977,N_8366);
xnor U10373 (N_10373,N_8498,N_7714);
and U10374 (N_10374,N_8110,N_8070);
nand U10375 (N_10375,N_8075,N_8804);
nand U10376 (N_10376,N_8389,N_7962);
nand U10377 (N_10377,N_7609,N_7896);
and U10378 (N_10378,N_8992,N_7527);
or U10379 (N_10379,N_7844,N_8831);
and U10380 (N_10380,N_7686,N_8897);
nor U10381 (N_10381,N_8107,N_8770);
or U10382 (N_10382,N_7679,N_7867);
and U10383 (N_10383,N_8901,N_8450);
nor U10384 (N_10384,N_8908,N_7549);
and U10385 (N_10385,N_8399,N_8179);
or U10386 (N_10386,N_8873,N_8793);
xnor U10387 (N_10387,N_8319,N_7779);
xnor U10388 (N_10388,N_8181,N_8325);
xor U10389 (N_10389,N_8681,N_8691);
nand U10390 (N_10390,N_8136,N_8169);
xnor U10391 (N_10391,N_7806,N_8327);
nor U10392 (N_10392,N_7727,N_8525);
nand U10393 (N_10393,N_8277,N_8887);
nand U10394 (N_10394,N_8514,N_8313);
nor U10395 (N_10395,N_8592,N_8799);
nor U10396 (N_10396,N_8124,N_8764);
and U10397 (N_10397,N_8807,N_8010);
xnor U10398 (N_10398,N_7793,N_7780);
xor U10399 (N_10399,N_8391,N_7980);
or U10400 (N_10400,N_7907,N_8059);
and U10401 (N_10401,N_8407,N_8672);
xnor U10402 (N_10402,N_8943,N_7558);
nor U10403 (N_10403,N_7946,N_7814);
xor U10404 (N_10404,N_8496,N_8035);
nand U10405 (N_10405,N_8907,N_8676);
nor U10406 (N_10406,N_8853,N_8623);
xnor U10407 (N_10407,N_8904,N_7726);
or U10408 (N_10408,N_8586,N_7636);
nor U10409 (N_10409,N_7565,N_8914);
and U10410 (N_10410,N_8074,N_8662);
nand U10411 (N_10411,N_7626,N_8871);
nor U10412 (N_10412,N_8406,N_8935);
nand U10413 (N_10413,N_7967,N_8687);
and U10414 (N_10414,N_7942,N_8291);
nor U10415 (N_10415,N_8899,N_8203);
xor U10416 (N_10416,N_8356,N_8858);
nand U10417 (N_10417,N_8043,N_7835);
or U10418 (N_10418,N_8785,N_8720);
nor U10419 (N_10419,N_8650,N_8392);
xnor U10420 (N_10420,N_7855,N_7645);
xnor U10421 (N_10421,N_7813,N_8029);
or U10422 (N_10422,N_7956,N_8205);
and U10423 (N_10423,N_7904,N_8902);
and U10424 (N_10424,N_8974,N_7646);
xor U10425 (N_10425,N_7669,N_8827);
nand U10426 (N_10426,N_8366,N_8401);
xor U10427 (N_10427,N_7611,N_8191);
nor U10428 (N_10428,N_7970,N_8998);
nand U10429 (N_10429,N_7879,N_8587);
or U10430 (N_10430,N_8148,N_7816);
nand U10431 (N_10431,N_8291,N_8962);
nor U10432 (N_10432,N_7853,N_8133);
nor U10433 (N_10433,N_8323,N_7946);
and U10434 (N_10434,N_8906,N_8528);
or U10435 (N_10435,N_8338,N_7808);
nor U10436 (N_10436,N_7689,N_8249);
and U10437 (N_10437,N_8815,N_8315);
nor U10438 (N_10438,N_7924,N_8766);
xor U10439 (N_10439,N_8539,N_7658);
or U10440 (N_10440,N_8642,N_8617);
or U10441 (N_10441,N_8197,N_7962);
nor U10442 (N_10442,N_7625,N_7785);
or U10443 (N_10443,N_7550,N_8029);
or U10444 (N_10444,N_8876,N_8496);
xnor U10445 (N_10445,N_8048,N_7848);
xnor U10446 (N_10446,N_8544,N_7927);
or U10447 (N_10447,N_8672,N_7930);
or U10448 (N_10448,N_8174,N_7762);
nand U10449 (N_10449,N_8517,N_8853);
nor U10450 (N_10450,N_7549,N_7922);
and U10451 (N_10451,N_8749,N_8137);
nor U10452 (N_10452,N_7603,N_8899);
xor U10453 (N_10453,N_8253,N_7991);
nor U10454 (N_10454,N_8048,N_8740);
xnor U10455 (N_10455,N_8180,N_8903);
xnor U10456 (N_10456,N_8065,N_8777);
xor U10457 (N_10457,N_8287,N_8400);
nand U10458 (N_10458,N_7778,N_7506);
nand U10459 (N_10459,N_7591,N_8327);
nand U10460 (N_10460,N_8115,N_7588);
nor U10461 (N_10461,N_8258,N_8562);
nand U10462 (N_10462,N_8353,N_8549);
or U10463 (N_10463,N_8070,N_8768);
and U10464 (N_10464,N_7822,N_8479);
or U10465 (N_10465,N_8898,N_8012);
and U10466 (N_10466,N_8794,N_8032);
nand U10467 (N_10467,N_8002,N_8024);
or U10468 (N_10468,N_8377,N_8308);
nand U10469 (N_10469,N_7594,N_8753);
or U10470 (N_10470,N_8592,N_8039);
and U10471 (N_10471,N_8752,N_8388);
and U10472 (N_10472,N_7932,N_8164);
and U10473 (N_10473,N_8330,N_8463);
nand U10474 (N_10474,N_8000,N_8248);
xor U10475 (N_10475,N_8974,N_8056);
nand U10476 (N_10476,N_8714,N_7887);
nand U10477 (N_10477,N_8964,N_8566);
or U10478 (N_10478,N_8186,N_8202);
and U10479 (N_10479,N_7599,N_8544);
and U10480 (N_10480,N_8758,N_7830);
xnor U10481 (N_10481,N_7976,N_7731);
and U10482 (N_10482,N_7802,N_7760);
nand U10483 (N_10483,N_8210,N_8574);
and U10484 (N_10484,N_8622,N_8576);
or U10485 (N_10485,N_8462,N_7646);
and U10486 (N_10486,N_8090,N_7859);
nor U10487 (N_10487,N_8184,N_7568);
nor U10488 (N_10488,N_8783,N_7736);
xor U10489 (N_10489,N_7692,N_8215);
nor U10490 (N_10490,N_7593,N_8185);
nor U10491 (N_10491,N_7670,N_7557);
and U10492 (N_10492,N_8057,N_8633);
nand U10493 (N_10493,N_7590,N_8724);
or U10494 (N_10494,N_8264,N_8621);
nand U10495 (N_10495,N_8001,N_7503);
or U10496 (N_10496,N_8847,N_7919);
nor U10497 (N_10497,N_7776,N_7669);
and U10498 (N_10498,N_7781,N_8548);
and U10499 (N_10499,N_7548,N_8456);
nand U10500 (N_10500,N_9606,N_9624);
nand U10501 (N_10501,N_10080,N_9349);
and U10502 (N_10502,N_9258,N_9456);
nor U10503 (N_10503,N_9806,N_10477);
and U10504 (N_10504,N_9556,N_9749);
nor U10505 (N_10505,N_10291,N_9306);
xor U10506 (N_10506,N_9681,N_9150);
and U10507 (N_10507,N_9940,N_10135);
or U10508 (N_10508,N_9555,N_9290);
nor U10509 (N_10509,N_10186,N_10497);
xnor U10510 (N_10510,N_9999,N_9305);
and U10511 (N_10511,N_9796,N_9830);
or U10512 (N_10512,N_10348,N_10173);
nand U10513 (N_10513,N_10161,N_9194);
xnor U10514 (N_10514,N_10391,N_9301);
nand U10515 (N_10515,N_9770,N_10101);
xor U10516 (N_10516,N_10312,N_10165);
nor U10517 (N_10517,N_10207,N_9615);
nand U10518 (N_10518,N_10462,N_10117);
nand U10519 (N_10519,N_9854,N_9472);
nor U10520 (N_10520,N_10199,N_9333);
or U10521 (N_10521,N_9224,N_9040);
nand U10522 (N_10522,N_9067,N_10150);
and U10523 (N_10523,N_10491,N_9804);
nor U10524 (N_10524,N_9761,N_9088);
nand U10525 (N_10525,N_9017,N_10012);
nor U10526 (N_10526,N_9044,N_9441);
or U10527 (N_10527,N_9825,N_10006);
nor U10528 (N_10528,N_9286,N_9664);
xnor U10529 (N_10529,N_9679,N_10263);
xor U10530 (N_10530,N_9449,N_9799);
nor U10531 (N_10531,N_10390,N_9170);
or U10532 (N_10532,N_9809,N_9880);
and U10533 (N_10533,N_9535,N_9543);
xnor U10534 (N_10534,N_9188,N_9596);
or U10535 (N_10535,N_9186,N_10028);
or U10536 (N_10536,N_9722,N_9317);
nor U10537 (N_10537,N_10473,N_9032);
or U10538 (N_10538,N_9402,N_10097);
or U10539 (N_10539,N_10287,N_10055);
or U10540 (N_10540,N_9148,N_9971);
nand U10541 (N_10541,N_9257,N_10131);
and U10542 (N_10542,N_9497,N_10201);
nor U10543 (N_10543,N_10014,N_9213);
xor U10544 (N_10544,N_9575,N_9523);
nand U10545 (N_10545,N_9812,N_9782);
xnor U10546 (N_10546,N_9878,N_9353);
xnor U10547 (N_10547,N_10400,N_9490);
or U10548 (N_10548,N_9862,N_10159);
and U10549 (N_10549,N_9502,N_10119);
or U10550 (N_10550,N_10399,N_9364);
xor U10551 (N_10551,N_10110,N_10032);
and U10552 (N_10552,N_9287,N_9611);
nor U10553 (N_10553,N_10375,N_10191);
or U10554 (N_10554,N_9656,N_10264);
or U10555 (N_10555,N_9025,N_9473);
nor U10556 (N_10556,N_9685,N_9351);
or U10557 (N_10557,N_10356,N_9002);
nand U10558 (N_10558,N_9215,N_10317);
or U10559 (N_10559,N_10449,N_9135);
nor U10560 (N_10560,N_9197,N_9289);
nand U10561 (N_10561,N_10351,N_10407);
nand U10562 (N_10562,N_10061,N_9597);
or U10563 (N_10563,N_10283,N_9807);
and U10564 (N_10564,N_9978,N_9553);
nor U10565 (N_10565,N_10498,N_9263);
and U10566 (N_10566,N_9089,N_9536);
xnor U10567 (N_10567,N_10451,N_10409);
or U10568 (N_10568,N_9193,N_9636);
or U10569 (N_10569,N_10043,N_9474);
nor U10570 (N_10570,N_9550,N_9237);
nor U10571 (N_10571,N_10084,N_9847);
or U10572 (N_10572,N_9779,N_9660);
or U10573 (N_10573,N_9871,N_10208);
nand U10574 (N_10574,N_10347,N_9525);
and U10575 (N_10575,N_9696,N_9166);
or U10576 (N_10576,N_9739,N_9266);
or U10577 (N_10577,N_10403,N_9683);
or U10578 (N_10578,N_10478,N_9726);
or U10579 (N_10579,N_9352,N_9600);
xor U10580 (N_10580,N_9203,N_9658);
xor U10581 (N_10581,N_9108,N_10001);
nor U10582 (N_10582,N_9835,N_9222);
nor U10583 (N_10583,N_9297,N_9922);
xnor U10584 (N_10584,N_9322,N_9250);
nand U10585 (N_10585,N_10321,N_9476);
and U10586 (N_10586,N_9813,N_9451);
nor U10587 (N_10587,N_9489,N_9443);
xor U10588 (N_10588,N_10248,N_9914);
nor U10589 (N_10589,N_9709,N_9657);
nor U10590 (N_10590,N_9540,N_9568);
nand U10591 (N_10591,N_9805,N_10083);
nand U10592 (N_10592,N_9665,N_9762);
or U10593 (N_10593,N_9817,N_9344);
nand U10594 (N_10594,N_9751,N_10433);
xor U10595 (N_10595,N_9917,N_10438);
xnor U10596 (N_10596,N_9050,N_9731);
or U10597 (N_10597,N_9243,N_9638);
nor U10598 (N_10598,N_10295,N_9339);
nand U10599 (N_10599,N_9926,N_9784);
nand U10600 (N_10600,N_10395,N_9220);
or U10601 (N_10601,N_9918,N_9792);
nor U10602 (N_10602,N_9292,N_10389);
and U10603 (N_10603,N_10034,N_10382);
xor U10604 (N_10604,N_10079,N_10422);
and U10605 (N_10605,N_9894,N_9533);
and U10606 (N_10606,N_9399,N_10410);
and U10607 (N_10607,N_10446,N_9617);
nand U10608 (N_10608,N_9732,N_10260);
and U10609 (N_10609,N_10194,N_9572);
and U10610 (N_10610,N_10171,N_9157);
or U10611 (N_10611,N_9361,N_9149);
nor U10612 (N_10612,N_9381,N_9702);
xnor U10613 (N_10613,N_10420,N_9299);
nor U10614 (N_10614,N_10257,N_10126);
nor U10615 (N_10615,N_10298,N_9013);
or U10616 (N_10616,N_9059,N_9569);
nor U10617 (N_10617,N_10481,N_9909);
or U10618 (N_10618,N_10387,N_9808);
xor U10619 (N_10619,N_9986,N_10058);
or U10620 (N_10620,N_10123,N_9628);
and U10621 (N_10621,N_9948,N_9652);
or U10622 (N_10622,N_9189,N_9057);
and U10623 (N_10623,N_9105,N_9083);
xor U10624 (N_10624,N_9358,N_9343);
xnor U10625 (N_10625,N_10251,N_9227);
nor U10626 (N_10626,N_9113,N_9255);
or U10627 (N_10627,N_10282,N_10447);
nand U10628 (N_10628,N_9532,N_9947);
and U10629 (N_10629,N_10211,N_9026);
nand U10630 (N_10630,N_10064,N_9637);
or U10631 (N_10631,N_9187,N_9405);
nor U10632 (N_10632,N_9336,N_10139);
or U10633 (N_10633,N_9527,N_10360);
xor U10634 (N_10634,N_9115,N_9750);
or U10635 (N_10635,N_10299,N_9642);
or U10636 (N_10636,N_9867,N_9695);
xor U10637 (N_10637,N_10279,N_9130);
nor U10638 (N_10638,N_10371,N_9863);
or U10639 (N_10639,N_9445,N_9071);
nand U10640 (N_10640,N_10378,N_9706);
or U10641 (N_10641,N_9435,N_9453);
nor U10642 (N_10642,N_9409,N_10175);
xnor U10643 (N_10643,N_9626,N_10411);
nand U10644 (N_10644,N_9654,N_9776);
nand U10645 (N_10645,N_9327,N_9162);
nor U10646 (N_10646,N_9531,N_10047);
nand U10647 (N_10647,N_9647,N_10326);
nand U10648 (N_10648,N_9547,N_9080);
and U10649 (N_10649,N_9946,N_10185);
and U10650 (N_10650,N_10346,N_9119);
nand U10651 (N_10651,N_9426,N_10107);
or U10652 (N_10652,N_9663,N_10322);
and U10653 (N_10653,N_9463,N_9646);
or U10654 (N_10654,N_9700,N_10294);
or U10655 (N_10655,N_10472,N_9365);
and U10656 (N_10656,N_9398,N_9114);
nor U10657 (N_10657,N_9885,N_9240);
nor U10658 (N_10658,N_9487,N_9325);
and U10659 (N_10659,N_9832,N_9068);
or U10660 (N_10660,N_9499,N_9980);
nand U10661 (N_10661,N_9208,N_10334);
or U10662 (N_10662,N_9753,N_9217);
or U10663 (N_10663,N_10457,N_10020);
nand U10664 (N_10664,N_9086,N_9455);
or U10665 (N_10665,N_10075,N_9640);
and U10666 (N_10666,N_9109,N_9414);
or U10667 (N_10667,N_9763,N_10431);
and U10668 (N_10668,N_10241,N_9406);
nor U10669 (N_10669,N_9842,N_10327);
or U10670 (N_10670,N_10417,N_9648);
nand U10671 (N_10671,N_9141,N_9676);
nand U10672 (N_10672,N_9586,N_10204);
nand U10673 (N_10673,N_10278,N_9239);
xor U10674 (N_10674,N_9356,N_9219);
nor U10675 (N_10675,N_10448,N_9641);
and U10676 (N_10676,N_10088,N_9493);
or U10677 (N_10677,N_9605,N_9697);
nand U10678 (N_10678,N_9147,N_10011);
nand U10679 (N_10679,N_9383,N_10373);
nor U10680 (N_10680,N_9350,N_10349);
and U10681 (N_10681,N_9524,N_9419);
and U10682 (N_10682,N_10179,N_10017);
and U10683 (N_10683,N_9171,N_9758);
xor U10684 (N_10684,N_10486,N_9688);
nand U10685 (N_10685,N_10316,N_10499);
xnor U10686 (N_10686,N_10189,N_9734);
nor U10687 (N_10687,N_10021,N_10000);
xor U10688 (N_10688,N_9639,N_9416);
nand U10689 (N_10689,N_9538,N_9400);
xor U10690 (N_10690,N_9081,N_10086);
nand U10691 (N_10691,N_10067,N_9016);
or U10692 (N_10692,N_10401,N_10377);
and U10693 (N_10693,N_9902,N_9049);
or U10694 (N_10694,N_9018,N_9466);
nor U10695 (N_10695,N_10015,N_10254);
or U10696 (N_10696,N_9727,N_9311);
nor U10697 (N_10697,N_9513,N_10070);
xnor U10698 (N_10698,N_9191,N_9201);
nor U10699 (N_10699,N_10217,N_9669);
or U10700 (N_10700,N_9315,N_9882);
nand U10701 (N_10701,N_9529,N_10030);
or U10702 (N_10702,N_10048,N_10138);
nor U10703 (N_10703,N_9632,N_9755);
xor U10704 (N_10704,N_10009,N_10104);
nand U10705 (N_10705,N_9460,N_9559);
xor U10706 (N_10706,N_10482,N_9142);
xor U10707 (N_10707,N_9843,N_10314);
and U10708 (N_10708,N_9877,N_9485);
or U10709 (N_10709,N_9376,N_10026);
and U10710 (N_10710,N_9670,N_9927);
and U10711 (N_10711,N_9504,N_9928);
nor U10712 (N_10712,N_10111,N_9587);
or U10713 (N_10713,N_10113,N_9087);
nor U10714 (N_10714,N_9342,N_10145);
nor U10715 (N_10715,N_9671,N_9833);
and U10716 (N_10716,N_10124,N_9649);
or U10717 (N_10717,N_10071,N_10464);
nand U10718 (N_10718,N_9300,N_10040);
and U10719 (N_10719,N_9552,N_10100);
xor U10720 (N_10720,N_9388,N_9477);
nand U10721 (N_10721,N_9438,N_9184);
xor U10722 (N_10722,N_9022,N_9881);
nor U10723 (N_10723,N_9936,N_9179);
nor U10724 (N_10724,N_9009,N_9218);
xnor U10725 (N_10725,N_9367,N_10225);
nor U10726 (N_10726,N_10151,N_9452);
nand U10727 (N_10727,N_9169,N_10008);
nand U10728 (N_10728,N_9124,N_10300);
xor U10729 (N_10729,N_9043,N_10495);
or U10730 (N_10730,N_9116,N_10042);
or U10731 (N_10731,N_9693,N_10418);
nand U10732 (N_10732,N_9053,N_9889);
nand U10733 (N_10733,N_9888,N_9372);
nand U10734 (N_10734,N_9037,N_10219);
xnor U10735 (N_10735,N_9030,N_9653);
xnor U10736 (N_10736,N_9848,N_9082);
xor U10737 (N_10737,N_9355,N_10428);
xor U10738 (N_10738,N_10484,N_10277);
nand U10739 (N_10739,N_9629,N_10181);
nor U10740 (N_10740,N_9394,N_9828);
or U10741 (N_10741,N_9613,N_10330);
or U10742 (N_10742,N_9713,N_10024);
or U10743 (N_10743,N_10333,N_10091);
xnor U10744 (N_10744,N_9982,N_9957);
xnor U10745 (N_10745,N_9964,N_9144);
nand U10746 (N_10746,N_9253,N_10213);
or U10747 (N_10747,N_9935,N_9512);
xor U10748 (N_10748,N_9873,N_9991);
xnor U10749 (N_10749,N_9977,N_9601);
nand U10750 (N_10750,N_10419,N_10023);
nor U10751 (N_10751,N_10053,N_9137);
nand U10752 (N_10752,N_9714,N_9506);
nand U10753 (N_10753,N_9181,N_9459);
and U10754 (N_10754,N_9915,N_10423);
xor U10755 (N_10755,N_10209,N_9786);
xnor U10756 (N_10756,N_9412,N_9246);
xor U10757 (N_10757,N_9987,N_10441);
and U10758 (N_10758,N_9816,N_10246);
nand U10759 (N_10759,N_9296,N_10466);
nor U10760 (N_10760,N_9974,N_10149);
or U10761 (N_10761,N_9158,N_9746);
nor U10762 (N_10762,N_9790,N_9844);
or U10763 (N_10763,N_10458,N_9682);
nor U10764 (N_10764,N_9276,N_9908);
xnor U10765 (N_10765,N_9103,N_10489);
and U10766 (N_10766,N_10002,N_10394);
and U10767 (N_10767,N_9427,N_10019);
nor U10768 (N_10768,N_9491,N_10049);
or U10769 (N_10769,N_9920,N_9967);
and U10770 (N_10770,N_9571,N_9185);
nand U10771 (N_10771,N_10013,N_9969);
and U10772 (N_10772,N_10154,N_9655);
xnor U10773 (N_10773,N_9274,N_9139);
nor U10774 (N_10774,N_9265,N_9096);
xnor U10775 (N_10775,N_10096,N_9836);
and U10776 (N_10776,N_10370,N_10365);
and U10777 (N_10777,N_9757,N_10092);
nand U10778 (N_10778,N_10271,N_10338);
or U10779 (N_10779,N_10483,N_9800);
or U10780 (N_10780,N_10054,N_10357);
nor U10781 (N_10781,N_9981,N_10052);
nor U10782 (N_10782,N_10041,N_9024);
nor U10783 (N_10783,N_9730,N_10465);
nor U10784 (N_10784,N_9737,N_9308);
and U10785 (N_10785,N_10276,N_9495);
or U10786 (N_10786,N_9341,N_9063);
nand U10787 (N_10787,N_10468,N_9846);
xor U10788 (N_10788,N_9937,N_9230);
xor U10789 (N_10789,N_9129,N_9318);
xor U10790 (N_10790,N_10308,N_9444);
or U10791 (N_10791,N_9360,N_9963);
xnor U10792 (N_10792,N_9277,N_9955);
xor U10793 (N_10793,N_9768,N_9033);
nand U10794 (N_10794,N_9408,N_9078);
and U10795 (N_10795,N_9202,N_9542);
nand U10796 (N_10796,N_9146,N_9269);
xor U10797 (N_10797,N_9397,N_9574);
or U10798 (N_10798,N_10331,N_10359);
and U10799 (N_10799,N_9074,N_9125);
nand U10800 (N_10800,N_9121,N_9905);
nand U10801 (N_10801,N_9772,N_10494);
or U10802 (N_10802,N_10436,N_9385);
nor U10803 (N_10803,N_9176,N_9012);
xnor U10804 (N_10804,N_9954,N_10073);
or U10805 (N_10805,N_9229,N_9519);
nor U10806 (N_10806,N_10060,N_9993);
xor U10807 (N_10807,N_10076,N_10228);
and U10808 (N_10808,N_9826,N_10218);
nor U10809 (N_10809,N_9155,N_9561);
nand U10810 (N_10810,N_10144,N_9190);
nand U10811 (N_10811,N_9959,N_10022);
xor U10812 (N_10812,N_9313,N_9590);
nand U10813 (N_10813,N_10461,N_9488);
nor U10814 (N_10814,N_9211,N_10339);
nand U10815 (N_10815,N_9284,N_10190);
xor U10816 (N_10816,N_9268,N_9212);
nor U10817 (N_10817,N_9968,N_10036);
or U10818 (N_10818,N_9055,N_9573);
nor U10819 (N_10819,N_9175,N_9038);
nand U10820 (N_10820,N_9686,N_9106);
xor U10821 (N_10821,N_10492,N_10141);
nor U10822 (N_10822,N_10450,N_9990);
nor U10823 (N_10823,N_10183,N_9780);
xor U10824 (N_10824,N_9324,N_10453);
nor U10825 (N_10825,N_10344,N_9966);
or U10826 (N_10826,N_9172,N_9484);
or U10827 (N_10827,N_10315,N_9764);
and U10828 (N_10828,N_9391,N_10142);
or U10829 (N_10829,N_10169,N_9973);
and U10830 (N_10830,N_9522,N_9164);
and U10831 (N_10831,N_9868,N_10031);
and U10832 (N_10832,N_9432,N_10487);
nand U10833 (N_10833,N_9478,N_10253);
nor U10834 (N_10834,N_9869,N_9410);
nand U10835 (N_10835,N_10247,N_10147);
nand U10836 (N_10836,N_10426,N_9811);
nand U10837 (N_10837,N_9235,N_10266);
nor U10838 (N_10838,N_9347,N_9395);
nand U10839 (N_10839,N_9960,N_9006);
nor U10840 (N_10840,N_10490,N_9595);
and U10841 (N_10841,N_9029,N_10098);
or U10842 (N_10842,N_9199,N_10106);
xor U10843 (N_10843,N_9956,N_9165);
nand U10844 (N_10844,N_9112,N_9430);
nor U10845 (N_10845,N_9226,N_9724);
and U10846 (N_10846,N_10078,N_9454);
xnor U10847 (N_10847,N_10429,N_9518);
nand U10848 (N_10848,N_9668,N_9994);
or U10849 (N_10849,N_9450,N_9421);
and U10850 (N_10850,N_10109,N_10252);
xor U10851 (N_10851,N_9934,N_9375);
and U10852 (N_10852,N_9879,N_10153);
and U10853 (N_10853,N_10474,N_9992);
nand U10854 (N_10854,N_9931,N_9008);
or U10855 (N_10855,N_9567,N_10146);
or U10856 (N_10856,N_9622,N_9797);
and U10857 (N_10857,N_9136,N_9072);
nor U10858 (N_10858,N_9717,N_9952);
nor U10859 (N_10859,N_9608,N_9810);
nand U10860 (N_10860,N_9077,N_9154);
xor U10861 (N_10861,N_10274,N_10444);
nand U10862 (N_10862,N_9035,N_9516);
nand U10863 (N_10863,N_9280,N_9330);
xor U10864 (N_10864,N_10004,N_9195);
or U10865 (N_10865,N_9890,N_9541);
nor U10866 (N_10866,N_9238,N_9769);
nand U10867 (N_10867,N_9126,N_10336);
nand U10868 (N_10868,N_10386,N_9442);
nor U10869 (N_10869,N_9924,N_10425);
nor U10870 (N_10870,N_10323,N_9446);
nor U10871 (N_10871,N_9584,N_9143);
xnor U10872 (N_10872,N_9962,N_9771);
or U10873 (N_10873,N_9910,N_10105);
or U10874 (N_10874,N_9396,N_9983);
xnor U10875 (N_10875,N_10259,N_10262);
and U10876 (N_10876,N_9895,N_9876);
nand U10877 (N_10877,N_10269,N_10280);
nand U10878 (N_10878,N_9241,N_9228);
or U10879 (N_10879,N_9675,N_9743);
nand U10880 (N_10880,N_9362,N_9643);
nor U10881 (N_10881,N_9778,N_9282);
nor U10882 (N_10882,N_10313,N_10116);
nor U10883 (N_10883,N_9036,N_10152);
or U10884 (N_10884,N_9363,N_9858);
or U10885 (N_10885,N_9845,N_9373);
and U10886 (N_10886,N_9598,N_10309);
xnor U10887 (N_10887,N_10227,N_10188);
nor U10888 (N_10888,N_10198,N_10235);
and U10889 (N_10889,N_9483,N_10035);
nor U10890 (N_10890,N_10268,N_10087);
and U10891 (N_10891,N_9509,N_9329);
nor U10892 (N_10892,N_9401,N_9505);
nor U10893 (N_10893,N_10214,N_9084);
or U10894 (N_10894,N_9929,N_9110);
nor U10895 (N_10895,N_9413,N_9995);
xor U10896 (N_10896,N_9650,N_9599);
nor U10897 (N_10897,N_9949,N_9554);
and U10898 (N_10898,N_9942,N_10362);
nand U10899 (N_10899,N_10454,N_9248);
xnor U10900 (N_10900,N_9591,N_10203);
nand U10901 (N_10901,N_10044,N_9581);
nand U10902 (N_10902,N_10258,N_9976);
nor U10903 (N_10903,N_9630,N_10305);
or U10904 (N_10904,N_9161,N_9687);
nand U10905 (N_10905,N_9680,N_10239);
xnor U10906 (N_10906,N_10121,N_10488);
and U10907 (N_10907,N_9851,N_9919);
and U10908 (N_10908,N_9699,N_10128);
nor U10909 (N_10909,N_10130,N_9251);
xnor U10910 (N_10910,N_9264,N_9837);
or U10911 (N_10911,N_9620,N_9625);
nor U10912 (N_10912,N_10281,N_10366);
nand U10913 (N_10913,N_9293,N_10493);
nor U10914 (N_10914,N_9386,N_9475);
or U10915 (N_10915,N_10112,N_9102);
nor U10916 (N_10916,N_9281,N_9609);
xnor U10917 (N_10917,N_9803,N_9874);
xor U10918 (N_10918,N_10379,N_10319);
nor U10919 (N_10919,N_9236,N_9298);
nor U10920 (N_10920,N_9131,N_9801);
or U10921 (N_10921,N_9859,N_9231);
and U10922 (N_10922,N_10158,N_9123);
nand U10923 (N_10923,N_9337,N_10414);
nor U10924 (N_10924,N_9777,N_9431);
nand U10925 (N_10925,N_10122,N_9100);
nor U10926 (N_10926,N_10289,N_9984);
and U10927 (N_10927,N_10063,N_10082);
nor U10928 (N_10928,N_9913,N_10430);
nand U10929 (N_10929,N_9511,N_10125);
nor U10930 (N_10930,N_9198,N_9133);
and U10931 (N_10931,N_9562,N_10220);
and U10932 (N_10932,N_9145,N_10270);
nor U10933 (N_10933,N_10232,N_10206);
xor U10934 (N_10934,N_10320,N_10345);
and U10935 (N_10935,N_9254,N_9719);
and U10936 (N_10936,N_9767,N_9965);
xor U10937 (N_10937,N_10479,N_9312);
nor U10938 (N_10938,N_9850,N_9612);
nor U10939 (N_10939,N_9214,N_9901);
nand U10940 (N_10940,N_10301,N_9010);
or U10941 (N_10941,N_9708,N_9689);
nor U10942 (N_10942,N_9046,N_9997);
xor U10943 (N_10943,N_9933,N_9062);
xnor U10944 (N_10944,N_9415,N_10195);
xnor U10945 (N_10945,N_9521,N_9517);
and U10946 (N_10946,N_9468,N_9140);
nand U10947 (N_10947,N_10434,N_10074);
and U10948 (N_10948,N_9206,N_9411);
nand U10949 (N_10949,N_9418,N_10212);
xnor U10950 (N_10950,N_9651,N_10196);
nand U10951 (N_10951,N_10396,N_10293);
xnor U10952 (N_10952,N_10475,N_9094);
nand U10953 (N_10953,N_10134,N_9823);
nor U10954 (N_10954,N_9093,N_9975);
xnor U10955 (N_10955,N_9793,N_9374);
and U10956 (N_10956,N_9501,N_9180);
nand U10957 (N_10957,N_10406,N_9610);
and U10958 (N_10958,N_9073,N_9701);
nor U10959 (N_10959,N_9721,N_9461);
and U10960 (N_10960,N_9548,N_9745);
or U10961 (N_10961,N_9303,N_9723);
nor U10962 (N_10962,N_9822,N_9530);
and U10963 (N_10963,N_10155,N_10455);
or U10964 (N_10964,N_10443,N_10255);
or U10965 (N_10965,N_10093,N_9849);
and U10966 (N_10966,N_9393,N_9633);
xor U10967 (N_10967,N_9285,N_10329);
or U10968 (N_10968,N_9659,N_9594);
nand U10969 (N_10969,N_9392,N_9005);
and U10970 (N_10970,N_10384,N_9423);
nor U10971 (N_10971,N_9950,N_9666);
nand U10972 (N_10972,N_9359,N_9467);
or U10973 (N_10973,N_9930,N_10230);
xnor U10974 (N_10974,N_9684,N_9748);
xnor U10975 (N_10975,N_9566,N_10480);
or U10976 (N_10976,N_10164,N_10413);
and U10977 (N_10977,N_10167,N_9703);
and U10978 (N_10978,N_9480,N_10292);
nor U10979 (N_10979,N_9672,N_9824);
nand U10980 (N_10980,N_9107,N_10467);
and U10981 (N_10981,N_10005,N_9883);
nor U10982 (N_10982,N_10069,N_9207);
nand U10983 (N_10983,N_9168,N_9773);
nor U10984 (N_10984,N_10355,N_9066);
nand U10985 (N_10985,N_10056,N_9326);
and U10986 (N_10986,N_9616,N_9234);
xnor U10987 (N_10987,N_10223,N_9134);
and U10988 (N_10988,N_10018,N_9316);
or U10989 (N_10989,N_10176,N_10140);
and U10990 (N_10990,N_9537,N_9526);
nand U10991 (N_10991,N_9494,N_9576);
nor U10992 (N_10992,N_9893,N_9334);
xnor U10993 (N_10993,N_9345,N_10421);
or U10994 (N_10994,N_9853,N_9906);
nor U10995 (N_10995,N_10470,N_10304);
or U10996 (N_10996,N_9787,N_10285);
xnor U10997 (N_10997,N_9802,N_10437);
nor U10998 (N_10998,N_9674,N_10148);
and U10999 (N_10999,N_9691,N_10376);
nor U11000 (N_11000,N_9321,N_10469);
xor U11001 (N_11001,N_9027,N_9335);
or U11002 (N_11002,N_9818,N_9623);
nor U11003 (N_11003,N_9514,N_9589);
nor U11004 (N_11004,N_9662,N_9865);
or U11005 (N_11005,N_10435,N_10306);
nand U11006 (N_11006,N_9607,N_9465);
nand U11007 (N_11007,N_9690,N_9961);
xnor U11008 (N_11008,N_10302,N_10416);
nand U11009 (N_11009,N_10335,N_9661);
and U11010 (N_11010,N_9733,N_9216);
nor U11011 (N_11011,N_10210,N_10234);
or U11012 (N_11012,N_9953,N_10231);
or U11013 (N_11013,N_10476,N_10233);
xor U11014 (N_11014,N_9271,N_9019);
nand U11015 (N_11015,N_9741,N_9378);
and U11016 (N_11016,N_10445,N_9247);
and U11017 (N_11017,N_9677,N_9970);
nand U11018 (N_11018,N_10068,N_10397);
or U11019 (N_11019,N_9544,N_9602);
xnor U11020 (N_11020,N_9943,N_9515);
nand U11021 (N_11021,N_9020,N_10310);
xnor U11022 (N_11022,N_9153,N_9099);
or U11023 (N_11023,N_9302,N_9331);
xnor U11024 (N_11024,N_9582,N_9380);
or U11025 (N_11025,N_9028,N_9420);
nand U11026 (N_11026,N_9998,N_9744);
xor U11027 (N_11027,N_10439,N_10129);
and U11028 (N_11028,N_10143,N_9132);
or U11029 (N_11029,N_9939,N_9896);
and U11030 (N_11030,N_10193,N_9437);
and U11031 (N_11031,N_10132,N_9945);
nor U11032 (N_11032,N_9644,N_9338);
or U11033 (N_11033,N_10393,N_10226);
and U11034 (N_11034,N_9256,N_9275);
xor U11035 (N_11035,N_9328,N_9056);
or U11036 (N_11036,N_9958,N_10261);
or U11037 (N_11037,N_9407,N_9716);
nand U11038 (N_11038,N_9482,N_9439);
nor U11039 (N_11039,N_9903,N_10374);
or U11040 (N_11040,N_10368,N_9041);
nand U11041 (N_11041,N_9756,N_10215);
or U11042 (N_11042,N_10415,N_10016);
nand U11043 (N_11043,N_10358,N_9004);
nor U11044 (N_11044,N_9560,N_10050);
xor U11045 (N_11045,N_9887,N_9794);
or U11046 (N_11046,N_10192,N_10077);
or U11047 (N_11047,N_10383,N_10388);
and U11048 (N_11048,N_9705,N_9127);
xnor U11049 (N_11049,N_9252,N_9320);
nor U11050 (N_11050,N_9163,N_10402);
xor U11051 (N_11051,N_10118,N_9583);
or U11052 (N_11052,N_9225,N_9852);
nor U11053 (N_11053,N_9481,N_9369);
or U11054 (N_11054,N_9923,N_9178);
and U11055 (N_11055,N_10200,N_9270);
and U11056 (N_11056,N_10243,N_9635);
or U11057 (N_11057,N_9736,N_10496);
nor U11058 (N_11058,N_9592,N_10102);
and U11059 (N_11059,N_9357,N_10156);
nor U11060 (N_11060,N_9838,N_10296);
nand U11061 (N_11061,N_9156,N_9972);
or U11062 (N_11062,N_10452,N_9051);
or U11063 (N_11063,N_10328,N_9384);
xor U11064 (N_11064,N_9278,N_10236);
nand U11065 (N_11065,N_10456,N_9619);
or U11066 (N_11066,N_9245,N_10010);
nand U11067 (N_11067,N_10363,N_9925);
nor U11068 (N_11068,N_10398,N_9340);
and U11069 (N_11069,N_10187,N_9204);
or U11070 (N_11070,N_9783,N_10350);
and U11071 (N_11071,N_10404,N_9045);
nand U11072 (N_11072,N_9534,N_9788);
and U11073 (N_11073,N_9814,N_9371);
nand U11074 (N_11074,N_9831,N_10242);
and U11075 (N_11075,N_9989,N_9921);
and U11076 (N_11076,N_9621,N_9173);
nand U11077 (N_11077,N_9507,N_9034);
and U11078 (N_11078,N_10137,N_10250);
nor U11079 (N_11079,N_9627,N_9047);
xor U11080 (N_11080,N_10120,N_10275);
nor U11081 (N_11081,N_9579,N_9604);
and U11082 (N_11082,N_10343,N_9122);
nor U11083 (N_11083,N_9578,N_9200);
nand U11084 (N_11084,N_9496,N_9259);
nand U11085 (N_11085,N_9052,N_10222);
or U11086 (N_11086,N_9897,N_9941);
or U11087 (N_11087,N_9159,N_10354);
and U11088 (N_11088,N_9738,N_9614);
xor U11089 (N_11089,N_9785,N_9307);
or U11090 (N_11090,N_10380,N_10272);
nand U11091 (N_11091,N_10288,N_9464);
or U11092 (N_11092,N_10229,N_9348);
and U11093 (N_11093,N_9283,N_9829);
xnor U11094 (N_11094,N_9711,N_9470);
nor U11095 (N_11095,N_9023,N_9434);
nand U11096 (N_11096,N_10157,N_9054);
nand U11097 (N_11097,N_9558,N_10202);
or U11098 (N_11098,N_9715,N_9152);
or U11099 (N_11099,N_9839,N_9209);
nand U11100 (N_11100,N_10440,N_9007);
nand U11101 (N_11101,N_9429,N_9428);
or U11102 (N_11102,N_9457,N_9042);
nor U11103 (N_11103,N_9260,N_9775);
nand U11104 (N_11104,N_10284,N_10361);
or U11105 (N_11105,N_9789,N_9210);
or U11106 (N_11106,N_9841,N_10381);
nand U11107 (N_11107,N_9916,N_9898);
xor U11108 (N_11108,N_9821,N_9907);
xor U11109 (N_11109,N_9551,N_9448);
nand U11110 (N_11110,N_10224,N_9712);
or U11111 (N_11111,N_10332,N_9479);
nor U11112 (N_11112,N_9075,N_9985);
nor U11113 (N_11113,N_9262,N_10045);
xor U11114 (N_11114,N_9798,N_9404);
or U11115 (N_11115,N_10460,N_10094);
nand U11116 (N_11116,N_9295,N_9174);
xnor U11117 (N_11117,N_10256,N_9498);
nand U11118 (N_11118,N_9160,N_9580);
nor U11119 (N_11119,N_10127,N_9382);
and U11120 (N_11120,N_9900,N_9692);
xnor U11121 (N_11121,N_10114,N_10364);
or U11122 (N_11122,N_9424,N_9031);
nand U11123 (N_11123,N_9310,N_9090);
nor U11124 (N_11124,N_9996,N_9065);
nor U11125 (N_11125,N_9151,N_10039);
nand U11126 (N_11126,N_9752,N_10216);
nand U11127 (N_11127,N_9766,N_9196);
nand U11128 (N_11128,N_10003,N_9855);
and U11129 (N_11129,N_9510,N_9003);
and U11130 (N_11130,N_9884,N_10340);
nor U11131 (N_11131,N_9631,N_9486);
nand U11132 (N_11132,N_9860,N_10424);
or U11133 (N_11133,N_9891,N_10318);
or U11134 (N_11134,N_9447,N_9323);
or U11135 (N_11135,N_9021,N_9001);
nor U11136 (N_11136,N_10367,N_9267);
and U11137 (N_11137,N_9440,N_10337);
nor U11138 (N_11138,N_9508,N_9549);
or U11139 (N_11139,N_9707,N_9436);
xor U11140 (N_11140,N_9857,N_9118);
nand U11141 (N_11141,N_10090,N_9061);
and U11142 (N_11142,N_9834,N_9718);
nand U11143 (N_11143,N_10463,N_9288);
nand U11144 (N_11144,N_10459,N_9354);
or U11145 (N_11145,N_10267,N_9725);
nor U11146 (N_11146,N_10273,N_9870);
nand U11147 (N_11147,N_9332,N_9742);
and U11148 (N_11148,N_9570,N_9872);
and U11149 (N_11149,N_10081,N_9720);
nor U11150 (N_11150,N_9564,N_9244);
nor U11151 (N_11151,N_10166,N_10037);
xnor U11152 (N_11152,N_10178,N_9076);
xnor U11153 (N_11153,N_9469,N_9232);
or U11154 (N_11154,N_9097,N_9389);
nand U11155 (N_11155,N_10369,N_9319);
nand U11156 (N_11156,N_9346,N_9698);
nor U11157 (N_11157,N_9425,N_9694);
nand U11158 (N_11158,N_10133,N_9273);
or U11159 (N_11159,N_9819,N_10342);
nand U11160 (N_11160,N_9177,N_10197);
and U11161 (N_11161,N_10182,N_9911);
and U11162 (N_11162,N_9634,N_10027);
xnor U11163 (N_11163,N_9223,N_9422);
and U11164 (N_11164,N_10303,N_9433);
and U11165 (N_11165,N_9892,N_9545);
and U11166 (N_11166,N_9886,N_9759);
and U11167 (N_11167,N_9912,N_9128);
nor U11168 (N_11168,N_9861,N_10038);
nand U11169 (N_11169,N_10372,N_10162);
nand U11170 (N_11170,N_9729,N_9138);
nand U11171 (N_11171,N_10290,N_10442);
nor U11172 (N_11172,N_10325,N_9979);
xnor U11173 (N_11173,N_9095,N_9557);
or U11174 (N_11174,N_10249,N_9403);
and U11175 (N_11175,N_9221,N_9528);
nor U11176 (N_11176,N_9520,N_10136);
nand U11177 (N_11177,N_10432,N_9205);
xnor U11178 (N_11178,N_9875,N_9563);
xnor U11179 (N_11179,N_9492,N_10353);
nor U11180 (N_11180,N_9091,N_10286);
and U11181 (N_11181,N_10471,N_10174);
nand U11182 (N_11182,N_9593,N_9048);
or U11183 (N_11183,N_9098,N_9740);
nor U11184 (N_11184,N_9603,N_10352);
xnor U11185 (N_11185,N_9774,N_9760);
nor U11186 (N_11186,N_10025,N_10244);
and U11187 (N_11187,N_9000,N_9101);
and U11188 (N_11188,N_9704,N_9192);
nor U11189 (N_11189,N_10221,N_10046);
or U11190 (N_11190,N_9899,N_9070);
xnor U11191 (N_11191,N_9366,N_10177);
nor U11192 (N_11192,N_9370,N_9014);
and U11193 (N_11193,N_9092,N_9944);
xor U11194 (N_11194,N_10099,N_9104);
nor U11195 (N_11195,N_9015,N_10170);
xor U11196 (N_11196,N_9747,N_10205);
nand U11197 (N_11197,N_10163,N_9673);
and U11198 (N_11198,N_10341,N_9791);
nor U11199 (N_11199,N_9577,N_10412);
nand U11200 (N_11200,N_10051,N_10307);
nand U11201 (N_11201,N_9309,N_9754);
and U11202 (N_11202,N_9645,N_10311);
nand U11203 (N_11203,N_9272,N_9820);
nor U11204 (N_11204,N_9039,N_9069);
and U11205 (N_11205,N_9294,N_9866);
nand U11206 (N_11206,N_9951,N_9167);
nor U11207 (N_11207,N_9471,N_10085);
or U11208 (N_11208,N_9678,N_9304);
nor U11209 (N_11209,N_10103,N_9291);
xor U11210 (N_11210,N_9815,N_10184);
nor U11211 (N_11211,N_10029,N_10297);
xor U11212 (N_11212,N_10062,N_10108);
nor U11213 (N_11213,N_9904,N_10066);
nor U11214 (N_11214,N_9932,N_9183);
nor U11215 (N_11215,N_10007,N_10265);
and U11216 (N_11216,N_9827,N_9500);
and U11217 (N_11217,N_10408,N_9390);
and U11218 (N_11218,N_9417,N_9781);
nor U11219 (N_11219,N_10089,N_9233);
xor U11220 (N_11220,N_9864,N_10427);
or U11221 (N_11221,N_10240,N_9728);
nor U11222 (N_11222,N_10160,N_9546);
nor U11223 (N_11223,N_9314,N_9182);
nor U11224 (N_11224,N_9242,N_9667);
or U11225 (N_11225,N_10324,N_9279);
and U11226 (N_11226,N_9565,N_10237);
nand U11227 (N_11227,N_10172,N_9064);
and U11228 (N_11228,N_9938,N_9840);
nand U11229 (N_11229,N_9060,N_9795);
or U11230 (N_11230,N_9249,N_9079);
nor U11231 (N_11231,N_9539,N_9710);
xor U11232 (N_11232,N_9765,N_9011);
xor U11233 (N_11233,N_10238,N_9120);
xnor U11234 (N_11234,N_9856,N_9462);
xnor U11235 (N_11235,N_9058,N_9379);
and U11236 (N_11236,N_10059,N_9458);
nor U11237 (N_11237,N_10033,N_10485);
nor U11238 (N_11238,N_10245,N_9117);
nand U11239 (N_11239,N_10072,N_9735);
nand U11240 (N_11240,N_10115,N_10057);
nand U11241 (N_11241,N_10392,N_9368);
and U11242 (N_11242,N_9085,N_10095);
and U11243 (N_11243,N_10405,N_9503);
xor U11244 (N_11244,N_10385,N_9387);
nand U11245 (N_11245,N_9111,N_9585);
nand U11246 (N_11246,N_9261,N_9988);
nand U11247 (N_11247,N_9588,N_10180);
or U11248 (N_11248,N_10065,N_9618);
nand U11249 (N_11249,N_10168,N_9377);
or U11250 (N_11250,N_10193,N_9081);
xor U11251 (N_11251,N_9550,N_10298);
nor U11252 (N_11252,N_10173,N_10391);
or U11253 (N_11253,N_9324,N_9462);
or U11254 (N_11254,N_10161,N_9701);
xnor U11255 (N_11255,N_9590,N_9037);
nand U11256 (N_11256,N_9668,N_10255);
nand U11257 (N_11257,N_10005,N_9931);
and U11258 (N_11258,N_10485,N_9663);
or U11259 (N_11259,N_10106,N_10107);
or U11260 (N_11260,N_10130,N_9994);
and U11261 (N_11261,N_10217,N_10239);
and U11262 (N_11262,N_9660,N_9103);
nor U11263 (N_11263,N_9252,N_10169);
or U11264 (N_11264,N_9007,N_9034);
and U11265 (N_11265,N_9902,N_9155);
or U11266 (N_11266,N_10079,N_10218);
nand U11267 (N_11267,N_9668,N_9611);
nand U11268 (N_11268,N_9374,N_9887);
nand U11269 (N_11269,N_10358,N_10333);
xor U11270 (N_11270,N_9104,N_10053);
or U11271 (N_11271,N_10061,N_9140);
nor U11272 (N_11272,N_9945,N_9633);
or U11273 (N_11273,N_9418,N_10291);
nor U11274 (N_11274,N_9477,N_9818);
and U11275 (N_11275,N_9065,N_9345);
and U11276 (N_11276,N_9957,N_10217);
and U11277 (N_11277,N_9393,N_9488);
nand U11278 (N_11278,N_9824,N_9577);
or U11279 (N_11279,N_9206,N_10248);
nor U11280 (N_11280,N_9488,N_10200);
nand U11281 (N_11281,N_9552,N_9766);
xor U11282 (N_11282,N_10301,N_9929);
xor U11283 (N_11283,N_9123,N_9878);
xnor U11284 (N_11284,N_9446,N_9622);
nand U11285 (N_11285,N_10293,N_9474);
or U11286 (N_11286,N_9730,N_9412);
xor U11287 (N_11287,N_9178,N_9530);
and U11288 (N_11288,N_9947,N_9732);
or U11289 (N_11289,N_10258,N_9518);
or U11290 (N_11290,N_9322,N_10272);
and U11291 (N_11291,N_9362,N_9966);
and U11292 (N_11292,N_10134,N_9113);
or U11293 (N_11293,N_10447,N_9141);
or U11294 (N_11294,N_9059,N_9318);
or U11295 (N_11295,N_9813,N_9527);
xnor U11296 (N_11296,N_9820,N_10486);
or U11297 (N_11297,N_10457,N_9441);
nand U11298 (N_11298,N_9684,N_9965);
or U11299 (N_11299,N_10352,N_10000);
xor U11300 (N_11300,N_10470,N_9216);
xnor U11301 (N_11301,N_9284,N_9783);
nand U11302 (N_11302,N_10248,N_9746);
nand U11303 (N_11303,N_9449,N_10346);
and U11304 (N_11304,N_10415,N_9705);
nor U11305 (N_11305,N_9823,N_10191);
nand U11306 (N_11306,N_10080,N_9597);
xnor U11307 (N_11307,N_9612,N_10463);
or U11308 (N_11308,N_9948,N_10497);
or U11309 (N_11309,N_9770,N_9756);
and U11310 (N_11310,N_9871,N_9404);
nor U11311 (N_11311,N_10004,N_9726);
nand U11312 (N_11312,N_10171,N_9648);
nand U11313 (N_11313,N_10130,N_9618);
nand U11314 (N_11314,N_9284,N_10068);
and U11315 (N_11315,N_9040,N_10084);
nor U11316 (N_11316,N_10090,N_10082);
or U11317 (N_11317,N_10040,N_10080);
nand U11318 (N_11318,N_9208,N_10066);
or U11319 (N_11319,N_9683,N_9392);
and U11320 (N_11320,N_9914,N_9504);
nand U11321 (N_11321,N_10468,N_10366);
or U11322 (N_11322,N_9145,N_9140);
and U11323 (N_11323,N_9106,N_9260);
nor U11324 (N_11324,N_9795,N_9617);
nor U11325 (N_11325,N_9393,N_9013);
and U11326 (N_11326,N_9593,N_10096);
or U11327 (N_11327,N_10135,N_10309);
and U11328 (N_11328,N_10038,N_9117);
xor U11329 (N_11329,N_9640,N_9251);
xor U11330 (N_11330,N_9125,N_10305);
nor U11331 (N_11331,N_9088,N_9805);
nand U11332 (N_11332,N_10436,N_10363);
nand U11333 (N_11333,N_10395,N_9649);
or U11334 (N_11334,N_9413,N_9153);
nand U11335 (N_11335,N_9763,N_9230);
or U11336 (N_11336,N_9218,N_9989);
and U11337 (N_11337,N_10411,N_10358);
and U11338 (N_11338,N_9371,N_10328);
nor U11339 (N_11339,N_10480,N_10184);
and U11340 (N_11340,N_9106,N_9002);
xor U11341 (N_11341,N_9488,N_9209);
and U11342 (N_11342,N_9684,N_9516);
nand U11343 (N_11343,N_9218,N_9437);
xor U11344 (N_11344,N_9547,N_9809);
nand U11345 (N_11345,N_9936,N_10228);
or U11346 (N_11346,N_10424,N_9569);
and U11347 (N_11347,N_9816,N_10229);
or U11348 (N_11348,N_10209,N_10337);
and U11349 (N_11349,N_10082,N_10473);
xor U11350 (N_11350,N_10318,N_10187);
nor U11351 (N_11351,N_10089,N_9342);
nor U11352 (N_11352,N_10070,N_9133);
xnor U11353 (N_11353,N_10415,N_9391);
nand U11354 (N_11354,N_10441,N_10203);
nor U11355 (N_11355,N_9487,N_9568);
nor U11356 (N_11356,N_9426,N_10309);
xnor U11357 (N_11357,N_9894,N_10279);
xnor U11358 (N_11358,N_9233,N_10352);
nor U11359 (N_11359,N_10399,N_10107);
nand U11360 (N_11360,N_9834,N_10079);
and U11361 (N_11361,N_9633,N_9150);
nand U11362 (N_11362,N_9605,N_9473);
nand U11363 (N_11363,N_9406,N_10132);
nand U11364 (N_11364,N_9622,N_10142);
xnor U11365 (N_11365,N_9471,N_9299);
and U11366 (N_11366,N_10422,N_9165);
nor U11367 (N_11367,N_9062,N_9158);
xor U11368 (N_11368,N_9036,N_10333);
nand U11369 (N_11369,N_9915,N_9818);
xor U11370 (N_11370,N_9306,N_9100);
and U11371 (N_11371,N_10230,N_10034);
or U11372 (N_11372,N_9007,N_10008);
nand U11373 (N_11373,N_10281,N_10040);
xor U11374 (N_11374,N_9401,N_10009);
or U11375 (N_11375,N_9942,N_9606);
nor U11376 (N_11376,N_10425,N_9062);
xnor U11377 (N_11377,N_9421,N_10438);
nor U11378 (N_11378,N_9563,N_9919);
nor U11379 (N_11379,N_10429,N_10404);
or U11380 (N_11380,N_10000,N_9765);
or U11381 (N_11381,N_10142,N_9145);
and U11382 (N_11382,N_9309,N_9345);
xnor U11383 (N_11383,N_9263,N_9059);
or U11384 (N_11384,N_9898,N_9007);
and U11385 (N_11385,N_10105,N_10053);
nand U11386 (N_11386,N_10462,N_9060);
and U11387 (N_11387,N_9395,N_9146);
xnor U11388 (N_11388,N_9488,N_9875);
or U11389 (N_11389,N_9611,N_10242);
and U11390 (N_11390,N_9446,N_9589);
xnor U11391 (N_11391,N_10411,N_9966);
xor U11392 (N_11392,N_9825,N_9970);
xor U11393 (N_11393,N_10438,N_9589);
or U11394 (N_11394,N_9869,N_9593);
nand U11395 (N_11395,N_9155,N_9465);
xor U11396 (N_11396,N_10218,N_10243);
xor U11397 (N_11397,N_10277,N_10020);
nand U11398 (N_11398,N_10099,N_9159);
nand U11399 (N_11399,N_10037,N_10358);
or U11400 (N_11400,N_9340,N_9124);
nor U11401 (N_11401,N_9754,N_9756);
or U11402 (N_11402,N_9927,N_9168);
xor U11403 (N_11403,N_10363,N_9541);
xnor U11404 (N_11404,N_10071,N_9034);
nand U11405 (N_11405,N_9903,N_10068);
nor U11406 (N_11406,N_10103,N_10222);
and U11407 (N_11407,N_9360,N_9397);
or U11408 (N_11408,N_10081,N_9481);
nor U11409 (N_11409,N_9843,N_10326);
xnor U11410 (N_11410,N_10366,N_9734);
nand U11411 (N_11411,N_9646,N_9636);
nor U11412 (N_11412,N_9939,N_10138);
xor U11413 (N_11413,N_9252,N_9710);
xnor U11414 (N_11414,N_9806,N_9127);
and U11415 (N_11415,N_9402,N_10406);
or U11416 (N_11416,N_10362,N_9694);
xor U11417 (N_11417,N_9516,N_9471);
or U11418 (N_11418,N_9596,N_9335);
nand U11419 (N_11419,N_10183,N_9577);
or U11420 (N_11420,N_10472,N_9524);
and U11421 (N_11421,N_9117,N_9236);
xor U11422 (N_11422,N_9239,N_10057);
nor U11423 (N_11423,N_9349,N_9680);
nor U11424 (N_11424,N_9534,N_9702);
or U11425 (N_11425,N_10152,N_9270);
nand U11426 (N_11426,N_10237,N_10189);
nor U11427 (N_11427,N_10025,N_10128);
nand U11428 (N_11428,N_9116,N_9372);
and U11429 (N_11429,N_9177,N_10150);
nor U11430 (N_11430,N_10113,N_10386);
nand U11431 (N_11431,N_9758,N_9361);
and U11432 (N_11432,N_9573,N_10426);
xor U11433 (N_11433,N_9830,N_10048);
or U11434 (N_11434,N_9947,N_9073);
nand U11435 (N_11435,N_9339,N_9640);
nor U11436 (N_11436,N_9759,N_10319);
xnor U11437 (N_11437,N_9666,N_9570);
or U11438 (N_11438,N_10427,N_10108);
nand U11439 (N_11439,N_9700,N_9402);
or U11440 (N_11440,N_10015,N_9797);
and U11441 (N_11441,N_9492,N_9683);
and U11442 (N_11442,N_10325,N_9311);
xor U11443 (N_11443,N_9090,N_9140);
or U11444 (N_11444,N_9652,N_9155);
nor U11445 (N_11445,N_9222,N_10134);
nor U11446 (N_11446,N_9738,N_9511);
or U11447 (N_11447,N_10148,N_9922);
xor U11448 (N_11448,N_9016,N_9101);
or U11449 (N_11449,N_9758,N_9348);
and U11450 (N_11450,N_9634,N_10356);
nor U11451 (N_11451,N_9226,N_9478);
nand U11452 (N_11452,N_10209,N_10424);
nor U11453 (N_11453,N_9003,N_10409);
nand U11454 (N_11454,N_9968,N_9260);
and U11455 (N_11455,N_9342,N_9678);
and U11456 (N_11456,N_9056,N_10490);
nor U11457 (N_11457,N_9517,N_10156);
xnor U11458 (N_11458,N_10092,N_9755);
and U11459 (N_11459,N_9504,N_9850);
nand U11460 (N_11460,N_9676,N_10255);
and U11461 (N_11461,N_10390,N_9322);
nor U11462 (N_11462,N_10376,N_9216);
nand U11463 (N_11463,N_10148,N_9630);
nand U11464 (N_11464,N_9626,N_9123);
xor U11465 (N_11465,N_10166,N_9501);
xor U11466 (N_11466,N_10463,N_10372);
nand U11467 (N_11467,N_9019,N_9445);
nor U11468 (N_11468,N_9676,N_10462);
nor U11469 (N_11469,N_9389,N_9555);
or U11470 (N_11470,N_10144,N_9777);
or U11471 (N_11471,N_10146,N_9901);
xor U11472 (N_11472,N_10491,N_9732);
nor U11473 (N_11473,N_9127,N_10179);
and U11474 (N_11474,N_9189,N_9937);
nor U11475 (N_11475,N_9056,N_10270);
nor U11476 (N_11476,N_9394,N_10340);
nand U11477 (N_11477,N_9713,N_9402);
nand U11478 (N_11478,N_9560,N_9018);
xor U11479 (N_11479,N_10148,N_9974);
xnor U11480 (N_11480,N_9496,N_10072);
nand U11481 (N_11481,N_9135,N_9446);
nor U11482 (N_11482,N_9015,N_9943);
nor U11483 (N_11483,N_9646,N_10320);
or U11484 (N_11484,N_9365,N_10186);
nand U11485 (N_11485,N_9028,N_9488);
xnor U11486 (N_11486,N_9027,N_10267);
nand U11487 (N_11487,N_10459,N_9725);
and U11488 (N_11488,N_9608,N_9548);
nor U11489 (N_11489,N_10434,N_9584);
xnor U11490 (N_11490,N_10054,N_9804);
and U11491 (N_11491,N_9990,N_10423);
nor U11492 (N_11492,N_9148,N_9481);
xnor U11493 (N_11493,N_10413,N_9451);
or U11494 (N_11494,N_10095,N_10346);
and U11495 (N_11495,N_9169,N_9226);
xnor U11496 (N_11496,N_9857,N_9574);
or U11497 (N_11497,N_9735,N_9784);
nor U11498 (N_11498,N_10438,N_9993);
nand U11499 (N_11499,N_10054,N_9491);
nor U11500 (N_11500,N_9629,N_9847);
nor U11501 (N_11501,N_9397,N_9815);
xor U11502 (N_11502,N_10163,N_9810);
and U11503 (N_11503,N_9739,N_10377);
xor U11504 (N_11504,N_9470,N_9713);
and U11505 (N_11505,N_10470,N_10393);
and U11506 (N_11506,N_10264,N_9134);
xnor U11507 (N_11507,N_9843,N_9464);
nand U11508 (N_11508,N_10002,N_9946);
nor U11509 (N_11509,N_10195,N_10435);
or U11510 (N_11510,N_9623,N_10366);
or U11511 (N_11511,N_9146,N_10365);
or U11512 (N_11512,N_10067,N_10035);
xnor U11513 (N_11513,N_9251,N_10151);
nor U11514 (N_11514,N_9582,N_9735);
or U11515 (N_11515,N_9331,N_9143);
or U11516 (N_11516,N_10074,N_9758);
nand U11517 (N_11517,N_10285,N_9020);
xor U11518 (N_11518,N_9675,N_10364);
xnor U11519 (N_11519,N_9042,N_9416);
nand U11520 (N_11520,N_10389,N_9848);
xnor U11521 (N_11521,N_9407,N_9382);
xor U11522 (N_11522,N_9065,N_10268);
or U11523 (N_11523,N_10105,N_9028);
nand U11524 (N_11524,N_9530,N_9023);
or U11525 (N_11525,N_9648,N_9100);
xor U11526 (N_11526,N_10398,N_9055);
or U11527 (N_11527,N_10088,N_10135);
and U11528 (N_11528,N_9873,N_10076);
xor U11529 (N_11529,N_9628,N_9230);
and U11530 (N_11530,N_9141,N_9899);
nor U11531 (N_11531,N_10201,N_10212);
nor U11532 (N_11532,N_10218,N_9411);
or U11533 (N_11533,N_10354,N_10243);
xnor U11534 (N_11534,N_10325,N_9317);
and U11535 (N_11535,N_10372,N_9394);
and U11536 (N_11536,N_9962,N_9215);
or U11537 (N_11537,N_9092,N_9327);
and U11538 (N_11538,N_10353,N_10431);
xnor U11539 (N_11539,N_9464,N_9588);
or U11540 (N_11540,N_10499,N_10157);
nor U11541 (N_11541,N_9688,N_9069);
or U11542 (N_11542,N_9529,N_9313);
nand U11543 (N_11543,N_9015,N_9688);
and U11544 (N_11544,N_10425,N_10378);
nor U11545 (N_11545,N_9149,N_9318);
and U11546 (N_11546,N_9548,N_10241);
nand U11547 (N_11547,N_9832,N_9250);
nor U11548 (N_11548,N_9777,N_9734);
nor U11549 (N_11549,N_10337,N_9560);
nor U11550 (N_11550,N_9421,N_9550);
nand U11551 (N_11551,N_9463,N_9149);
or U11552 (N_11552,N_10055,N_9612);
xor U11553 (N_11553,N_9196,N_10443);
xor U11554 (N_11554,N_10343,N_9096);
nand U11555 (N_11555,N_9722,N_9809);
xnor U11556 (N_11556,N_10274,N_9003);
nor U11557 (N_11557,N_9359,N_9867);
xnor U11558 (N_11558,N_9997,N_10417);
or U11559 (N_11559,N_9851,N_9457);
and U11560 (N_11560,N_9564,N_9548);
and U11561 (N_11561,N_10392,N_10202);
nand U11562 (N_11562,N_10139,N_9417);
nor U11563 (N_11563,N_10028,N_10479);
xor U11564 (N_11564,N_9824,N_9458);
nor U11565 (N_11565,N_10077,N_9581);
and U11566 (N_11566,N_9029,N_9020);
and U11567 (N_11567,N_10483,N_9093);
or U11568 (N_11568,N_9752,N_9239);
or U11569 (N_11569,N_10219,N_9938);
or U11570 (N_11570,N_10099,N_9234);
or U11571 (N_11571,N_9469,N_9077);
nand U11572 (N_11572,N_9013,N_9883);
or U11573 (N_11573,N_10479,N_9345);
xor U11574 (N_11574,N_9738,N_10022);
xor U11575 (N_11575,N_9129,N_9124);
or U11576 (N_11576,N_9151,N_9733);
xnor U11577 (N_11577,N_9345,N_10224);
and U11578 (N_11578,N_9197,N_10400);
nor U11579 (N_11579,N_9506,N_10233);
xnor U11580 (N_11580,N_10319,N_9976);
and U11581 (N_11581,N_10315,N_9156);
or U11582 (N_11582,N_9389,N_9051);
and U11583 (N_11583,N_9197,N_9428);
nand U11584 (N_11584,N_9115,N_9925);
nand U11585 (N_11585,N_9226,N_10047);
xor U11586 (N_11586,N_10368,N_10163);
nand U11587 (N_11587,N_10248,N_10442);
and U11588 (N_11588,N_9147,N_10087);
and U11589 (N_11589,N_10045,N_9686);
xor U11590 (N_11590,N_9336,N_9711);
or U11591 (N_11591,N_9160,N_10015);
and U11592 (N_11592,N_9116,N_9730);
nor U11593 (N_11593,N_9064,N_9827);
xor U11594 (N_11594,N_10075,N_9165);
or U11595 (N_11595,N_10446,N_9490);
nand U11596 (N_11596,N_10164,N_9467);
nand U11597 (N_11597,N_9274,N_9138);
nor U11598 (N_11598,N_9700,N_9985);
xnor U11599 (N_11599,N_9871,N_9753);
and U11600 (N_11600,N_9867,N_9727);
or U11601 (N_11601,N_9261,N_9129);
nand U11602 (N_11602,N_9043,N_10009);
xor U11603 (N_11603,N_10342,N_10089);
nor U11604 (N_11604,N_9404,N_9208);
nand U11605 (N_11605,N_9932,N_10098);
and U11606 (N_11606,N_9069,N_10279);
xor U11607 (N_11607,N_9593,N_9257);
xnor U11608 (N_11608,N_9657,N_10150);
or U11609 (N_11609,N_9217,N_9257);
nand U11610 (N_11610,N_9031,N_9554);
xnor U11611 (N_11611,N_9059,N_9843);
nand U11612 (N_11612,N_9677,N_9414);
nor U11613 (N_11613,N_9118,N_10457);
nor U11614 (N_11614,N_9575,N_9439);
nor U11615 (N_11615,N_9207,N_9948);
and U11616 (N_11616,N_10131,N_9894);
nor U11617 (N_11617,N_9704,N_10453);
and U11618 (N_11618,N_10327,N_10499);
nand U11619 (N_11619,N_9899,N_9693);
xor U11620 (N_11620,N_9020,N_9108);
or U11621 (N_11621,N_9024,N_9482);
xor U11622 (N_11622,N_9781,N_9426);
and U11623 (N_11623,N_9864,N_9472);
and U11624 (N_11624,N_10192,N_9086);
or U11625 (N_11625,N_9521,N_9648);
and U11626 (N_11626,N_10238,N_10185);
nor U11627 (N_11627,N_9205,N_9448);
or U11628 (N_11628,N_9816,N_9748);
nor U11629 (N_11629,N_9203,N_9488);
xor U11630 (N_11630,N_9305,N_10342);
xor U11631 (N_11631,N_9405,N_9778);
xnor U11632 (N_11632,N_10484,N_9982);
nor U11633 (N_11633,N_9735,N_9254);
nand U11634 (N_11634,N_10491,N_9901);
xor U11635 (N_11635,N_9613,N_9302);
nor U11636 (N_11636,N_9351,N_9643);
or U11637 (N_11637,N_10107,N_9102);
or U11638 (N_11638,N_9191,N_9252);
nor U11639 (N_11639,N_10330,N_9554);
or U11640 (N_11640,N_10273,N_9223);
or U11641 (N_11641,N_10146,N_9818);
xnor U11642 (N_11642,N_9665,N_10202);
or U11643 (N_11643,N_9031,N_9998);
and U11644 (N_11644,N_9776,N_10360);
xnor U11645 (N_11645,N_10340,N_9799);
and U11646 (N_11646,N_10329,N_9636);
nor U11647 (N_11647,N_9175,N_10494);
nand U11648 (N_11648,N_9547,N_10063);
or U11649 (N_11649,N_9168,N_9983);
nor U11650 (N_11650,N_9063,N_10369);
nor U11651 (N_11651,N_10215,N_9152);
nor U11652 (N_11652,N_10149,N_9167);
nor U11653 (N_11653,N_9601,N_10041);
and U11654 (N_11654,N_10401,N_9241);
or U11655 (N_11655,N_10121,N_9832);
or U11656 (N_11656,N_9243,N_10206);
and U11657 (N_11657,N_10429,N_10257);
or U11658 (N_11658,N_10437,N_9241);
or U11659 (N_11659,N_10365,N_9090);
nor U11660 (N_11660,N_10005,N_9980);
and U11661 (N_11661,N_9604,N_10054);
nor U11662 (N_11662,N_10063,N_9801);
xor U11663 (N_11663,N_9940,N_9137);
xnor U11664 (N_11664,N_10036,N_9166);
nor U11665 (N_11665,N_9114,N_10175);
nor U11666 (N_11666,N_9413,N_10250);
and U11667 (N_11667,N_9742,N_9060);
and U11668 (N_11668,N_9725,N_9331);
xnor U11669 (N_11669,N_10219,N_9091);
nand U11670 (N_11670,N_9108,N_9557);
or U11671 (N_11671,N_9432,N_10185);
nand U11672 (N_11672,N_9200,N_10428);
xnor U11673 (N_11673,N_9783,N_10406);
nor U11674 (N_11674,N_9702,N_10112);
and U11675 (N_11675,N_10267,N_9935);
xor U11676 (N_11676,N_9433,N_9780);
nor U11677 (N_11677,N_9593,N_9244);
nand U11678 (N_11678,N_9821,N_9807);
xor U11679 (N_11679,N_9340,N_9087);
nor U11680 (N_11680,N_10368,N_9643);
nand U11681 (N_11681,N_9450,N_9973);
or U11682 (N_11682,N_10058,N_9869);
or U11683 (N_11683,N_9139,N_9363);
xnor U11684 (N_11684,N_9671,N_9090);
nor U11685 (N_11685,N_10198,N_9708);
or U11686 (N_11686,N_9772,N_10145);
nand U11687 (N_11687,N_10060,N_9534);
and U11688 (N_11688,N_9333,N_10396);
or U11689 (N_11689,N_10492,N_9145);
xor U11690 (N_11690,N_9436,N_10185);
and U11691 (N_11691,N_10366,N_9545);
and U11692 (N_11692,N_9579,N_9177);
nand U11693 (N_11693,N_9748,N_10484);
and U11694 (N_11694,N_10268,N_9327);
nor U11695 (N_11695,N_9326,N_9981);
nand U11696 (N_11696,N_9529,N_10162);
nor U11697 (N_11697,N_9662,N_10117);
nand U11698 (N_11698,N_9774,N_9844);
or U11699 (N_11699,N_10332,N_9884);
xnor U11700 (N_11700,N_9120,N_10122);
nor U11701 (N_11701,N_9078,N_10459);
nor U11702 (N_11702,N_10217,N_9393);
nand U11703 (N_11703,N_9585,N_9072);
nand U11704 (N_11704,N_9825,N_10160);
and U11705 (N_11705,N_9861,N_9101);
or U11706 (N_11706,N_9365,N_9052);
nor U11707 (N_11707,N_9008,N_10335);
and U11708 (N_11708,N_10308,N_9090);
xnor U11709 (N_11709,N_9503,N_9176);
and U11710 (N_11710,N_9368,N_9555);
nor U11711 (N_11711,N_10436,N_10205);
xor U11712 (N_11712,N_9869,N_10436);
or U11713 (N_11713,N_9758,N_9882);
xor U11714 (N_11714,N_9112,N_10479);
xnor U11715 (N_11715,N_9641,N_9235);
xor U11716 (N_11716,N_10269,N_9593);
xor U11717 (N_11717,N_10078,N_10060);
xor U11718 (N_11718,N_9435,N_10161);
nand U11719 (N_11719,N_9315,N_9029);
or U11720 (N_11720,N_9132,N_9468);
nor U11721 (N_11721,N_10175,N_9284);
xor U11722 (N_11722,N_10197,N_9916);
nand U11723 (N_11723,N_10140,N_9313);
and U11724 (N_11724,N_9376,N_9489);
or U11725 (N_11725,N_9154,N_9035);
nor U11726 (N_11726,N_9125,N_10041);
nand U11727 (N_11727,N_9322,N_9262);
nand U11728 (N_11728,N_9595,N_10148);
and U11729 (N_11729,N_9851,N_10137);
nor U11730 (N_11730,N_9175,N_10077);
xor U11731 (N_11731,N_9897,N_9840);
nand U11732 (N_11732,N_9979,N_10257);
and U11733 (N_11733,N_10096,N_9402);
and U11734 (N_11734,N_10478,N_9457);
and U11735 (N_11735,N_9589,N_9569);
nand U11736 (N_11736,N_9534,N_9225);
or U11737 (N_11737,N_9545,N_9672);
xnor U11738 (N_11738,N_9956,N_9453);
and U11739 (N_11739,N_10217,N_9929);
and U11740 (N_11740,N_9249,N_9353);
and U11741 (N_11741,N_10407,N_9311);
or U11742 (N_11742,N_9692,N_9075);
nor U11743 (N_11743,N_9612,N_9759);
nor U11744 (N_11744,N_9240,N_10305);
and U11745 (N_11745,N_10040,N_9208);
nor U11746 (N_11746,N_9044,N_10315);
nor U11747 (N_11747,N_10010,N_9867);
nor U11748 (N_11748,N_9211,N_9722);
and U11749 (N_11749,N_9435,N_9457);
and U11750 (N_11750,N_9658,N_10106);
nor U11751 (N_11751,N_10318,N_10009);
nor U11752 (N_11752,N_10419,N_9798);
nand U11753 (N_11753,N_9172,N_10123);
nor U11754 (N_11754,N_9110,N_9530);
nand U11755 (N_11755,N_9885,N_9701);
nand U11756 (N_11756,N_9220,N_9717);
and U11757 (N_11757,N_9117,N_10029);
xor U11758 (N_11758,N_9013,N_9966);
and U11759 (N_11759,N_9581,N_10195);
or U11760 (N_11760,N_9736,N_9496);
xor U11761 (N_11761,N_9694,N_9588);
xnor U11762 (N_11762,N_9726,N_9007);
nand U11763 (N_11763,N_9939,N_9772);
xnor U11764 (N_11764,N_10060,N_9235);
nor U11765 (N_11765,N_10306,N_9892);
nor U11766 (N_11766,N_9419,N_9377);
nand U11767 (N_11767,N_9947,N_10026);
nand U11768 (N_11768,N_9907,N_9490);
nand U11769 (N_11769,N_10230,N_9479);
nor U11770 (N_11770,N_9839,N_9353);
nand U11771 (N_11771,N_9477,N_9377);
nand U11772 (N_11772,N_10042,N_10278);
nor U11773 (N_11773,N_9576,N_9147);
xnor U11774 (N_11774,N_9343,N_9961);
xor U11775 (N_11775,N_10381,N_10432);
nand U11776 (N_11776,N_9730,N_9530);
nor U11777 (N_11777,N_10298,N_9043);
xor U11778 (N_11778,N_10480,N_9274);
and U11779 (N_11779,N_9654,N_9733);
and U11780 (N_11780,N_9204,N_9925);
or U11781 (N_11781,N_9631,N_9916);
nand U11782 (N_11782,N_9885,N_9363);
nor U11783 (N_11783,N_9316,N_9946);
nand U11784 (N_11784,N_10471,N_9675);
nand U11785 (N_11785,N_9971,N_9424);
nor U11786 (N_11786,N_9258,N_10357);
nand U11787 (N_11787,N_9874,N_9196);
or U11788 (N_11788,N_10012,N_10354);
nor U11789 (N_11789,N_10495,N_10196);
and U11790 (N_11790,N_9959,N_9301);
or U11791 (N_11791,N_10244,N_9749);
and U11792 (N_11792,N_9514,N_9407);
nor U11793 (N_11793,N_9045,N_9854);
xnor U11794 (N_11794,N_10267,N_10132);
xor U11795 (N_11795,N_9579,N_9997);
xor U11796 (N_11796,N_9375,N_10333);
and U11797 (N_11797,N_9429,N_9784);
nand U11798 (N_11798,N_9333,N_9125);
or U11799 (N_11799,N_9109,N_9572);
nor U11800 (N_11800,N_9966,N_9474);
xnor U11801 (N_11801,N_10281,N_9319);
nand U11802 (N_11802,N_9595,N_9201);
nor U11803 (N_11803,N_9409,N_9290);
xor U11804 (N_11804,N_10209,N_9281);
xor U11805 (N_11805,N_10392,N_9466);
nand U11806 (N_11806,N_9351,N_10356);
nand U11807 (N_11807,N_9142,N_9510);
xor U11808 (N_11808,N_9117,N_9433);
and U11809 (N_11809,N_10470,N_9653);
xor U11810 (N_11810,N_9499,N_9240);
nor U11811 (N_11811,N_10491,N_9981);
xnor U11812 (N_11812,N_9377,N_10463);
and U11813 (N_11813,N_9452,N_9747);
xnor U11814 (N_11814,N_9194,N_10206);
xnor U11815 (N_11815,N_10035,N_9239);
nor U11816 (N_11816,N_9651,N_10460);
nor U11817 (N_11817,N_9686,N_9906);
and U11818 (N_11818,N_9769,N_9506);
xor U11819 (N_11819,N_9711,N_9656);
and U11820 (N_11820,N_9985,N_9363);
or U11821 (N_11821,N_9005,N_10334);
or U11822 (N_11822,N_9240,N_9536);
nor U11823 (N_11823,N_9892,N_9085);
nand U11824 (N_11824,N_9113,N_10120);
nor U11825 (N_11825,N_9577,N_9489);
and U11826 (N_11826,N_9693,N_10205);
nor U11827 (N_11827,N_9138,N_9071);
and U11828 (N_11828,N_10066,N_9319);
xor U11829 (N_11829,N_9184,N_10477);
nand U11830 (N_11830,N_9271,N_10430);
and U11831 (N_11831,N_10412,N_10378);
and U11832 (N_11832,N_10025,N_10088);
or U11833 (N_11833,N_9119,N_10351);
xor U11834 (N_11834,N_10270,N_9545);
nand U11835 (N_11835,N_9001,N_10126);
xnor U11836 (N_11836,N_10419,N_9732);
or U11837 (N_11837,N_10334,N_10164);
or U11838 (N_11838,N_9358,N_10364);
xnor U11839 (N_11839,N_9848,N_9864);
or U11840 (N_11840,N_10259,N_9853);
and U11841 (N_11841,N_10198,N_9648);
nor U11842 (N_11842,N_9237,N_10047);
and U11843 (N_11843,N_9234,N_10209);
xnor U11844 (N_11844,N_10010,N_10226);
xor U11845 (N_11845,N_9716,N_10026);
xor U11846 (N_11846,N_9631,N_10091);
xnor U11847 (N_11847,N_10303,N_9516);
xnor U11848 (N_11848,N_9553,N_9589);
or U11849 (N_11849,N_9423,N_10202);
xor U11850 (N_11850,N_9319,N_10233);
nor U11851 (N_11851,N_10235,N_10283);
nor U11852 (N_11852,N_9497,N_9526);
nand U11853 (N_11853,N_10019,N_10283);
nor U11854 (N_11854,N_10336,N_10288);
xor U11855 (N_11855,N_9077,N_9478);
nor U11856 (N_11856,N_9662,N_9694);
nand U11857 (N_11857,N_9489,N_10041);
nand U11858 (N_11858,N_10305,N_9577);
nand U11859 (N_11859,N_10125,N_9887);
nor U11860 (N_11860,N_9730,N_9580);
and U11861 (N_11861,N_9296,N_10114);
and U11862 (N_11862,N_10144,N_10446);
and U11863 (N_11863,N_9714,N_10273);
xnor U11864 (N_11864,N_9064,N_9509);
nand U11865 (N_11865,N_9424,N_9490);
nor U11866 (N_11866,N_9769,N_9935);
or U11867 (N_11867,N_9896,N_9261);
and U11868 (N_11868,N_9371,N_9441);
xor U11869 (N_11869,N_9297,N_10006);
or U11870 (N_11870,N_9496,N_9859);
nand U11871 (N_11871,N_9939,N_9124);
and U11872 (N_11872,N_9829,N_10065);
or U11873 (N_11873,N_9044,N_10172);
xnor U11874 (N_11874,N_9317,N_10174);
and U11875 (N_11875,N_9062,N_10161);
nor U11876 (N_11876,N_10201,N_10006);
and U11877 (N_11877,N_10002,N_9492);
nor U11878 (N_11878,N_9891,N_9397);
or U11879 (N_11879,N_9049,N_10112);
nand U11880 (N_11880,N_9522,N_9958);
or U11881 (N_11881,N_10174,N_10499);
and U11882 (N_11882,N_9841,N_9304);
or U11883 (N_11883,N_10481,N_9746);
xnor U11884 (N_11884,N_9863,N_9173);
nor U11885 (N_11885,N_9131,N_9336);
and U11886 (N_11886,N_9678,N_9521);
or U11887 (N_11887,N_10024,N_9305);
xnor U11888 (N_11888,N_9420,N_9807);
and U11889 (N_11889,N_9685,N_10412);
or U11890 (N_11890,N_9110,N_9202);
nor U11891 (N_11891,N_10297,N_10102);
nand U11892 (N_11892,N_10210,N_9163);
nand U11893 (N_11893,N_10216,N_10345);
and U11894 (N_11894,N_9555,N_9412);
and U11895 (N_11895,N_9537,N_9897);
nor U11896 (N_11896,N_9887,N_10214);
and U11897 (N_11897,N_9038,N_10305);
nor U11898 (N_11898,N_9056,N_10486);
nor U11899 (N_11899,N_10094,N_10383);
nor U11900 (N_11900,N_10195,N_10455);
and U11901 (N_11901,N_9893,N_9071);
nand U11902 (N_11902,N_9300,N_9536);
nor U11903 (N_11903,N_10456,N_10080);
xnor U11904 (N_11904,N_9428,N_9175);
nand U11905 (N_11905,N_10387,N_10007);
nor U11906 (N_11906,N_9185,N_9269);
nor U11907 (N_11907,N_9908,N_10073);
or U11908 (N_11908,N_9848,N_9633);
nor U11909 (N_11909,N_10092,N_10197);
nand U11910 (N_11910,N_9520,N_9618);
and U11911 (N_11911,N_9181,N_10492);
nand U11912 (N_11912,N_9029,N_9934);
nand U11913 (N_11913,N_9798,N_10135);
xor U11914 (N_11914,N_9521,N_9280);
nor U11915 (N_11915,N_10331,N_10305);
xnor U11916 (N_11916,N_9187,N_9831);
and U11917 (N_11917,N_9716,N_9847);
nor U11918 (N_11918,N_9831,N_10404);
nand U11919 (N_11919,N_9921,N_9952);
nor U11920 (N_11920,N_10337,N_9962);
nand U11921 (N_11921,N_9092,N_10047);
nand U11922 (N_11922,N_9337,N_9676);
nand U11923 (N_11923,N_9461,N_9061);
nand U11924 (N_11924,N_9292,N_9806);
or U11925 (N_11925,N_9736,N_9322);
and U11926 (N_11926,N_10089,N_9399);
nand U11927 (N_11927,N_9327,N_9111);
and U11928 (N_11928,N_9038,N_10475);
xnor U11929 (N_11929,N_9548,N_9641);
xor U11930 (N_11930,N_10279,N_9886);
nand U11931 (N_11931,N_9544,N_9252);
or U11932 (N_11932,N_9811,N_9790);
or U11933 (N_11933,N_9190,N_9828);
nor U11934 (N_11934,N_9650,N_10443);
nand U11935 (N_11935,N_10289,N_9480);
nand U11936 (N_11936,N_9539,N_9639);
nor U11937 (N_11937,N_10360,N_9278);
xnor U11938 (N_11938,N_10097,N_9570);
xor U11939 (N_11939,N_9146,N_9360);
and U11940 (N_11940,N_9865,N_9745);
nor U11941 (N_11941,N_10064,N_10112);
or U11942 (N_11942,N_10333,N_9687);
and U11943 (N_11943,N_9630,N_9865);
and U11944 (N_11944,N_10136,N_9996);
or U11945 (N_11945,N_9480,N_10409);
nand U11946 (N_11946,N_10199,N_10013);
xnor U11947 (N_11947,N_9876,N_9646);
and U11948 (N_11948,N_9434,N_10152);
or U11949 (N_11949,N_9697,N_9459);
xnor U11950 (N_11950,N_10215,N_10139);
and U11951 (N_11951,N_9162,N_9482);
or U11952 (N_11952,N_9176,N_9096);
nor U11953 (N_11953,N_9458,N_9257);
and U11954 (N_11954,N_9324,N_9202);
or U11955 (N_11955,N_9551,N_9726);
nor U11956 (N_11956,N_9800,N_9426);
or U11957 (N_11957,N_9479,N_10188);
and U11958 (N_11958,N_10274,N_9102);
xor U11959 (N_11959,N_9442,N_9505);
or U11960 (N_11960,N_9895,N_10071);
nand U11961 (N_11961,N_9069,N_10039);
and U11962 (N_11962,N_9342,N_9129);
or U11963 (N_11963,N_9380,N_9868);
xor U11964 (N_11964,N_9125,N_10255);
or U11965 (N_11965,N_9622,N_10112);
nand U11966 (N_11966,N_9406,N_10126);
and U11967 (N_11967,N_9955,N_9792);
and U11968 (N_11968,N_9627,N_9199);
or U11969 (N_11969,N_9469,N_9742);
and U11970 (N_11970,N_9191,N_9478);
nand U11971 (N_11971,N_9127,N_9695);
nand U11972 (N_11972,N_9423,N_9341);
xnor U11973 (N_11973,N_9523,N_10113);
nand U11974 (N_11974,N_10186,N_9740);
xor U11975 (N_11975,N_10482,N_9291);
or U11976 (N_11976,N_10011,N_10472);
xor U11977 (N_11977,N_9685,N_9151);
xnor U11978 (N_11978,N_9111,N_9196);
nand U11979 (N_11979,N_9486,N_9416);
xor U11980 (N_11980,N_9051,N_9225);
nand U11981 (N_11981,N_9446,N_10272);
nor U11982 (N_11982,N_9159,N_9475);
and U11983 (N_11983,N_9598,N_10162);
nand U11984 (N_11984,N_9009,N_9173);
and U11985 (N_11985,N_9431,N_9595);
and U11986 (N_11986,N_9554,N_9313);
or U11987 (N_11987,N_9639,N_9940);
nor U11988 (N_11988,N_10489,N_9920);
and U11989 (N_11989,N_10416,N_9706);
or U11990 (N_11990,N_10306,N_9079);
xnor U11991 (N_11991,N_9295,N_9549);
and U11992 (N_11992,N_10097,N_9136);
nand U11993 (N_11993,N_9217,N_9159);
xnor U11994 (N_11994,N_9401,N_9025);
nor U11995 (N_11995,N_9085,N_9627);
or U11996 (N_11996,N_9801,N_9155);
nor U11997 (N_11997,N_9103,N_9330);
nor U11998 (N_11998,N_10443,N_9216);
xor U11999 (N_11999,N_10347,N_10093);
nor U12000 (N_12000,N_11870,N_11650);
nor U12001 (N_12001,N_11043,N_11471);
nand U12002 (N_12002,N_11366,N_10878);
xor U12003 (N_12003,N_11249,N_11268);
nand U12004 (N_12004,N_10981,N_10687);
and U12005 (N_12005,N_11240,N_11474);
nand U12006 (N_12006,N_11913,N_11824);
nor U12007 (N_12007,N_11964,N_11382);
nor U12008 (N_12008,N_11620,N_11588);
nand U12009 (N_12009,N_10931,N_11244);
nand U12010 (N_12010,N_10753,N_11879);
and U12011 (N_12011,N_10983,N_11123);
xor U12012 (N_12012,N_11888,N_11355);
or U12013 (N_12013,N_10596,N_11832);
and U12014 (N_12014,N_10590,N_11267);
xnor U12015 (N_12015,N_10782,N_11018);
xnor U12016 (N_12016,N_10679,N_11279);
nand U12017 (N_12017,N_11393,N_11220);
nand U12018 (N_12018,N_10885,N_11531);
xor U12019 (N_12019,N_11633,N_10555);
xor U12020 (N_12020,N_10853,N_11954);
nand U12021 (N_12021,N_11016,N_11993);
xor U12022 (N_12022,N_11166,N_11768);
nor U12023 (N_12023,N_10593,N_11770);
nand U12024 (N_12024,N_11945,N_10938);
xnor U12025 (N_12025,N_11276,N_11014);
xnor U12026 (N_12026,N_10867,N_11872);
or U12027 (N_12027,N_11097,N_11373);
or U12028 (N_12028,N_10940,N_10559);
nor U12029 (N_12029,N_10714,N_10866);
nor U12030 (N_12030,N_10979,N_11419);
nand U12031 (N_12031,N_11789,N_11417);
nand U12032 (N_12032,N_11710,N_11414);
or U12033 (N_12033,N_11013,N_11804);
and U12034 (N_12034,N_11970,N_11568);
or U12035 (N_12035,N_11010,N_11165);
and U12036 (N_12036,N_10550,N_11085);
nand U12037 (N_12037,N_10810,N_10846);
nor U12038 (N_12038,N_10901,N_11863);
nand U12039 (N_12039,N_11904,N_11918);
nand U12040 (N_12040,N_11066,N_10951);
or U12041 (N_12041,N_11444,N_10727);
or U12042 (N_12042,N_11708,N_11684);
nor U12043 (N_12043,N_11337,N_10992);
and U12044 (N_12044,N_11101,N_11562);
nor U12045 (N_12045,N_10614,N_11113);
and U12046 (N_12046,N_10883,N_10584);
xnor U12047 (N_12047,N_11692,N_10793);
xor U12048 (N_12048,N_11928,N_11490);
and U12049 (N_12049,N_11180,N_11374);
nand U12050 (N_12050,N_11302,N_10795);
xor U12051 (N_12051,N_11813,N_11963);
xnor U12052 (N_12052,N_11527,N_11231);
or U12053 (N_12053,N_11916,N_11186);
nor U12054 (N_12054,N_11111,N_11732);
nor U12055 (N_12055,N_11184,N_11545);
nand U12056 (N_12056,N_10710,N_10513);
nor U12057 (N_12057,N_11228,N_10798);
or U12058 (N_12058,N_11570,N_11183);
nor U12059 (N_12059,N_11925,N_10953);
xnor U12060 (N_12060,N_11936,N_11537);
nand U12061 (N_12061,N_11323,N_10703);
xor U12062 (N_12062,N_11286,N_11901);
or U12063 (N_12063,N_11195,N_11460);
nor U12064 (N_12064,N_11528,N_10778);
nand U12065 (N_12065,N_11896,N_11478);
and U12066 (N_12066,N_10632,N_10926);
nand U12067 (N_12067,N_10959,N_10945);
and U12068 (N_12068,N_11283,N_11274);
nor U12069 (N_12069,N_11818,N_11724);
and U12070 (N_12070,N_11681,N_11668);
or U12071 (N_12071,N_11775,N_11644);
nand U12072 (N_12072,N_11536,N_10543);
nor U12073 (N_12073,N_11859,N_11674);
and U12074 (N_12074,N_10569,N_10923);
xor U12075 (N_12075,N_11887,N_11764);
nand U12076 (N_12076,N_10964,N_11773);
or U12077 (N_12077,N_10807,N_11981);
and U12078 (N_12078,N_10948,N_11222);
nand U12079 (N_12079,N_11593,N_11217);
xnor U12080 (N_12080,N_10823,N_10527);
and U12081 (N_12081,N_11574,N_10505);
and U12082 (N_12082,N_11951,N_11608);
nand U12083 (N_12083,N_10877,N_10654);
nand U12084 (N_12084,N_11680,N_11080);
and U12085 (N_12085,N_11455,N_11696);
or U12086 (N_12086,N_11045,N_11172);
nand U12087 (N_12087,N_11740,N_11157);
nor U12088 (N_12088,N_11598,N_11573);
or U12089 (N_12089,N_10644,N_11483);
and U12090 (N_12090,N_11495,N_10652);
nor U12091 (N_12091,N_10561,N_11299);
xor U12092 (N_12092,N_11623,N_10939);
and U12093 (N_12093,N_11575,N_11445);
nor U12094 (N_12094,N_11966,N_11513);
or U12095 (N_12095,N_11838,N_11930);
xor U12096 (N_12096,N_11814,N_11019);
or U12097 (N_12097,N_11731,N_11008);
nor U12098 (N_12098,N_11007,N_11200);
and U12099 (N_12099,N_11163,N_11194);
xnor U12100 (N_12100,N_11224,N_11233);
xor U12101 (N_12101,N_11336,N_10726);
xor U12102 (N_12102,N_10743,N_10766);
and U12103 (N_12103,N_11505,N_11516);
nand U12104 (N_12104,N_11778,N_10733);
nand U12105 (N_12105,N_10967,N_11169);
xor U12106 (N_12106,N_11895,N_11409);
nand U12107 (N_12107,N_10749,N_10787);
and U12108 (N_12108,N_11144,N_10740);
or U12109 (N_12109,N_11726,N_11304);
nor U12110 (N_12110,N_10755,N_10560);
nand U12111 (N_12111,N_11785,N_11462);
or U12112 (N_12112,N_11796,N_10512);
and U12113 (N_12113,N_10845,N_10500);
or U12114 (N_12114,N_11050,N_11329);
or U12115 (N_12115,N_10974,N_11990);
nor U12116 (N_12116,N_11703,N_10977);
xnor U12117 (N_12117,N_10768,N_10902);
nor U12118 (N_12118,N_11852,N_11754);
nor U12119 (N_12119,N_11864,N_10635);
nor U12120 (N_12120,N_10792,N_11994);
and U12121 (N_12121,N_10683,N_10913);
nor U12122 (N_12122,N_10628,N_11324);
nor U12123 (N_12123,N_10690,N_11952);
nand U12124 (N_12124,N_11004,N_10738);
nand U12125 (N_12125,N_11563,N_11525);
xor U12126 (N_12126,N_11844,N_10579);
xor U12127 (N_12127,N_11027,N_11346);
nor U12128 (N_12128,N_11907,N_10697);
or U12129 (N_12129,N_10562,N_10578);
xnor U12130 (N_12130,N_11430,N_11421);
and U12131 (N_12131,N_11160,N_11858);
and U12132 (N_12132,N_11903,N_11151);
or U12133 (N_12133,N_10581,N_11629);
nand U12134 (N_12134,N_11874,N_10589);
xor U12135 (N_12135,N_11368,N_10709);
nor U12136 (N_12136,N_11214,N_11091);
or U12137 (N_12137,N_11108,N_11883);
nand U12138 (N_12138,N_11170,N_10580);
nor U12139 (N_12139,N_11543,N_11320);
nor U12140 (N_12140,N_11877,N_11557);
or U12141 (N_12141,N_10761,N_11362);
nand U12142 (N_12142,N_11853,N_11225);
xor U12143 (N_12143,N_11875,N_11847);
and U12144 (N_12144,N_11028,N_11552);
nor U12145 (N_12145,N_11198,N_11248);
nor U12146 (N_12146,N_10636,N_11783);
nand U12147 (N_12147,N_11950,N_10919);
nand U12148 (N_12148,N_11640,N_11694);
nor U12149 (N_12149,N_11216,N_10676);
nand U12150 (N_12150,N_11797,N_11148);
and U12151 (N_12151,N_11638,N_10600);
xnor U12152 (N_12152,N_11415,N_10594);
or U12153 (N_12153,N_10634,N_11475);
xnor U12154 (N_12154,N_10972,N_11912);
nor U12155 (N_12155,N_11071,N_11618);
and U12156 (N_12156,N_10587,N_10924);
nand U12157 (N_12157,N_10642,N_11012);
xnor U12158 (N_12158,N_11520,N_10980);
nor U12159 (N_12159,N_11985,N_11688);
xnor U12160 (N_12160,N_11539,N_10597);
nand U12161 (N_12161,N_11564,N_11816);
xor U12162 (N_12162,N_11940,N_11514);
nor U12163 (N_12163,N_11300,N_11499);
or U12164 (N_12164,N_11529,N_11866);
and U12165 (N_12165,N_11882,N_11017);
nor U12166 (N_12166,N_10801,N_11295);
and U12167 (N_12167,N_10789,N_11745);
nand U12168 (N_12168,N_11992,N_11182);
nor U12169 (N_12169,N_11141,N_11817);
xor U12170 (N_12170,N_11153,N_11069);
nor U12171 (N_12171,N_10520,N_11094);
nor U12172 (N_12172,N_10701,N_11728);
or U12173 (N_12173,N_11188,N_11743);
nor U12174 (N_12174,N_10618,N_11048);
nand U12175 (N_12175,N_11058,N_11278);
and U12176 (N_12176,N_11805,N_10888);
xor U12177 (N_12177,N_11892,N_11118);
nor U12178 (N_12178,N_10833,N_11693);
nand U12179 (N_12179,N_10721,N_10706);
xnor U12180 (N_12180,N_11512,N_11943);
nor U12181 (N_12181,N_11931,N_11597);
nand U12182 (N_12182,N_10835,N_11342);
nand U12183 (N_12183,N_11860,N_10582);
xor U12184 (N_12184,N_11034,N_11837);
nor U12185 (N_12185,N_10704,N_10884);
nand U12186 (N_12186,N_11841,N_10524);
xnor U12187 (N_12187,N_10758,N_11929);
nand U12188 (N_12188,N_11917,N_10640);
or U12189 (N_12189,N_11470,N_11894);
nor U12190 (N_12190,N_11707,N_11594);
nand U12191 (N_12191,N_11481,N_11026);
nor U12192 (N_12192,N_10966,N_11130);
xnor U12193 (N_12193,N_10803,N_10925);
nor U12194 (N_12194,N_11193,N_11654);
nand U12195 (N_12195,N_10626,N_11482);
nor U12196 (N_12196,N_10754,N_11155);
nor U12197 (N_12197,N_11236,N_11635);
or U12198 (N_12198,N_11944,N_11103);
or U12199 (N_12199,N_11345,N_11310);
and U12200 (N_12200,N_11765,N_10765);
or U12201 (N_12201,N_11766,N_11744);
nor U12202 (N_12202,N_11908,N_10598);
or U12203 (N_12203,N_11721,N_11697);
and U12204 (N_12204,N_10851,N_10759);
or U12205 (N_12205,N_11582,N_11352);
and U12206 (N_12206,N_11507,N_11054);
and U12207 (N_12207,N_11698,N_10741);
and U12208 (N_12208,N_11297,N_11578);
and U12209 (N_12209,N_10824,N_11689);
xnor U12210 (N_12210,N_11639,N_11973);
or U12211 (N_12211,N_11534,N_10645);
or U12212 (N_12212,N_11843,N_11029);
nand U12213 (N_12213,N_11658,N_11659);
and U12214 (N_12214,N_11965,N_11987);
or U12215 (N_12215,N_11363,N_11828);
xnor U12216 (N_12216,N_10944,N_11404);
and U12217 (N_12217,N_10954,N_11653);
nor U12218 (N_12218,N_11571,N_11255);
nand U12219 (N_12219,N_10804,N_11104);
and U12220 (N_12220,N_11530,N_10523);
nor U12221 (N_12221,N_11344,N_10941);
nand U12222 (N_12222,N_10568,N_11424);
and U12223 (N_12223,N_11391,N_10860);
nor U12224 (N_12224,N_11603,N_11319);
xnor U12225 (N_12225,N_11042,N_11434);
nor U12226 (N_12226,N_11713,N_11939);
or U12227 (N_12227,N_11230,N_10763);
nor U12228 (N_12228,N_11815,N_10933);
nand U12229 (N_12229,N_10889,N_11712);
or U12230 (N_12230,N_11187,N_11282);
and U12231 (N_12231,N_11755,N_10760);
nand U12232 (N_12232,N_11289,N_11932);
and U12233 (N_12233,N_11347,N_11110);
xor U12234 (N_12234,N_10750,N_11736);
nor U12235 (N_12235,N_11955,N_11269);
xor U12236 (N_12236,N_10825,N_11669);
or U12237 (N_12237,N_10519,N_11072);
nor U12238 (N_12238,N_11695,N_11384);
and U12239 (N_12239,N_11836,N_11999);
or U12240 (N_12240,N_11567,N_11447);
xor U12241 (N_12241,N_11227,N_11308);
and U12242 (N_12242,N_11760,N_10570);
nand U12243 (N_12243,N_11957,N_10665);
xor U12244 (N_12244,N_10928,N_11395);
nand U12245 (N_12245,N_10712,N_11122);
nand U12246 (N_12246,N_11910,N_11839);
and U12247 (N_12247,N_10842,N_11208);
nor U12248 (N_12248,N_11077,N_10747);
nor U12249 (N_12249,N_11159,N_11211);
nor U12250 (N_12250,N_11825,N_11834);
nand U12251 (N_12251,N_11995,N_11833);
xor U12252 (N_12252,N_11702,N_11114);
xnor U12253 (N_12253,N_11651,N_10657);
and U12254 (N_12254,N_11284,N_10854);
nand U12255 (N_12255,N_11009,N_10605);
or U12256 (N_12256,N_10912,N_10836);
or U12257 (N_12257,N_11400,N_11306);
nor U12258 (N_12258,N_11387,N_11138);
nand U12259 (N_12259,N_11020,N_11035);
or U12260 (N_12260,N_11742,N_11241);
nor U12261 (N_12261,N_11243,N_11664);
or U12262 (N_12262,N_11519,N_10748);
or U12263 (N_12263,N_11041,N_10893);
and U12264 (N_12264,N_11254,N_11919);
xor U12265 (N_12265,N_11780,N_10610);
xnor U12266 (N_12266,N_11672,N_10988);
xor U12267 (N_12267,N_11162,N_11673);
nand U12268 (N_12268,N_11037,N_11370);
and U12269 (N_12269,N_11354,N_10908);
and U12270 (N_12270,N_10502,N_11142);
or U12271 (N_12271,N_11022,N_10751);
xor U12272 (N_12272,N_11011,N_11496);
nor U12273 (N_12273,N_11585,N_11835);
or U12274 (N_12274,N_10847,N_11823);
xnor U12275 (N_12275,N_11532,N_10631);
or U12276 (N_12276,N_11427,N_11466);
nand U12277 (N_12277,N_11178,N_10918);
xor U12278 (N_12278,N_11518,N_10973);
nand U12279 (N_12279,N_10936,N_11105);
xor U12280 (N_12280,N_11686,N_10985);
or U12281 (N_12281,N_10622,N_11472);
or U12282 (N_12282,N_11806,N_11542);
and U12283 (N_12283,N_10869,N_11364);
and U12284 (N_12284,N_11605,N_11508);
nand U12285 (N_12285,N_11491,N_11622);
or U12286 (N_12286,N_10950,N_10564);
nand U12287 (N_12287,N_11587,N_11185);
and U12288 (N_12288,N_10872,N_11733);
or U12289 (N_12289,N_11260,N_11949);
xor U12290 (N_12290,N_11579,N_10909);
nor U12291 (N_12291,N_11328,N_11660);
xnor U12292 (N_12292,N_11106,N_11005);
nor U12293 (N_12293,N_10557,N_10968);
nand U12294 (N_12294,N_11088,N_11869);
or U12295 (N_12295,N_11506,N_11596);
or U12296 (N_12296,N_11868,N_11782);
xor U12297 (N_12297,N_10526,N_11318);
nand U12298 (N_12298,N_10999,N_11209);
nand U12299 (N_12299,N_11889,N_11422);
nor U12300 (N_12300,N_11880,N_11706);
xor U12301 (N_12301,N_11924,N_11270);
nand U12302 (N_12302,N_11645,N_11790);
xnor U12303 (N_12303,N_10781,N_10556);
and U12304 (N_12304,N_10831,N_11049);
or U12305 (N_12305,N_10688,N_11972);
nor U12306 (N_12306,N_11353,N_11365);
xnor U12307 (N_12307,N_11792,N_11060);
xnor U12308 (N_12308,N_11920,N_10935);
nor U12309 (N_12309,N_11357,N_11546);
nor U12310 (N_12310,N_11411,N_11959);
and U12311 (N_12311,N_11497,N_11607);
nand U12312 (N_12312,N_10623,N_11207);
nand U12313 (N_12313,N_11914,N_11139);
and U12314 (N_12314,N_10887,N_10814);
nand U12315 (N_12315,N_10828,N_11641);
and U12316 (N_12316,N_11649,N_11038);
nand U12317 (N_12317,N_11379,N_10509);
nand U12318 (N_12318,N_11070,N_11339);
nor U12319 (N_12319,N_11033,N_11601);
nand U12320 (N_12320,N_11126,N_11937);
or U12321 (N_12321,N_11277,N_10678);
nor U12322 (N_12322,N_10525,N_10599);
nand U12323 (N_12323,N_11290,N_11052);
nand U12324 (N_12324,N_11135,N_10879);
nand U12325 (N_12325,N_10708,N_11750);
xnor U12326 (N_12326,N_11886,N_11662);
or U12327 (N_12327,N_10773,N_11458);
nand U12328 (N_12328,N_11425,N_11465);
nand U12329 (N_12329,N_10800,N_11002);
nor U12330 (N_12330,N_11156,N_11192);
and U12331 (N_12331,N_10535,N_11509);
xor U12332 (N_12332,N_11372,N_10563);
or U12333 (N_12333,N_10890,N_11909);
nor U12334 (N_12334,N_11087,N_10834);
or U12335 (N_12335,N_10819,N_10895);
or U12336 (N_12336,N_11386,N_10677);
nand U12337 (N_12337,N_11210,N_11331);
xor U12338 (N_12338,N_11627,N_11281);
xnor U12339 (N_12339,N_11566,N_11565);
nand U12340 (N_12340,N_11309,N_11469);
and U12341 (N_12341,N_11068,N_11991);
nor U12342 (N_12342,N_11456,N_11642);
nand U12343 (N_12343,N_11367,N_11643);
nor U12344 (N_12344,N_11377,N_11493);
nand U12345 (N_12345,N_11793,N_11338);
nor U12346 (N_12346,N_11544,N_11583);
nand U12347 (N_12347,N_11501,N_11341);
or U12348 (N_12348,N_11962,N_10822);
nand U12349 (N_12349,N_10920,N_11855);
xor U12350 (N_12350,N_11271,N_11121);
and U12351 (N_12351,N_10583,N_10648);
or U12352 (N_12352,N_10521,N_11047);
xor U12353 (N_12353,N_10558,N_10670);
nand U12354 (N_12354,N_11794,N_10547);
or U12355 (N_12355,N_11389,N_11885);
or U12356 (N_12356,N_11390,N_11416);
nand U12357 (N_12357,N_11238,N_10855);
or U12358 (N_12358,N_10987,N_10522);
xor U12359 (N_12359,N_11967,N_10881);
nand U12360 (N_12360,N_11715,N_10608);
and U12361 (N_12361,N_11753,N_10989);
or U12362 (N_12362,N_10691,N_10573);
nor U12363 (N_12363,N_11436,N_11779);
nand U12364 (N_12364,N_11891,N_10903);
xnor U12365 (N_12365,N_11759,N_11001);
and U12366 (N_12366,N_10906,N_10894);
and U12367 (N_12367,N_10715,N_11751);
nand U12368 (N_12368,N_11448,N_11921);
xnor U12369 (N_12369,N_10711,N_11849);
and U12370 (N_12370,N_11055,N_11609);
xor U12371 (N_12371,N_11258,N_10651);
xnor U12372 (N_12372,N_10553,N_10791);
nand U12373 (N_12373,N_11203,N_10947);
nand U12374 (N_12374,N_11468,N_10790);
nand U12375 (N_12375,N_10529,N_11443);
nand U12376 (N_12376,N_11092,N_11763);
or U12377 (N_12377,N_11250,N_11535);
xnor U12378 (N_12378,N_10997,N_10886);
nor U12379 (N_12379,N_10699,N_11485);
and U12380 (N_12380,N_11840,N_11305);
nor U12381 (N_12381,N_11734,N_10776);
nor U12382 (N_12382,N_11560,N_11676);
or U12383 (N_12383,N_11061,N_11062);
and U12384 (N_12384,N_10943,N_11046);
nor U12385 (N_12385,N_11065,N_10737);
or U12386 (N_12386,N_11705,N_11812);
xnor U12387 (N_12387,N_10639,N_11915);
nand U12388 (N_12388,N_10732,N_11861);
xnor U12389 (N_12389,N_11667,N_11761);
and U12390 (N_12390,N_11854,N_11376);
and U12391 (N_12391,N_10829,N_10694);
nor U12392 (N_12392,N_10510,N_10840);
or U12393 (N_12393,N_11292,N_11719);
or U12394 (N_12394,N_11489,N_10856);
nand U12395 (N_12395,N_11934,N_11510);
nand U12396 (N_12396,N_11558,N_11086);
xnor U12397 (N_12397,N_11827,N_11850);
and U12398 (N_12398,N_11221,N_10850);
xor U12399 (N_12399,N_11191,N_10692);
nor U12400 (N_12400,N_11730,N_11577);
nand U12401 (N_12401,N_10857,N_11787);
or U12402 (N_12402,N_11399,N_11599);
nand U12403 (N_12403,N_11540,N_11624);
or U12404 (N_12404,N_10716,N_11361);
xnor U12405 (N_12405,N_11158,N_11846);
nand U12406 (N_12406,N_11677,N_10832);
or U12407 (N_12407,N_11067,N_11032);
and U12408 (N_12408,N_10899,N_10976);
xor U12409 (N_12409,N_11056,N_11413);
nand U12410 (N_12410,N_10577,N_10960);
or U12411 (N_12411,N_10629,N_10772);
and U12412 (N_12412,N_11079,N_11125);
nor U12413 (N_12413,N_11219,N_11500);
nor U12414 (N_12414,N_11251,N_11360);
nand U12415 (N_12415,N_10544,N_10813);
or U12416 (N_12416,N_11439,N_10916);
nor U12417 (N_12417,N_10859,N_11821);
or U12418 (N_12418,N_11589,N_11757);
xnor U12419 (N_12419,N_11205,N_11590);
and U12420 (N_12420,N_10917,N_10602);
and U12421 (N_12421,N_11451,N_11722);
or U12422 (N_12422,N_11926,N_10551);
nor U12423 (N_12423,N_11176,N_10796);
nor U12424 (N_12424,N_11871,N_10952);
and U12425 (N_12425,N_11625,N_11723);
xor U12426 (N_12426,N_11647,N_11147);
xnor U12427 (N_12427,N_11700,N_11729);
or U12428 (N_12428,N_11661,N_11524);
and U12429 (N_12429,N_11498,N_11177);
nand U12430 (N_12430,N_11408,N_10794);
xnor U12431 (N_12431,N_11388,N_10870);
nand U12432 (N_12432,N_10680,N_11115);
or U12433 (N_12433,N_11477,N_11829);
and U12434 (N_12434,N_10830,N_11906);
nand U12435 (N_12435,N_10686,N_11884);
and U12436 (N_12436,N_11977,N_10506);
or U12437 (N_12437,N_11898,N_11212);
or U12438 (N_12438,N_11714,N_11982);
nand U12439 (N_12439,N_11246,N_10817);
nor U12440 (N_12440,N_11044,N_11392);
and U12441 (N_12441,N_11800,N_11772);
nand U12442 (N_12442,N_11340,N_11741);
and U12443 (N_12443,N_11989,N_11922);
nor U12444 (N_12444,N_11533,N_11820);
and U12445 (N_12445,N_10864,N_10868);
or U12446 (N_12446,N_10638,N_11810);
nand U12447 (N_12447,N_11412,N_10821);
nor U12448 (N_12448,N_11264,N_11636);
xor U12449 (N_12449,N_10735,N_10720);
and U12450 (N_12450,N_11876,N_11396);
or U12451 (N_12451,N_10606,N_10546);
and U12452 (N_12452,N_11717,N_11407);
nand U12453 (N_12453,N_10533,N_10900);
nand U12454 (N_12454,N_11167,N_11383);
and U12455 (N_12455,N_11976,N_11801);
nand U12456 (N_12456,N_10730,N_11547);
nand U12457 (N_12457,N_11437,N_11819);
xor U12458 (N_12458,N_10669,N_11867);
or U12459 (N_12459,N_11090,N_10849);
nand U12460 (N_12460,N_11725,N_10507);
or U12461 (N_12461,N_10611,N_10719);
nor U12462 (N_12462,N_10752,N_11541);
xor U12463 (N_12463,N_11146,N_11381);
xnor U12464 (N_12464,N_10880,N_11202);
or U12465 (N_12465,N_11682,N_11515);
xnor U12466 (N_12466,N_11663,N_11933);
nor U12467 (N_12467,N_10892,N_11610);
or U12468 (N_12468,N_11315,N_10565);
nand U12469 (N_12469,N_11795,N_10998);
and U12470 (N_12470,N_11616,N_11762);
nand U12471 (N_12471,N_11776,N_11288);
nand U12472 (N_12472,N_11997,N_10724);
xnor U12473 (N_12473,N_10996,N_11401);
or U12474 (N_12474,N_11581,N_11040);
or U12475 (N_12475,N_10536,N_10962);
and U12476 (N_12476,N_10514,N_10707);
nor U12477 (N_12477,N_10612,N_11441);
and U12478 (N_12478,N_11348,N_11971);
or U12479 (N_12479,N_11665,N_10530);
and U12480 (N_12480,N_10588,N_11064);
nand U12481 (N_12481,N_10861,N_11078);
nor U12482 (N_12482,N_11612,N_10745);
nand U12483 (N_12483,N_11215,N_11199);
or U12484 (N_12484,N_11057,N_11911);
xnor U12485 (N_12485,N_10844,N_11201);
nand U12486 (N_12486,N_11133,N_11280);
and U12487 (N_12487,N_11272,N_11927);
and U12488 (N_12488,N_11611,N_10874);
and U12489 (N_12489,N_11486,N_11025);
and U12490 (N_12490,N_11727,N_10591);
nor U12491 (N_12491,N_11397,N_10656);
or U12492 (N_12492,N_10620,N_11856);
xor U12493 (N_12493,N_11015,N_11418);
nor U12494 (N_12494,N_11332,N_11735);
nor U12495 (N_12495,N_11747,N_10643);
nor U12496 (N_12496,N_11137,N_10875);
nand U12497 (N_12497,N_11375,N_11204);
and U12498 (N_12498,N_11628,N_11093);
and U12499 (N_12499,N_11648,N_10542);
and U12500 (N_12500,N_11670,N_11960);
or U12501 (N_12501,N_10876,N_10921);
nor U12502 (N_12502,N_11406,N_11613);
nand U12503 (N_12503,N_11197,N_10723);
or U12504 (N_12504,N_10698,N_11938);
nand U12505 (N_12505,N_11826,N_11956);
nor U12506 (N_12506,N_11398,N_10837);
and U12507 (N_12507,N_10615,N_11082);
nor U12508 (N_12508,N_10771,N_11737);
and U12509 (N_12509,N_10970,N_10673);
xnor U12510 (N_12510,N_10827,N_11983);
nand U12511 (N_12511,N_10971,N_10646);
nand U12512 (N_12512,N_11784,N_11857);
xor U12513 (N_12513,N_10958,N_10575);
nand U12514 (N_12514,N_11378,N_10641);
or U12515 (N_12515,N_10808,N_10508);
xnor U12516 (N_12516,N_10797,N_11143);
and U12517 (N_12517,N_11223,N_11652);
and U12518 (N_12518,N_11235,N_11556);
or U12519 (N_12519,N_11394,N_11189);
xor U12520 (N_12520,N_10649,N_10922);
and U12521 (N_12521,N_11678,N_11656);
or U12522 (N_12522,N_11709,N_11523);
nor U12523 (N_12523,N_10865,N_10934);
xor U12524 (N_12524,N_10725,N_11494);
or U12525 (N_12525,N_11675,N_10567);
nor U12526 (N_12526,N_10503,N_11808);
and U12527 (N_12527,N_10650,N_10769);
xnor U12528 (N_12528,N_11316,N_11322);
or U12529 (N_12529,N_11655,N_11830);
nand U12530 (N_12530,N_11953,N_11239);
and U12531 (N_12531,N_11798,N_11081);
nor U12532 (N_12532,N_11548,N_11873);
nand U12533 (N_12533,N_10982,N_11591);
or U12534 (N_12534,N_11559,N_11538);
nor U12535 (N_12535,N_11600,N_11426);
xnor U12536 (N_12536,N_11429,N_11181);
nand U12537 (N_12537,N_10898,N_11941);
and U12538 (N_12538,N_11473,N_10826);
xor U12539 (N_12539,N_11602,N_10991);
or U12540 (N_12540,N_10969,N_10666);
xor U12541 (N_12541,N_11380,N_11132);
xor U12542 (N_12542,N_11317,N_10780);
nand U12543 (N_12543,N_11371,N_10986);
or U12544 (N_12544,N_11423,N_10871);
or U12545 (N_12545,N_11107,N_11958);
or U12546 (N_12546,N_10839,N_11758);
xor U12547 (N_12547,N_11059,N_11102);
and U12548 (N_12548,N_10537,N_10734);
and U12549 (N_12549,N_10965,N_10538);
and U12550 (N_12550,N_10619,N_11333);
xnor U12551 (N_12551,N_11988,N_11774);
or U12552 (N_12552,N_11595,N_10504);
xnor U12553 (N_12553,N_11164,N_11173);
xnor U12554 (N_12554,N_10915,N_10929);
xor U12555 (N_12555,N_10805,N_10621);
nor U12556 (N_12556,N_10515,N_11576);
and U12557 (N_12557,N_11890,N_10684);
nand U12558 (N_12558,N_10722,N_11402);
nand U12559 (N_12559,N_11614,N_10862);
nand U12560 (N_12560,N_11767,N_11511);
or U12561 (N_12561,N_10742,N_11234);
nor U12562 (N_12562,N_10625,N_11428);
nor U12563 (N_12563,N_10774,N_10777);
nor U12564 (N_12564,N_11074,N_11311);
xnor U12565 (N_12565,N_11807,N_10882);
nor U12566 (N_12566,N_10984,N_10757);
and U12567 (N_12567,N_11334,N_11095);
or U12568 (N_12568,N_11484,N_11604);
nand U12569 (N_12569,N_10930,N_11136);
nor U12570 (N_12570,N_11076,N_11974);
nor U12571 (N_12571,N_10627,N_11247);
or U12572 (N_12572,N_11343,N_10511);
nand U12573 (N_12573,N_10910,N_11657);
and U12574 (N_12574,N_10539,N_10518);
or U12575 (N_12575,N_11947,N_11961);
or U12576 (N_12576,N_10674,N_11036);
nor U12577 (N_12577,N_10762,N_10820);
and U12578 (N_12578,N_10994,N_11196);
and U12579 (N_12579,N_11213,N_11021);
and U12580 (N_12580,N_11161,N_11263);
or U12581 (N_12581,N_11504,N_10545);
nor U12582 (N_12582,N_10609,N_10731);
nor U12583 (N_12583,N_11454,N_11720);
and U12584 (N_12584,N_11127,N_11449);
xnor U12585 (N_12585,N_11799,N_11948);
nand U12586 (N_12586,N_11549,N_11083);
xor U12587 (N_12587,N_10660,N_11120);
nand U12588 (N_12588,N_10667,N_10552);
nor U12589 (N_12589,N_10891,N_10516);
nand U12590 (N_12590,N_11502,N_10995);
or U12591 (N_12591,N_11555,N_11626);
and U12592 (N_12592,N_11786,N_11432);
nor U12593 (N_12593,N_11756,N_11503);
nor U12594 (N_12594,N_11803,N_10540);
xor U12595 (N_12595,N_10574,N_11487);
nand U12596 (N_12596,N_10576,N_10566);
xnor U12597 (N_12597,N_10658,N_11273);
or U12598 (N_12598,N_11586,N_11802);
nand U12599 (N_12599,N_11256,N_10955);
nor U12600 (N_12600,N_11124,N_11229);
nor U12601 (N_12601,N_10783,N_11986);
nor U12602 (N_12602,N_11980,N_11718);
xor U12603 (N_12603,N_10630,N_10961);
or U12604 (N_12604,N_11606,N_11356);
nor U12605 (N_12605,N_11327,N_11897);
xor U12606 (N_12606,N_11550,N_11298);
nor U12607 (N_12607,N_10756,N_11492);
and U12608 (N_12608,N_10956,N_10927);
xnor U12609 (N_12609,N_11084,N_11584);
nor U12610 (N_12610,N_11738,N_11580);
nand U12611 (N_12611,N_11100,N_11621);
or U12612 (N_12612,N_10764,N_10802);
and U12613 (N_12613,N_11438,N_10897);
and U12614 (N_12614,N_10843,N_10815);
and U12615 (N_12615,N_11096,N_11285);
nor U12616 (N_12616,N_10816,N_10607);
nand U12617 (N_12617,N_11517,N_11174);
or U12618 (N_12618,N_10501,N_11572);
nor U12619 (N_12619,N_11003,N_11592);
nor U12620 (N_12620,N_11253,N_11433);
xnor U12621 (N_12621,N_11112,N_11701);
nand U12622 (N_12622,N_10571,N_11350);
nor U12623 (N_12623,N_10770,N_11632);
nor U12624 (N_12624,N_11242,N_10528);
and U12625 (N_12625,N_11553,N_10914);
nor U12626 (N_12626,N_11526,N_10613);
and U12627 (N_12627,N_11457,N_10601);
nor U12628 (N_12628,N_11881,N_10695);
nand U12629 (N_12629,N_11788,N_10541);
nand U12630 (N_12630,N_10718,N_11551);
and U12631 (N_12631,N_11467,N_10841);
xor U12632 (N_12632,N_10905,N_10617);
nor U12633 (N_12633,N_11358,N_11522);
nand U12634 (N_12634,N_10784,N_10942);
xor U12635 (N_12635,N_11781,N_11446);
nand U12636 (N_12636,N_11615,N_11257);
and U12637 (N_12637,N_10647,N_10812);
nor U12638 (N_12638,N_10904,N_11206);
xor U12639 (N_12639,N_11359,N_11218);
and U12640 (N_12640,N_10767,N_10775);
or U12641 (N_12641,N_11063,N_11811);
nand U12642 (N_12642,N_10963,N_11129);
xor U12643 (N_12643,N_11294,N_11984);
and U12644 (N_12644,N_10729,N_11307);
nor U12645 (N_12645,N_10653,N_10549);
nor U12646 (N_12646,N_10744,N_10949);
nor U12647 (N_12647,N_10548,N_11942);
xor U12648 (N_12648,N_11175,N_10534);
nor U12649 (N_12649,N_11226,N_11459);
and U12650 (N_12650,N_10681,N_11746);
and U12651 (N_12651,N_11691,N_11561);
and U12652 (N_12652,N_11979,N_11154);
nor U12653 (N_12653,N_11969,N_10517);
and U12654 (N_12654,N_11039,N_11119);
xnor U12655 (N_12655,N_11666,N_11865);
nand U12656 (N_12656,N_11739,N_11330);
nor U12657 (N_12657,N_10993,N_10788);
nand U12658 (N_12658,N_10978,N_10717);
or U12659 (N_12659,N_11245,N_11935);
and U12660 (N_12660,N_10911,N_11410);
nor U12661 (N_12661,N_10672,N_11630);
nor U12662 (N_12662,N_11179,N_11646);
xor U12663 (N_12663,N_11099,N_11435);
nand U12664 (N_12664,N_11140,N_11312);
nand U12665 (N_12665,N_11685,N_10655);
xor U12666 (N_12666,N_10585,N_11420);
and U12667 (N_12667,N_11634,N_10531);
nor U12668 (N_12668,N_10809,N_11349);
xnor U12669 (N_12669,N_11569,N_11716);
and U12670 (N_12670,N_11899,N_11385);
nor U12671 (N_12671,N_10671,N_11314);
xor U12672 (N_12672,N_11452,N_11403);
and U12673 (N_12673,N_10572,N_11946);
xnor U12674 (N_12674,N_11023,N_10661);
and U12675 (N_12675,N_10785,N_11024);
nor U12676 (N_12676,N_11521,N_11480);
or U12677 (N_12677,N_11905,N_11150);
or U12678 (N_12678,N_10637,N_11266);
nor U12679 (N_12679,N_11291,N_11321);
nor U12680 (N_12680,N_11152,N_10592);
nor U12681 (N_12681,N_11301,N_11862);
or U12682 (N_12682,N_11752,N_11326);
nand U12683 (N_12683,N_11335,N_10586);
or U12684 (N_12684,N_10682,N_11978);
and U12685 (N_12685,N_11996,N_11171);
nor U12686 (N_12686,N_11450,N_10685);
xor U12687 (N_12687,N_11109,N_11748);
nand U12688 (N_12688,N_11631,N_10702);
or U12689 (N_12689,N_10736,N_10624);
and U12690 (N_12690,N_10603,N_11232);
nor U12691 (N_12691,N_10932,N_10946);
nand U12692 (N_12692,N_10700,N_11476);
xor U12693 (N_12693,N_10696,N_10693);
or U12694 (N_12694,N_11237,N_11442);
and U12695 (N_12695,N_10957,N_10728);
or U12696 (N_12696,N_11116,N_11619);
nand U12697 (N_12697,N_11453,N_11554);
xor U12698 (N_12698,N_11488,N_10907);
nor U12699 (N_12699,N_10633,N_11968);
and U12700 (N_12700,N_10858,N_10689);
and U12701 (N_12701,N_10604,N_11145);
or U12702 (N_12702,N_11848,N_11704);
or U12703 (N_12703,N_11325,N_10848);
or U12704 (N_12704,N_10739,N_11369);
or U12705 (N_12705,N_11893,N_11671);
or U12706 (N_12706,N_11464,N_11431);
and U12707 (N_12707,N_10664,N_10818);
and U12708 (N_12708,N_11053,N_11679);
nor U12709 (N_12709,N_10713,N_10896);
xnor U12710 (N_12710,N_10705,N_11822);
xnor U12711 (N_12711,N_11075,N_10873);
and U12712 (N_12712,N_11259,N_11031);
or U12713 (N_12713,N_11351,N_11711);
nand U12714 (N_12714,N_11073,N_10838);
nor U12715 (N_12715,N_11637,N_11117);
nor U12716 (N_12716,N_11051,N_10663);
xnor U12717 (N_12717,N_11303,N_10554);
and U12718 (N_12718,N_11791,N_11902);
and U12719 (N_12719,N_11975,N_10975);
and U12720 (N_12720,N_11261,N_11769);
nand U12721 (N_12721,N_11265,N_11190);
nand U12722 (N_12722,N_11006,N_10786);
or U12723 (N_12723,N_11134,N_11777);
or U12724 (N_12724,N_11089,N_11131);
and U12725 (N_12725,N_10811,N_11479);
and U12726 (N_12726,N_11000,N_11878);
nor U12727 (N_12727,N_11461,N_10659);
nor U12728 (N_12728,N_11923,N_10595);
xnor U12729 (N_12729,N_11699,N_11851);
or U12730 (N_12730,N_10675,N_10990);
xnor U12731 (N_12731,N_10863,N_11683);
nand U12732 (N_12732,N_11313,N_11831);
xor U12733 (N_12733,N_10937,N_11440);
or U12734 (N_12734,N_10799,N_10746);
nand U12735 (N_12735,N_11098,N_10852);
xnor U12736 (N_12736,N_11842,N_11749);
or U12737 (N_12737,N_10806,N_11771);
nand U12738 (N_12738,N_11275,N_11900);
nor U12739 (N_12739,N_11617,N_11168);
nand U12740 (N_12740,N_11809,N_10662);
nor U12741 (N_12741,N_11690,N_11998);
nand U12742 (N_12742,N_11030,N_11128);
nand U12743 (N_12743,N_11262,N_11287);
and U12744 (N_12744,N_10616,N_11845);
nor U12745 (N_12745,N_10779,N_11463);
xor U12746 (N_12746,N_11687,N_11405);
xnor U12747 (N_12747,N_10668,N_11296);
nor U12748 (N_12748,N_11293,N_11252);
and U12749 (N_12749,N_10532,N_11149);
nand U12750 (N_12750,N_11208,N_11565);
nor U12751 (N_12751,N_11633,N_10665);
or U12752 (N_12752,N_10864,N_11449);
xor U12753 (N_12753,N_11131,N_11368);
xor U12754 (N_12754,N_11420,N_10785);
nor U12755 (N_12755,N_10925,N_11423);
xnor U12756 (N_12756,N_10589,N_11713);
and U12757 (N_12757,N_11377,N_11869);
and U12758 (N_12758,N_10753,N_10791);
nand U12759 (N_12759,N_11560,N_11069);
nor U12760 (N_12760,N_11412,N_11874);
xnor U12761 (N_12761,N_10917,N_11999);
nor U12762 (N_12762,N_11018,N_11993);
or U12763 (N_12763,N_11209,N_11812);
or U12764 (N_12764,N_11377,N_11708);
xnor U12765 (N_12765,N_11882,N_11018);
xnor U12766 (N_12766,N_10956,N_11276);
and U12767 (N_12767,N_11498,N_11973);
and U12768 (N_12768,N_10837,N_11223);
xnor U12769 (N_12769,N_11574,N_11789);
xor U12770 (N_12770,N_11927,N_11723);
nand U12771 (N_12771,N_10624,N_10677);
and U12772 (N_12772,N_11320,N_11214);
xnor U12773 (N_12773,N_11772,N_11028);
nand U12774 (N_12774,N_11124,N_11435);
nand U12775 (N_12775,N_11474,N_11590);
nor U12776 (N_12776,N_11642,N_11421);
xnor U12777 (N_12777,N_11518,N_11945);
xnor U12778 (N_12778,N_11109,N_11638);
nor U12779 (N_12779,N_10619,N_11198);
nor U12780 (N_12780,N_11279,N_11826);
and U12781 (N_12781,N_11482,N_11997);
nand U12782 (N_12782,N_11677,N_11264);
xnor U12783 (N_12783,N_11966,N_11899);
xor U12784 (N_12784,N_11583,N_11337);
nor U12785 (N_12785,N_11385,N_11013);
nand U12786 (N_12786,N_11205,N_11555);
xnor U12787 (N_12787,N_10781,N_11221);
nor U12788 (N_12788,N_11785,N_10570);
or U12789 (N_12789,N_10718,N_11508);
xor U12790 (N_12790,N_11665,N_11844);
nand U12791 (N_12791,N_10625,N_10933);
nand U12792 (N_12792,N_11487,N_10733);
nor U12793 (N_12793,N_11786,N_10794);
xor U12794 (N_12794,N_10853,N_11843);
and U12795 (N_12795,N_11237,N_11885);
nor U12796 (N_12796,N_11040,N_10569);
xor U12797 (N_12797,N_10940,N_10589);
or U12798 (N_12798,N_10538,N_11876);
and U12799 (N_12799,N_10997,N_11796);
nor U12800 (N_12800,N_10755,N_11046);
and U12801 (N_12801,N_11778,N_11541);
and U12802 (N_12802,N_11171,N_11840);
nor U12803 (N_12803,N_11440,N_10530);
and U12804 (N_12804,N_11098,N_11538);
nor U12805 (N_12805,N_11425,N_11548);
xor U12806 (N_12806,N_11264,N_10902);
or U12807 (N_12807,N_10887,N_11765);
xor U12808 (N_12808,N_11446,N_11350);
or U12809 (N_12809,N_11674,N_11178);
or U12810 (N_12810,N_11805,N_11071);
nor U12811 (N_12811,N_10770,N_11982);
or U12812 (N_12812,N_10722,N_11775);
nand U12813 (N_12813,N_11448,N_11882);
xnor U12814 (N_12814,N_10670,N_11909);
or U12815 (N_12815,N_10515,N_11065);
xnor U12816 (N_12816,N_10886,N_10558);
xor U12817 (N_12817,N_10797,N_11480);
nor U12818 (N_12818,N_11616,N_11134);
nand U12819 (N_12819,N_11879,N_10592);
xnor U12820 (N_12820,N_11297,N_11372);
or U12821 (N_12821,N_11896,N_11659);
nand U12822 (N_12822,N_10507,N_10662);
nand U12823 (N_12823,N_11656,N_11418);
nor U12824 (N_12824,N_11259,N_11660);
xnor U12825 (N_12825,N_10828,N_11562);
xnor U12826 (N_12826,N_10601,N_11276);
and U12827 (N_12827,N_10573,N_11100);
and U12828 (N_12828,N_11297,N_11474);
and U12829 (N_12829,N_11622,N_11748);
and U12830 (N_12830,N_11975,N_11398);
or U12831 (N_12831,N_11372,N_11388);
xor U12832 (N_12832,N_11572,N_10878);
xor U12833 (N_12833,N_11280,N_11283);
nand U12834 (N_12834,N_11376,N_10958);
or U12835 (N_12835,N_10503,N_10761);
and U12836 (N_12836,N_11025,N_11059);
or U12837 (N_12837,N_10508,N_11403);
and U12838 (N_12838,N_11172,N_11487);
and U12839 (N_12839,N_11767,N_11940);
or U12840 (N_12840,N_11338,N_11629);
or U12841 (N_12841,N_10652,N_10894);
and U12842 (N_12842,N_11190,N_11938);
and U12843 (N_12843,N_10682,N_10510);
nand U12844 (N_12844,N_11715,N_10716);
or U12845 (N_12845,N_10526,N_10595);
and U12846 (N_12846,N_11879,N_10691);
xnor U12847 (N_12847,N_11118,N_11094);
or U12848 (N_12848,N_11470,N_11316);
or U12849 (N_12849,N_10638,N_11052);
or U12850 (N_12850,N_11138,N_11279);
xor U12851 (N_12851,N_11422,N_11642);
nor U12852 (N_12852,N_10620,N_11637);
xnor U12853 (N_12853,N_11673,N_11799);
and U12854 (N_12854,N_11330,N_11911);
nand U12855 (N_12855,N_11313,N_10611);
or U12856 (N_12856,N_11793,N_11797);
nor U12857 (N_12857,N_11322,N_11400);
and U12858 (N_12858,N_10974,N_11951);
nor U12859 (N_12859,N_11152,N_10758);
nor U12860 (N_12860,N_10846,N_10976);
or U12861 (N_12861,N_11964,N_11024);
xor U12862 (N_12862,N_10878,N_10963);
nand U12863 (N_12863,N_11055,N_11117);
nand U12864 (N_12864,N_11882,N_11419);
or U12865 (N_12865,N_11278,N_11155);
or U12866 (N_12866,N_11415,N_11601);
xnor U12867 (N_12867,N_11869,N_10840);
nand U12868 (N_12868,N_11055,N_11113);
and U12869 (N_12869,N_11640,N_11393);
nor U12870 (N_12870,N_10971,N_11844);
and U12871 (N_12871,N_11419,N_11218);
or U12872 (N_12872,N_11568,N_11692);
or U12873 (N_12873,N_11712,N_11878);
nand U12874 (N_12874,N_10968,N_11297);
nand U12875 (N_12875,N_11524,N_11571);
nor U12876 (N_12876,N_11379,N_11419);
or U12877 (N_12877,N_10536,N_10615);
nand U12878 (N_12878,N_11427,N_11342);
nand U12879 (N_12879,N_10935,N_11505);
nor U12880 (N_12880,N_11802,N_11309);
nor U12881 (N_12881,N_10643,N_11229);
or U12882 (N_12882,N_11298,N_10849);
or U12883 (N_12883,N_11884,N_11085);
xnor U12884 (N_12884,N_11565,N_11698);
nor U12885 (N_12885,N_11712,N_11760);
xnor U12886 (N_12886,N_10920,N_11623);
xor U12887 (N_12887,N_11697,N_11762);
nor U12888 (N_12888,N_10809,N_11751);
or U12889 (N_12889,N_10992,N_11525);
nor U12890 (N_12890,N_11268,N_10501);
or U12891 (N_12891,N_11911,N_11152);
or U12892 (N_12892,N_10623,N_11172);
or U12893 (N_12893,N_11661,N_11294);
and U12894 (N_12894,N_10794,N_10767);
nor U12895 (N_12895,N_11238,N_11957);
or U12896 (N_12896,N_11673,N_11400);
nor U12897 (N_12897,N_11508,N_11513);
nor U12898 (N_12898,N_10545,N_11564);
xor U12899 (N_12899,N_10678,N_11241);
xnor U12900 (N_12900,N_11919,N_11389);
and U12901 (N_12901,N_11721,N_11318);
xnor U12902 (N_12902,N_10678,N_10861);
xor U12903 (N_12903,N_10710,N_11360);
xor U12904 (N_12904,N_11145,N_10599);
xor U12905 (N_12905,N_10500,N_10706);
nand U12906 (N_12906,N_11796,N_11532);
nor U12907 (N_12907,N_11403,N_11596);
nand U12908 (N_12908,N_11389,N_11767);
nand U12909 (N_12909,N_11164,N_11532);
xor U12910 (N_12910,N_11006,N_11609);
and U12911 (N_12911,N_11723,N_11066);
nand U12912 (N_12912,N_11368,N_10967);
xnor U12913 (N_12913,N_11184,N_10525);
nand U12914 (N_12914,N_11118,N_11730);
or U12915 (N_12915,N_11621,N_11873);
xor U12916 (N_12916,N_10667,N_11615);
nor U12917 (N_12917,N_11283,N_10654);
xnor U12918 (N_12918,N_11957,N_11580);
and U12919 (N_12919,N_11234,N_10647);
nand U12920 (N_12920,N_10810,N_11245);
nor U12921 (N_12921,N_11626,N_10742);
xor U12922 (N_12922,N_11583,N_11013);
or U12923 (N_12923,N_11433,N_11162);
xor U12924 (N_12924,N_11875,N_11127);
nand U12925 (N_12925,N_11808,N_11270);
or U12926 (N_12926,N_10831,N_11457);
nor U12927 (N_12927,N_11792,N_11982);
nor U12928 (N_12928,N_11212,N_11859);
nor U12929 (N_12929,N_11677,N_11601);
nand U12930 (N_12930,N_10797,N_11660);
and U12931 (N_12931,N_10648,N_11545);
nand U12932 (N_12932,N_10785,N_11010);
and U12933 (N_12933,N_11277,N_11486);
nand U12934 (N_12934,N_11730,N_11262);
xnor U12935 (N_12935,N_11194,N_11252);
nand U12936 (N_12936,N_11656,N_10851);
or U12937 (N_12937,N_10719,N_10783);
or U12938 (N_12938,N_11461,N_11349);
or U12939 (N_12939,N_11827,N_10968);
nand U12940 (N_12940,N_10709,N_11582);
nand U12941 (N_12941,N_10651,N_11142);
and U12942 (N_12942,N_11699,N_11089);
xnor U12943 (N_12943,N_10726,N_11867);
xnor U12944 (N_12944,N_11679,N_11615);
nor U12945 (N_12945,N_11382,N_10931);
and U12946 (N_12946,N_11882,N_11441);
and U12947 (N_12947,N_10642,N_11379);
xnor U12948 (N_12948,N_11821,N_10787);
xor U12949 (N_12949,N_11600,N_11718);
or U12950 (N_12950,N_11679,N_10981);
or U12951 (N_12951,N_10836,N_11179);
and U12952 (N_12952,N_11530,N_11125);
or U12953 (N_12953,N_11425,N_10873);
nand U12954 (N_12954,N_11236,N_11891);
nor U12955 (N_12955,N_10910,N_11805);
xor U12956 (N_12956,N_10507,N_11884);
or U12957 (N_12957,N_10709,N_11292);
xor U12958 (N_12958,N_11629,N_10549);
or U12959 (N_12959,N_11205,N_11365);
and U12960 (N_12960,N_11738,N_11263);
xnor U12961 (N_12961,N_10511,N_11978);
xor U12962 (N_12962,N_11981,N_10545);
and U12963 (N_12963,N_11226,N_11624);
nand U12964 (N_12964,N_11436,N_10812);
xnor U12965 (N_12965,N_10650,N_11502);
and U12966 (N_12966,N_10637,N_10556);
or U12967 (N_12967,N_10655,N_10762);
xnor U12968 (N_12968,N_10636,N_11850);
xnor U12969 (N_12969,N_11444,N_10542);
nand U12970 (N_12970,N_11213,N_11791);
nand U12971 (N_12971,N_11902,N_11098);
and U12972 (N_12972,N_10858,N_10998);
nand U12973 (N_12973,N_11498,N_11584);
and U12974 (N_12974,N_10563,N_11143);
and U12975 (N_12975,N_10518,N_11487);
nand U12976 (N_12976,N_10624,N_11278);
nor U12977 (N_12977,N_11542,N_11844);
xor U12978 (N_12978,N_10843,N_11403);
nor U12979 (N_12979,N_11142,N_11030);
or U12980 (N_12980,N_10838,N_10531);
nor U12981 (N_12981,N_11441,N_11824);
or U12982 (N_12982,N_11054,N_11521);
or U12983 (N_12983,N_10984,N_10912);
or U12984 (N_12984,N_10943,N_11109);
or U12985 (N_12985,N_11529,N_10600);
nand U12986 (N_12986,N_10889,N_11870);
nor U12987 (N_12987,N_11517,N_10523);
xor U12988 (N_12988,N_10763,N_10783);
nor U12989 (N_12989,N_11325,N_10704);
xnor U12990 (N_12990,N_10874,N_11722);
xnor U12991 (N_12991,N_10915,N_11921);
xor U12992 (N_12992,N_11127,N_10895);
nor U12993 (N_12993,N_10986,N_10578);
nor U12994 (N_12994,N_10848,N_11664);
and U12995 (N_12995,N_10615,N_11346);
and U12996 (N_12996,N_11170,N_10747);
nand U12997 (N_12997,N_10520,N_11621);
and U12998 (N_12998,N_10775,N_11378);
xnor U12999 (N_12999,N_10567,N_10995);
xor U13000 (N_13000,N_11906,N_11208);
or U13001 (N_13001,N_10957,N_10741);
and U13002 (N_13002,N_11917,N_11520);
or U13003 (N_13003,N_10961,N_11718);
nand U13004 (N_13004,N_11909,N_11850);
xor U13005 (N_13005,N_10783,N_11869);
nand U13006 (N_13006,N_11251,N_11626);
and U13007 (N_13007,N_10553,N_11706);
nand U13008 (N_13008,N_11491,N_11706);
or U13009 (N_13009,N_10836,N_11409);
nor U13010 (N_13010,N_10615,N_10991);
nor U13011 (N_13011,N_10916,N_11765);
xnor U13012 (N_13012,N_10790,N_11667);
nor U13013 (N_13013,N_11476,N_10864);
nor U13014 (N_13014,N_10861,N_11266);
or U13015 (N_13015,N_11734,N_11091);
nand U13016 (N_13016,N_11298,N_11459);
nand U13017 (N_13017,N_11084,N_10569);
nand U13018 (N_13018,N_11643,N_11579);
nand U13019 (N_13019,N_11125,N_10930);
or U13020 (N_13020,N_10824,N_10516);
nand U13021 (N_13021,N_11374,N_10909);
nor U13022 (N_13022,N_11063,N_11385);
and U13023 (N_13023,N_11470,N_10908);
xor U13024 (N_13024,N_11479,N_11207);
nor U13025 (N_13025,N_11258,N_11540);
or U13026 (N_13026,N_11516,N_10518);
or U13027 (N_13027,N_10956,N_10902);
nor U13028 (N_13028,N_10587,N_11481);
xor U13029 (N_13029,N_11522,N_11264);
nor U13030 (N_13030,N_10870,N_11949);
or U13031 (N_13031,N_10861,N_11823);
nand U13032 (N_13032,N_10716,N_11113);
and U13033 (N_13033,N_11311,N_11690);
and U13034 (N_13034,N_10543,N_11062);
or U13035 (N_13035,N_10954,N_11251);
nor U13036 (N_13036,N_11481,N_11354);
and U13037 (N_13037,N_10621,N_11447);
nor U13038 (N_13038,N_11262,N_11080);
nor U13039 (N_13039,N_11147,N_11224);
and U13040 (N_13040,N_10926,N_10940);
or U13041 (N_13041,N_11819,N_10731);
or U13042 (N_13042,N_11305,N_11035);
nor U13043 (N_13043,N_11852,N_10928);
and U13044 (N_13044,N_11179,N_11545);
and U13045 (N_13045,N_11784,N_11933);
xnor U13046 (N_13046,N_11881,N_11942);
xor U13047 (N_13047,N_10807,N_10604);
and U13048 (N_13048,N_10989,N_11219);
nand U13049 (N_13049,N_10719,N_10813);
nor U13050 (N_13050,N_10614,N_10515);
and U13051 (N_13051,N_11341,N_10680);
nor U13052 (N_13052,N_11101,N_11988);
xnor U13053 (N_13053,N_11715,N_11316);
and U13054 (N_13054,N_11098,N_10513);
and U13055 (N_13055,N_10743,N_11807);
nor U13056 (N_13056,N_10899,N_11183);
nand U13057 (N_13057,N_10782,N_10835);
nand U13058 (N_13058,N_10941,N_11555);
nand U13059 (N_13059,N_11423,N_11985);
and U13060 (N_13060,N_11233,N_11323);
nand U13061 (N_13061,N_10630,N_11522);
and U13062 (N_13062,N_11929,N_11394);
and U13063 (N_13063,N_11602,N_11105);
nor U13064 (N_13064,N_10929,N_11886);
nor U13065 (N_13065,N_10603,N_10532);
or U13066 (N_13066,N_11871,N_10574);
xor U13067 (N_13067,N_11330,N_10766);
or U13068 (N_13068,N_11810,N_11139);
nor U13069 (N_13069,N_11249,N_10973);
xor U13070 (N_13070,N_11200,N_11742);
nor U13071 (N_13071,N_11140,N_10869);
or U13072 (N_13072,N_11905,N_10714);
xor U13073 (N_13073,N_10754,N_10595);
xor U13074 (N_13074,N_10844,N_10699);
nand U13075 (N_13075,N_10808,N_10556);
xnor U13076 (N_13076,N_11253,N_11917);
nand U13077 (N_13077,N_11347,N_11409);
nor U13078 (N_13078,N_10901,N_10841);
and U13079 (N_13079,N_10888,N_10934);
nor U13080 (N_13080,N_10866,N_11541);
nand U13081 (N_13081,N_10504,N_10514);
or U13082 (N_13082,N_10958,N_11722);
xnor U13083 (N_13083,N_11039,N_10664);
and U13084 (N_13084,N_11047,N_11102);
and U13085 (N_13085,N_10842,N_11466);
nand U13086 (N_13086,N_10903,N_11502);
nand U13087 (N_13087,N_11452,N_10642);
xnor U13088 (N_13088,N_11483,N_11712);
and U13089 (N_13089,N_11940,N_10875);
nand U13090 (N_13090,N_11551,N_11593);
or U13091 (N_13091,N_11436,N_11764);
nor U13092 (N_13092,N_10674,N_11654);
or U13093 (N_13093,N_11948,N_11435);
nand U13094 (N_13094,N_11244,N_11811);
nor U13095 (N_13095,N_11146,N_11980);
nor U13096 (N_13096,N_10752,N_11417);
or U13097 (N_13097,N_11562,N_10629);
nor U13098 (N_13098,N_11408,N_10589);
or U13099 (N_13099,N_11466,N_11871);
nand U13100 (N_13100,N_11681,N_11119);
or U13101 (N_13101,N_10823,N_10560);
nand U13102 (N_13102,N_11033,N_11008);
nand U13103 (N_13103,N_11616,N_10986);
xor U13104 (N_13104,N_11518,N_11575);
and U13105 (N_13105,N_11919,N_11243);
and U13106 (N_13106,N_11260,N_10808);
and U13107 (N_13107,N_11325,N_11476);
nor U13108 (N_13108,N_10556,N_11006);
and U13109 (N_13109,N_11712,N_11934);
or U13110 (N_13110,N_11333,N_11052);
nand U13111 (N_13111,N_11474,N_11285);
nor U13112 (N_13112,N_11996,N_11411);
nor U13113 (N_13113,N_11897,N_10575);
nand U13114 (N_13114,N_10804,N_10761);
and U13115 (N_13115,N_11455,N_10953);
nand U13116 (N_13116,N_11409,N_10880);
nand U13117 (N_13117,N_11110,N_11757);
and U13118 (N_13118,N_10966,N_11717);
or U13119 (N_13119,N_10535,N_11827);
and U13120 (N_13120,N_11821,N_11003);
or U13121 (N_13121,N_10879,N_10950);
nor U13122 (N_13122,N_10647,N_11250);
or U13123 (N_13123,N_10631,N_10761);
and U13124 (N_13124,N_11856,N_11514);
and U13125 (N_13125,N_11560,N_11487);
or U13126 (N_13126,N_10911,N_11970);
or U13127 (N_13127,N_11955,N_10618);
or U13128 (N_13128,N_10634,N_10832);
nor U13129 (N_13129,N_11023,N_11744);
and U13130 (N_13130,N_11146,N_10684);
and U13131 (N_13131,N_11545,N_11359);
or U13132 (N_13132,N_10719,N_10630);
and U13133 (N_13133,N_11667,N_10657);
nand U13134 (N_13134,N_10612,N_10604);
nand U13135 (N_13135,N_11463,N_11280);
nor U13136 (N_13136,N_11052,N_11690);
and U13137 (N_13137,N_10722,N_11606);
or U13138 (N_13138,N_10813,N_11769);
nor U13139 (N_13139,N_11345,N_10659);
xnor U13140 (N_13140,N_11493,N_10926);
nand U13141 (N_13141,N_11402,N_11073);
nand U13142 (N_13142,N_11644,N_11610);
xor U13143 (N_13143,N_11065,N_11688);
and U13144 (N_13144,N_11626,N_11634);
and U13145 (N_13145,N_11594,N_11921);
nor U13146 (N_13146,N_11262,N_11127);
nor U13147 (N_13147,N_10888,N_10640);
nor U13148 (N_13148,N_10640,N_11320);
xor U13149 (N_13149,N_10940,N_11183);
nor U13150 (N_13150,N_11124,N_10683);
or U13151 (N_13151,N_11231,N_10602);
and U13152 (N_13152,N_11202,N_11166);
or U13153 (N_13153,N_11970,N_11128);
and U13154 (N_13154,N_11801,N_10759);
xor U13155 (N_13155,N_11257,N_11873);
and U13156 (N_13156,N_10593,N_11566);
nand U13157 (N_13157,N_11045,N_10929);
nand U13158 (N_13158,N_11286,N_11019);
nor U13159 (N_13159,N_11017,N_11256);
or U13160 (N_13160,N_11218,N_11354);
nor U13161 (N_13161,N_11076,N_11260);
nand U13162 (N_13162,N_11621,N_11874);
nand U13163 (N_13163,N_10986,N_11414);
nand U13164 (N_13164,N_11688,N_11949);
nor U13165 (N_13165,N_11233,N_11101);
nand U13166 (N_13166,N_11409,N_11384);
and U13167 (N_13167,N_11622,N_11099);
and U13168 (N_13168,N_11053,N_11046);
xor U13169 (N_13169,N_11277,N_10661);
nor U13170 (N_13170,N_11889,N_10880);
xnor U13171 (N_13171,N_11215,N_10590);
nand U13172 (N_13172,N_11658,N_11046);
nor U13173 (N_13173,N_11030,N_10981);
and U13174 (N_13174,N_10840,N_11536);
or U13175 (N_13175,N_11911,N_11136);
and U13176 (N_13176,N_10691,N_11742);
or U13177 (N_13177,N_11419,N_10584);
and U13178 (N_13178,N_11778,N_11542);
nand U13179 (N_13179,N_11056,N_11579);
nor U13180 (N_13180,N_10631,N_11652);
or U13181 (N_13181,N_11965,N_10606);
nand U13182 (N_13182,N_11007,N_11317);
nand U13183 (N_13183,N_11988,N_11830);
or U13184 (N_13184,N_11770,N_10616);
nor U13185 (N_13185,N_11196,N_11676);
or U13186 (N_13186,N_11349,N_10661);
nor U13187 (N_13187,N_10974,N_10630);
xnor U13188 (N_13188,N_11975,N_10860);
xor U13189 (N_13189,N_10739,N_11471);
and U13190 (N_13190,N_10725,N_10807);
and U13191 (N_13191,N_10653,N_11531);
nor U13192 (N_13192,N_11747,N_11982);
nand U13193 (N_13193,N_10522,N_11021);
nor U13194 (N_13194,N_11407,N_11334);
xnor U13195 (N_13195,N_11042,N_11438);
and U13196 (N_13196,N_11435,N_11154);
nor U13197 (N_13197,N_10896,N_10783);
nand U13198 (N_13198,N_11108,N_10929);
nor U13199 (N_13199,N_11714,N_11526);
and U13200 (N_13200,N_11395,N_11190);
or U13201 (N_13201,N_10770,N_11823);
and U13202 (N_13202,N_11275,N_11098);
or U13203 (N_13203,N_11503,N_11105);
nand U13204 (N_13204,N_10757,N_11455);
or U13205 (N_13205,N_10929,N_11000);
nor U13206 (N_13206,N_11008,N_11937);
xor U13207 (N_13207,N_11818,N_11824);
or U13208 (N_13208,N_11953,N_11155);
nand U13209 (N_13209,N_10549,N_11181);
and U13210 (N_13210,N_10572,N_11214);
nand U13211 (N_13211,N_11742,N_10723);
nand U13212 (N_13212,N_11799,N_11261);
or U13213 (N_13213,N_10942,N_11016);
nor U13214 (N_13214,N_11848,N_11130);
and U13215 (N_13215,N_11712,N_11911);
nor U13216 (N_13216,N_10737,N_11072);
and U13217 (N_13217,N_11494,N_10697);
or U13218 (N_13218,N_11388,N_11385);
or U13219 (N_13219,N_11303,N_10953);
nor U13220 (N_13220,N_11386,N_11302);
xnor U13221 (N_13221,N_11753,N_10835);
or U13222 (N_13222,N_11719,N_11333);
xnor U13223 (N_13223,N_10795,N_10737);
nor U13224 (N_13224,N_10724,N_11506);
and U13225 (N_13225,N_10797,N_10735);
xor U13226 (N_13226,N_11035,N_11588);
xor U13227 (N_13227,N_10909,N_10823);
and U13228 (N_13228,N_11018,N_11986);
and U13229 (N_13229,N_11566,N_11961);
nor U13230 (N_13230,N_11651,N_10946);
nand U13231 (N_13231,N_10593,N_11852);
nand U13232 (N_13232,N_11225,N_10935);
and U13233 (N_13233,N_11604,N_11904);
xor U13234 (N_13234,N_11043,N_11841);
and U13235 (N_13235,N_11115,N_11092);
nor U13236 (N_13236,N_11256,N_11844);
xnor U13237 (N_13237,N_11720,N_11521);
xor U13238 (N_13238,N_11918,N_10604);
nand U13239 (N_13239,N_10730,N_11121);
or U13240 (N_13240,N_11777,N_11048);
nor U13241 (N_13241,N_10520,N_11146);
xor U13242 (N_13242,N_10927,N_10639);
nand U13243 (N_13243,N_11130,N_11245);
nand U13244 (N_13244,N_10966,N_10834);
or U13245 (N_13245,N_11227,N_11742);
nor U13246 (N_13246,N_10529,N_11963);
nand U13247 (N_13247,N_11236,N_11080);
and U13248 (N_13248,N_11736,N_10723);
and U13249 (N_13249,N_11416,N_11283);
xnor U13250 (N_13250,N_11429,N_11080);
xor U13251 (N_13251,N_11237,N_10684);
nor U13252 (N_13252,N_11550,N_11525);
nor U13253 (N_13253,N_10736,N_11358);
and U13254 (N_13254,N_11452,N_10652);
and U13255 (N_13255,N_11184,N_11995);
and U13256 (N_13256,N_11333,N_11537);
nor U13257 (N_13257,N_11072,N_11906);
nand U13258 (N_13258,N_11981,N_11027);
or U13259 (N_13259,N_11709,N_11615);
nand U13260 (N_13260,N_11547,N_10674);
and U13261 (N_13261,N_10671,N_11481);
or U13262 (N_13262,N_11288,N_10861);
or U13263 (N_13263,N_11069,N_10633);
or U13264 (N_13264,N_11358,N_11508);
or U13265 (N_13265,N_11052,N_10791);
nand U13266 (N_13266,N_11044,N_11778);
nor U13267 (N_13267,N_11702,N_11487);
and U13268 (N_13268,N_10710,N_11610);
nand U13269 (N_13269,N_11799,N_10534);
and U13270 (N_13270,N_11799,N_11130);
or U13271 (N_13271,N_10890,N_11595);
nor U13272 (N_13272,N_11982,N_10555);
nand U13273 (N_13273,N_10798,N_11854);
nor U13274 (N_13274,N_11817,N_11608);
nand U13275 (N_13275,N_10656,N_10768);
nand U13276 (N_13276,N_11378,N_11575);
nand U13277 (N_13277,N_11262,N_11931);
xor U13278 (N_13278,N_10880,N_10658);
nand U13279 (N_13279,N_10757,N_11258);
nor U13280 (N_13280,N_11097,N_11165);
xor U13281 (N_13281,N_10696,N_10739);
nor U13282 (N_13282,N_11755,N_11764);
xor U13283 (N_13283,N_11972,N_10588);
or U13284 (N_13284,N_11300,N_11445);
and U13285 (N_13285,N_10803,N_11361);
or U13286 (N_13286,N_10744,N_10575);
nor U13287 (N_13287,N_10993,N_11601);
nand U13288 (N_13288,N_11744,N_10593);
and U13289 (N_13289,N_11119,N_11540);
or U13290 (N_13290,N_11910,N_10948);
and U13291 (N_13291,N_10898,N_11326);
nor U13292 (N_13292,N_11985,N_10749);
nand U13293 (N_13293,N_10684,N_11785);
and U13294 (N_13294,N_11506,N_10734);
nand U13295 (N_13295,N_11195,N_11647);
xor U13296 (N_13296,N_11942,N_11660);
xnor U13297 (N_13297,N_10568,N_10553);
nor U13298 (N_13298,N_11549,N_11503);
nand U13299 (N_13299,N_11991,N_10613);
xnor U13300 (N_13300,N_10667,N_11106);
xnor U13301 (N_13301,N_11800,N_10552);
or U13302 (N_13302,N_11617,N_11218);
nor U13303 (N_13303,N_11052,N_11145);
nand U13304 (N_13304,N_11671,N_11447);
nand U13305 (N_13305,N_10932,N_10877);
nor U13306 (N_13306,N_11984,N_10649);
or U13307 (N_13307,N_10606,N_11657);
and U13308 (N_13308,N_11595,N_11520);
xnor U13309 (N_13309,N_11833,N_11924);
nor U13310 (N_13310,N_11229,N_11732);
nor U13311 (N_13311,N_11054,N_10877);
nor U13312 (N_13312,N_11576,N_11284);
and U13313 (N_13313,N_11139,N_11747);
and U13314 (N_13314,N_10648,N_11141);
nand U13315 (N_13315,N_11255,N_11672);
xor U13316 (N_13316,N_11922,N_11591);
xor U13317 (N_13317,N_11348,N_11759);
xnor U13318 (N_13318,N_11801,N_10961);
and U13319 (N_13319,N_10575,N_11367);
nand U13320 (N_13320,N_11027,N_10694);
nand U13321 (N_13321,N_11978,N_11220);
and U13322 (N_13322,N_11291,N_11793);
or U13323 (N_13323,N_11884,N_10722);
nor U13324 (N_13324,N_11189,N_10715);
xor U13325 (N_13325,N_11586,N_11098);
nor U13326 (N_13326,N_10954,N_11385);
nand U13327 (N_13327,N_10852,N_11427);
nand U13328 (N_13328,N_11265,N_10718);
xnor U13329 (N_13329,N_11297,N_10965);
xnor U13330 (N_13330,N_11834,N_10960);
and U13331 (N_13331,N_11410,N_10585);
xor U13332 (N_13332,N_11400,N_11717);
xnor U13333 (N_13333,N_11193,N_11722);
xor U13334 (N_13334,N_10551,N_11286);
or U13335 (N_13335,N_10916,N_11964);
xnor U13336 (N_13336,N_10737,N_10965);
and U13337 (N_13337,N_11075,N_11281);
nand U13338 (N_13338,N_11404,N_11992);
xor U13339 (N_13339,N_10877,N_11434);
nor U13340 (N_13340,N_11397,N_11424);
nor U13341 (N_13341,N_11624,N_11119);
xnor U13342 (N_13342,N_10889,N_10817);
nand U13343 (N_13343,N_11361,N_11259);
nand U13344 (N_13344,N_10950,N_10757);
and U13345 (N_13345,N_10644,N_11513);
or U13346 (N_13346,N_11295,N_10921);
and U13347 (N_13347,N_11810,N_11660);
nor U13348 (N_13348,N_11846,N_11533);
nor U13349 (N_13349,N_11795,N_10808);
and U13350 (N_13350,N_11053,N_11236);
xor U13351 (N_13351,N_11172,N_10545);
nor U13352 (N_13352,N_11932,N_10984);
or U13353 (N_13353,N_11825,N_11915);
nand U13354 (N_13354,N_11247,N_11507);
nor U13355 (N_13355,N_10654,N_11146);
nand U13356 (N_13356,N_10934,N_11499);
nor U13357 (N_13357,N_10533,N_11354);
or U13358 (N_13358,N_11569,N_10729);
xnor U13359 (N_13359,N_10966,N_11501);
and U13360 (N_13360,N_11348,N_10640);
or U13361 (N_13361,N_11410,N_11253);
or U13362 (N_13362,N_11762,N_10709);
and U13363 (N_13363,N_10946,N_11680);
xor U13364 (N_13364,N_11665,N_10886);
nor U13365 (N_13365,N_11202,N_10690);
nor U13366 (N_13366,N_11136,N_11065);
or U13367 (N_13367,N_11435,N_11165);
nor U13368 (N_13368,N_11262,N_11172);
and U13369 (N_13369,N_11666,N_11222);
or U13370 (N_13370,N_10631,N_10651);
nand U13371 (N_13371,N_11509,N_11360);
nor U13372 (N_13372,N_11000,N_11712);
nand U13373 (N_13373,N_11638,N_11277);
or U13374 (N_13374,N_11560,N_11985);
or U13375 (N_13375,N_11355,N_11243);
or U13376 (N_13376,N_10601,N_11627);
nor U13377 (N_13377,N_10863,N_11357);
and U13378 (N_13378,N_11413,N_10514);
or U13379 (N_13379,N_10587,N_10974);
or U13380 (N_13380,N_10620,N_10920);
nand U13381 (N_13381,N_11775,N_10763);
nand U13382 (N_13382,N_10809,N_11428);
xor U13383 (N_13383,N_11084,N_10583);
nor U13384 (N_13384,N_10968,N_11500);
and U13385 (N_13385,N_10902,N_11272);
nor U13386 (N_13386,N_10582,N_10692);
or U13387 (N_13387,N_10788,N_10990);
nand U13388 (N_13388,N_11845,N_11238);
and U13389 (N_13389,N_11513,N_11424);
or U13390 (N_13390,N_10600,N_10904);
and U13391 (N_13391,N_10968,N_11619);
xor U13392 (N_13392,N_11163,N_10990);
nand U13393 (N_13393,N_10669,N_11334);
xnor U13394 (N_13394,N_11750,N_11202);
nor U13395 (N_13395,N_11541,N_11723);
and U13396 (N_13396,N_11453,N_11093);
and U13397 (N_13397,N_11429,N_10678);
xor U13398 (N_13398,N_10681,N_11180);
nor U13399 (N_13399,N_11737,N_11334);
nand U13400 (N_13400,N_11144,N_11645);
nor U13401 (N_13401,N_11107,N_11541);
and U13402 (N_13402,N_10634,N_11221);
or U13403 (N_13403,N_10617,N_11793);
or U13404 (N_13404,N_11100,N_10738);
nand U13405 (N_13405,N_11463,N_11075);
xnor U13406 (N_13406,N_11231,N_11866);
and U13407 (N_13407,N_10837,N_11310);
and U13408 (N_13408,N_11875,N_10713);
nor U13409 (N_13409,N_11480,N_10736);
or U13410 (N_13410,N_10718,N_11306);
or U13411 (N_13411,N_10865,N_11465);
or U13412 (N_13412,N_10688,N_10923);
or U13413 (N_13413,N_10946,N_11498);
xor U13414 (N_13414,N_10846,N_10537);
xnor U13415 (N_13415,N_10852,N_11136);
xnor U13416 (N_13416,N_10568,N_10738);
nor U13417 (N_13417,N_11869,N_10811);
xor U13418 (N_13418,N_11482,N_10798);
and U13419 (N_13419,N_11879,N_11358);
nand U13420 (N_13420,N_10519,N_10825);
and U13421 (N_13421,N_11708,N_10727);
or U13422 (N_13422,N_11101,N_10995);
or U13423 (N_13423,N_11037,N_10660);
nor U13424 (N_13424,N_11209,N_10532);
nand U13425 (N_13425,N_11325,N_11596);
nor U13426 (N_13426,N_10542,N_11269);
or U13427 (N_13427,N_11567,N_11216);
or U13428 (N_13428,N_11329,N_11171);
xnor U13429 (N_13429,N_11251,N_11761);
nand U13430 (N_13430,N_11703,N_10611);
nor U13431 (N_13431,N_11088,N_10740);
xor U13432 (N_13432,N_11639,N_11223);
xor U13433 (N_13433,N_11125,N_11687);
nand U13434 (N_13434,N_11492,N_10806);
or U13435 (N_13435,N_11372,N_11191);
xnor U13436 (N_13436,N_11230,N_11065);
nor U13437 (N_13437,N_10753,N_11227);
or U13438 (N_13438,N_11321,N_10553);
nand U13439 (N_13439,N_11429,N_10513);
and U13440 (N_13440,N_11238,N_10914);
or U13441 (N_13441,N_10966,N_11020);
nor U13442 (N_13442,N_11136,N_11151);
or U13443 (N_13443,N_11626,N_11035);
or U13444 (N_13444,N_11352,N_10932);
nor U13445 (N_13445,N_11193,N_10627);
nand U13446 (N_13446,N_10965,N_11580);
nor U13447 (N_13447,N_10946,N_10777);
xor U13448 (N_13448,N_11744,N_11696);
or U13449 (N_13449,N_10938,N_10820);
nor U13450 (N_13450,N_10606,N_11855);
and U13451 (N_13451,N_10876,N_10547);
nor U13452 (N_13452,N_11883,N_11408);
and U13453 (N_13453,N_11310,N_11769);
or U13454 (N_13454,N_11968,N_10969);
nor U13455 (N_13455,N_11462,N_11015);
xor U13456 (N_13456,N_11343,N_10716);
and U13457 (N_13457,N_11300,N_11000);
nor U13458 (N_13458,N_11119,N_11868);
nand U13459 (N_13459,N_11702,N_11851);
and U13460 (N_13460,N_10848,N_11450);
nor U13461 (N_13461,N_11023,N_10731);
xor U13462 (N_13462,N_11027,N_11199);
nor U13463 (N_13463,N_11196,N_11958);
and U13464 (N_13464,N_10637,N_11020);
nand U13465 (N_13465,N_10500,N_10812);
nor U13466 (N_13466,N_10668,N_11336);
and U13467 (N_13467,N_11124,N_11871);
or U13468 (N_13468,N_11797,N_11512);
and U13469 (N_13469,N_11596,N_10721);
nor U13470 (N_13470,N_10753,N_10942);
nor U13471 (N_13471,N_11300,N_11088);
xor U13472 (N_13472,N_10685,N_10829);
xnor U13473 (N_13473,N_11433,N_11857);
nor U13474 (N_13474,N_11838,N_11776);
and U13475 (N_13475,N_11454,N_11106);
xor U13476 (N_13476,N_11152,N_11924);
nor U13477 (N_13477,N_11839,N_11420);
or U13478 (N_13478,N_11292,N_11338);
nor U13479 (N_13479,N_11050,N_11103);
and U13480 (N_13480,N_11351,N_11759);
nor U13481 (N_13481,N_10659,N_11788);
and U13482 (N_13482,N_10702,N_10922);
or U13483 (N_13483,N_11207,N_11109);
and U13484 (N_13484,N_11662,N_11272);
nand U13485 (N_13485,N_11221,N_11189);
xnor U13486 (N_13486,N_11095,N_10746);
xor U13487 (N_13487,N_11533,N_10765);
and U13488 (N_13488,N_11935,N_10671);
nor U13489 (N_13489,N_10633,N_10971);
and U13490 (N_13490,N_11140,N_10929);
or U13491 (N_13491,N_11673,N_11127);
nand U13492 (N_13492,N_10713,N_10586);
and U13493 (N_13493,N_11266,N_11582);
xnor U13494 (N_13494,N_10591,N_11870);
nand U13495 (N_13495,N_10766,N_10719);
or U13496 (N_13496,N_11462,N_10589);
nand U13497 (N_13497,N_11271,N_11475);
xor U13498 (N_13498,N_11526,N_11849);
or U13499 (N_13499,N_11979,N_11652);
nand U13500 (N_13500,N_13114,N_12564);
nor U13501 (N_13501,N_12818,N_12924);
xnor U13502 (N_13502,N_13397,N_13310);
nor U13503 (N_13503,N_13041,N_12788);
and U13504 (N_13504,N_13147,N_12215);
xor U13505 (N_13505,N_12599,N_12542);
or U13506 (N_13506,N_13103,N_13115);
nor U13507 (N_13507,N_13472,N_12834);
xor U13508 (N_13508,N_12546,N_12668);
xnor U13509 (N_13509,N_12034,N_13182);
nor U13510 (N_13510,N_12868,N_12961);
or U13511 (N_13511,N_12429,N_12410);
xor U13512 (N_13512,N_13307,N_12880);
nand U13513 (N_13513,N_13411,N_12044);
nand U13514 (N_13514,N_12396,N_13415);
nor U13515 (N_13515,N_12799,N_12297);
and U13516 (N_13516,N_12979,N_13269);
nor U13517 (N_13517,N_13490,N_12060);
nand U13518 (N_13518,N_12755,N_12790);
nor U13519 (N_13519,N_12512,N_13420);
nor U13520 (N_13520,N_13018,N_12246);
nand U13521 (N_13521,N_12813,N_13121);
or U13522 (N_13522,N_13130,N_12758);
nand U13523 (N_13523,N_12761,N_12481);
or U13524 (N_13524,N_13061,N_12404);
or U13525 (N_13525,N_13045,N_12915);
and U13526 (N_13526,N_13488,N_12837);
nor U13527 (N_13527,N_12316,N_12814);
nand U13528 (N_13528,N_13142,N_13006);
nand U13529 (N_13529,N_13199,N_12402);
nand U13530 (N_13530,N_12858,N_13205);
and U13531 (N_13531,N_12072,N_13025);
and U13532 (N_13532,N_13227,N_13403);
and U13533 (N_13533,N_12738,N_12647);
nand U13534 (N_13534,N_13105,N_12077);
xnor U13535 (N_13535,N_13438,N_12025);
xnor U13536 (N_13536,N_13470,N_12553);
or U13537 (N_13537,N_13497,N_12812);
and U13538 (N_13538,N_12832,N_13391);
nand U13539 (N_13539,N_13418,N_12590);
or U13540 (N_13540,N_13172,N_13480);
xor U13541 (N_13541,N_12145,N_12888);
nor U13542 (N_13542,N_12510,N_12356);
nor U13543 (N_13543,N_12259,N_12796);
or U13544 (N_13544,N_12664,N_12511);
and U13545 (N_13545,N_13355,N_12539);
nor U13546 (N_13546,N_12482,N_13020);
and U13547 (N_13547,N_12754,N_12719);
and U13548 (N_13548,N_13184,N_12631);
nand U13549 (N_13549,N_12211,N_12384);
or U13550 (N_13550,N_13486,N_13186);
and U13551 (N_13551,N_12919,N_13311);
nor U13552 (N_13552,N_12112,N_12596);
nand U13553 (N_13553,N_13487,N_12697);
and U13554 (N_13554,N_12670,N_12896);
nand U13555 (N_13555,N_13316,N_12008);
or U13556 (N_13556,N_13251,N_13402);
or U13557 (N_13557,N_13027,N_13323);
nor U13558 (N_13558,N_12016,N_12760);
xnor U13559 (N_13559,N_12126,N_13209);
nor U13560 (N_13560,N_13382,N_12020);
and U13561 (N_13561,N_12945,N_13279);
xnor U13562 (N_13562,N_12521,N_13240);
nor U13563 (N_13563,N_12375,N_13309);
nand U13564 (N_13564,N_13318,N_12161);
nand U13565 (N_13565,N_12256,N_12274);
and U13566 (N_13566,N_12809,N_13445);
nor U13567 (N_13567,N_12932,N_12684);
or U13568 (N_13568,N_13262,N_13000);
nand U13569 (N_13569,N_12492,N_12759);
or U13570 (N_13570,N_12876,N_12844);
xnor U13571 (N_13571,N_13482,N_12966);
nor U13572 (N_13572,N_12476,N_12420);
xor U13573 (N_13573,N_12214,N_12722);
nor U13574 (N_13574,N_12720,N_12323);
or U13575 (N_13575,N_12373,N_13484);
nor U13576 (N_13576,N_13376,N_13293);
and U13577 (N_13577,N_13417,N_13428);
nor U13578 (N_13578,N_13167,N_13283);
nand U13579 (N_13579,N_12332,N_12107);
and U13580 (N_13580,N_12391,N_12672);
nor U13581 (N_13581,N_13166,N_13008);
or U13582 (N_13582,N_12886,N_12456);
nand U13583 (N_13583,N_13052,N_13434);
or U13584 (N_13584,N_12347,N_13195);
xor U13585 (N_13585,N_13098,N_12284);
xnor U13586 (N_13586,N_12475,N_12007);
nand U13587 (N_13587,N_13222,N_12643);
nor U13588 (N_13588,N_12198,N_12047);
nand U13589 (N_13589,N_12645,N_12383);
xnor U13590 (N_13590,N_13196,N_13270);
or U13591 (N_13591,N_13046,N_12787);
nand U13592 (N_13592,N_12341,N_12368);
and U13593 (N_13593,N_12207,N_12298);
and U13594 (N_13594,N_13230,N_12073);
nand U13595 (N_13595,N_12202,N_13327);
nand U13596 (N_13596,N_12319,N_12763);
nand U13597 (N_13597,N_12312,N_13024);
nand U13598 (N_13598,N_13254,N_13232);
and U13599 (N_13599,N_12301,N_12851);
and U13600 (N_13600,N_12270,N_12946);
nand U13601 (N_13601,N_12650,N_12639);
xnor U13602 (N_13602,N_12432,N_12150);
nand U13603 (N_13603,N_12283,N_12750);
nand U13604 (N_13604,N_13469,N_12694);
nor U13605 (N_13605,N_13449,N_13407);
and U13606 (N_13606,N_12223,N_12955);
xor U13607 (N_13607,N_12495,N_12068);
xor U13608 (N_13608,N_12351,N_13109);
nor U13609 (N_13609,N_13285,N_12209);
xnor U13610 (N_13610,N_13080,N_13120);
or U13611 (N_13611,N_12033,N_13248);
nand U13612 (N_13612,N_12716,N_13009);
and U13613 (N_13613,N_12773,N_12948);
and U13614 (N_13614,N_12582,N_12499);
or U13615 (N_13615,N_13047,N_12522);
nand U13616 (N_13616,N_12036,N_12300);
nand U13617 (N_13617,N_12046,N_12914);
and U13618 (N_13618,N_12290,N_12556);
and U13619 (N_13619,N_13463,N_12620);
and U13620 (N_13620,N_12305,N_13335);
or U13621 (N_13621,N_12689,N_12731);
or U13622 (N_13622,N_13341,N_13457);
nor U13623 (N_13623,N_12823,N_12504);
nor U13624 (N_13624,N_13298,N_12792);
nand U13625 (N_13625,N_13158,N_12137);
nor U13626 (N_13626,N_12217,N_12528);
or U13627 (N_13627,N_13042,N_12062);
xnor U13628 (N_13628,N_12767,N_12882);
nand U13629 (N_13629,N_12050,N_12236);
xnor U13630 (N_13630,N_12573,N_12286);
or U13631 (N_13631,N_12142,N_12359);
and U13632 (N_13632,N_12221,N_12729);
nor U13633 (N_13633,N_12540,N_12218);
and U13634 (N_13634,N_12801,N_12369);
xnor U13635 (N_13635,N_12533,N_12588);
nor U13636 (N_13636,N_12996,N_13342);
nor U13637 (N_13637,N_12190,N_13108);
nand U13638 (N_13638,N_12013,N_12193);
nor U13639 (N_13639,N_12224,N_13149);
and U13640 (N_13640,N_12904,N_12635);
nor U13641 (N_13641,N_13243,N_13221);
nor U13642 (N_13642,N_12802,N_12695);
xnor U13643 (N_13643,N_12313,N_13344);
nand U13644 (N_13644,N_13040,N_13371);
or U13645 (N_13645,N_12155,N_12531);
nor U13646 (N_13646,N_12096,N_12632);
nand U13647 (N_13647,N_12944,N_12345);
xor U13648 (N_13648,N_13078,N_12029);
xnor U13649 (N_13649,N_13125,N_13067);
xnor U13650 (N_13650,N_12774,N_12417);
and U13651 (N_13651,N_13264,N_13494);
nor U13652 (N_13652,N_12600,N_12080);
or U13653 (N_13653,N_12192,N_12976);
nand U13654 (N_13654,N_13132,N_12387);
or U13655 (N_13655,N_12304,N_13295);
and U13656 (N_13656,N_12999,N_13016);
and U13657 (N_13657,N_12881,N_13198);
nor U13658 (N_13658,N_12199,N_12532);
nor U13659 (N_13659,N_13441,N_12690);
nor U13660 (N_13660,N_13287,N_13225);
nor U13661 (N_13661,N_13328,N_13276);
nand U13662 (N_13662,N_12120,N_12807);
nor U13663 (N_13663,N_12901,N_13210);
and U13664 (N_13664,N_12595,N_12965);
nor U13665 (N_13665,N_12674,N_12343);
and U13666 (N_13666,N_12163,N_12705);
or U13667 (N_13667,N_12435,N_12905);
and U13668 (N_13668,N_13259,N_12929);
or U13669 (N_13669,N_13477,N_12831);
xnor U13670 (N_13670,N_12365,N_12213);
nor U13671 (N_13671,N_12841,N_12865);
nand U13672 (N_13672,N_12032,N_13357);
or U13673 (N_13673,N_12911,N_13206);
or U13674 (N_13674,N_12744,N_13267);
and U13675 (N_13675,N_13491,N_13346);
nand U13676 (N_13676,N_12430,N_12717);
xnor U13677 (N_13677,N_12870,N_13272);
nand U13678 (N_13678,N_12361,N_12793);
and U13679 (N_13679,N_12201,N_13003);
and U13680 (N_13680,N_12418,N_12503);
and U13681 (N_13681,N_13011,N_13313);
xnor U13682 (N_13682,N_12994,N_13076);
xnor U13683 (N_13683,N_12604,N_13385);
xor U13684 (N_13684,N_13197,N_12266);
nor U13685 (N_13685,N_12083,N_13324);
or U13686 (N_13686,N_12063,N_12415);
and U13687 (N_13687,N_12940,N_13127);
nand U13688 (N_13688,N_12395,N_13292);
nand U13689 (N_13689,N_13116,N_13029);
xnor U13690 (N_13690,N_12655,N_12459);
or U13691 (N_13691,N_12329,N_12835);
xor U13692 (N_13692,N_12562,N_12017);
nor U13693 (N_13693,N_12607,N_12644);
nand U13694 (N_13694,N_12977,N_12254);
or U13695 (N_13695,N_12115,N_12464);
or U13696 (N_13696,N_13348,N_13201);
nor U13697 (N_13697,N_13155,N_13377);
nand U13698 (N_13698,N_12563,N_12339);
nor U13699 (N_13699,N_12200,N_12229);
nor U13700 (N_13700,N_13375,N_12331);
xor U13701 (N_13701,N_13413,N_12815);
xnor U13702 (N_13702,N_13455,N_12354);
and U13703 (N_13703,N_13202,N_12134);
nand U13704 (N_13704,N_12446,N_12125);
and U13705 (N_13705,N_12123,N_13162);
nand U13706 (N_13706,N_12276,N_13138);
nor U13707 (N_13707,N_12678,N_12405);
or U13708 (N_13708,N_13352,N_12959);
xnor U13709 (N_13709,N_12550,N_12687);
or U13710 (N_13710,N_13414,N_13366);
nor U13711 (N_13711,N_12751,N_12691);
or U13712 (N_13712,N_13361,N_12450);
nor U13713 (N_13713,N_12916,N_13070);
or U13714 (N_13714,N_12637,N_12660);
or U13715 (N_13715,N_12547,N_13440);
and U13716 (N_13716,N_13235,N_12983);
nand U13717 (N_13717,N_12514,N_12900);
and U13718 (N_13718,N_13213,N_13435);
xor U13719 (N_13719,N_12930,N_12657);
and U13720 (N_13720,N_13443,N_12220);
nor U13721 (N_13721,N_13444,N_13056);
xnor U13722 (N_13722,N_13427,N_12454);
nand U13723 (N_13723,N_12838,N_12043);
or U13724 (N_13724,N_13203,N_13485);
and U13725 (N_13725,N_12128,N_13218);
or U13726 (N_13726,N_13333,N_12106);
nand U13727 (N_13727,N_12549,N_12537);
xor U13728 (N_13728,N_12167,N_13063);
nand U13729 (N_13729,N_12001,N_12127);
and U13730 (N_13730,N_13176,N_13146);
xnor U13731 (N_13731,N_12129,N_13296);
and U13732 (N_13732,N_12669,N_13388);
and U13733 (N_13733,N_12232,N_13392);
and U13734 (N_13734,N_12183,N_12548);
or U13735 (N_13735,N_13302,N_12421);
nor U13736 (N_13736,N_12673,N_13356);
nor U13737 (N_13737,N_12084,N_13161);
and U13738 (N_13738,N_12101,N_12640);
xnor U13739 (N_13739,N_12377,N_12071);
nand U13740 (N_13740,N_12749,N_13019);
nor U13741 (N_13741,N_12413,N_13153);
and U13742 (N_13742,N_13447,N_12656);
xor U13743 (N_13743,N_12642,N_12109);
and U13744 (N_13744,N_13073,N_12839);
nand U13745 (N_13745,N_12970,N_12630);
or U13746 (N_13746,N_12140,N_12988);
nor U13747 (N_13747,N_12285,N_12820);
nor U13748 (N_13748,N_12500,N_12295);
xor U13749 (N_13749,N_12936,N_12114);
nor U13750 (N_13750,N_12912,N_12544);
xor U13751 (N_13751,N_12189,N_12090);
xnor U13752 (N_13752,N_12560,N_13256);
xnor U13753 (N_13753,N_13462,N_13014);
xor U13754 (N_13754,N_13100,N_12765);
or U13755 (N_13755,N_13017,N_13107);
or U13756 (N_13756,N_13173,N_13087);
nor U13757 (N_13757,N_12682,N_12272);
nand U13758 (N_13758,N_12381,N_12156);
or U13759 (N_13759,N_12349,N_13265);
nand U13760 (N_13760,N_12055,N_12899);
or U13761 (N_13761,N_12181,N_13345);
nor U13762 (N_13762,N_13096,N_13060);
and U13763 (N_13763,N_12978,N_13277);
xor U13764 (N_13764,N_13223,N_13126);
nor U13765 (N_13765,N_13159,N_12350);
nor U13766 (N_13766,N_12121,N_12419);
and U13767 (N_13767,N_12177,N_12455);
xor U13768 (N_13768,N_13113,N_12724);
or U13769 (N_13769,N_13004,N_12095);
nand U13770 (N_13770,N_12808,N_12424);
nor U13771 (N_13771,N_12484,N_13079);
nand U13772 (N_13772,N_12160,N_12408);
nand U13773 (N_13773,N_13372,N_12263);
or U13774 (N_13774,N_12583,N_12742);
xor U13775 (N_13775,N_12525,N_12367);
and U13776 (N_13776,N_13390,N_13317);
nor U13777 (N_13777,N_13257,N_13300);
or U13778 (N_13778,N_13093,N_13325);
xnor U13779 (N_13779,N_13048,N_12718);
and U13780 (N_13780,N_12176,N_12412);
and U13781 (N_13781,N_12594,N_12661);
nor U13782 (N_13782,N_12920,N_12348);
nor U13783 (N_13783,N_12089,N_13340);
or U13784 (N_13784,N_12058,N_13124);
and U13785 (N_13785,N_13141,N_12825);
xor U13786 (N_13786,N_12288,N_12781);
and U13787 (N_13787,N_12108,N_13021);
or U13788 (N_13788,N_12676,N_13406);
and U13789 (N_13789,N_13399,N_12061);
and U13790 (N_13790,N_12993,N_13074);
nand U13791 (N_13791,N_13204,N_12997);
and U13792 (N_13792,N_13102,N_12049);
and U13793 (N_13793,N_12649,N_13266);
nor U13794 (N_13794,N_13358,N_13091);
or U13795 (N_13795,N_13465,N_13422);
and U13796 (N_13796,N_12529,N_13305);
or U13797 (N_13797,N_12516,N_12757);
xnor U13798 (N_13798,N_13170,N_12141);
xnor U13799 (N_13799,N_13038,N_12592);
nor U13800 (N_13800,N_12182,N_13245);
xor U13801 (N_13801,N_13145,N_13291);
nand U13802 (N_13802,N_12518,N_12960);
xor U13803 (N_13803,N_12986,N_13249);
or U13804 (N_13804,N_13495,N_13253);
xor U13805 (N_13805,N_12015,N_13036);
xnor U13806 (N_13806,N_12099,N_12238);
and U13807 (N_13807,N_12784,N_13104);
and U13808 (N_13808,N_12299,N_12989);
nor U13809 (N_13809,N_12398,N_12478);
and U13810 (N_13810,N_12162,N_12364);
nor U13811 (N_13811,N_12703,N_13099);
xor U13812 (N_13812,N_12507,N_12735);
and U13813 (N_13813,N_12292,N_12241);
nor U13814 (N_13814,N_12289,N_13442);
or U13815 (N_13815,N_13174,N_13478);
xnor U13816 (N_13816,N_12712,N_13331);
xnor U13817 (N_13817,N_12505,N_12064);
nor U13818 (N_13818,N_13007,N_12279);
or U13819 (N_13819,N_13072,N_12386);
xor U13820 (N_13820,N_12371,N_12038);
nor U13821 (N_13821,N_12752,N_12196);
or U13822 (N_13822,N_12308,N_12119);
nor U13823 (N_13823,N_13466,N_12235);
and U13824 (N_13824,N_12311,N_12554);
or U13825 (N_13825,N_13089,N_12938);
or U13826 (N_13826,N_12337,N_13189);
nor U13827 (N_13827,N_13150,N_12219);
xnor U13828 (N_13828,N_12513,N_12216);
nor U13829 (N_13829,N_12616,N_13321);
or U13830 (N_13830,N_12857,N_13054);
xnor U13831 (N_13831,N_12496,N_12242);
nand U13832 (N_13832,N_12093,N_12042);
nand U13833 (N_13833,N_12833,N_12654);
xnor U13834 (N_13834,N_12804,N_12023);
nor U13835 (N_13835,N_12863,N_12949);
xor U13836 (N_13836,N_12580,N_12471);
nand U13837 (N_13837,N_12428,N_13412);
nand U13838 (N_13838,N_12702,N_13133);
or U13839 (N_13839,N_12249,N_13252);
nand U13840 (N_13840,N_12928,N_13471);
or U13841 (N_13841,N_13123,N_12909);
nor U13842 (N_13842,N_12700,N_12489);
nand U13843 (N_13843,N_12185,N_13171);
nand U13844 (N_13844,N_12461,N_13334);
nand U13845 (N_13845,N_13062,N_12449);
xor U13846 (N_13846,N_12037,N_12667);
nand U13847 (N_13847,N_12538,N_13424);
xor U13848 (N_13848,N_12075,N_12414);
and U13849 (N_13849,N_13084,N_12598);
nand U13850 (N_13850,N_13128,N_13479);
or U13851 (N_13851,N_13446,N_12617);
xor U13852 (N_13852,N_12927,N_13131);
and U13853 (N_13853,N_12205,N_12953);
or U13854 (N_13854,N_13339,N_12974);
xnor U13855 (N_13855,N_12954,N_12338);
nor U13856 (N_13856,N_12467,N_12030);
or U13857 (N_13857,N_13398,N_12097);
nor U13858 (N_13858,N_13448,N_12004);
xnor U13859 (N_13859,N_13404,N_12665);
nor U13860 (N_13860,N_12470,N_12585);
or U13861 (N_13861,N_12895,N_12204);
nand U13862 (N_13862,N_12378,N_13005);
nor U13863 (N_13863,N_12764,N_13168);
nor U13864 (N_13864,N_13432,N_13112);
and U13865 (N_13865,N_12726,N_12252);
or U13866 (N_13866,N_12747,N_12842);
nand U13867 (N_13867,N_12278,N_12769);
nand U13868 (N_13868,N_13299,N_12610);
nand U13869 (N_13869,N_12302,N_12853);
nand U13870 (N_13870,N_12445,N_13364);
or U13871 (N_13871,N_13026,N_12618);
nand U13872 (N_13872,N_13304,N_12231);
xnor U13873 (N_13873,N_12855,N_13044);
or U13874 (N_13874,N_12626,N_12591);
and U13875 (N_13875,N_13453,N_13139);
nor U13876 (N_13876,N_12878,N_12170);
xnor U13877 (N_13877,N_12225,N_12621);
nor U13878 (N_13878,N_12984,N_12164);
nand U13879 (N_13879,N_12791,N_12091);
xnor U13880 (N_13880,N_12506,N_13483);
nand U13881 (N_13881,N_13499,N_13436);
xor U13882 (N_13882,N_12575,N_13387);
nand U13883 (N_13883,N_12152,N_13338);
nor U13884 (N_13884,N_12964,N_12143);
nor U13885 (N_13885,N_12054,N_12326);
and U13886 (N_13886,N_12245,N_13274);
xnor U13887 (N_13887,N_12158,N_13476);
or U13888 (N_13888,N_12179,N_12541);
and U13889 (N_13889,N_13135,N_13134);
nor U13890 (N_13890,N_13034,N_13181);
nand U13891 (N_13891,N_13492,N_12658);
nand U13892 (N_13892,N_12951,N_12934);
xor U13893 (N_13893,N_12869,N_12982);
nand U13894 (N_13894,N_12859,N_12102);
nand U13895 (N_13895,N_12407,N_13315);
nor U13896 (N_13896,N_12486,N_12733);
and U13897 (N_13897,N_13258,N_12309);
xnor U13898 (N_13898,N_12031,N_12730);
xor U13899 (N_13899,N_12233,N_12366);
or U13900 (N_13900,N_13247,N_12146);
xnor U13901 (N_13901,N_12732,N_12612);
nand U13902 (N_13902,N_12374,N_13129);
xnor U13903 (N_13903,N_12795,N_12426);
nand U13904 (N_13904,N_12191,N_12133);
or U13905 (N_13905,N_12014,N_13237);
or U13906 (N_13906,N_12203,N_13347);
nor U13907 (N_13907,N_12536,N_12973);
xor U13908 (N_13908,N_12234,N_12138);
xor U13909 (N_13909,N_13092,N_12836);
or U13910 (N_13910,N_12330,N_13244);
or U13911 (N_13911,N_13363,N_12889);
and U13912 (N_13912,N_12762,N_12258);
nand U13913 (N_13913,N_12609,N_13066);
and U13914 (N_13914,N_12466,N_12257);
xor U13915 (N_13915,N_12543,N_13489);
xnor U13916 (N_13916,N_12498,N_13282);
nand U13917 (N_13917,N_12570,N_12494);
nor U13918 (N_13918,N_13421,N_12867);
nor U13919 (N_13919,N_13106,N_12452);
or U13920 (N_13920,N_12971,N_13360);
or U13921 (N_13921,N_13242,N_13308);
nand U13922 (N_13922,N_13330,N_12082);
nor U13923 (N_13923,N_12826,N_13286);
or U13924 (N_13924,N_13231,N_12910);
nor U13925 (N_13925,N_12315,N_13459);
nand U13926 (N_13926,N_13001,N_12041);
xnor U13927 (N_13927,N_12956,N_12178);
xor U13928 (N_13928,N_12406,N_13023);
or U13929 (N_13929,N_13059,N_12069);
nand U13930 (N_13930,N_13157,N_13143);
or U13931 (N_13931,N_12022,N_12727);
nor U13932 (N_13932,N_12753,N_12741);
nor U13933 (N_13933,N_13426,N_12962);
and U13934 (N_13934,N_12397,N_13433);
and U13935 (N_13935,N_13454,N_12433);
nor U13936 (N_13936,N_13368,N_12006);
xnor U13937 (N_13937,N_13410,N_12625);
and U13938 (N_13938,N_13263,N_12891);
xor U13939 (N_13939,N_12324,N_12389);
nand U13940 (N_13940,N_13090,N_12462);
nor U13941 (N_13941,N_13187,N_12646);
nand U13942 (N_13942,N_13163,N_12416);
nand U13943 (N_13943,N_13301,N_13343);
or U13944 (N_13944,N_12437,N_13030);
and U13945 (N_13945,N_12824,N_12045);
nand U13946 (N_13946,N_13160,N_12144);
and U13947 (N_13947,N_12866,N_12587);
nor U13948 (N_13948,N_13393,N_12698);
nor U13949 (N_13949,N_13362,N_12699);
or U13950 (N_13950,N_12624,N_12713);
and U13951 (N_13951,N_12453,N_12883);
or U13952 (N_13952,N_12088,N_13053);
nor U13953 (N_13953,N_12057,N_13278);
or U13954 (N_13954,N_12636,N_12666);
nor U13955 (N_13955,N_12056,N_12659);
nor U13956 (N_13956,N_13200,N_12746);
and U13957 (N_13957,N_12987,N_12222);
xor U13958 (N_13958,N_12443,N_12282);
nand U13959 (N_13959,N_12567,N_12872);
or U13960 (N_13960,N_13320,N_13294);
xnor U13961 (N_13961,N_13303,N_12611);
nand U13962 (N_13962,N_12711,N_12493);
and U13963 (N_13963,N_13228,N_12985);
xnor U13964 (N_13964,N_13033,N_12287);
and U13965 (N_13965,N_12508,N_12376);
or U13966 (N_13966,N_12362,N_12728);
nand U13967 (N_13967,N_12800,N_12425);
nor U13968 (N_13968,N_12314,N_12469);
nor U13969 (N_13969,N_12725,N_13071);
and U13970 (N_13970,N_12370,N_13241);
xnor U13971 (N_13971,N_12680,N_12816);
or U13972 (N_13972,N_13261,N_12104);
xor U13973 (N_13973,N_12307,N_12334);
and U13974 (N_13974,N_12963,N_12265);
nor U13975 (N_13975,N_12817,N_12465);
nor U13976 (N_13976,N_12171,N_12188);
nor U13977 (N_13977,N_13405,N_12401);
and U13978 (N_13978,N_13164,N_12704);
nor U13979 (N_13979,N_13329,N_13430);
nor U13980 (N_13980,N_12797,N_13015);
and U13981 (N_13981,N_13178,N_12390);
or U13982 (N_13982,N_12686,N_13086);
and U13983 (N_13983,N_12677,N_13049);
nand U13984 (N_13984,N_13193,N_12923);
nand U13985 (N_13985,N_13369,N_13367);
xor U13986 (N_13986,N_13475,N_12777);
nor U13987 (N_13987,N_13437,N_12614);
or U13988 (N_13988,N_12555,N_12662);
or U13989 (N_13989,N_12622,N_12322);
nor U13990 (N_13990,N_12002,N_12081);
and U13991 (N_13991,N_13394,N_12709);
or U13992 (N_13992,N_12879,N_12363);
xnor U13993 (N_13993,N_12967,N_12785);
nor U13994 (N_13994,N_12151,N_12076);
or U13995 (N_13995,N_12388,N_12551);
xor U13996 (N_13996,N_12184,N_13152);
nand U13997 (N_13997,N_12439,N_12586);
nor U13998 (N_13998,N_12803,N_12501);
xnor U13999 (N_13999,N_12360,N_12281);
or U14000 (N_14000,N_12124,N_12154);
nor U14001 (N_14001,N_12078,N_13493);
nand U14002 (N_14002,N_12372,N_12688);
xnor U14003 (N_14003,N_12576,N_13207);
nor U14004 (N_14004,N_13013,N_13010);
or U14005 (N_14005,N_12990,N_13075);
nand U14006 (N_14006,N_12821,N_12786);
or U14007 (N_14007,N_12444,N_12488);
nand U14008 (N_14008,N_13383,N_12685);
xor U14009 (N_14009,N_12706,N_12251);
xor U14010 (N_14010,N_12094,N_12110);
nand U14011 (N_14011,N_13032,N_13220);
and U14012 (N_14012,N_12244,N_12675);
or U14013 (N_14013,N_12606,N_12782);
xor U14014 (N_14014,N_12427,N_12264);
or U14015 (N_14015,N_12357,N_13456);
or U14016 (N_14016,N_12597,N_12652);
nand U14017 (N_14017,N_13425,N_13260);
and U14018 (N_14018,N_13065,N_13095);
nor U14019 (N_14019,N_13306,N_13088);
or U14020 (N_14020,N_13239,N_12113);
nor U14021 (N_14021,N_12066,N_12559);
or U14022 (N_14022,N_12603,N_12903);
or U14023 (N_14023,N_12577,N_13043);
xor U14024 (N_14024,N_13050,N_13273);
or U14025 (N_14025,N_13035,N_12906);
or U14026 (N_14026,N_12210,N_12227);
and U14027 (N_14027,N_13268,N_12394);
nand U14028 (N_14028,N_12840,N_12681);
or U14029 (N_14029,N_12926,N_12874);
nor U14030 (N_14030,N_12778,N_13288);
xnor U14031 (N_14031,N_13461,N_12019);
or U14032 (N_14032,N_12355,N_13349);
or U14033 (N_14033,N_13165,N_12601);
xor U14034 (N_14034,N_13233,N_12111);
xor U14035 (N_14035,N_12187,N_12228);
or U14036 (N_14036,N_13498,N_13496);
xnor U14037 (N_14037,N_12132,N_12707);
nor U14038 (N_14038,N_12310,N_12515);
or U14039 (N_14039,N_12561,N_12186);
nand U14040 (N_14040,N_12085,N_12981);
or U14041 (N_14041,N_12380,N_13055);
nor U14042 (N_14042,N_12783,N_12074);
nor U14043 (N_14043,N_13022,N_12619);
nor U14044 (N_14044,N_12848,N_13234);
and U14045 (N_14045,N_12458,N_13378);
or U14046 (N_14046,N_12487,N_13380);
xnor U14047 (N_14047,N_12136,N_12018);
nand U14048 (N_14048,N_12441,N_12422);
nand U14049 (N_14049,N_12766,N_12230);
xor U14050 (N_14050,N_12291,N_12165);
xor U14051 (N_14051,N_12400,N_13077);
and U14052 (N_14052,N_13154,N_12892);
nor U14053 (N_14053,N_12572,N_12497);
or U14054 (N_14054,N_12530,N_12627);
or U14055 (N_14055,N_12519,N_12860);
or U14056 (N_14056,N_12819,N_12320);
nand U14057 (N_14057,N_13284,N_13224);
and U14058 (N_14058,N_13401,N_13137);
xor U14059 (N_14059,N_12696,N_13177);
nor U14060 (N_14060,N_12431,N_12340);
and U14061 (N_14061,N_12527,N_12502);
nand U14062 (N_14062,N_12756,N_12629);
xor U14063 (N_14063,N_12237,N_13354);
xor U14064 (N_14064,N_12552,N_12358);
and U14065 (N_14065,N_12296,N_12884);
nor U14066 (N_14066,N_13226,N_12648);
xnor U14067 (N_14067,N_12827,N_13314);
or U14068 (N_14068,N_13175,N_12000);
nand U14069 (N_14069,N_12255,N_12885);
and U14070 (N_14070,N_12887,N_13151);
or U14071 (N_14071,N_12862,N_13332);
and U14072 (N_14072,N_12921,N_12169);
or U14073 (N_14073,N_12931,N_12328);
xnor U14074 (N_14074,N_12480,N_12040);
nand U14075 (N_14075,N_12980,N_12262);
xnor U14076 (N_14076,N_12776,N_13416);
nand U14077 (N_14077,N_12943,N_12770);
xnor U14078 (N_14078,N_12995,N_13281);
nand U14079 (N_14079,N_12180,N_12092);
and U14080 (N_14080,N_12798,N_12890);
and U14081 (N_14081,N_12897,N_12135);
nor U14082 (N_14082,N_13094,N_12399);
and U14083 (N_14083,N_12208,N_12893);
nor U14084 (N_14084,N_13337,N_12490);
nand U14085 (N_14085,N_12535,N_12861);
nor U14086 (N_14086,N_13037,N_12992);
nor U14087 (N_14087,N_12239,N_12557);
nand U14088 (N_14088,N_13460,N_12873);
nand U14089 (N_14089,N_12269,N_13212);
nand U14090 (N_14090,N_12472,N_13322);
nand U14091 (N_14091,N_12615,N_12411);
nand U14092 (N_14092,N_12710,N_12130);
nor U14093 (N_14093,N_12558,N_12534);
or U14094 (N_14094,N_13350,N_12852);
or U14095 (N_14095,N_12335,N_12253);
and U14096 (N_14096,N_12721,N_12325);
nand U14097 (N_14097,N_13081,N_12275);
xnor U14098 (N_14098,N_12952,N_13384);
nor U14099 (N_14099,N_13409,N_13185);
nand U14100 (N_14100,N_12477,N_12157);
and U14101 (N_14101,N_13379,N_12247);
xnor U14102 (N_14102,N_12633,N_13118);
or U14103 (N_14103,N_13419,N_12448);
xnor U14104 (N_14104,N_12991,N_12027);
or U14105 (N_14105,N_12159,N_13208);
nor U14106 (N_14106,N_12035,N_13188);
or U14107 (N_14107,N_13057,N_12344);
nand U14108 (N_14108,N_12197,N_12771);
nand U14109 (N_14109,N_12212,N_13229);
or U14110 (N_14110,N_12174,N_12321);
nand U14111 (N_14111,N_13012,N_12303);
nand U14112 (N_14112,N_12671,N_12250);
or U14113 (N_14113,N_12474,N_13386);
or U14114 (N_14114,N_12473,N_12608);
nand U14115 (N_14115,N_12052,N_12070);
xor U14116 (N_14116,N_12922,N_13031);
and U14117 (N_14117,N_13215,N_12568);
xor U14118 (N_14118,N_13169,N_12306);
xnor U14119 (N_14119,N_13464,N_12173);
and U14120 (N_14120,N_12342,N_12051);
nand U14121 (N_14121,N_13068,N_13474);
and U14122 (N_14122,N_13085,N_13381);
nand U14123 (N_14123,N_13028,N_12830);
xor U14124 (N_14124,N_12745,N_12195);
or U14125 (N_14125,N_12118,N_12854);
or U14126 (N_14126,N_12913,N_12545);
nor U14127 (N_14127,N_13326,N_13097);
nand U14128 (N_14128,N_12613,N_12149);
and U14129 (N_14129,N_12261,N_12382);
or U14130 (N_14130,N_13122,N_12248);
and U14131 (N_14131,N_12485,N_12122);
xor U14132 (N_14132,N_12723,N_12353);
nand U14133 (N_14133,N_12794,N_13191);
xnor U14134 (N_14134,N_12327,N_13156);
and U14135 (N_14135,N_13117,N_12907);
nor U14136 (N_14136,N_12087,N_12226);
or U14137 (N_14137,N_13312,N_12021);
xor U14138 (N_14138,N_12828,N_12740);
nand U14139 (N_14139,N_12438,N_12011);
and U14140 (N_14140,N_12273,N_12409);
or U14141 (N_14141,N_12268,N_12957);
and U14142 (N_14142,N_12902,N_12939);
nand U14143 (N_14143,N_12969,N_13250);
or U14144 (N_14144,N_12845,N_12918);
nor U14145 (N_14145,N_13365,N_13370);
and U14146 (N_14146,N_13246,N_12148);
nand U14147 (N_14147,N_12294,N_12005);
and U14148 (N_14148,N_12692,N_12168);
and U14149 (N_14149,N_12581,N_13373);
nand U14150 (N_14150,N_13082,N_13280);
or U14151 (N_14151,N_12849,N_12423);
nand U14152 (N_14152,N_12243,N_13217);
nor U14153 (N_14153,N_13148,N_12277);
xnor U14154 (N_14154,N_12693,N_12651);
and U14155 (N_14155,N_13450,N_13389);
nand U14156 (N_14156,N_12634,N_12950);
nor U14157 (N_14157,N_12937,N_12569);
and U14158 (N_14158,N_12628,N_12864);
nand U14159 (N_14159,N_12194,N_12172);
nand U14160 (N_14160,N_12779,N_13289);
xor U14161 (N_14161,N_13452,N_13423);
and U14162 (N_14162,N_12385,N_12780);
nand U14163 (N_14163,N_12175,N_12491);
or U14164 (N_14164,N_13183,N_13194);
or U14165 (N_14165,N_12067,N_12526);
or U14166 (N_14166,N_12403,N_13473);
nand U14167 (N_14167,N_12877,N_13144);
and U14168 (N_14168,N_12942,N_12003);
and U14169 (N_14169,N_12336,N_12024);
nand U14170 (N_14170,N_13458,N_13400);
and U14171 (N_14171,N_13216,N_12968);
and U14172 (N_14172,N_12941,N_12958);
nand U14173 (N_14173,N_12772,N_12975);
nand U14174 (N_14174,N_12623,N_13319);
nand U14175 (N_14175,N_13111,N_12947);
nand U14176 (N_14176,N_13179,N_13374);
xor U14177 (N_14177,N_12768,N_12240);
and U14178 (N_14178,N_12898,N_12053);
xor U14179 (N_14179,N_13468,N_12260);
xor U14180 (N_14180,N_12166,N_12679);
nand U14181 (N_14181,N_13353,N_12908);
and U14182 (N_14182,N_12748,N_13351);
and U14183 (N_14183,N_12483,N_12116);
or U14184 (N_14184,N_12810,N_12447);
xor U14185 (N_14185,N_12998,N_13271);
or U14186 (N_14186,N_12280,N_13192);
and U14187 (N_14187,N_13136,N_12743);
and U14188 (N_14188,N_12012,N_12153);
or U14189 (N_14189,N_12850,N_12856);
and U14190 (N_14190,N_13101,N_12972);
nor U14191 (N_14191,N_13083,N_12805);
xor U14192 (N_14192,N_13451,N_12775);
and U14193 (N_14193,N_12440,N_12789);
nand U14194 (N_14194,N_13439,N_12451);
and U14195 (N_14195,N_12715,N_12653);
xor U14196 (N_14196,N_12917,N_13396);
and U14197 (N_14197,N_13211,N_12318);
nor U14198 (N_14198,N_12039,N_13336);
nand U14199 (N_14199,N_13429,N_13214);
xnor U14200 (N_14200,N_13180,N_12708);
or U14201 (N_14201,N_12811,N_13119);
and U14202 (N_14202,N_12641,N_12059);
nor U14203 (N_14203,N_12714,N_12520);
nand U14204 (N_14204,N_12460,N_12086);
and U14205 (N_14205,N_13219,N_12442);
and U14206 (N_14206,N_12293,N_12566);
nor U14207 (N_14207,N_12875,N_12048);
or U14208 (N_14208,N_13069,N_13238);
nand U14209 (N_14209,N_12028,N_12829);
and U14210 (N_14210,N_12935,N_12847);
nor U14211 (N_14211,N_12463,N_12434);
xnor U14212 (N_14212,N_12663,N_12267);
nand U14213 (N_14213,N_12317,N_12436);
xnor U14214 (N_14214,N_12117,N_12457);
or U14215 (N_14215,N_13058,N_12524);
nand U14216 (N_14216,N_13297,N_13359);
xnor U14217 (N_14217,N_12584,N_12103);
nor U14218 (N_14218,N_13140,N_13255);
or U14219 (N_14219,N_12571,N_13051);
nand U14220 (N_14220,N_12509,N_12605);
and U14221 (N_14221,N_12393,N_12105);
or U14222 (N_14222,N_13467,N_12593);
and U14223 (N_14223,N_12392,N_12638);
and U14224 (N_14224,N_12578,N_12701);
xor U14225 (N_14225,N_12468,N_13395);
nor U14226 (N_14226,N_12079,N_13290);
and U14227 (N_14227,N_12479,N_13002);
nor U14228 (N_14228,N_12010,N_12523);
xnor U14229 (N_14229,N_13190,N_12871);
and U14230 (N_14230,N_12739,N_12065);
and U14231 (N_14231,N_12352,N_13275);
or U14232 (N_14232,N_12843,N_13236);
and U14233 (N_14233,N_13039,N_12589);
xor U14234 (N_14234,N_13431,N_12333);
nand U14235 (N_14235,N_12131,N_12806);
nand U14236 (N_14236,N_12271,N_13064);
nand U14237 (N_14237,N_13408,N_12894);
nand U14238 (N_14238,N_12026,N_12565);
and U14239 (N_14239,N_12925,N_12602);
xor U14240 (N_14240,N_12683,N_12379);
nand U14241 (N_14241,N_12346,N_12139);
xor U14242 (N_14242,N_12100,N_13481);
or U14243 (N_14243,N_12009,N_12737);
nand U14244 (N_14244,N_12579,N_13110);
nand U14245 (N_14245,N_12098,N_12734);
nor U14246 (N_14246,N_12574,N_12822);
xor U14247 (N_14247,N_12517,N_12206);
and U14248 (N_14248,N_12736,N_12933);
nor U14249 (N_14249,N_12846,N_12147);
nand U14250 (N_14250,N_12224,N_12165);
nand U14251 (N_14251,N_12208,N_12394);
nor U14252 (N_14252,N_13224,N_13058);
nor U14253 (N_14253,N_13437,N_12094);
xnor U14254 (N_14254,N_13182,N_13194);
nand U14255 (N_14255,N_12961,N_12198);
or U14256 (N_14256,N_12632,N_12845);
and U14257 (N_14257,N_12360,N_13049);
or U14258 (N_14258,N_12729,N_12514);
xnor U14259 (N_14259,N_12884,N_12478);
or U14260 (N_14260,N_12460,N_12100);
or U14261 (N_14261,N_12309,N_13452);
or U14262 (N_14262,N_12893,N_12539);
xor U14263 (N_14263,N_12297,N_12820);
and U14264 (N_14264,N_12035,N_12289);
xor U14265 (N_14265,N_12016,N_12612);
nor U14266 (N_14266,N_13144,N_12985);
and U14267 (N_14267,N_12012,N_13235);
xor U14268 (N_14268,N_12401,N_12963);
nand U14269 (N_14269,N_12420,N_12355);
nor U14270 (N_14270,N_12331,N_12725);
nor U14271 (N_14271,N_12448,N_13493);
nor U14272 (N_14272,N_13152,N_12802);
xor U14273 (N_14273,N_13117,N_13187);
nor U14274 (N_14274,N_13141,N_12747);
nand U14275 (N_14275,N_12370,N_12784);
or U14276 (N_14276,N_13179,N_13255);
xnor U14277 (N_14277,N_12279,N_12659);
nand U14278 (N_14278,N_12858,N_13174);
xnor U14279 (N_14279,N_13360,N_13381);
xor U14280 (N_14280,N_12977,N_12933);
xor U14281 (N_14281,N_12951,N_13300);
or U14282 (N_14282,N_12058,N_13444);
nand U14283 (N_14283,N_12484,N_13135);
xor U14284 (N_14284,N_13163,N_12871);
xor U14285 (N_14285,N_13141,N_12314);
nor U14286 (N_14286,N_12562,N_13115);
xor U14287 (N_14287,N_12862,N_12296);
nor U14288 (N_14288,N_13449,N_13470);
and U14289 (N_14289,N_12175,N_12085);
nand U14290 (N_14290,N_12952,N_12283);
nor U14291 (N_14291,N_12519,N_12807);
and U14292 (N_14292,N_12386,N_12099);
nand U14293 (N_14293,N_12572,N_12564);
nor U14294 (N_14294,N_13273,N_12256);
nand U14295 (N_14295,N_13492,N_13225);
and U14296 (N_14296,N_13091,N_13328);
or U14297 (N_14297,N_13475,N_12436);
and U14298 (N_14298,N_12094,N_12350);
or U14299 (N_14299,N_13356,N_13107);
nand U14300 (N_14300,N_13475,N_13207);
or U14301 (N_14301,N_13265,N_12363);
and U14302 (N_14302,N_12997,N_13271);
xor U14303 (N_14303,N_12745,N_12512);
nor U14304 (N_14304,N_13302,N_12766);
and U14305 (N_14305,N_13331,N_13193);
nor U14306 (N_14306,N_12410,N_13084);
nand U14307 (N_14307,N_13141,N_13288);
or U14308 (N_14308,N_12202,N_12698);
xor U14309 (N_14309,N_12067,N_13299);
xor U14310 (N_14310,N_12031,N_12588);
xor U14311 (N_14311,N_13397,N_13040);
xnor U14312 (N_14312,N_12853,N_12115);
nand U14313 (N_14313,N_12838,N_12210);
or U14314 (N_14314,N_13260,N_12203);
or U14315 (N_14315,N_13150,N_12747);
or U14316 (N_14316,N_13306,N_12511);
or U14317 (N_14317,N_12719,N_12864);
and U14318 (N_14318,N_12702,N_12477);
nor U14319 (N_14319,N_12179,N_13232);
nor U14320 (N_14320,N_13413,N_13024);
nand U14321 (N_14321,N_13398,N_12337);
or U14322 (N_14322,N_12255,N_13308);
and U14323 (N_14323,N_12200,N_12698);
and U14324 (N_14324,N_12960,N_12847);
xor U14325 (N_14325,N_13094,N_12575);
and U14326 (N_14326,N_12902,N_13242);
nand U14327 (N_14327,N_12509,N_13220);
or U14328 (N_14328,N_12147,N_13198);
and U14329 (N_14329,N_12636,N_13488);
or U14330 (N_14330,N_12534,N_12628);
nand U14331 (N_14331,N_12509,N_12526);
and U14332 (N_14332,N_12243,N_12233);
nor U14333 (N_14333,N_12309,N_13103);
xor U14334 (N_14334,N_12140,N_13485);
xnor U14335 (N_14335,N_13027,N_12057);
xor U14336 (N_14336,N_12555,N_13387);
nand U14337 (N_14337,N_12471,N_12260);
xnor U14338 (N_14338,N_12676,N_12703);
xnor U14339 (N_14339,N_13116,N_12484);
xnor U14340 (N_14340,N_12581,N_12686);
nor U14341 (N_14341,N_13394,N_13262);
or U14342 (N_14342,N_13202,N_12843);
nand U14343 (N_14343,N_12540,N_12902);
nor U14344 (N_14344,N_12820,N_13401);
nand U14345 (N_14345,N_12310,N_13415);
and U14346 (N_14346,N_13188,N_12561);
nand U14347 (N_14347,N_12449,N_12620);
nand U14348 (N_14348,N_13419,N_12498);
and U14349 (N_14349,N_13473,N_13067);
xor U14350 (N_14350,N_12845,N_13302);
or U14351 (N_14351,N_12063,N_12906);
xor U14352 (N_14352,N_12527,N_12667);
xnor U14353 (N_14353,N_12064,N_12489);
nand U14354 (N_14354,N_12061,N_12088);
nor U14355 (N_14355,N_13332,N_12316);
or U14356 (N_14356,N_12634,N_12338);
xor U14357 (N_14357,N_12589,N_12375);
and U14358 (N_14358,N_12372,N_12202);
or U14359 (N_14359,N_13340,N_12302);
xor U14360 (N_14360,N_13482,N_13056);
nor U14361 (N_14361,N_12005,N_13103);
xor U14362 (N_14362,N_13267,N_12492);
nor U14363 (N_14363,N_12395,N_13444);
xor U14364 (N_14364,N_12051,N_13127);
xor U14365 (N_14365,N_12033,N_12445);
nand U14366 (N_14366,N_12986,N_13387);
or U14367 (N_14367,N_12610,N_13079);
or U14368 (N_14368,N_12385,N_12972);
nor U14369 (N_14369,N_12757,N_13485);
nor U14370 (N_14370,N_12379,N_12933);
xor U14371 (N_14371,N_12663,N_12550);
nand U14372 (N_14372,N_12168,N_12695);
xnor U14373 (N_14373,N_12430,N_12493);
xor U14374 (N_14374,N_13349,N_12509);
or U14375 (N_14375,N_12496,N_12823);
xnor U14376 (N_14376,N_13352,N_13153);
or U14377 (N_14377,N_12215,N_12947);
nand U14378 (N_14378,N_12488,N_12738);
and U14379 (N_14379,N_12526,N_12241);
nor U14380 (N_14380,N_12483,N_12178);
nand U14381 (N_14381,N_13222,N_12691);
and U14382 (N_14382,N_13065,N_12761);
nor U14383 (N_14383,N_12679,N_12379);
nor U14384 (N_14384,N_12285,N_12303);
and U14385 (N_14385,N_12437,N_13006);
xor U14386 (N_14386,N_12994,N_12508);
or U14387 (N_14387,N_12468,N_13388);
and U14388 (N_14388,N_12148,N_12904);
or U14389 (N_14389,N_12205,N_12950);
xnor U14390 (N_14390,N_12970,N_13216);
and U14391 (N_14391,N_13043,N_13046);
xnor U14392 (N_14392,N_12821,N_12569);
and U14393 (N_14393,N_12705,N_13203);
xnor U14394 (N_14394,N_12122,N_13443);
nor U14395 (N_14395,N_12371,N_12753);
xor U14396 (N_14396,N_12854,N_13297);
xor U14397 (N_14397,N_12992,N_13181);
and U14398 (N_14398,N_12913,N_13067);
and U14399 (N_14399,N_12723,N_13475);
or U14400 (N_14400,N_12924,N_13206);
xnor U14401 (N_14401,N_12097,N_13243);
nand U14402 (N_14402,N_13489,N_13199);
xnor U14403 (N_14403,N_13287,N_13404);
nor U14404 (N_14404,N_12994,N_12440);
or U14405 (N_14405,N_12715,N_12646);
or U14406 (N_14406,N_12897,N_12779);
and U14407 (N_14407,N_13267,N_13185);
nand U14408 (N_14408,N_13026,N_13483);
nand U14409 (N_14409,N_12584,N_13293);
nor U14410 (N_14410,N_13306,N_12868);
and U14411 (N_14411,N_12504,N_13065);
xor U14412 (N_14412,N_12686,N_12217);
nor U14413 (N_14413,N_12449,N_12477);
nor U14414 (N_14414,N_12870,N_13033);
and U14415 (N_14415,N_13179,N_13351);
nor U14416 (N_14416,N_12140,N_12660);
nor U14417 (N_14417,N_12694,N_13055);
or U14418 (N_14418,N_12036,N_12583);
or U14419 (N_14419,N_13097,N_13029);
or U14420 (N_14420,N_13179,N_13283);
or U14421 (N_14421,N_12964,N_13275);
nand U14422 (N_14422,N_12974,N_12527);
or U14423 (N_14423,N_12626,N_13460);
xnor U14424 (N_14424,N_13020,N_13012);
or U14425 (N_14425,N_12031,N_12148);
or U14426 (N_14426,N_12176,N_12609);
or U14427 (N_14427,N_12041,N_13174);
and U14428 (N_14428,N_13078,N_13441);
nor U14429 (N_14429,N_13077,N_13432);
and U14430 (N_14430,N_12668,N_12957);
or U14431 (N_14431,N_12518,N_12474);
nor U14432 (N_14432,N_12540,N_13139);
nor U14433 (N_14433,N_13169,N_13427);
nor U14434 (N_14434,N_12133,N_12811);
and U14435 (N_14435,N_13334,N_12913);
and U14436 (N_14436,N_12499,N_12349);
or U14437 (N_14437,N_12627,N_12135);
and U14438 (N_14438,N_12375,N_12681);
nand U14439 (N_14439,N_12332,N_12634);
or U14440 (N_14440,N_12832,N_13076);
and U14441 (N_14441,N_12034,N_12000);
xor U14442 (N_14442,N_13429,N_13167);
and U14443 (N_14443,N_12623,N_13404);
and U14444 (N_14444,N_13420,N_12029);
nor U14445 (N_14445,N_12300,N_12601);
xnor U14446 (N_14446,N_12913,N_12112);
nor U14447 (N_14447,N_12161,N_12241);
or U14448 (N_14448,N_13494,N_12574);
nand U14449 (N_14449,N_13215,N_13104);
xor U14450 (N_14450,N_13092,N_12340);
and U14451 (N_14451,N_13124,N_12865);
nand U14452 (N_14452,N_12114,N_12518);
xnor U14453 (N_14453,N_12801,N_13141);
and U14454 (N_14454,N_12652,N_13125);
nor U14455 (N_14455,N_12782,N_13198);
nand U14456 (N_14456,N_13349,N_12889);
and U14457 (N_14457,N_12464,N_12915);
and U14458 (N_14458,N_13310,N_13449);
xor U14459 (N_14459,N_13149,N_12875);
or U14460 (N_14460,N_12806,N_13451);
xnor U14461 (N_14461,N_12437,N_12856);
nand U14462 (N_14462,N_12091,N_12534);
and U14463 (N_14463,N_12809,N_12698);
or U14464 (N_14464,N_12325,N_12104);
nand U14465 (N_14465,N_12691,N_12366);
nor U14466 (N_14466,N_12930,N_13335);
nor U14467 (N_14467,N_12668,N_12976);
nor U14468 (N_14468,N_12145,N_13059);
or U14469 (N_14469,N_12565,N_13220);
or U14470 (N_14470,N_12396,N_13093);
or U14471 (N_14471,N_13159,N_12043);
and U14472 (N_14472,N_12185,N_12444);
and U14473 (N_14473,N_12076,N_12149);
nor U14474 (N_14474,N_12681,N_13037);
xor U14475 (N_14475,N_13068,N_13418);
xor U14476 (N_14476,N_13199,N_12303);
and U14477 (N_14477,N_12849,N_12939);
and U14478 (N_14478,N_12262,N_13297);
or U14479 (N_14479,N_13474,N_12833);
nand U14480 (N_14480,N_12410,N_12999);
or U14481 (N_14481,N_13284,N_12404);
nor U14482 (N_14482,N_12852,N_12776);
xnor U14483 (N_14483,N_13086,N_12544);
nand U14484 (N_14484,N_12575,N_13223);
or U14485 (N_14485,N_12329,N_12485);
nand U14486 (N_14486,N_12923,N_12410);
xor U14487 (N_14487,N_12963,N_13410);
nor U14488 (N_14488,N_13360,N_12967);
nand U14489 (N_14489,N_13493,N_12450);
and U14490 (N_14490,N_12547,N_13291);
xor U14491 (N_14491,N_12541,N_12066);
or U14492 (N_14492,N_13411,N_13000);
nand U14493 (N_14493,N_12531,N_12215);
xor U14494 (N_14494,N_13053,N_13414);
xnor U14495 (N_14495,N_12549,N_13136);
nor U14496 (N_14496,N_12891,N_13347);
and U14497 (N_14497,N_12705,N_13177);
xnor U14498 (N_14498,N_12279,N_12466);
nor U14499 (N_14499,N_13437,N_13383);
or U14500 (N_14500,N_12321,N_13301);
nor U14501 (N_14501,N_13157,N_13350);
nand U14502 (N_14502,N_12268,N_12395);
xnor U14503 (N_14503,N_12812,N_12349);
nand U14504 (N_14504,N_12469,N_13153);
and U14505 (N_14505,N_12529,N_12253);
or U14506 (N_14506,N_12245,N_12638);
or U14507 (N_14507,N_13008,N_12618);
xor U14508 (N_14508,N_12691,N_13329);
or U14509 (N_14509,N_13098,N_13356);
or U14510 (N_14510,N_12033,N_12563);
nand U14511 (N_14511,N_12656,N_13144);
nor U14512 (N_14512,N_12884,N_13317);
and U14513 (N_14513,N_12566,N_12130);
nor U14514 (N_14514,N_12518,N_12418);
nand U14515 (N_14515,N_13396,N_12445);
xor U14516 (N_14516,N_13139,N_12754);
or U14517 (N_14517,N_12000,N_12311);
or U14518 (N_14518,N_13130,N_13480);
or U14519 (N_14519,N_12590,N_12971);
nand U14520 (N_14520,N_12616,N_12590);
and U14521 (N_14521,N_12360,N_12645);
xor U14522 (N_14522,N_12681,N_12760);
xor U14523 (N_14523,N_12510,N_13025);
nor U14524 (N_14524,N_12120,N_12458);
nor U14525 (N_14525,N_12620,N_12454);
and U14526 (N_14526,N_12174,N_13315);
xor U14527 (N_14527,N_13306,N_12326);
nor U14528 (N_14528,N_12888,N_12087);
or U14529 (N_14529,N_12891,N_12442);
nand U14530 (N_14530,N_13266,N_12613);
xnor U14531 (N_14531,N_12001,N_12803);
nand U14532 (N_14532,N_12879,N_12826);
nor U14533 (N_14533,N_13350,N_13136);
nor U14534 (N_14534,N_12439,N_12324);
xor U14535 (N_14535,N_12350,N_12972);
or U14536 (N_14536,N_12667,N_13305);
xnor U14537 (N_14537,N_12075,N_12591);
or U14538 (N_14538,N_13086,N_12216);
nor U14539 (N_14539,N_13131,N_12517);
xnor U14540 (N_14540,N_12578,N_13486);
or U14541 (N_14541,N_13341,N_13198);
xnor U14542 (N_14542,N_12729,N_13372);
xor U14543 (N_14543,N_13046,N_13260);
and U14544 (N_14544,N_12081,N_12350);
xor U14545 (N_14545,N_12813,N_12667);
xor U14546 (N_14546,N_13294,N_12815);
nor U14547 (N_14547,N_12646,N_12931);
and U14548 (N_14548,N_13137,N_12515);
and U14549 (N_14549,N_12607,N_12594);
nand U14550 (N_14550,N_13427,N_12027);
nor U14551 (N_14551,N_12183,N_13364);
and U14552 (N_14552,N_13150,N_13486);
nand U14553 (N_14553,N_12039,N_13279);
nand U14554 (N_14554,N_12698,N_12156);
xor U14555 (N_14555,N_12370,N_12112);
nor U14556 (N_14556,N_12858,N_12537);
and U14557 (N_14557,N_12317,N_12693);
and U14558 (N_14558,N_13015,N_13363);
and U14559 (N_14559,N_12537,N_13171);
or U14560 (N_14560,N_12450,N_13443);
xnor U14561 (N_14561,N_13489,N_13183);
nor U14562 (N_14562,N_12176,N_12429);
nand U14563 (N_14563,N_12277,N_12951);
xnor U14564 (N_14564,N_13108,N_12120);
xor U14565 (N_14565,N_12733,N_13211);
or U14566 (N_14566,N_12528,N_12776);
nor U14567 (N_14567,N_12684,N_12002);
or U14568 (N_14568,N_12963,N_12671);
xnor U14569 (N_14569,N_13281,N_12855);
and U14570 (N_14570,N_13383,N_12214);
and U14571 (N_14571,N_12830,N_12466);
or U14572 (N_14572,N_13313,N_13190);
or U14573 (N_14573,N_13222,N_13196);
xnor U14574 (N_14574,N_12385,N_13438);
and U14575 (N_14575,N_12494,N_12606);
xor U14576 (N_14576,N_12030,N_12572);
nand U14577 (N_14577,N_13214,N_13234);
xnor U14578 (N_14578,N_13493,N_13208);
nor U14579 (N_14579,N_13089,N_13139);
nor U14580 (N_14580,N_12187,N_12780);
nand U14581 (N_14581,N_13039,N_13436);
xnor U14582 (N_14582,N_13393,N_12084);
and U14583 (N_14583,N_12347,N_12250);
nand U14584 (N_14584,N_12779,N_12671);
nand U14585 (N_14585,N_13432,N_12374);
nor U14586 (N_14586,N_12690,N_13420);
and U14587 (N_14587,N_12879,N_12946);
xnor U14588 (N_14588,N_13095,N_12897);
or U14589 (N_14589,N_13267,N_12831);
nand U14590 (N_14590,N_12030,N_12214);
xnor U14591 (N_14591,N_13348,N_13279);
and U14592 (N_14592,N_12337,N_13042);
and U14593 (N_14593,N_12087,N_12124);
nand U14594 (N_14594,N_13472,N_12367);
nor U14595 (N_14595,N_13156,N_13387);
xnor U14596 (N_14596,N_12805,N_12506);
nand U14597 (N_14597,N_13170,N_12666);
nand U14598 (N_14598,N_12214,N_12060);
or U14599 (N_14599,N_12734,N_12893);
nand U14600 (N_14600,N_12612,N_12382);
and U14601 (N_14601,N_12296,N_12199);
nor U14602 (N_14602,N_12070,N_12373);
nor U14603 (N_14603,N_12784,N_12033);
nor U14604 (N_14604,N_12424,N_13142);
nor U14605 (N_14605,N_13154,N_13278);
and U14606 (N_14606,N_12787,N_12995);
nor U14607 (N_14607,N_13391,N_12024);
nor U14608 (N_14608,N_12421,N_12962);
xnor U14609 (N_14609,N_12006,N_12290);
nor U14610 (N_14610,N_13442,N_12146);
nor U14611 (N_14611,N_13355,N_12768);
nor U14612 (N_14612,N_13121,N_12078);
xor U14613 (N_14613,N_13051,N_12598);
xnor U14614 (N_14614,N_12303,N_12126);
xnor U14615 (N_14615,N_13129,N_12855);
nand U14616 (N_14616,N_12475,N_13172);
nor U14617 (N_14617,N_12942,N_13225);
or U14618 (N_14618,N_12465,N_12346);
nand U14619 (N_14619,N_12764,N_12360);
nor U14620 (N_14620,N_13305,N_13465);
or U14621 (N_14621,N_13206,N_12430);
nor U14622 (N_14622,N_12303,N_13453);
and U14623 (N_14623,N_12316,N_13192);
nand U14624 (N_14624,N_13447,N_12763);
nor U14625 (N_14625,N_13421,N_12651);
and U14626 (N_14626,N_12560,N_12315);
nor U14627 (N_14627,N_12342,N_12766);
or U14628 (N_14628,N_13443,N_12762);
or U14629 (N_14629,N_12006,N_13346);
nor U14630 (N_14630,N_13271,N_12135);
xnor U14631 (N_14631,N_12752,N_12531);
nor U14632 (N_14632,N_12681,N_12129);
nor U14633 (N_14633,N_13206,N_12137);
nor U14634 (N_14634,N_13034,N_12609);
or U14635 (N_14635,N_13083,N_12500);
xor U14636 (N_14636,N_13183,N_13165);
nand U14637 (N_14637,N_12088,N_13119);
and U14638 (N_14638,N_12022,N_12652);
nor U14639 (N_14639,N_12582,N_12557);
nor U14640 (N_14640,N_12024,N_12151);
xnor U14641 (N_14641,N_12869,N_12467);
and U14642 (N_14642,N_13024,N_12338);
or U14643 (N_14643,N_12806,N_12644);
nor U14644 (N_14644,N_12866,N_12981);
nor U14645 (N_14645,N_13382,N_12674);
nor U14646 (N_14646,N_12090,N_13459);
or U14647 (N_14647,N_12028,N_12764);
or U14648 (N_14648,N_13291,N_13364);
and U14649 (N_14649,N_12364,N_12501);
nor U14650 (N_14650,N_12996,N_12226);
xor U14651 (N_14651,N_12086,N_13468);
and U14652 (N_14652,N_13033,N_12240);
or U14653 (N_14653,N_12686,N_13112);
nand U14654 (N_14654,N_12437,N_13437);
and U14655 (N_14655,N_12626,N_12055);
nor U14656 (N_14656,N_12495,N_12125);
or U14657 (N_14657,N_12720,N_12582);
and U14658 (N_14658,N_12626,N_12722);
nand U14659 (N_14659,N_12220,N_12597);
and U14660 (N_14660,N_13440,N_13192);
nor U14661 (N_14661,N_12804,N_12619);
or U14662 (N_14662,N_12146,N_12105);
nand U14663 (N_14663,N_12636,N_12541);
or U14664 (N_14664,N_12137,N_13277);
nand U14665 (N_14665,N_12203,N_12207);
nor U14666 (N_14666,N_12487,N_12943);
nor U14667 (N_14667,N_12028,N_13219);
nor U14668 (N_14668,N_12967,N_13213);
nor U14669 (N_14669,N_13063,N_12763);
xor U14670 (N_14670,N_12297,N_13284);
or U14671 (N_14671,N_12104,N_12006);
nand U14672 (N_14672,N_13158,N_12958);
and U14673 (N_14673,N_12741,N_13299);
xor U14674 (N_14674,N_12018,N_13470);
and U14675 (N_14675,N_13304,N_12688);
nand U14676 (N_14676,N_13488,N_12392);
xor U14677 (N_14677,N_12030,N_12347);
nor U14678 (N_14678,N_12806,N_13167);
or U14679 (N_14679,N_12983,N_13409);
nand U14680 (N_14680,N_12436,N_12841);
xnor U14681 (N_14681,N_13285,N_12073);
nand U14682 (N_14682,N_13140,N_12029);
nand U14683 (N_14683,N_12342,N_13061);
nand U14684 (N_14684,N_12103,N_12727);
nand U14685 (N_14685,N_12410,N_13337);
xnor U14686 (N_14686,N_13053,N_13249);
xor U14687 (N_14687,N_12039,N_13134);
or U14688 (N_14688,N_13278,N_12473);
nand U14689 (N_14689,N_12092,N_12600);
nand U14690 (N_14690,N_13455,N_12754);
or U14691 (N_14691,N_13288,N_12550);
or U14692 (N_14692,N_13398,N_12884);
nor U14693 (N_14693,N_12469,N_12863);
xnor U14694 (N_14694,N_12445,N_13331);
xor U14695 (N_14695,N_12464,N_12426);
xor U14696 (N_14696,N_13380,N_12037);
xor U14697 (N_14697,N_13453,N_12449);
nor U14698 (N_14698,N_12611,N_13310);
and U14699 (N_14699,N_13493,N_12295);
or U14700 (N_14700,N_13114,N_12027);
nand U14701 (N_14701,N_12547,N_13310);
nand U14702 (N_14702,N_12100,N_12444);
nand U14703 (N_14703,N_12502,N_13370);
nor U14704 (N_14704,N_13473,N_12954);
or U14705 (N_14705,N_12700,N_12549);
xnor U14706 (N_14706,N_13019,N_12959);
nor U14707 (N_14707,N_13389,N_12922);
xnor U14708 (N_14708,N_12455,N_12607);
nor U14709 (N_14709,N_13416,N_12719);
or U14710 (N_14710,N_12773,N_12274);
or U14711 (N_14711,N_12170,N_13017);
nand U14712 (N_14712,N_12351,N_12648);
xor U14713 (N_14713,N_12953,N_13031);
nor U14714 (N_14714,N_12461,N_12154);
nand U14715 (N_14715,N_12606,N_13496);
and U14716 (N_14716,N_12443,N_12764);
nand U14717 (N_14717,N_12411,N_13489);
or U14718 (N_14718,N_12757,N_13274);
xnor U14719 (N_14719,N_12318,N_12065);
nand U14720 (N_14720,N_13382,N_12594);
or U14721 (N_14721,N_13291,N_13004);
and U14722 (N_14722,N_13450,N_13337);
and U14723 (N_14723,N_13353,N_12363);
xor U14724 (N_14724,N_12354,N_13282);
nand U14725 (N_14725,N_12060,N_13408);
xnor U14726 (N_14726,N_12804,N_12093);
or U14727 (N_14727,N_13361,N_12494);
or U14728 (N_14728,N_12783,N_12111);
and U14729 (N_14729,N_13363,N_12598);
nor U14730 (N_14730,N_12529,N_13232);
and U14731 (N_14731,N_12733,N_12030);
nand U14732 (N_14732,N_12299,N_12719);
nor U14733 (N_14733,N_12394,N_12811);
nand U14734 (N_14734,N_12554,N_12188);
and U14735 (N_14735,N_12047,N_12665);
and U14736 (N_14736,N_12289,N_13354);
nand U14737 (N_14737,N_12086,N_13418);
xor U14738 (N_14738,N_12655,N_13356);
or U14739 (N_14739,N_12576,N_12150);
nor U14740 (N_14740,N_12050,N_12951);
nor U14741 (N_14741,N_12099,N_13427);
nand U14742 (N_14742,N_12410,N_12229);
and U14743 (N_14743,N_12862,N_13467);
xnor U14744 (N_14744,N_12198,N_12901);
xor U14745 (N_14745,N_12752,N_12898);
or U14746 (N_14746,N_12438,N_13340);
nand U14747 (N_14747,N_13369,N_12786);
xnor U14748 (N_14748,N_12872,N_13461);
xnor U14749 (N_14749,N_12319,N_12064);
xor U14750 (N_14750,N_12151,N_12922);
and U14751 (N_14751,N_13033,N_12830);
xor U14752 (N_14752,N_13016,N_12981);
nand U14753 (N_14753,N_12006,N_13172);
and U14754 (N_14754,N_12491,N_12613);
xor U14755 (N_14755,N_13032,N_12016);
nand U14756 (N_14756,N_13300,N_13400);
or U14757 (N_14757,N_13254,N_12870);
and U14758 (N_14758,N_13372,N_13403);
or U14759 (N_14759,N_12793,N_12758);
nand U14760 (N_14760,N_13381,N_12224);
nand U14761 (N_14761,N_12661,N_12452);
nand U14762 (N_14762,N_12905,N_12793);
nor U14763 (N_14763,N_12120,N_12163);
and U14764 (N_14764,N_12013,N_12135);
or U14765 (N_14765,N_12943,N_13133);
or U14766 (N_14766,N_13476,N_12023);
nand U14767 (N_14767,N_12810,N_12760);
nand U14768 (N_14768,N_13420,N_13092);
xnor U14769 (N_14769,N_13369,N_12851);
and U14770 (N_14770,N_13348,N_12364);
or U14771 (N_14771,N_12419,N_12473);
or U14772 (N_14772,N_12111,N_12505);
nor U14773 (N_14773,N_13387,N_12149);
and U14774 (N_14774,N_13040,N_13072);
and U14775 (N_14775,N_12167,N_12330);
xor U14776 (N_14776,N_12500,N_13433);
nand U14777 (N_14777,N_12165,N_12387);
or U14778 (N_14778,N_12572,N_12088);
nor U14779 (N_14779,N_12477,N_13243);
nor U14780 (N_14780,N_13139,N_12656);
or U14781 (N_14781,N_13162,N_12003);
nor U14782 (N_14782,N_12892,N_12036);
nand U14783 (N_14783,N_12683,N_12306);
nand U14784 (N_14784,N_13252,N_13364);
and U14785 (N_14785,N_12028,N_13292);
nor U14786 (N_14786,N_13065,N_12302);
nand U14787 (N_14787,N_12939,N_12679);
nand U14788 (N_14788,N_12312,N_12702);
and U14789 (N_14789,N_13476,N_12458);
or U14790 (N_14790,N_13320,N_12236);
nor U14791 (N_14791,N_12415,N_13035);
nor U14792 (N_14792,N_12446,N_12408);
nand U14793 (N_14793,N_12621,N_13395);
nor U14794 (N_14794,N_12750,N_12254);
xnor U14795 (N_14795,N_12972,N_13463);
xor U14796 (N_14796,N_13283,N_12898);
xnor U14797 (N_14797,N_13286,N_12360);
nand U14798 (N_14798,N_12359,N_12825);
nor U14799 (N_14799,N_13126,N_12246);
and U14800 (N_14800,N_13292,N_12088);
or U14801 (N_14801,N_12912,N_12080);
nand U14802 (N_14802,N_12800,N_12228);
and U14803 (N_14803,N_13364,N_12733);
or U14804 (N_14804,N_13302,N_12797);
xor U14805 (N_14805,N_12298,N_12803);
and U14806 (N_14806,N_12294,N_12837);
nor U14807 (N_14807,N_13403,N_12152);
nor U14808 (N_14808,N_12950,N_13085);
nor U14809 (N_14809,N_12546,N_12364);
nand U14810 (N_14810,N_12322,N_13334);
or U14811 (N_14811,N_12719,N_12268);
or U14812 (N_14812,N_13211,N_13088);
nor U14813 (N_14813,N_12728,N_12593);
and U14814 (N_14814,N_12636,N_12500);
xnor U14815 (N_14815,N_12759,N_12310);
nand U14816 (N_14816,N_12223,N_12722);
xor U14817 (N_14817,N_12915,N_12025);
or U14818 (N_14818,N_12089,N_12985);
nor U14819 (N_14819,N_13151,N_13489);
nor U14820 (N_14820,N_13209,N_13162);
xor U14821 (N_14821,N_13476,N_12125);
nand U14822 (N_14822,N_12073,N_12064);
xor U14823 (N_14823,N_12959,N_12405);
or U14824 (N_14824,N_12259,N_12574);
and U14825 (N_14825,N_13294,N_12181);
nor U14826 (N_14826,N_12309,N_12473);
nand U14827 (N_14827,N_12830,N_12135);
nor U14828 (N_14828,N_13422,N_13262);
and U14829 (N_14829,N_13208,N_12834);
xnor U14830 (N_14830,N_13450,N_13350);
xnor U14831 (N_14831,N_12546,N_12467);
nor U14832 (N_14832,N_12405,N_13024);
nor U14833 (N_14833,N_12523,N_12709);
xnor U14834 (N_14834,N_12852,N_13460);
nor U14835 (N_14835,N_12763,N_12126);
or U14836 (N_14836,N_12039,N_12206);
xnor U14837 (N_14837,N_12174,N_12157);
xor U14838 (N_14838,N_12159,N_12075);
nand U14839 (N_14839,N_12422,N_12447);
and U14840 (N_14840,N_12027,N_13446);
and U14841 (N_14841,N_13282,N_13171);
or U14842 (N_14842,N_12298,N_12643);
nand U14843 (N_14843,N_12338,N_13269);
and U14844 (N_14844,N_13447,N_13376);
or U14845 (N_14845,N_12820,N_12463);
and U14846 (N_14846,N_13419,N_12878);
and U14847 (N_14847,N_12176,N_12701);
and U14848 (N_14848,N_12421,N_12523);
or U14849 (N_14849,N_13193,N_12859);
nand U14850 (N_14850,N_13270,N_12332);
or U14851 (N_14851,N_13199,N_12421);
or U14852 (N_14852,N_13260,N_12540);
xor U14853 (N_14853,N_12607,N_12658);
xor U14854 (N_14854,N_13116,N_13432);
nor U14855 (N_14855,N_12415,N_13146);
and U14856 (N_14856,N_12046,N_12100);
or U14857 (N_14857,N_13198,N_12904);
nand U14858 (N_14858,N_13100,N_12766);
nor U14859 (N_14859,N_13360,N_12767);
and U14860 (N_14860,N_13176,N_12700);
or U14861 (N_14861,N_13333,N_12526);
xor U14862 (N_14862,N_13498,N_13325);
and U14863 (N_14863,N_13234,N_13150);
nor U14864 (N_14864,N_12521,N_13121);
xor U14865 (N_14865,N_13027,N_12257);
nand U14866 (N_14866,N_12220,N_12092);
nand U14867 (N_14867,N_12523,N_12178);
or U14868 (N_14868,N_13353,N_12962);
nor U14869 (N_14869,N_13400,N_12535);
or U14870 (N_14870,N_13041,N_12838);
nand U14871 (N_14871,N_12715,N_12959);
or U14872 (N_14872,N_12983,N_12807);
or U14873 (N_14873,N_13045,N_12950);
and U14874 (N_14874,N_12636,N_12902);
nand U14875 (N_14875,N_12068,N_12391);
nor U14876 (N_14876,N_12626,N_13050);
xor U14877 (N_14877,N_12011,N_12609);
nand U14878 (N_14878,N_12848,N_12459);
xor U14879 (N_14879,N_12794,N_12978);
xnor U14880 (N_14880,N_12570,N_12981);
or U14881 (N_14881,N_13071,N_13444);
and U14882 (N_14882,N_13465,N_12388);
nor U14883 (N_14883,N_13122,N_13142);
nand U14884 (N_14884,N_12886,N_13052);
and U14885 (N_14885,N_12657,N_12062);
and U14886 (N_14886,N_13267,N_12966);
or U14887 (N_14887,N_12290,N_13406);
xor U14888 (N_14888,N_12826,N_12043);
nor U14889 (N_14889,N_12286,N_12592);
and U14890 (N_14890,N_12740,N_13175);
xor U14891 (N_14891,N_12617,N_12241);
and U14892 (N_14892,N_12243,N_12206);
or U14893 (N_14893,N_13169,N_12180);
and U14894 (N_14894,N_12134,N_13026);
nor U14895 (N_14895,N_12268,N_13345);
xnor U14896 (N_14896,N_12630,N_12902);
and U14897 (N_14897,N_12108,N_12285);
or U14898 (N_14898,N_12543,N_13112);
xnor U14899 (N_14899,N_12284,N_12042);
nor U14900 (N_14900,N_12003,N_12054);
nand U14901 (N_14901,N_13244,N_12169);
nor U14902 (N_14902,N_12006,N_12950);
and U14903 (N_14903,N_12411,N_12281);
nand U14904 (N_14904,N_13306,N_12394);
nor U14905 (N_14905,N_13303,N_12297);
nor U14906 (N_14906,N_12434,N_13103);
and U14907 (N_14907,N_12848,N_13320);
and U14908 (N_14908,N_12693,N_12774);
and U14909 (N_14909,N_12993,N_12649);
nor U14910 (N_14910,N_12320,N_12269);
xnor U14911 (N_14911,N_12340,N_12456);
nand U14912 (N_14912,N_12052,N_12002);
and U14913 (N_14913,N_12523,N_12092);
or U14914 (N_14914,N_13202,N_13193);
xnor U14915 (N_14915,N_12608,N_12531);
xnor U14916 (N_14916,N_12027,N_12788);
nor U14917 (N_14917,N_12343,N_12913);
xnor U14918 (N_14918,N_12554,N_13354);
nor U14919 (N_14919,N_12471,N_12839);
or U14920 (N_14920,N_13363,N_13445);
or U14921 (N_14921,N_13322,N_12147);
nor U14922 (N_14922,N_12701,N_13434);
nor U14923 (N_14923,N_13285,N_12682);
and U14924 (N_14924,N_13335,N_12861);
and U14925 (N_14925,N_12221,N_12377);
or U14926 (N_14926,N_12625,N_13375);
and U14927 (N_14927,N_12459,N_12123);
xnor U14928 (N_14928,N_12261,N_13175);
xnor U14929 (N_14929,N_12729,N_12725);
xnor U14930 (N_14930,N_12779,N_12927);
or U14931 (N_14931,N_12104,N_12256);
nand U14932 (N_14932,N_12444,N_12624);
nand U14933 (N_14933,N_12471,N_12676);
nand U14934 (N_14934,N_12631,N_12420);
and U14935 (N_14935,N_12784,N_12681);
and U14936 (N_14936,N_12256,N_13306);
and U14937 (N_14937,N_12198,N_13234);
nor U14938 (N_14938,N_12243,N_13074);
or U14939 (N_14939,N_13170,N_13409);
xor U14940 (N_14940,N_12528,N_12199);
nand U14941 (N_14941,N_12240,N_12467);
xnor U14942 (N_14942,N_13373,N_13262);
xor U14943 (N_14943,N_13460,N_12309);
xnor U14944 (N_14944,N_12070,N_13100);
nand U14945 (N_14945,N_13477,N_12772);
or U14946 (N_14946,N_12631,N_12415);
nor U14947 (N_14947,N_13474,N_12266);
or U14948 (N_14948,N_12510,N_13353);
xnor U14949 (N_14949,N_13379,N_12836);
nor U14950 (N_14950,N_12756,N_12094);
and U14951 (N_14951,N_12648,N_13196);
xnor U14952 (N_14952,N_13414,N_12591);
xnor U14953 (N_14953,N_13270,N_12502);
xor U14954 (N_14954,N_13285,N_12559);
nor U14955 (N_14955,N_12925,N_12107);
xnor U14956 (N_14956,N_12752,N_13019);
and U14957 (N_14957,N_12311,N_13367);
or U14958 (N_14958,N_12799,N_12645);
and U14959 (N_14959,N_13197,N_13017);
or U14960 (N_14960,N_12795,N_13072);
and U14961 (N_14961,N_12385,N_12353);
nand U14962 (N_14962,N_12373,N_12926);
and U14963 (N_14963,N_13446,N_12855);
nor U14964 (N_14964,N_12269,N_12374);
nor U14965 (N_14965,N_12899,N_12248);
and U14966 (N_14966,N_12054,N_13266);
or U14967 (N_14967,N_13286,N_12705);
or U14968 (N_14968,N_12751,N_12202);
nor U14969 (N_14969,N_12526,N_12033);
and U14970 (N_14970,N_12228,N_13485);
or U14971 (N_14971,N_12270,N_12576);
nor U14972 (N_14972,N_12698,N_13362);
and U14973 (N_14973,N_12743,N_12670);
and U14974 (N_14974,N_13412,N_12478);
and U14975 (N_14975,N_13310,N_12659);
and U14976 (N_14976,N_12349,N_12615);
or U14977 (N_14977,N_13340,N_12135);
nor U14978 (N_14978,N_12449,N_12744);
or U14979 (N_14979,N_13109,N_13205);
nand U14980 (N_14980,N_13326,N_13159);
xor U14981 (N_14981,N_13333,N_12989);
and U14982 (N_14982,N_12849,N_12235);
xnor U14983 (N_14983,N_12528,N_13031);
or U14984 (N_14984,N_12867,N_12131);
xor U14985 (N_14985,N_12013,N_12072);
and U14986 (N_14986,N_12178,N_12139);
nand U14987 (N_14987,N_12026,N_12221);
xnor U14988 (N_14988,N_13217,N_13105);
nand U14989 (N_14989,N_12768,N_13135);
xor U14990 (N_14990,N_13485,N_12462);
nand U14991 (N_14991,N_12931,N_12756);
nand U14992 (N_14992,N_13113,N_12686);
and U14993 (N_14993,N_12324,N_12817);
or U14994 (N_14994,N_12435,N_12529);
or U14995 (N_14995,N_13483,N_12355);
or U14996 (N_14996,N_12596,N_12911);
nor U14997 (N_14997,N_12202,N_12794);
xor U14998 (N_14998,N_13052,N_13178);
xor U14999 (N_14999,N_12957,N_12527);
nor U15000 (N_15000,N_14401,N_13590);
nor U15001 (N_15001,N_14066,N_13874);
nand U15002 (N_15002,N_14676,N_14684);
nand U15003 (N_15003,N_14866,N_13789);
or U15004 (N_15004,N_14240,N_14029);
xor U15005 (N_15005,N_14476,N_14126);
or U15006 (N_15006,N_13885,N_14856);
and U15007 (N_15007,N_14209,N_14742);
nand U15008 (N_15008,N_14148,N_13866);
nand U15009 (N_15009,N_14344,N_14728);
and U15010 (N_15010,N_14058,N_14767);
and U15011 (N_15011,N_14446,N_13548);
xor U15012 (N_15012,N_14818,N_13762);
xor U15013 (N_15013,N_14044,N_14501);
nand U15014 (N_15014,N_14068,N_13618);
nor U15015 (N_15015,N_13586,N_14153);
or U15016 (N_15016,N_14226,N_14549);
xnor U15017 (N_15017,N_14535,N_14933);
nor U15018 (N_15018,N_14995,N_13985);
nor U15019 (N_15019,N_13931,N_14237);
or U15020 (N_15020,N_14613,N_14335);
and U15021 (N_15021,N_13938,N_14521);
or U15022 (N_15022,N_14439,N_13587);
nor U15023 (N_15023,N_14248,N_14449);
nor U15024 (N_15024,N_14485,N_13783);
or U15025 (N_15025,N_14729,N_13860);
nand U15026 (N_15026,N_13830,N_13663);
nand U15027 (N_15027,N_14942,N_13514);
nor U15028 (N_15028,N_13792,N_14215);
or U15029 (N_15029,N_13575,N_14940);
xor U15030 (N_15030,N_14218,N_14991);
or U15031 (N_15031,N_14482,N_13650);
nand U15032 (N_15032,N_13827,N_13956);
and U15033 (N_15033,N_13670,N_13883);
nand U15034 (N_15034,N_14494,N_14517);
and U15035 (N_15035,N_14574,N_13741);
nor U15036 (N_15036,N_14046,N_13601);
xnor U15037 (N_15037,N_13527,N_13844);
nand U15038 (N_15038,N_13731,N_13542);
xor U15039 (N_15039,N_13612,N_14602);
and U15040 (N_15040,N_13683,N_14558);
xor U15041 (N_15041,N_14496,N_13773);
xnor U15042 (N_15042,N_13732,N_14430);
or U15043 (N_15043,N_13609,N_14853);
nand U15044 (N_15044,N_14758,N_13557);
nor U15045 (N_15045,N_14698,N_14421);
nor U15046 (N_15046,N_14817,N_14487);
or U15047 (N_15047,N_13721,N_14162);
nor U15048 (N_15048,N_13843,N_14263);
xnor U15049 (N_15049,N_14834,N_14082);
nand U15050 (N_15050,N_14099,N_13686);
nand U15051 (N_15051,N_14718,N_13564);
xor U15052 (N_15052,N_14376,N_14552);
or U15053 (N_15053,N_14310,N_14125);
and U15054 (N_15054,N_14318,N_14283);
nand U15055 (N_15055,N_14929,N_14025);
or U15056 (N_15056,N_14909,N_14720);
nor U15057 (N_15057,N_14147,N_14726);
or U15058 (N_15058,N_14217,N_14682);
xor U15059 (N_15059,N_13616,N_13652);
nor U15060 (N_15060,N_13972,N_14548);
or U15061 (N_15061,N_13727,N_13513);
nand U15062 (N_15062,N_14403,N_14631);
xnor U15063 (N_15063,N_13695,N_14806);
and U15064 (N_15064,N_14087,N_14234);
xor U15065 (N_15065,N_14298,N_14073);
xnor U15066 (N_15066,N_14898,N_13770);
xor U15067 (N_15067,N_13978,N_13791);
and U15068 (N_15068,N_13696,N_14183);
nand U15069 (N_15069,N_14400,N_13822);
xor U15070 (N_15070,N_14832,N_14406);
nand U15071 (N_15071,N_14170,N_14792);
nor U15072 (N_15072,N_14712,N_14737);
nor U15073 (N_15073,N_14645,N_14634);
nor U15074 (N_15074,N_13636,N_13966);
and U15075 (N_15075,N_14269,N_13999);
nor U15076 (N_15076,N_14803,N_13613);
nand U15077 (N_15077,N_14828,N_13880);
nor U15078 (N_15078,N_14708,N_14661);
nand U15079 (N_15079,N_14242,N_14716);
or U15080 (N_15080,N_13908,N_14724);
xnor U15081 (N_15081,N_14876,N_14700);
xnor U15082 (N_15082,N_14197,N_14214);
nor U15083 (N_15083,N_13918,N_14247);
or U15084 (N_15084,N_14951,N_14090);
or U15085 (N_15085,N_14561,N_14470);
nor U15086 (N_15086,N_14241,N_14659);
nand U15087 (N_15087,N_14596,N_13550);
or U15088 (N_15088,N_14727,N_14789);
nand U15089 (N_15089,N_14911,N_14765);
and U15090 (N_15090,N_14685,N_14220);
nor U15091 (N_15091,N_13664,N_13976);
nor U15092 (N_15092,N_13647,N_13506);
nor U15093 (N_15093,N_14831,N_14670);
or U15094 (N_15094,N_13625,N_13904);
xnor U15095 (N_15095,N_14469,N_14748);
nor U15096 (N_15096,N_13697,N_14976);
or U15097 (N_15097,N_13814,N_14041);
or U15098 (N_15098,N_13558,N_14287);
nor U15099 (N_15099,N_13679,N_14018);
xnor U15100 (N_15100,N_14925,N_14489);
nor U15101 (N_15101,N_14594,N_14711);
or U15102 (N_15102,N_13848,N_14175);
or U15103 (N_15103,N_13975,N_14761);
nor U15104 (N_15104,N_14683,N_13782);
xnor U15105 (N_15105,N_14134,N_14585);
or U15106 (N_15106,N_14580,N_14579);
nand U15107 (N_15107,N_14363,N_13617);
nand U15108 (N_15108,N_13855,N_14352);
nor U15109 (N_15109,N_14045,N_14979);
nor U15110 (N_15110,N_14042,N_13959);
nor U15111 (N_15111,N_14502,N_14905);
nand U15112 (N_15112,N_14703,N_13882);
nand U15113 (N_15113,N_14477,N_14719);
or U15114 (N_15114,N_14405,N_14907);
xnor U15115 (N_15115,N_14842,N_14709);
xnor U15116 (N_15116,N_14130,N_14691);
and U15117 (N_15117,N_14650,N_14349);
nand U15118 (N_15118,N_13559,N_13933);
nor U15119 (N_15119,N_13740,N_13632);
nor U15120 (N_15120,N_14358,N_13736);
nor U15121 (N_15121,N_14837,N_13849);
and U15122 (N_15122,N_14902,N_13797);
or U15123 (N_15123,N_14397,N_14393);
xor U15124 (N_15124,N_13940,N_13535);
nor U15125 (N_15125,N_13593,N_14394);
nor U15126 (N_15126,N_13911,N_13547);
and U15127 (N_15127,N_14395,N_13622);
xnor U15128 (N_15128,N_13929,N_14739);
and U15129 (N_15129,N_13517,N_13716);
nor U15130 (N_15130,N_13605,N_13501);
nor U15131 (N_15131,N_14434,N_13944);
nor U15132 (N_15132,N_13749,N_14428);
or U15133 (N_15133,N_14623,N_14048);
or U15134 (N_15134,N_14009,N_14576);
and U15135 (N_15135,N_14480,N_14996);
xnor U15136 (N_15136,N_14111,N_13901);
xor U15137 (N_15137,N_14507,N_14939);
nor U15138 (N_15138,N_13539,N_14355);
nand U15139 (N_15139,N_13812,N_14267);
or U15140 (N_15140,N_14696,N_14776);
nand U15141 (N_15141,N_14014,N_14182);
nor U15142 (N_15142,N_14750,N_14144);
and U15143 (N_15143,N_13576,N_14367);
nor U15144 (N_15144,N_14591,N_14997);
or U15145 (N_15145,N_13896,N_13687);
nand U15146 (N_15146,N_13841,N_14740);
or U15147 (N_15147,N_14804,N_14903);
and U15148 (N_15148,N_13536,N_14096);
and U15149 (N_15149,N_13873,N_14266);
nor U15150 (N_15150,N_14201,N_13832);
or U15151 (N_15151,N_14338,N_14589);
nand U15152 (N_15152,N_14086,N_14398);
and U15153 (N_15153,N_13853,N_14999);
xor U15154 (N_15154,N_14163,N_13596);
or U15155 (N_15155,N_14302,N_14990);
and U15156 (N_15156,N_14199,N_14968);
and U15157 (N_15157,N_13733,N_14923);
or U15158 (N_15158,N_14347,N_14833);
or U15159 (N_15159,N_13916,N_13977);
nand U15160 (N_15160,N_14206,N_14190);
nor U15161 (N_15161,N_14080,N_14305);
nor U15162 (N_15162,N_14572,N_14402);
xor U15163 (N_15163,N_13724,N_13584);
nor U15164 (N_15164,N_13953,N_14440);
nor U15165 (N_15165,N_14910,N_13910);
nor U15166 (N_15166,N_14284,N_14205);
nor U15167 (N_15167,N_14020,N_13702);
nor U15168 (N_15168,N_13598,N_14345);
xnor U15169 (N_15169,N_14459,N_14760);
or U15170 (N_15170,N_14513,N_14464);
nor U15171 (N_15171,N_14076,N_14953);
xor U15172 (N_15172,N_14644,N_13546);
nand U15173 (N_15173,N_14977,N_14294);
and U15174 (N_15174,N_14889,N_14187);
or U15175 (N_15175,N_13989,N_13756);
or U15176 (N_15176,N_14617,N_14555);
and U15177 (N_15177,N_14749,N_14260);
or U15178 (N_15178,N_13681,N_14836);
nor U15179 (N_15179,N_14427,N_14523);
nor U15180 (N_15180,N_14895,N_14559);
and U15181 (N_15181,N_13656,N_14094);
nor U15182 (N_15182,N_13665,N_14825);
nor U15183 (N_15183,N_14114,N_13788);
nor U15184 (N_15184,N_14551,N_14830);
nor U15185 (N_15185,N_14000,N_13766);
nand U15186 (N_15186,N_14746,N_13887);
nand U15187 (N_15187,N_14871,N_14787);
nor U15188 (N_15188,N_13675,N_14004);
or U15189 (N_15189,N_14541,N_13942);
nor U15190 (N_15190,N_14462,N_13745);
xor U15191 (N_15191,N_14587,N_13599);
nand U15192 (N_15192,N_14669,N_14678);
nand U15193 (N_15193,N_14992,N_13932);
and U15194 (N_15194,N_14515,N_14178);
and U15195 (N_15195,N_14962,N_14304);
nor U15196 (N_15196,N_14544,N_14736);
nand U15197 (N_15197,N_13723,N_14658);
nand U15198 (N_15198,N_14584,N_13754);
or U15199 (N_15199,N_13893,N_14475);
xor U15200 (N_15200,N_13804,N_13962);
and U15201 (N_15201,N_13528,N_14067);
nand U15202 (N_15202,N_13748,N_14961);
xor U15203 (N_15203,N_14447,N_13631);
and U15204 (N_15204,N_14132,N_14399);
or U15205 (N_15205,N_14754,N_14875);
nor U15206 (N_15206,N_13961,N_14829);
and U15207 (N_15207,N_14486,N_14627);
nand U15208 (N_15208,N_13900,N_13897);
xnor U15209 (N_15209,N_14966,N_14822);
nor U15210 (N_15210,N_14200,N_14981);
xor U15211 (N_15211,N_14024,N_13921);
and U15212 (N_15212,N_14371,N_13560);
and U15213 (N_15213,N_14801,N_13825);
nand U15214 (N_15214,N_14835,N_14137);
and U15215 (N_15215,N_13694,N_14954);
nor U15216 (N_15216,N_14180,N_14495);
or U15217 (N_15217,N_14013,N_14612);
nor U15218 (N_15218,N_14914,N_13820);
xor U15219 (N_15219,N_13516,N_13951);
and U15220 (N_15220,N_14624,N_14500);
nand U15221 (N_15221,N_14191,N_14564);
nand U15222 (N_15222,N_14978,N_14693);
nor U15223 (N_15223,N_14243,N_14504);
nor U15224 (N_15224,N_14770,N_14662);
xor U15225 (N_15225,N_14257,N_13693);
nand U15226 (N_15226,N_14780,N_14651);
xor U15227 (N_15227,N_14356,N_14880);
or U15228 (N_15228,N_13668,N_13915);
or U15229 (N_15229,N_14531,N_14643);
or U15230 (N_15230,N_14797,N_14926);
nand U15231 (N_15231,N_13705,N_14100);
and U15232 (N_15232,N_14415,N_14616);
or U15233 (N_15233,N_14568,N_14556);
xnor U15234 (N_15234,N_13523,N_14275);
nand U15235 (N_15235,N_13597,N_14619);
xnor U15236 (N_15236,N_14106,N_13717);
and U15237 (N_15237,N_14692,N_14854);
xor U15238 (N_15238,N_14849,N_14844);
or U15239 (N_15239,N_13997,N_14117);
nand U15240 (N_15240,N_13917,N_14107);
or U15241 (N_15241,N_14103,N_14941);
nor U15242 (N_15242,N_14127,N_14581);
and U15243 (N_15243,N_14276,N_14823);
and U15244 (N_15244,N_13872,N_14033);
nand U15245 (N_15245,N_13864,N_14625);
nor U15246 (N_15246,N_13980,N_14814);
or U15247 (N_15247,N_14472,N_13753);
nor U15248 (N_15248,N_14173,N_13595);
nand U15249 (N_15249,N_14306,N_13785);
or U15250 (N_15250,N_14286,N_14229);
or U15251 (N_15251,N_14799,N_13569);
nor U15252 (N_15252,N_13658,N_13919);
xnor U15253 (N_15253,N_13868,N_14769);
or U15254 (N_15254,N_14262,N_13905);
and U15255 (N_15255,N_14189,N_14537);
or U15256 (N_15256,N_13660,N_13769);
xor U15257 (N_15257,N_14956,N_14289);
nand U15258 (N_15258,N_13798,N_14845);
nor U15259 (N_15259,N_14618,N_14037);
nand U15260 (N_15260,N_14034,N_14946);
and U15261 (N_15261,N_13993,N_13881);
xnor U15262 (N_15262,N_14630,N_14960);
nor U15263 (N_15263,N_14164,N_14679);
or U15264 (N_15264,N_13774,N_13676);
nand U15265 (N_15265,N_14341,N_14988);
xor U15266 (N_15266,N_13592,N_14936);
or U15267 (N_15267,N_13643,N_13579);
xnor U15268 (N_15268,N_13509,N_14320);
nor U15269 (N_15269,N_14563,N_13570);
xnor U15270 (N_15270,N_14340,N_14158);
or U15271 (N_15271,N_14809,N_14453);
and U15272 (N_15272,N_14391,N_13699);
nand U15273 (N_15273,N_13817,N_14115);
nand U15274 (N_15274,N_14900,N_13903);
and U15275 (N_15275,N_14062,N_13790);
or U15276 (N_15276,N_14204,N_14466);
nand U15277 (N_15277,N_14455,N_13674);
nand U15278 (N_15278,N_13779,N_14641);
xnor U15279 (N_15279,N_13898,N_13627);
xor U15280 (N_15280,N_13979,N_14882);
nor U15281 (N_15281,N_14343,N_13588);
nand U15282 (N_15282,N_14874,N_14802);
and U15283 (N_15283,N_13994,N_14293);
xnor U15284 (N_15284,N_14075,N_14438);
or U15285 (N_15285,N_13713,N_14649);
or U15286 (N_15286,N_14252,N_14974);
and U15287 (N_15287,N_13553,N_13886);
and U15288 (N_15288,N_14884,N_14141);
or U15289 (N_15289,N_14852,N_14223);
xor U15290 (N_15290,N_14723,N_14943);
xnor U15291 (N_15291,N_14138,N_13525);
and U15292 (N_15292,N_13837,N_14983);
or U15293 (N_15293,N_14697,N_14931);
nor U15294 (N_15294,N_14721,N_14534);
or U15295 (N_15295,N_14969,N_13854);
nand U15296 (N_15296,N_14963,N_13765);
or U15297 (N_15297,N_13718,N_13661);
or U15298 (N_15298,N_14733,N_14586);
nand U15299 (N_15299,N_13786,N_14151);
and U15300 (N_15300,N_14605,N_14256);
nand U15301 (N_15301,N_14744,N_13628);
nor U15302 (N_15302,N_14278,N_14878);
xor U15303 (N_15303,N_14553,N_13920);
xnor U15304 (N_15304,N_13761,N_14411);
xor U15305 (N_15305,N_13698,N_14674);
nor U15306 (N_15306,N_13710,N_13706);
and U15307 (N_15307,N_14764,N_14575);
nor U15308 (N_15308,N_13682,N_13534);
nand U15309 (N_15309,N_14881,N_14311);
and U15310 (N_15310,N_13906,N_14527);
nand U15311 (N_15311,N_14493,N_13651);
nor U15312 (N_15312,N_14509,N_14407);
xnor U15313 (N_15313,N_13899,N_13971);
nor U15314 (N_15314,N_14277,N_14506);
xnor U15315 (N_15315,N_13737,N_14379);
nor U15316 (N_15316,N_13839,N_14689);
and U15317 (N_15317,N_14143,N_14443);
nand U15318 (N_15318,N_13757,N_13891);
and U15319 (N_15319,N_13970,N_13521);
xnor U15320 (N_15320,N_14543,N_14353);
nand U15321 (N_15321,N_14285,N_14657);
nand U15322 (N_15322,N_13680,N_14303);
and U15323 (N_15323,N_13561,N_13730);
or U15324 (N_15324,N_14361,N_14867);
nand U15325 (N_15325,N_14414,N_13955);
nand U15326 (N_15326,N_13811,N_13585);
and U15327 (N_15327,N_13568,N_13799);
and U15328 (N_15328,N_14452,N_14827);
xor U15329 (N_15329,N_13793,N_14036);
or U15330 (N_15330,N_13573,N_14920);
or U15331 (N_15331,N_14412,N_14597);
or U15332 (N_15332,N_14364,N_13505);
or U15333 (N_15333,N_13946,N_14308);
and U15334 (N_15334,N_13943,N_14167);
xnor U15335 (N_15335,N_14694,N_14794);
nor U15336 (N_15336,N_13728,N_14927);
nand U15337 (N_15337,N_13987,N_13764);
nor U15338 (N_15338,N_13986,N_14047);
nor U15339 (N_15339,N_14957,N_14639);
and U15340 (N_15340,N_13644,N_13602);
or U15341 (N_15341,N_13889,N_14425);
nor U15342 (N_15342,N_13771,N_13642);
or U15343 (N_15343,N_13875,N_14840);
nor U15344 (N_15344,N_13563,N_14265);
nand U15345 (N_15345,N_13815,N_13934);
nand U15346 (N_15346,N_14457,N_14959);
or U15347 (N_15347,N_13842,N_14342);
xnor U15348 (N_15348,N_14530,N_14172);
or U15349 (N_15349,N_13857,N_14213);
nor U15350 (N_15350,N_13930,N_14088);
xnor U15351 (N_15351,N_14777,N_14264);
or U15352 (N_15352,N_14897,N_14588);
or U15353 (N_15353,N_14741,N_13522);
or U15354 (N_15354,N_14196,N_14307);
nor U15355 (N_15355,N_13935,N_14993);
nor U15356 (N_15356,N_13649,N_14811);
or U15357 (N_15357,N_14194,N_13809);
or U15358 (N_15358,N_14301,N_14653);
nand U15359 (N_15359,N_14860,N_13800);
xor U15360 (N_15360,N_14442,N_14052);
and U15361 (N_15361,N_14177,N_14707);
xor U15362 (N_15362,N_14410,N_13600);
and U15363 (N_15363,N_14065,N_14539);
and U15364 (N_15364,N_14005,N_14757);
or U15365 (N_15365,N_14017,N_13512);
nor U15366 (N_15366,N_13531,N_14784);
nor U15367 (N_15367,N_14258,N_14893);
or U15368 (N_15368,N_14747,N_14686);
or U15369 (N_15369,N_14069,N_13719);
or U15370 (N_15370,N_14971,N_14778);
or U15371 (N_15371,N_14031,N_13926);
or U15372 (N_15372,N_14525,N_13856);
or U15373 (N_15373,N_14774,N_14230);
nand U15374 (N_15374,N_14948,N_13924);
and U15375 (N_15375,N_13876,N_14437);
nor U15376 (N_15376,N_14102,N_14077);
and U15377 (N_15377,N_13807,N_14635);
or U15378 (N_15378,N_13715,N_14505);
or U15379 (N_15379,N_14016,N_14015);
or U15380 (N_15380,N_13968,N_14123);
or U15381 (N_15381,N_14224,N_14296);
and U15382 (N_15382,N_14484,N_14660);
xnor U15383 (N_15383,N_13519,N_14595);
nand U15384 (N_15384,N_13928,N_13577);
nor U15385 (N_15385,N_13510,N_14498);
nor U15386 (N_15386,N_13655,N_14753);
nand U15387 (N_15387,N_14917,N_14314);
xor U15388 (N_15388,N_14492,N_13678);
or U15389 (N_15389,N_13677,N_14465);
or U15390 (N_15390,N_14348,N_13974);
nor U15391 (N_15391,N_14851,N_13796);
xnor U15392 (N_15392,N_13768,N_14611);
nor U15393 (N_15393,N_13801,N_13562);
or U15394 (N_15394,N_14432,N_14687);
xor U15395 (N_15395,N_14947,N_13692);
nand U15396 (N_15396,N_14300,N_14323);
nand U15397 (N_15397,N_14336,N_13673);
nand U15398 (N_15398,N_14628,N_14174);
xnor U15399 (N_15399,N_14456,N_14642);
or U15400 (N_15400,N_14710,N_14193);
nand U15401 (N_15401,N_14858,N_14629);
nand U15402 (N_15402,N_13795,N_14478);
and U15403 (N_15403,N_14357,N_14816);
xor U15404 (N_15404,N_13508,N_14848);
nand U15405 (N_15405,N_14212,N_13818);
or U15406 (N_15406,N_14652,N_14070);
nand U15407 (N_15407,N_14725,N_14610);
or U15408 (N_15408,N_13758,N_14176);
or U15409 (N_15409,N_14821,N_14445);
and U15410 (N_15410,N_14186,N_13549);
and U15411 (N_15411,N_14759,N_13688);
and U15412 (N_15412,N_13672,N_14673);
nor U15413 (N_15413,N_14423,N_14636);
or U15414 (N_15414,N_14565,N_14188);
nor U15415 (N_15415,N_14280,N_13529);
nor U15416 (N_15416,N_14524,N_14566);
nor U15417 (N_15417,N_14120,N_13626);
nor U15418 (N_15418,N_14731,N_14124);
and U15419 (N_15419,N_13998,N_13996);
and U15420 (N_15420,N_14315,N_14250);
nand U15421 (N_15421,N_14715,N_14781);
or U15422 (N_15422,N_14532,N_14608);
nand U15423 (N_15423,N_13635,N_14664);
nand U15424 (N_15424,N_14989,N_13530);
nand U15425 (N_15425,N_14582,N_14675);
or U15426 (N_15426,N_14150,N_14074);
or U15427 (N_15427,N_14609,N_14413);
or U15428 (N_15428,N_13925,N_14026);
or U15429 (N_15429,N_13895,N_13892);
nand U15430 (N_15430,N_13709,N_14329);
or U15431 (N_15431,N_14743,N_14236);
xor U15432 (N_15432,N_13828,N_14228);
and U15433 (N_15433,N_14987,N_13594);
nor U15434 (N_15434,N_14488,N_13954);
nand U15435 (N_15435,N_14104,N_14637);
nor U15436 (N_15436,N_13991,N_14454);
or U15437 (N_15437,N_13888,N_14131);
xor U15438 (N_15438,N_14392,N_14665);
nand U15439 (N_15439,N_13615,N_14093);
nand U15440 (N_15440,N_14688,N_14035);
or U15441 (N_15441,N_14370,N_14444);
and U15442 (N_15442,N_13772,N_14672);
and U15443 (N_15443,N_14570,N_14159);
and U15444 (N_15444,N_14762,N_14557);
and U15445 (N_15445,N_13614,N_14771);
xnor U15446 (N_15446,N_13545,N_14598);
and U15447 (N_15447,N_14497,N_14601);
or U15448 (N_15448,N_13816,N_13850);
nand U15449 (N_15449,N_14288,N_13927);
and U15450 (N_15450,N_14385,N_14232);
or U15451 (N_15451,N_14334,N_14207);
nor U15452 (N_15452,N_14061,N_13750);
nor U15453 (N_15453,N_14824,N_13781);
xor U15454 (N_15454,N_14049,N_14592);
nor U15455 (N_15455,N_13633,N_14192);
nand U15456 (N_15456,N_13566,N_13852);
nand U15457 (N_15457,N_14377,N_14239);
or U15458 (N_15458,N_14779,N_14663);
nand U15459 (N_15459,N_14820,N_14313);
and U15460 (N_15460,N_14451,N_13912);
xor U15461 (N_15461,N_14246,N_14529);
or U15462 (N_15462,N_14873,N_14021);
and U15463 (N_15463,N_14322,N_14896);
nor U15464 (N_15464,N_13623,N_14560);
and U15465 (N_15465,N_14038,N_14540);
and U15466 (N_15466,N_14547,N_14108);
or U15467 (N_15467,N_14632,N_13950);
nand U15468 (N_15468,N_13707,N_14463);
nand U15469 (N_15469,N_13701,N_14417);
or U15470 (N_15470,N_14928,N_14857);
or U15471 (N_15471,N_14508,N_13810);
or U15472 (N_15472,N_13725,N_13567);
nand U15473 (N_15473,N_13639,N_14503);
nor U15474 (N_15474,N_14590,N_14695);
nand U15475 (N_15475,N_14766,N_13540);
or U15476 (N_15476,N_14059,N_13823);
xnor U15477 (N_15477,N_13544,N_13836);
nor U15478 (N_15478,N_13541,N_13580);
nor U15479 (N_15479,N_13829,N_13981);
nor U15480 (N_15480,N_13787,N_14967);
nor U15481 (N_15481,N_14154,N_13657);
or U15482 (N_15482,N_14161,N_14906);
and U15483 (N_15483,N_14290,N_13640);
or U15484 (N_15484,N_14350,N_14089);
or U15485 (N_15485,N_14129,N_14095);
or U15486 (N_15486,N_13805,N_14975);
or U15487 (N_15487,N_14460,N_14118);
xor U15488 (N_15488,N_14324,N_14056);
and U15489 (N_15489,N_14846,N_14003);
and U15490 (N_15490,N_14885,N_14790);
or U15491 (N_15491,N_14222,N_13964);
nor U15492 (N_15492,N_14467,N_14225);
or U15493 (N_15493,N_14435,N_14755);
and U15494 (N_15494,N_14116,N_13708);
nor U15495 (N_15495,N_14921,N_14812);
and U15496 (N_15496,N_14932,N_14119);
xor U15497 (N_15497,N_14359,N_14360);
xnor U15498 (N_15498,N_14145,N_14011);
xor U15499 (N_15499,N_14337,N_13936);
and U15500 (N_15500,N_14795,N_14964);
xnor U15501 (N_15501,N_14550,N_14972);
or U15502 (N_15502,N_14615,N_14491);
and U15503 (N_15503,N_14690,N_14773);
xor U15504 (N_15504,N_13983,N_14429);
and U15505 (N_15505,N_14772,N_14063);
and U15506 (N_15506,N_14332,N_13834);
nor U15507 (N_15507,N_14573,N_14751);
nand U15508 (N_15508,N_13591,N_13990);
and U15509 (N_15509,N_14892,N_13747);
or U15510 (N_15510,N_14272,N_14368);
xnor U15511 (N_15511,N_14519,N_14448);
nor U15512 (N_15512,N_13503,N_14254);
xnor U15513 (N_15513,N_13552,N_13952);
nor U15514 (N_15514,N_13729,N_14312);
nand U15515 (N_15515,N_14404,N_14887);
or U15516 (N_15516,N_14622,N_14538);
or U15517 (N_15517,N_14373,N_13862);
or U15518 (N_15518,N_14146,N_13879);
nand U15519 (N_15519,N_13826,N_14808);
or U15520 (N_15520,N_14886,N_14841);
xnor U15521 (N_15521,N_14219,N_14919);
xor U15522 (N_15522,N_13846,N_13583);
or U15523 (N_15523,N_14899,N_14481);
xnor U15524 (N_15524,N_14950,N_14092);
xnor U15525 (N_15525,N_14791,N_13755);
nor U15526 (N_15526,N_14701,N_13641);
and U15527 (N_15527,N_14546,N_13526);
nor U15528 (N_15528,N_14937,N_13775);
xnor U15529 (N_15529,N_13965,N_13565);
nor U15530 (N_15530,N_14862,N_13813);
and U15531 (N_15531,N_13859,N_14390);
and U15532 (N_15532,N_14383,N_14606);
or U15533 (N_15533,N_14384,N_13957);
xnor U15534 (N_15534,N_13877,N_13507);
nand U15535 (N_15535,N_14677,N_14621);
and U15536 (N_15536,N_14600,N_14577);
or U15537 (N_15537,N_13637,N_13659);
nand U15538 (N_15538,N_14273,N_14043);
xor U15539 (N_15539,N_14139,N_14211);
or U15540 (N_15540,N_14471,N_13778);
xor U15541 (N_15541,N_13907,N_13831);
and U15542 (N_15542,N_14734,N_14528);
or U15543 (N_15543,N_13949,N_14958);
and U15544 (N_15544,N_14374,N_14520);
or U15545 (N_15545,N_14922,N_14441);
xnor U15546 (N_15546,N_14667,N_14654);
xor U15547 (N_15547,N_13941,N_14533);
nor U15548 (N_15548,N_14526,N_14952);
nand U15549 (N_15549,N_14918,N_14105);
or U15550 (N_15550,N_13603,N_14083);
and U15551 (N_15551,N_14051,N_13621);
or U15552 (N_15552,N_14419,N_13515);
xor U15553 (N_15553,N_14965,N_13638);
and U15554 (N_15554,N_14949,N_13863);
nor U15555 (N_15555,N_13902,N_14261);
xnor U15556 (N_15556,N_13776,N_14915);
nand U15557 (N_15557,N_13645,N_13870);
and U15558 (N_15558,N_14319,N_13524);
xnor U15559 (N_15559,N_14891,N_13835);
nand U15560 (N_15560,N_14388,N_13711);
or U15561 (N_15561,N_14717,N_13690);
and U15562 (N_15562,N_14297,N_14567);
xnor U15563 (N_15563,N_13784,N_14868);
nor U15564 (N_15564,N_13923,N_14160);
or U15565 (N_15565,N_13984,N_14877);
nor U15566 (N_15566,N_14128,N_13607);
or U15567 (N_15567,N_14253,N_14012);
nand U15568 (N_15568,N_14783,N_14039);
and U15569 (N_15569,N_14179,N_14387);
and U15570 (N_15570,N_13861,N_14571);
nand U15571 (N_15571,N_14461,N_14354);
and U15572 (N_15572,N_14512,N_14198);
and U15573 (N_15573,N_13704,N_13726);
or U15574 (N_15574,N_14317,N_14578);
xnor U15575 (N_15575,N_14064,N_14483);
nand U15576 (N_15576,N_13604,N_13858);
and U15577 (N_15577,N_13739,N_13909);
and U15578 (N_15578,N_14149,N_13894);
nand U15579 (N_15579,N_14863,N_14879);
xor U15580 (N_15580,N_14800,N_14850);
or U15581 (N_15581,N_14081,N_14745);
and U15582 (N_15582,N_13808,N_13845);
and U15583 (N_15583,N_14562,N_14326);
xor U15584 (N_15584,N_14133,N_13520);
nand U15585 (N_15585,N_13802,N_14155);
xnor U15586 (N_15586,N_13806,N_14810);
xor U15587 (N_15587,N_13865,N_14666);
and U15588 (N_15588,N_13556,N_14195);
xor U15589 (N_15589,N_14259,N_14839);
or U15590 (N_15590,N_14210,N_13767);
and U15591 (N_15591,N_14168,N_14706);
xnor U15592 (N_15592,N_14604,N_13945);
or U15593 (N_15593,N_13620,N_14714);
nor U15594 (N_15594,N_14295,N_14372);
nand U15595 (N_15595,N_13634,N_13578);
and U15596 (N_15596,N_14788,N_14752);
nor U15597 (N_15597,N_14735,N_14450);
and U15598 (N_15598,N_14010,N_14647);
xor U15599 (N_15599,N_14362,N_14112);
nor U15600 (N_15600,N_14730,N_14416);
or U15601 (N_15601,N_14378,N_13960);
xnor U15602 (N_15602,N_13629,N_14208);
and U15603 (N_15603,N_14518,N_14136);
or U15604 (N_15604,N_14202,N_13574);
nor U15605 (N_15605,N_14732,N_14101);
xor U15606 (N_15606,N_13537,N_14904);
nand U15607 (N_15607,N_14522,N_14913);
nor U15608 (N_15608,N_13763,N_14235);
nand U15609 (N_15609,N_14511,N_13780);
and U15610 (N_15610,N_14980,N_14426);
nand U15611 (N_15611,N_14861,N_14274);
xor U15612 (N_15612,N_14815,N_14474);
nor U15613 (N_15613,N_13691,N_14055);
xor U15614 (N_15614,N_13992,N_14050);
or U15615 (N_15615,N_14333,N_14510);
or U15616 (N_15616,N_13669,N_13500);
or U15617 (N_15617,N_14973,N_13744);
or U15618 (N_15618,N_13884,N_13869);
or U15619 (N_15619,N_14022,N_14027);
xor U15620 (N_15620,N_14542,N_14536);
and U15621 (N_15621,N_14331,N_14768);
and U15622 (N_15622,N_14912,N_14365);
and U15623 (N_15623,N_14514,N_14847);
nand U15624 (N_15624,N_13610,N_13684);
nand U15625 (N_15625,N_14569,N_13619);
or U15626 (N_15626,N_14671,N_13646);
nand U15627 (N_15627,N_14872,N_13571);
nor U15628 (N_15628,N_13939,N_14620);
nand U15629 (N_15629,N_14227,N_14152);
nand U15630 (N_15630,N_13689,N_14375);
and U15631 (N_15631,N_13700,N_14986);
or U15632 (N_15632,N_13511,N_14245);
nand U15633 (N_15633,N_13824,N_13819);
nor U15634 (N_15634,N_14807,N_14894);
and U15635 (N_15635,N_13555,N_14380);
xor U15636 (N_15636,N_14626,N_14113);
or U15637 (N_15637,N_13838,N_14763);
and U15638 (N_15638,N_13589,N_14249);
xor U15639 (N_15639,N_14216,N_14185);
nand U15640 (N_15640,N_14169,N_14458);
nor U15641 (N_15641,N_13840,N_13958);
nor U15642 (N_15642,N_14468,N_13648);
xor U15643 (N_15643,N_14431,N_13914);
nand U15644 (N_15644,N_14473,N_14424);
or U15645 (N_15645,N_14826,N_14171);
and U15646 (N_15646,N_14382,N_14433);
nor U15647 (N_15647,N_14079,N_14648);
nor U15648 (N_15648,N_13532,N_14071);
nor U15649 (N_15649,N_14327,N_14203);
nand U15650 (N_15650,N_13666,N_14409);
nor U15651 (N_15651,N_14057,N_14381);
or U15652 (N_15652,N_13922,N_14330);
nand U15653 (N_15653,N_13878,N_14389);
xor U15654 (N_15654,N_14268,N_14545);
nand U15655 (N_15655,N_14864,N_14422);
and U15656 (N_15656,N_13738,N_14053);
or U15657 (N_15657,N_14924,N_13712);
or U15658 (N_15658,N_14756,N_13502);
xnor U15659 (N_15659,N_13890,N_14140);
xor U15660 (N_15660,N_13988,N_14030);
nor U15661 (N_15661,N_14028,N_14955);
or U15662 (N_15662,N_13504,N_14346);
nand U15663 (N_15663,N_14233,N_14985);
or U15664 (N_15664,N_14554,N_13685);
or U15665 (N_15665,N_13630,N_13967);
nand U15666 (N_15666,N_14798,N_13671);
nor U15667 (N_15667,N_13624,N_14078);
xnor U15668 (N_15668,N_14040,N_14157);
xnor U15669 (N_15669,N_14583,N_14001);
nor U15670 (N_15670,N_14369,N_14640);
nand U15671 (N_15671,N_13746,N_14396);
and U15672 (N_15672,N_14984,N_14002);
nor U15673 (N_15673,N_14890,N_13608);
and U15674 (N_15674,N_14516,N_14142);
nand U15675 (N_15675,N_14281,N_14231);
or U15676 (N_15676,N_14699,N_13963);
nand U15677 (N_15677,N_13735,N_14166);
or U15678 (N_15678,N_14865,N_14436);
nand U15679 (N_15679,N_13851,N_14184);
xnor U15680 (N_15680,N_13937,N_14366);
xor U15681 (N_15681,N_14479,N_13821);
nor U15682 (N_15682,N_13722,N_14843);
and U15683 (N_15683,N_13533,N_14238);
nor U15684 (N_15684,N_14908,N_14813);
nand U15685 (N_15685,N_13582,N_13847);
nor U15686 (N_15686,N_14603,N_14702);
and U15687 (N_15687,N_14386,N_14888);
nand U15688 (N_15688,N_14084,N_14785);
nand U15689 (N_15689,N_14793,N_14085);
or U15690 (N_15690,N_14599,N_13662);
nor U15691 (N_15691,N_14982,N_13760);
nor U15692 (N_15692,N_14007,N_14244);
nand U15693 (N_15693,N_14072,N_14646);
xnor U15694 (N_15694,N_13538,N_14499);
nor U15695 (N_15695,N_13734,N_13654);
xor U15696 (N_15696,N_14819,N_14328);
or U15697 (N_15697,N_14054,N_14060);
and U15698 (N_15698,N_14859,N_14418);
or U15699 (N_15699,N_14994,N_14181);
and U15700 (N_15700,N_14291,N_14023);
and U15701 (N_15701,N_14490,N_14722);
nand U15702 (N_15702,N_13982,N_14668);
nand U15703 (N_15703,N_14408,N_14122);
nor U15704 (N_15704,N_14638,N_13743);
nor U15705 (N_15705,N_14339,N_14938);
or U15706 (N_15706,N_14614,N_14420);
xor U15707 (N_15707,N_14934,N_14110);
nor U15708 (N_15708,N_14838,N_13948);
xor U15709 (N_15709,N_14299,N_14713);
and U15710 (N_15710,N_14019,N_14681);
and U15711 (N_15711,N_14870,N_14270);
or U15712 (N_15712,N_14292,N_14869);
and U15713 (N_15713,N_14935,N_14321);
and U15714 (N_15714,N_13833,N_14970);
xnor U15715 (N_15715,N_13581,N_13714);
nand U15716 (N_15716,N_14916,N_14738);
and U15717 (N_15717,N_13794,N_13611);
nor U15718 (N_15718,N_13759,N_13777);
nand U15719 (N_15719,N_13871,N_14656);
xor U15720 (N_15720,N_14156,N_13995);
and U15721 (N_15721,N_14098,N_14607);
xor U15722 (N_15722,N_14165,N_14279);
or U15723 (N_15723,N_13653,N_13973);
and U15724 (N_15724,N_13947,N_13572);
xnor U15725 (N_15725,N_13606,N_13742);
and U15726 (N_15726,N_14782,N_14680);
and U15727 (N_15727,N_14282,N_14930);
nand U15728 (N_15728,N_14097,N_14325);
nor U15729 (N_15729,N_14309,N_13551);
nor U15730 (N_15730,N_14796,N_14316);
or U15731 (N_15731,N_14945,N_13703);
and U15732 (N_15732,N_14121,N_14901);
and U15733 (N_15733,N_14351,N_13720);
and U15734 (N_15734,N_14006,N_13518);
xnor U15735 (N_15735,N_14032,N_13913);
nand U15736 (N_15736,N_14091,N_14704);
xor U15737 (N_15737,N_14633,N_13751);
xnor U15738 (N_15738,N_13969,N_13803);
and U15739 (N_15739,N_14221,N_14008);
and U15740 (N_15740,N_13667,N_14251);
and U15741 (N_15741,N_14593,N_14944);
nand U15742 (N_15742,N_14109,N_14775);
xor U15743 (N_15743,N_13867,N_14271);
or U15744 (N_15744,N_14655,N_14883);
xor U15745 (N_15745,N_14998,N_14786);
and U15746 (N_15746,N_13543,N_14705);
xnor U15747 (N_15747,N_14805,N_14855);
and U15748 (N_15748,N_14255,N_13554);
or U15749 (N_15749,N_14135,N_13752);
nand U15750 (N_15750,N_14986,N_14833);
and U15751 (N_15751,N_14255,N_14324);
nand U15752 (N_15752,N_14368,N_14718);
xor U15753 (N_15753,N_14734,N_13682);
nor U15754 (N_15754,N_14582,N_14384);
nor U15755 (N_15755,N_13694,N_14141);
nand U15756 (N_15756,N_13739,N_13599);
or U15757 (N_15757,N_14900,N_13934);
nor U15758 (N_15758,N_14403,N_13874);
xnor U15759 (N_15759,N_13695,N_14243);
nor U15760 (N_15760,N_14102,N_13677);
and U15761 (N_15761,N_14286,N_14278);
and U15762 (N_15762,N_13841,N_14596);
xor U15763 (N_15763,N_13931,N_14960);
xnor U15764 (N_15764,N_14439,N_13555);
or U15765 (N_15765,N_14668,N_14600);
and U15766 (N_15766,N_13609,N_14196);
and U15767 (N_15767,N_14338,N_13549);
or U15768 (N_15768,N_13628,N_14454);
nor U15769 (N_15769,N_14032,N_14748);
or U15770 (N_15770,N_14215,N_14993);
nor U15771 (N_15771,N_14601,N_13764);
xor U15772 (N_15772,N_14610,N_14511);
xor U15773 (N_15773,N_14627,N_14177);
and U15774 (N_15774,N_14600,N_14752);
or U15775 (N_15775,N_13728,N_14576);
or U15776 (N_15776,N_13645,N_14727);
xnor U15777 (N_15777,N_14736,N_14250);
and U15778 (N_15778,N_13701,N_14771);
and U15779 (N_15779,N_14273,N_14441);
or U15780 (N_15780,N_14677,N_14525);
and U15781 (N_15781,N_14083,N_13555);
or U15782 (N_15782,N_13813,N_14576);
nand U15783 (N_15783,N_14084,N_13887);
xor U15784 (N_15784,N_14606,N_14695);
and U15785 (N_15785,N_13699,N_14376);
or U15786 (N_15786,N_14100,N_14062);
nand U15787 (N_15787,N_14549,N_13757);
xnor U15788 (N_15788,N_13651,N_14500);
or U15789 (N_15789,N_14208,N_14813);
nor U15790 (N_15790,N_13708,N_13797);
or U15791 (N_15791,N_13582,N_13855);
or U15792 (N_15792,N_14642,N_14481);
and U15793 (N_15793,N_13798,N_13846);
nor U15794 (N_15794,N_14580,N_13718);
nor U15795 (N_15795,N_14830,N_14520);
nor U15796 (N_15796,N_14608,N_14155);
and U15797 (N_15797,N_13507,N_13976);
nor U15798 (N_15798,N_14065,N_14695);
or U15799 (N_15799,N_14340,N_13503);
nand U15800 (N_15800,N_14439,N_14542);
nor U15801 (N_15801,N_14689,N_14927);
or U15802 (N_15802,N_13897,N_14965);
and U15803 (N_15803,N_14569,N_14401);
nand U15804 (N_15804,N_14927,N_13581);
nand U15805 (N_15805,N_14102,N_14459);
nand U15806 (N_15806,N_14690,N_14212);
or U15807 (N_15807,N_14488,N_14691);
or U15808 (N_15808,N_13920,N_14376);
and U15809 (N_15809,N_14751,N_13686);
xor U15810 (N_15810,N_14786,N_13849);
nor U15811 (N_15811,N_14694,N_13770);
and U15812 (N_15812,N_13660,N_13874);
or U15813 (N_15813,N_14974,N_14547);
xnor U15814 (N_15814,N_13788,N_13678);
or U15815 (N_15815,N_14616,N_13729);
xnor U15816 (N_15816,N_13934,N_14293);
and U15817 (N_15817,N_13829,N_14735);
nor U15818 (N_15818,N_13549,N_14657);
and U15819 (N_15819,N_14567,N_14039);
nand U15820 (N_15820,N_14506,N_13900);
xnor U15821 (N_15821,N_14022,N_14145);
or U15822 (N_15822,N_13984,N_13972);
xor U15823 (N_15823,N_13876,N_14059);
nor U15824 (N_15824,N_13794,N_14276);
nor U15825 (N_15825,N_13944,N_13894);
nand U15826 (N_15826,N_14787,N_14706);
nor U15827 (N_15827,N_14821,N_13746);
nor U15828 (N_15828,N_14007,N_13727);
or U15829 (N_15829,N_14185,N_13649);
nand U15830 (N_15830,N_13554,N_13756);
and U15831 (N_15831,N_14854,N_14824);
nand U15832 (N_15832,N_13802,N_14260);
and U15833 (N_15833,N_13915,N_13627);
nand U15834 (N_15834,N_14247,N_13721);
and U15835 (N_15835,N_14218,N_14026);
and U15836 (N_15836,N_14804,N_14754);
xnor U15837 (N_15837,N_14515,N_14938);
or U15838 (N_15838,N_14864,N_14902);
xnor U15839 (N_15839,N_14754,N_14278);
or U15840 (N_15840,N_14958,N_13759);
nor U15841 (N_15841,N_14366,N_14050);
or U15842 (N_15842,N_14583,N_14692);
xnor U15843 (N_15843,N_14138,N_14980);
and U15844 (N_15844,N_13889,N_13609);
xnor U15845 (N_15845,N_14814,N_13668);
nor U15846 (N_15846,N_14235,N_14139);
nand U15847 (N_15847,N_13907,N_14125);
xnor U15848 (N_15848,N_13847,N_14738);
nand U15849 (N_15849,N_14406,N_14283);
nor U15850 (N_15850,N_13848,N_14472);
nand U15851 (N_15851,N_14401,N_14408);
nor U15852 (N_15852,N_14843,N_14628);
or U15853 (N_15853,N_14622,N_14908);
xor U15854 (N_15854,N_14957,N_13502);
xor U15855 (N_15855,N_14932,N_14701);
and U15856 (N_15856,N_14306,N_14981);
and U15857 (N_15857,N_14119,N_13888);
xnor U15858 (N_15858,N_13720,N_13610);
and U15859 (N_15859,N_14181,N_14330);
nor U15860 (N_15860,N_14503,N_13586);
nor U15861 (N_15861,N_14499,N_13568);
or U15862 (N_15862,N_14903,N_14505);
nand U15863 (N_15863,N_13523,N_14371);
xnor U15864 (N_15864,N_13985,N_14303);
and U15865 (N_15865,N_13614,N_14350);
or U15866 (N_15866,N_14214,N_14396);
nor U15867 (N_15867,N_14517,N_13543);
xnor U15868 (N_15868,N_13589,N_14520);
nand U15869 (N_15869,N_14163,N_14077);
and U15870 (N_15870,N_14665,N_14761);
and U15871 (N_15871,N_13995,N_14388);
nand U15872 (N_15872,N_14003,N_13887);
or U15873 (N_15873,N_14433,N_14829);
nor U15874 (N_15874,N_14319,N_14223);
xnor U15875 (N_15875,N_14073,N_14940);
xor U15876 (N_15876,N_14751,N_14936);
or U15877 (N_15877,N_14599,N_13962);
xor U15878 (N_15878,N_14499,N_13974);
nand U15879 (N_15879,N_14373,N_13858);
nand U15880 (N_15880,N_13791,N_14184);
nor U15881 (N_15881,N_13872,N_14831);
xor U15882 (N_15882,N_13842,N_14148);
nand U15883 (N_15883,N_13709,N_13889);
nor U15884 (N_15884,N_13831,N_14105);
and U15885 (N_15885,N_13843,N_14132);
nand U15886 (N_15886,N_14500,N_14098);
nor U15887 (N_15887,N_13952,N_14503);
nand U15888 (N_15888,N_14633,N_13684);
nor U15889 (N_15889,N_13947,N_14506);
and U15890 (N_15890,N_14652,N_14374);
and U15891 (N_15891,N_14259,N_13772);
or U15892 (N_15892,N_14091,N_14619);
nor U15893 (N_15893,N_13955,N_14982);
or U15894 (N_15894,N_14423,N_13635);
xnor U15895 (N_15895,N_14859,N_13829);
nand U15896 (N_15896,N_14356,N_14889);
xor U15897 (N_15897,N_14258,N_14749);
nor U15898 (N_15898,N_13989,N_13559);
nand U15899 (N_15899,N_14005,N_14341);
and U15900 (N_15900,N_14141,N_14205);
and U15901 (N_15901,N_13655,N_14202);
nand U15902 (N_15902,N_14679,N_13595);
or U15903 (N_15903,N_14222,N_14987);
xnor U15904 (N_15904,N_13641,N_14888);
xor U15905 (N_15905,N_14996,N_13990);
xnor U15906 (N_15906,N_14115,N_13770);
nor U15907 (N_15907,N_14556,N_14014);
or U15908 (N_15908,N_14036,N_13927);
nand U15909 (N_15909,N_14069,N_14507);
or U15910 (N_15910,N_14473,N_13559);
nand U15911 (N_15911,N_14492,N_14108);
xor U15912 (N_15912,N_14861,N_14425);
nor U15913 (N_15913,N_13802,N_14148);
and U15914 (N_15914,N_13508,N_13961);
nand U15915 (N_15915,N_14253,N_14463);
and U15916 (N_15916,N_14538,N_14396);
xor U15917 (N_15917,N_13920,N_13998);
or U15918 (N_15918,N_14533,N_13886);
or U15919 (N_15919,N_14074,N_14693);
nor U15920 (N_15920,N_14265,N_14103);
or U15921 (N_15921,N_13937,N_14560);
nand U15922 (N_15922,N_13684,N_14604);
or U15923 (N_15923,N_14326,N_14300);
xnor U15924 (N_15924,N_14635,N_14205);
and U15925 (N_15925,N_13897,N_14831);
and U15926 (N_15926,N_13848,N_13692);
or U15927 (N_15927,N_14695,N_13905);
and U15928 (N_15928,N_14539,N_14781);
or U15929 (N_15929,N_14381,N_13626);
and U15930 (N_15930,N_13893,N_14353);
xnor U15931 (N_15931,N_13882,N_14440);
and U15932 (N_15932,N_14115,N_13572);
nand U15933 (N_15933,N_14979,N_13629);
nor U15934 (N_15934,N_14713,N_14572);
nor U15935 (N_15935,N_14615,N_14071);
nor U15936 (N_15936,N_14338,N_13892);
or U15937 (N_15937,N_13941,N_14840);
or U15938 (N_15938,N_14014,N_14664);
and U15939 (N_15939,N_14805,N_13652);
nand U15940 (N_15940,N_14469,N_14325);
xor U15941 (N_15941,N_13876,N_14110);
nand U15942 (N_15942,N_14191,N_14636);
nand U15943 (N_15943,N_14762,N_13634);
nor U15944 (N_15944,N_14558,N_13759);
and U15945 (N_15945,N_14208,N_14421);
xor U15946 (N_15946,N_13728,N_13901);
or U15947 (N_15947,N_13576,N_13557);
xnor U15948 (N_15948,N_13962,N_14474);
nand U15949 (N_15949,N_14106,N_13956);
nand U15950 (N_15950,N_13885,N_14497);
xnor U15951 (N_15951,N_14695,N_14155);
nand U15952 (N_15952,N_14039,N_13590);
nand U15953 (N_15953,N_13803,N_14244);
xor U15954 (N_15954,N_14550,N_13517);
nand U15955 (N_15955,N_13638,N_13878);
nand U15956 (N_15956,N_14948,N_14212);
nand U15957 (N_15957,N_14955,N_14884);
nand U15958 (N_15958,N_14294,N_14904);
nand U15959 (N_15959,N_14795,N_13874);
or U15960 (N_15960,N_13946,N_13646);
nand U15961 (N_15961,N_14396,N_14884);
xnor U15962 (N_15962,N_14319,N_14536);
or U15963 (N_15963,N_14052,N_14482);
nor U15964 (N_15964,N_13775,N_13681);
or U15965 (N_15965,N_13527,N_14819);
nor U15966 (N_15966,N_13541,N_14255);
and U15967 (N_15967,N_14158,N_14446);
nor U15968 (N_15968,N_14147,N_13592);
and U15969 (N_15969,N_14697,N_14122);
or U15970 (N_15970,N_14058,N_14304);
xor U15971 (N_15971,N_14216,N_14982);
or U15972 (N_15972,N_14792,N_13648);
nand U15973 (N_15973,N_14564,N_14706);
nand U15974 (N_15974,N_14409,N_14666);
nand U15975 (N_15975,N_13632,N_13734);
nor U15976 (N_15976,N_14854,N_13983);
xor U15977 (N_15977,N_13866,N_14265);
nor U15978 (N_15978,N_13903,N_14750);
xor U15979 (N_15979,N_14521,N_13775);
and U15980 (N_15980,N_13609,N_14031);
and U15981 (N_15981,N_14229,N_14366);
nand U15982 (N_15982,N_13997,N_14197);
nor U15983 (N_15983,N_14370,N_13639);
nand U15984 (N_15984,N_14435,N_14523);
xor U15985 (N_15985,N_14919,N_14536);
and U15986 (N_15986,N_13651,N_14085);
or U15987 (N_15987,N_14212,N_13813);
nor U15988 (N_15988,N_13905,N_13787);
xnor U15989 (N_15989,N_13673,N_14433);
xor U15990 (N_15990,N_13543,N_14212);
and U15991 (N_15991,N_14586,N_14746);
nor U15992 (N_15992,N_13580,N_13801);
and U15993 (N_15993,N_14428,N_14348);
or U15994 (N_15994,N_14538,N_14945);
nand U15995 (N_15995,N_14210,N_13893);
xor U15996 (N_15996,N_14234,N_14341);
and U15997 (N_15997,N_14661,N_14627);
nor U15998 (N_15998,N_13954,N_13647);
or U15999 (N_15999,N_13895,N_13728);
or U16000 (N_16000,N_14521,N_14799);
nor U16001 (N_16001,N_14226,N_14102);
or U16002 (N_16002,N_14298,N_13745);
or U16003 (N_16003,N_14807,N_14421);
nand U16004 (N_16004,N_14097,N_14800);
xor U16005 (N_16005,N_14532,N_14780);
nor U16006 (N_16006,N_14249,N_14439);
nand U16007 (N_16007,N_14861,N_14726);
and U16008 (N_16008,N_13778,N_13788);
xor U16009 (N_16009,N_14057,N_14918);
xnor U16010 (N_16010,N_13952,N_14259);
xor U16011 (N_16011,N_14353,N_13761);
and U16012 (N_16012,N_14628,N_14811);
nand U16013 (N_16013,N_14614,N_14644);
nor U16014 (N_16014,N_14912,N_14371);
or U16015 (N_16015,N_13903,N_14699);
nand U16016 (N_16016,N_13899,N_13681);
nand U16017 (N_16017,N_14255,N_14942);
nand U16018 (N_16018,N_13514,N_14199);
and U16019 (N_16019,N_14585,N_14880);
xnor U16020 (N_16020,N_14509,N_14276);
nand U16021 (N_16021,N_14420,N_14856);
xor U16022 (N_16022,N_14652,N_14190);
or U16023 (N_16023,N_14482,N_14675);
nor U16024 (N_16024,N_14633,N_14413);
or U16025 (N_16025,N_13841,N_14588);
and U16026 (N_16026,N_14858,N_13818);
and U16027 (N_16027,N_13652,N_13758);
nand U16028 (N_16028,N_14837,N_14767);
or U16029 (N_16029,N_14224,N_14679);
nand U16030 (N_16030,N_14488,N_14659);
and U16031 (N_16031,N_13577,N_14321);
xnor U16032 (N_16032,N_14755,N_14429);
nand U16033 (N_16033,N_14514,N_14090);
xnor U16034 (N_16034,N_13657,N_13807);
nor U16035 (N_16035,N_14004,N_14036);
nand U16036 (N_16036,N_14559,N_14953);
or U16037 (N_16037,N_13701,N_14132);
or U16038 (N_16038,N_13793,N_13986);
and U16039 (N_16039,N_14858,N_14197);
nor U16040 (N_16040,N_13532,N_14625);
or U16041 (N_16041,N_13744,N_14525);
and U16042 (N_16042,N_14656,N_14924);
nor U16043 (N_16043,N_14986,N_14046);
and U16044 (N_16044,N_14375,N_14589);
nor U16045 (N_16045,N_13900,N_14799);
or U16046 (N_16046,N_14686,N_13869);
and U16047 (N_16047,N_14116,N_14528);
xnor U16048 (N_16048,N_13822,N_14866);
nor U16049 (N_16049,N_14262,N_14624);
nand U16050 (N_16050,N_14110,N_13705);
nor U16051 (N_16051,N_14790,N_14706);
nor U16052 (N_16052,N_14251,N_13684);
nor U16053 (N_16053,N_13645,N_13998);
and U16054 (N_16054,N_14927,N_14604);
and U16055 (N_16055,N_13723,N_14286);
or U16056 (N_16056,N_14988,N_14902);
and U16057 (N_16057,N_14896,N_13752);
nand U16058 (N_16058,N_14622,N_13849);
and U16059 (N_16059,N_13959,N_13729);
xor U16060 (N_16060,N_13575,N_13773);
or U16061 (N_16061,N_14716,N_14066);
nand U16062 (N_16062,N_13785,N_14913);
nand U16063 (N_16063,N_13760,N_14753);
nor U16064 (N_16064,N_14137,N_14429);
nor U16065 (N_16065,N_14674,N_13516);
and U16066 (N_16066,N_13656,N_14969);
or U16067 (N_16067,N_14572,N_13562);
nand U16068 (N_16068,N_14470,N_14571);
and U16069 (N_16069,N_13513,N_14894);
or U16070 (N_16070,N_14969,N_14382);
nand U16071 (N_16071,N_13905,N_14598);
or U16072 (N_16072,N_13523,N_14703);
or U16073 (N_16073,N_14843,N_14442);
nor U16074 (N_16074,N_14900,N_14893);
xor U16075 (N_16075,N_13615,N_13792);
and U16076 (N_16076,N_13577,N_13778);
nand U16077 (N_16077,N_13624,N_14907);
nand U16078 (N_16078,N_13973,N_14329);
nor U16079 (N_16079,N_14667,N_14296);
or U16080 (N_16080,N_13580,N_14235);
or U16081 (N_16081,N_14665,N_14947);
and U16082 (N_16082,N_14261,N_14725);
nand U16083 (N_16083,N_13639,N_13787);
nand U16084 (N_16084,N_13822,N_13980);
nor U16085 (N_16085,N_13938,N_13697);
nand U16086 (N_16086,N_14372,N_14134);
and U16087 (N_16087,N_13590,N_14430);
nor U16088 (N_16088,N_14125,N_14415);
nor U16089 (N_16089,N_13743,N_13827);
and U16090 (N_16090,N_14565,N_13863);
or U16091 (N_16091,N_13897,N_14874);
nand U16092 (N_16092,N_13583,N_14269);
nand U16093 (N_16093,N_14473,N_14976);
nand U16094 (N_16094,N_14089,N_14924);
nor U16095 (N_16095,N_14362,N_14791);
xnor U16096 (N_16096,N_14607,N_14497);
nor U16097 (N_16097,N_13616,N_14594);
nand U16098 (N_16098,N_13778,N_13705);
xnor U16099 (N_16099,N_14518,N_13664);
or U16100 (N_16100,N_14828,N_14024);
nor U16101 (N_16101,N_14973,N_14786);
or U16102 (N_16102,N_14756,N_14492);
nand U16103 (N_16103,N_14244,N_14342);
nand U16104 (N_16104,N_13908,N_14449);
xor U16105 (N_16105,N_14562,N_13913);
and U16106 (N_16106,N_14722,N_14560);
and U16107 (N_16107,N_14300,N_14587);
nor U16108 (N_16108,N_13915,N_14687);
nand U16109 (N_16109,N_14110,N_13670);
nor U16110 (N_16110,N_14485,N_14107);
xnor U16111 (N_16111,N_14361,N_14532);
and U16112 (N_16112,N_13811,N_14299);
or U16113 (N_16113,N_14338,N_14954);
or U16114 (N_16114,N_13780,N_14382);
nor U16115 (N_16115,N_14476,N_14095);
or U16116 (N_16116,N_14223,N_14978);
nor U16117 (N_16117,N_14847,N_13939);
nor U16118 (N_16118,N_13508,N_13678);
xnor U16119 (N_16119,N_14874,N_13754);
or U16120 (N_16120,N_14573,N_14205);
and U16121 (N_16121,N_14790,N_13951);
xor U16122 (N_16122,N_13590,N_13730);
and U16123 (N_16123,N_14687,N_13511);
or U16124 (N_16124,N_13685,N_14674);
nor U16125 (N_16125,N_14581,N_13787);
and U16126 (N_16126,N_14820,N_14768);
or U16127 (N_16127,N_14088,N_13736);
nand U16128 (N_16128,N_13732,N_14904);
and U16129 (N_16129,N_14513,N_13666);
nor U16130 (N_16130,N_14017,N_14678);
xnor U16131 (N_16131,N_14250,N_13521);
xnor U16132 (N_16132,N_14976,N_13595);
nor U16133 (N_16133,N_14557,N_13567);
or U16134 (N_16134,N_14745,N_13545);
or U16135 (N_16135,N_14262,N_14381);
and U16136 (N_16136,N_13889,N_14008);
and U16137 (N_16137,N_13518,N_14678);
xnor U16138 (N_16138,N_14224,N_14635);
or U16139 (N_16139,N_14435,N_14429);
nor U16140 (N_16140,N_14942,N_13508);
and U16141 (N_16141,N_14479,N_13873);
and U16142 (N_16142,N_14719,N_14170);
or U16143 (N_16143,N_14357,N_14856);
nor U16144 (N_16144,N_14956,N_14740);
nand U16145 (N_16145,N_14923,N_13889);
and U16146 (N_16146,N_13786,N_14079);
and U16147 (N_16147,N_14099,N_13963);
xor U16148 (N_16148,N_14238,N_14169);
xnor U16149 (N_16149,N_14522,N_14926);
and U16150 (N_16150,N_14757,N_14525);
nand U16151 (N_16151,N_14011,N_14891);
or U16152 (N_16152,N_14593,N_14956);
nor U16153 (N_16153,N_14466,N_14480);
nor U16154 (N_16154,N_14868,N_14097);
nor U16155 (N_16155,N_14528,N_13870);
and U16156 (N_16156,N_14286,N_14051);
or U16157 (N_16157,N_14211,N_13771);
nor U16158 (N_16158,N_14662,N_14341);
or U16159 (N_16159,N_14936,N_14526);
xnor U16160 (N_16160,N_14015,N_13675);
xnor U16161 (N_16161,N_14234,N_14845);
nor U16162 (N_16162,N_13590,N_14511);
and U16163 (N_16163,N_14165,N_14013);
nor U16164 (N_16164,N_13508,N_13631);
and U16165 (N_16165,N_14627,N_14581);
nand U16166 (N_16166,N_14941,N_13880);
xor U16167 (N_16167,N_14910,N_14286);
nor U16168 (N_16168,N_13576,N_14085);
nand U16169 (N_16169,N_14798,N_13895);
xor U16170 (N_16170,N_13630,N_14803);
or U16171 (N_16171,N_14271,N_14144);
nor U16172 (N_16172,N_14120,N_14836);
nor U16173 (N_16173,N_14970,N_14257);
nand U16174 (N_16174,N_14506,N_14202);
nand U16175 (N_16175,N_14067,N_13656);
xnor U16176 (N_16176,N_13543,N_14740);
and U16177 (N_16177,N_14822,N_14256);
or U16178 (N_16178,N_14702,N_14827);
xnor U16179 (N_16179,N_14276,N_14190);
nand U16180 (N_16180,N_13643,N_14241);
nor U16181 (N_16181,N_14485,N_14501);
or U16182 (N_16182,N_13730,N_14770);
xnor U16183 (N_16183,N_14877,N_14147);
nand U16184 (N_16184,N_13902,N_13690);
or U16185 (N_16185,N_14594,N_14494);
xor U16186 (N_16186,N_14785,N_14927);
and U16187 (N_16187,N_14153,N_14859);
or U16188 (N_16188,N_14621,N_14929);
nor U16189 (N_16189,N_13966,N_14181);
and U16190 (N_16190,N_14583,N_14084);
nor U16191 (N_16191,N_14194,N_13756);
xor U16192 (N_16192,N_13665,N_14498);
nor U16193 (N_16193,N_14146,N_13701);
or U16194 (N_16194,N_14749,N_13562);
or U16195 (N_16195,N_14512,N_14962);
and U16196 (N_16196,N_14057,N_14513);
or U16197 (N_16197,N_13636,N_14939);
and U16198 (N_16198,N_13602,N_13679);
or U16199 (N_16199,N_14208,N_13682);
xnor U16200 (N_16200,N_13801,N_14850);
xnor U16201 (N_16201,N_14740,N_14395);
nor U16202 (N_16202,N_14315,N_13851);
and U16203 (N_16203,N_14088,N_14081);
and U16204 (N_16204,N_14290,N_14147);
nand U16205 (N_16205,N_14205,N_14770);
xnor U16206 (N_16206,N_14193,N_14339);
nor U16207 (N_16207,N_14346,N_14918);
or U16208 (N_16208,N_14268,N_14290);
xor U16209 (N_16209,N_14226,N_14622);
xor U16210 (N_16210,N_14770,N_14152);
or U16211 (N_16211,N_13649,N_14526);
xnor U16212 (N_16212,N_14478,N_14783);
nor U16213 (N_16213,N_13641,N_13900);
xnor U16214 (N_16214,N_14399,N_13924);
or U16215 (N_16215,N_14272,N_14216);
nand U16216 (N_16216,N_14522,N_14908);
xnor U16217 (N_16217,N_14866,N_14413);
nor U16218 (N_16218,N_14410,N_14987);
xor U16219 (N_16219,N_14578,N_14107);
nand U16220 (N_16220,N_14129,N_13951);
and U16221 (N_16221,N_13719,N_14948);
xnor U16222 (N_16222,N_14680,N_13927);
nor U16223 (N_16223,N_13724,N_14871);
nand U16224 (N_16224,N_14220,N_13680);
nor U16225 (N_16225,N_13573,N_14393);
nand U16226 (N_16226,N_13799,N_13547);
nand U16227 (N_16227,N_14616,N_14468);
or U16228 (N_16228,N_14798,N_13699);
nand U16229 (N_16229,N_13918,N_13603);
nor U16230 (N_16230,N_14443,N_13733);
xor U16231 (N_16231,N_14282,N_13717);
nand U16232 (N_16232,N_14902,N_14097);
nor U16233 (N_16233,N_14340,N_13901);
or U16234 (N_16234,N_14966,N_13533);
or U16235 (N_16235,N_13713,N_14990);
xnor U16236 (N_16236,N_14192,N_14642);
and U16237 (N_16237,N_14770,N_14747);
nor U16238 (N_16238,N_13783,N_14274);
or U16239 (N_16239,N_14297,N_14963);
or U16240 (N_16240,N_14738,N_14255);
or U16241 (N_16241,N_14720,N_14740);
nor U16242 (N_16242,N_14028,N_14912);
nand U16243 (N_16243,N_13995,N_13684);
and U16244 (N_16244,N_13509,N_14648);
or U16245 (N_16245,N_13804,N_14988);
and U16246 (N_16246,N_14932,N_14618);
nor U16247 (N_16247,N_14464,N_14585);
or U16248 (N_16248,N_13965,N_13923);
nor U16249 (N_16249,N_14489,N_14311);
xor U16250 (N_16250,N_14888,N_13796);
xor U16251 (N_16251,N_13845,N_13507);
xor U16252 (N_16252,N_14160,N_13715);
nand U16253 (N_16253,N_14936,N_13751);
and U16254 (N_16254,N_13557,N_13924);
nor U16255 (N_16255,N_14443,N_14870);
xnor U16256 (N_16256,N_13948,N_13757);
nand U16257 (N_16257,N_13595,N_13852);
nor U16258 (N_16258,N_13926,N_13679);
xor U16259 (N_16259,N_13790,N_14682);
or U16260 (N_16260,N_14886,N_13562);
and U16261 (N_16261,N_14410,N_13877);
or U16262 (N_16262,N_13961,N_13683);
nor U16263 (N_16263,N_14501,N_14656);
or U16264 (N_16264,N_14877,N_13735);
nor U16265 (N_16265,N_14627,N_14260);
and U16266 (N_16266,N_13553,N_14837);
nand U16267 (N_16267,N_14314,N_13534);
and U16268 (N_16268,N_14303,N_14351);
nor U16269 (N_16269,N_14346,N_13686);
and U16270 (N_16270,N_13900,N_14327);
xor U16271 (N_16271,N_13583,N_13749);
and U16272 (N_16272,N_13802,N_14038);
and U16273 (N_16273,N_14799,N_14697);
or U16274 (N_16274,N_14514,N_13773);
and U16275 (N_16275,N_14086,N_14011);
nor U16276 (N_16276,N_14916,N_13956);
and U16277 (N_16277,N_14602,N_14171);
xnor U16278 (N_16278,N_13568,N_14727);
xor U16279 (N_16279,N_14352,N_13810);
nand U16280 (N_16280,N_14021,N_14553);
nor U16281 (N_16281,N_14788,N_14357);
nand U16282 (N_16282,N_14027,N_13850);
nor U16283 (N_16283,N_13881,N_14454);
and U16284 (N_16284,N_13645,N_14111);
and U16285 (N_16285,N_14598,N_14034);
nand U16286 (N_16286,N_13538,N_14259);
nand U16287 (N_16287,N_14499,N_14934);
nand U16288 (N_16288,N_13517,N_13911);
and U16289 (N_16289,N_14255,N_14591);
nand U16290 (N_16290,N_13974,N_13772);
nand U16291 (N_16291,N_13865,N_14824);
nand U16292 (N_16292,N_13562,N_13602);
nand U16293 (N_16293,N_14706,N_14444);
nor U16294 (N_16294,N_13686,N_14848);
xor U16295 (N_16295,N_14415,N_13637);
nand U16296 (N_16296,N_14267,N_14404);
xnor U16297 (N_16297,N_14200,N_13956);
nor U16298 (N_16298,N_13976,N_14899);
and U16299 (N_16299,N_13642,N_14316);
or U16300 (N_16300,N_14888,N_14327);
nand U16301 (N_16301,N_14839,N_13888);
or U16302 (N_16302,N_13605,N_13855);
or U16303 (N_16303,N_13897,N_13513);
nor U16304 (N_16304,N_13520,N_14680);
xnor U16305 (N_16305,N_14235,N_13794);
nor U16306 (N_16306,N_13954,N_14435);
nand U16307 (N_16307,N_14425,N_14036);
xnor U16308 (N_16308,N_14936,N_13561);
xnor U16309 (N_16309,N_14431,N_14175);
nand U16310 (N_16310,N_13996,N_14190);
and U16311 (N_16311,N_14892,N_14893);
or U16312 (N_16312,N_13775,N_14038);
or U16313 (N_16313,N_14683,N_14763);
and U16314 (N_16314,N_14811,N_14079);
or U16315 (N_16315,N_14685,N_14335);
xor U16316 (N_16316,N_14766,N_14532);
or U16317 (N_16317,N_13563,N_13626);
and U16318 (N_16318,N_13551,N_14304);
and U16319 (N_16319,N_14959,N_14223);
nor U16320 (N_16320,N_14572,N_13706);
nor U16321 (N_16321,N_14161,N_13769);
nand U16322 (N_16322,N_13625,N_14003);
or U16323 (N_16323,N_14369,N_14053);
or U16324 (N_16324,N_14415,N_14861);
nand U16325 (N_16325,N_13621,N_13689);
or U16326 (N_16326,N_14940,N_13580);
or U16327 (N_16327,N_14619,N_14138);
nand U16328 (N_16328,N_13715,N_14777);
nor U16329 (N_16329,N_13875,N_14379);
xor U16330 (N_16330,N_14886,N_14706);
nand U16331 (N_16331,N_14841,N_14792);
or U16332 (N_16332,N_13982,N_14837);
or U16333 (N_16333,N_13547,N_13961);
nor U16334 (N_16334,N_14302,N_14435);
nor U16335 (N_16335,N_13555,N_14777);
xnor U16336 (N_16336,N_13659,N_14565);
xnor U16337 (N_16337,N_13803,N_14665);
or U16338 (N_16338,N_14627,N_13579);
nand U16339 (N_16339,N_14444,N_14576);
xor U16340 (N_16340,N_14130,N_13583);
or U16341 (N_16341,N_13895,N_13785);
nand U16342 (N_16342,N_14608,N_13773);
or U16343 (N_16343,N_14357,N_13837);
or U16344 (N_16344,N_13929,N_13742);
and U16345 (N_16345,N_14920,N_13897);
xnor U16346 (N_16346,N_13954,N_14327);
nor U16347 (N_16347,N_14197,N_13870);
xor U16348 (N_16348,N_14242,N_13599);
nand U16349 (N_16349,N_14315,N_14638);
nor U16350 (N_16350,N_14844,N_14634);
nor U16351 (N_16351,N_13941,N_14076);
nor U16352 (N_16352,N_14542,N_13642);
nor U16353 (N_16353,N_14830,N_13778);
nor U16354 (N_16354,N_14217,N_13931);
nor U16355 (N_16355,N_13761,N_14258);
nor U16356 (N_16356,N_14728,N_14025);
and U16357 (N_16357,N_14895,N_14800);
nor U16358 (N_16358,N_13606,N_14436);
nor U16359 (N_16359,N_13674,N_14075);
or U16360 (N_16360,N_13745,N_14321);
nor U16361 (N_16361,N_14018,N_14953);
nor U16362 (N_16362,N_14692,N_14908);
or U16363 (N_16363,N_14325,N_14414);
and U16364 (N_16364,N_14692,N_14375);
nor U16365 (N_16365,N_13595,N_13845);
xor U16366 (N_16366,N_14083,N_14972);
xnor U16367 (N_16367,N_14001,N_13644);
or U16368 (N_16368,N_14533,N_14653);
xor U16369 (N_16369,N_14980,N_13609);
and U16370 (N_16370,N_13663,N_14522);
nand U16371 (N_16371,N_14136,N_13831);
nor U16372 (N_16372,N_14040,N_14075);
nor U16373 (N_16373,N_13923,N_13733);
xnor U16374 (N_16374,N_14355,N_13762);
nor U16375 (N_16375,N_13660,N_14975);
nand U16376 (N_16376,N_14819,N_13984);
nand U16377 (N_16377,N_14265,N_13557);
nand U16378 (N_16378,N_13882,N_14848);
xnor U16379 (N_16379,N_14087,N_13826);
nand U16380 (N_16380,N_14323,N_14115);
or U16381 (N_16381,N_14168,N_13741);
or U16382 (N_16382,N_14398,N_13890);
xnor U16383 (N_16383,N_14626,N_13830);
nor U16384 (N_16384,N_14222,N_14449);
xnor U16385 (N_16385,N_14352,N_14934);
xor U16386 (N_16386,N_14106,N_13899);
nor U16387 (N_16387,N_14086,N_13783);
and U16388 (N_16388,N_14485,N_13776);
or U16389 (N_16389,N_14488,N_14471);
nand U16390 (N_16390,N_14951,N_14514);
nor U16391 (N_16391,N_14461,N_14255);
xor U16392 (N_16392,N_14824,N_14500);
nand U16393 (N_16393,N_14967,N_14195);
nand U16394 (N_16394,N_14855,N_14872);
xnor U16395 (N_16395,N_13744,N_14059);
or U16396 (N_16396,N_13847,N_13763);
xor U16397 (N_16397,N_13972,N_13883);
nand U16398 (N_16398,N_13946,N_14158);
nand U16399 (N_16399,N_14672,N_14967);
nand U16400 (N_16400,N_14552,N_13570);
nand U16401 (N_16401,N_13652,N_14398);
nand U16402 (N_16402,N_13822,N_14673);
or U16403 (N_16403,N_14505,N_14149);
nor U16404 (N_16404,N_13932,N_14192);
nor U16405 (N_16405,N_14714,N_13789);
and U16406 (N_16406,N_14081,N_14504);
nand U16407 (N_16407,N_14477,N_13785);
xnor U16408 (N_16408,N_14689,N_14845);
and U16409 (N_16409,N_13880,N_14053);
or U16410 (N_16410,N_14745,N_14568);
nor U16411 (N_16411,N_14775,N_13607);
or U16412 (N_16412,N_14856,N_13834);
nand U16413 (N_16413,N_14486,N_14721);
nor U16414 (N_16414,N_13922,N_14766);
xnor U16415 (N_16415,N_14484,N_13507);
xnor U16416 (N_16416,N_14684,N_13673);
xor U16417 (N_16417,N_13537,N_14045);
or U16418 (N_16418,N_14778,N_13772);
xor U16419 (N_16419,N_14899,N_14308);
xor U16420 (N_16420,N_14282,N_14339);
and U16421 (N_16421,N_14905,N_14427);
nand U16422 (N_16422,N_14996,N_14325);
or U16423 (N_16423,N_13519,N_14517);
nand U16424 (N_16424,N_14216,N_14124);
and U16425 (N_16425,N_14327,N_14898);
xnor U16426 (N_16426,N_14681,N_13844);
nor U16427 (N_16427,N_14611,N_14851);
or U16428 (N_16428,N_14926,N_13987);
or U16429 (N_16429,N_13580,N_14322);
nand U16430 (N_16430,N_14627,N_14384);
or U16431 (N_16431,N_14296,N_14200);
and U16432 (N_16432,N_13859,N_14913);
xor U16433 (N_16433,N_14056,N_14127);
nor U16434 (N_16434,N_13552,N_13741);
xnor U16435 (N_16435,N_14085,N_14000);
nand U16436 (N_16436,N_14338,N_13975);
xnor U16437 (N_16437,N_14588,N_14439);
xnor U16438 (N_16438,N_14742,N_13705);
or U16439 (N_16439,N_14087,N_14394);
nor U16440 (N_16440,N_13792,N_13856);
or U16441 (N_16441,N_13553,N_13892);
nor U16442 (N_16442,N_14079,N_14244);
xnor U16443 (N_16443,N_13716,N_14726);
or U16444 (N_16444,N_14041,N_13839);
and U16445 (N_16445,N_14294,N_14671);
nand U16446 (N_16446,N_13954,N_14861);
and U16447 (N_16447,N_14560,N_14307);
xor U16448 (N_16448,N_14282,N_14731);
nor U16449 (N_16449,N_14772,N_14508);
nand U16450 (N_16450,N_14357,N_14980);
xor U16451 (N_16451,N_14963,N_14597);
nand U16452 (N_16452,N_14285,N_14916);
xor U16453 (N_16453,N_14061,N_14583);
and U16454 (N_16454,N_14828,N_14215);
and U16455 (N_16455,N_14392,N_14586);
and U16456 (N_16456,N_14126,N_14487);
xor U16457 (N_16457,N_13605,N_13933);
and U16458 (N_16458,N_14365,N_14161);
xor U16459 (N_16459,N_13627,N_14566);
or U16460 (N_16460,N_13711,N_14301);
nand U16461 (N_16461,N_13568,N_13527);
nor U16462 (N_16462,N_13585,N_13573);
nor U16463 (N_16463,N_13643,N_14304);
nand U16464 (N_16464,N_13587,N_13570);
or U16465 (N_16465,N_14383,N_14348);
nand U16466 (N_16466,N_14213,N_13567);
or U16467 (N_16467,N_13524,N_14090);
and U16468 (N_16468,N_14852,N_14505);
xor U16469 (N_16469,N_13889,N_14826);
and U16470 (N_16470,N_14120,N_13766);
nand U16471 (N_16471,N_14112,N_14577);
xnor U16472 (N_16472,N_14760,N_14405);
xnor U16473 (N_16473,N_14809,N_13728);
or U16474 (N_16474,N_14610,N_14791);
or U16475 (N_16475,N_13538,N_14506);
and U16476 (N_16476,N_14734,N_13519);
nand U16477 (N_16477,N_13610,N_14048);
nor U16478 (N_16478,N_13741,N_13577);
nand U16479 (N_16479,N_14214,N_14639);
or U16480 (N_16480,N_14340,N_14005);
nor U16481 (N_16481,N_14789,N_14997);
or U16482 (N_16482,N_14190,N_14803);
or U16483 (N_16483,N_14053,N_14293);
xor U16484 (N_16484,N_14775,N_13602);
or U16485 (N_16485,N_14902,N_14523);
xnor U16486 (N_16486,N_14319,N_14279);
and U16487 (N_16487,N_14142,N_13699);
and U16488 (N_16488,N_14018,N_14913);
xor U16489 (N_16489,N_14735,N_14305);
or U16490 (N_16490,N_14667,N_13953);
xnor U16491 (N_16491,N_14797,N_14576);
and U16492 (N_16492,N_14279,N_13547);
nor U16493 (N_16493,N_14579,N_14775);
xnor U16494 (N_16494,N_14648,N_13701);
and U16495 (N_16495,N_13849,N_13898);
and U16496 (N_16496,N_13822,N_14823);
nor U16497 (N_16497,N_14261,N_13885);
nor U16498 (N_16498,N_13993,N_14395);
and U16499 (N_16499,N_14695,N_14662);
nor U16500 (N_16500,N_15727,N_15895);
xor U16501 (N_16501,N_15398,N_16109);
xnor U16502 (N_16502,N_16419,N_15259);
xnor U16503 (N_16503,N_15699,N_15902);
nand U16504 (N_16504,N_15276,N_15011);
nor U16505 (N_16505,N_16336,N_15362);
or U16506 (N_16506,N_15364,N_16120);
and U16507 (N_16507,N_16104,N_15549);
xor U16508 (N_16508,N_16192,N_15838);
xor U16509 (N_16509,N_15719,N_15649);
nor U16510 (N_16510,N_15056,N_16086);
nand U16511 (N_16511,N_15129,N_16289);
xnor U16512 (N_16512,N_16191,N_16110);
nor U16513 (N_16513,N_16448,N_16445);
and U16514 (N_16514,N_15973,N_16487);
xnor U16515 (N_16515,N_16429,N_16058);
nor U16516 (N_16516,N_15655,N_16034);
or U16517 (N_16517,N_16428,N_16490);
nor U16518 (N_16518,N_15892,N_15706);
xor U16519 (N_16519,N_15277,N_15758);
nand U16520 (N_16520,N_15370,N_16303);
or U16521 (N_16521,N_15726,N_15438);
or U16522 (N_16522,N_15076,N_15921);
xor U16523 (N_16523,N_16117,N_15609);
nand U16524 (N_16524,N_15185,N_15877);
nand U16525 (N_16525,N_15216,N_15426);
and U16526 (N_16526,N_16122,N_15809);
and U16527 (N_16527,N_15115,N_16290);
and U16528 (N_16528,N_15763,N_15712);
nand U16529 (N_16529,N_16276,N_15485);
xnor U16530 (N_16530,N_15837,N_15095);
and U16531 (N_16531,N_16468,N_16296);
and U16532 (N_16532,N_15596,N_16147);
nor U16533 (N_16533,N_16033,N_15860);
and U16534 (N_16534,N_16000,N_16301);
nor U16535 (N_16535,N_16411,N_16321);
nand U16536 (N_16536,N_16111,N_16157);
nor U16537 (N_16537,N_15691,N_15698);
nor U16538 (N_16538,N_16295,N_15529);
nand U16539 (N_16539,N_15540,N_15832);
nor U16540 (N_16540,N_16356,N_15608);
xor U16541 (N_16541,N_16227,N_15483);
nand U16542 (N_16542,N_15054,N_15964);
or U16543 (N_16543,N_15998,N_15330);
or U16544 (N_16544,N_15887,N_16377);
or U16545 (N_16545,N_15700,N_15530);
nand U16546 (N_16546,N_15612,N_16374);
and U16547 (N_16547,N_15231,N_15177);
xor U16548 (N_16548,N_15855,N_15792);
and U16549 (N_16549,N_15939,N_15573);
nor U16550 (N_16550,N_16386,N_15825);
or U16551 (N_16551,N_15894,N_15842);
or U16552 (N_16552,N_15215,N_15948);
and U16553 (N_16553,N_16202,N_16119);
nand U16554 (N_16554,N_15790,N_16491);
xnor U16555 (N_16555,N_15603,N_15203);
xor U16556 (N_16556,N_16248,N_16348);
xnor U16557 (N_16557,N_16354,N_15085);
or U16558 (N_16558,N_16352,N_15339);
nand U16559 (N_16559,N_15724,N_15545);
nand U16560 (N_16560,N_15965,N_16341);
nor U16561 (N_16561,N_15361,N_15197);
and U16562 (N_16562,N_16071,N_15909);
and U16563 (N_16563,N_15123,N_16394);
nor U16564 (N_16564,N_16010,N_15447);
nor U16565 (N_16565,N_15641,N_16262);
nand U16566 (N_16566,N_16112,N_15968);
nand U16567 (N_16567,N_16218,N_15774);
and U16568 (N_16568,N_16068,N_15273);
or U16569 (N_16569,N_16275,N_16249);
or U16570 (N_16570,N_15025,N_15158);
nand U16571 (N_16571,N_16049,N_16298);
and U16572 (N_16572,N_15335,N_16399);
xor U16573 (N_16573,N_15289,N_16153);
xnor U16574 (N_16574,N_15082,N_16063);
xnor U16575 (N_16575,N_15086,N_16201);
nand U16576 (N_16576,N_16114,N_15263);
or U16577 (N_16577,N_15850,N_15280);
or U16578 (N_16578,N_16257,N_15249);
and U16579 (N_16579,N_15637,N_16042);
nor U16580 (N_16580,N_15214,N_15118);
nand U16581 (N_16581,N_15788,N_15898);
nor U16582 (N_16582,N_15652,N_15754);
xnor U16583 (N_16583,N_16362,N_15507);
nor U16584 (N_16584,N_15879,N_16162);
or U16585 (N_16585,N_15552,N_16170);
nand U16586 (N_16586,N_16494,N_16477);
or U16587 (N_16587,N_15930,N_15681);
nor U16588 (N_16588,N_15765,N_15728);
or U16589 (N_16589,N_15924,N_15105);
xor U16590 (N_16590,N_16047,N_16219);
and U16591 (N_16591,N_15599,N_15200);
nand U16592 (N_16592,N_15382,N_15949);
xor U16593 (N_16593,N_15816,N_15759);
xnor U16594 (N_16594,N_16233,N_15291);
or U16595 (N_16595,N_15081,N_16138);
nor U16596 (N_16596,N_15099,N_16172);
and U16597 (N_16597,N_15631,N_16409);
and U16598 (N_16598,N_15650,N_15802);
nor U16599 (N_16599,N_16451,N_16200);
xor U16600 (N_16600,N_16217,N_15640);
nor U16601 (N_16601,N_15154,N_15668);
xor U16602 (N_16602,N_15069,N_16496);
or U16603 (N_16603,N_15854,N_15334);
or U16604 (N_16604,N_15675,N_16361);
xor U16605 (N_16605,N_15340,N_15153);
nor U16606 (N_16606,N_15161,N_16417);
xnor U16607 (N_16607,N_16018,N_15981);
xor U16608 (N_16608,N_16072,N_16273);
nand U16609 (N_16609,N_15164,N_15421);
nand U16610 (N_16610,N_16251,N_15532);
xor U16611 (N_16611,N_15635,N_15394);
xor U16612 (N_16612,N_15418,N_15481);
and U16613 (N_16613,N_15567,N_15270);
nand U16614 (N_16614,N_16323,N_15392);
xnor U16615 (N_16615,N_16091,N_15793);
and U16616 (N_16616,N_15680,N_15477);
nand U16617 (N_16617,N_16467,N_15536);
and U16618 (N_16618,N_15862,N_16061);
xor U16619 (N_16619,N_16267,N_16366);
nand U16620 (N_16620,N_16213,N_16133);
and U16621 (N_16621,N_15414,N_15278);
xor U16622 (N_16622,N_15120,N_16315);
or U16623 (N_16623,N_15302,N_16163);
or U16624 (N_16624,N_15296,N_16476);
nor U16625 (N_16625,N_15046,N_15119);
xor U16626 (N_16626,N_15987,N_16032);
nand U16627 (N_16627,N_15893,N_15142);
xnor U16628 (N_16628,N_16343,N_15366);
or U16629 (N_16629,N_15137,N_15749);
nand U16630 (N_16630,N_16064,N_15441);
or U16631 (N_16631,N_16441,N_15646);
and U16632 (N_16632,N_15172,N_16272);
nand U16633 (N_16633,N_16115,N_15138);
nand U16634 (N_16634,N_15254,N_16196);
xor U16635 (N_16635,N_15328,N_15840);
nand U16636 (N_16636,N_15791,N_16055);
xor U16637 (N_16637,N_15386,N_16472);
xnor U16638 (N_16638,N_15055,N_16353);
nand U16639 (N_16639,N_16479,N_15610);
nand U16640 (N_16640,N_15126,N_16141);
and U16641 (N_16641,N_15569,N_15692);
xnor U16642 (N_16642,N_15799,N_15733);
nor U16643 (N_16643,N_16039,N_15400);
xnor U16644 (N_16644,N_15482,N_15347);
or U16645 (N_16645,N_15236,N_16132);
and U16646 (N_16646,N_16131,N_16384);
or U16647 (N_16647,N_16370,N_15527);
nand U16648 (N_16648,N_15885,N_15807);
or U16649 (N_16649,N_15678,N_16378);
and U16650 (N_16650,N_16422,N_15248);
nor U16651 (N_16651,N_15494,N_15146);
or U16652 (N_16652,N_16087,N_15720);
nor U16653 (N_16653,N_16439,N_15408);
nor U16654 (N_16654,N_15217,N_15794);
or U16655 (N_16655,N_15204,N_15562);
nor U16656 (N_16656,N_16212,N_15570);
nand U16657 (N_16657,N_15133,N_16434);
nand U16658 (N_16658,N_16221,N_15354);
nand U16659 (N_16659,N_15260,N_15342);
nand U16660 (N_16660,N_16449,N_15967);
nor U16661 (N_16661,N_16349,N_15053);
or U16662 (N_16662,N_15104,N_15311);
xor U16663 (N_16663,N_16299,N_16358);
nor U16664 (N_16664,N_16407,N_15677);
or U16665 (N_16665,N_15566,N_15982);
and U16666 (N_16666,N_15778,N_15616);
and U16667 (N_16667,N_16266,N_15232);
or U16668 (N_16668,N_16012,N_16339);
and U16669 (N_16669,N_15420,N_15518);
xnor U16670 (N_16670,N_15308,N_15595);
or U16671 (N_16671,N_16327,N_16440);
xnor U16672 (N_16672,N_16139,N_15316);
xor U16673 (N_16673,N_15456,N_15935);
xnor U16674 (N_16674,N_15384,N_16169);
or U16675 (N_16675,N_16195,N_16264);
and U16676 (N_16676,N_16329,N_16204);
nand U16677 (N_16677,N_15001,N_15294);
nor U16678 (N_16678,N_15100,N_15206);
and U16679 (N_16679,N_16392,N_15828);
xor U16680 (N_16680,N_15159,N_15522);
and U16681 (N_16681,N_15078,N_15615);
nand U16682 (N_16682,N_15397,N_16060);
xor U16683 (N_16683,N_15723,N_16046);
nand U16684 (N_16684,N_15525,N_16176);
xor U16685 (N_16685,N_15365,N_15149);
nand U16686 (N_16686,N_15410,N_15090);
xnor U16687 (N_16687,N_15002,N_16216);
or U16688 (N_16688,N_16402,N_15600);
nor U16689 (N_16689,N_15008,N_15568);
nor U16690 (N_16690,N_16453,N_16181);
nor U16691 (N_16691,N_16076,N_15089);
or U16692 (N_16692,N_15623,N_15238);
xor U16693 (N_16693,N_15240,N_15849);
xor U16694 (N_16694,N_16474,N_16395);
nand U16695 (N_16695,N_15509,N_15049);
xnor U16696 (N_16696,N_16475,N_16263);
and U16697 (N_16697,N_16148,N_15601);
and U16698 (N_16698,N_16178,N_15017);
xnor U16699 (N_16699,N_15343,N_15437);
and U16700 (N_16700,N_16461,N_15212);
xnor U16701 (N_16701,N_16226,N_16433);
xor U16702 (N_16702,N_15404,N_16238);
nand U16703 (N_16703,N_16415,N_15521);
nand U16704 (N_16704,N_15127,N_16035);
xor U16705 (N_16705,N_15381,N_15312);
and U16706 (N_16706,N_15274,N_15554);
or U16707 (N_16707,N_15506,N_15432);
or U16708 (N_16708,N_15564,N_15586);
nand U16709 (N_16709,N_15150,N_16067);
nor U16710 (N_16710,N_15593,N_16306);
xnor U16711 (N_16711,N_16123,N_16156);
nor U16712 (N_16712,N_16137,N_15766);
nand U16713 (N_16713,N_16432,N_15590);
xor U16714 (N_16714,N_16258,N_15288);
xnor U16715 (N_16715,N_15314,N_16319);
and U16716 (N_16716,N_15209,N_15945);
and U16717 (N_16717,N_15777,N_15062);
nor U16718 (N_16718,N_16281,N_15472);
nor U16719 (N_16719,N_15018,N_16292);
nand U16720 (N_16720,N_16335,N_15951);
xor U16721 (N_16721,N_15210,N_15369);
nand U16722 (N_16722,N_16090,N_15304);
nand U16723 (N_16723,N_15391,N_15764);
nor U16724 (N_16724,N_15351,N_16426);
xnor U16725 (N_16725,N_16317,N_15747);
nor U16726 (N_16726,N_15870,N_16245);
nand U16727 (N_16727,N_15189,N_15975);
nor U16728 (N_16728,N_15092,N_15102);
and U16729 (N_16729,N_15143,N_15242);
nand U16730 (N_16730,N_15136,N_16084);
nand U16731 (N_16731,N_16359,N_15901);
or U16732 (N_16732,N_15088,N_16239);
nand U16733 (N_16733,N_15332,N_15972);
xor U16734 (N_16734,N_15106,N_15041);
nand U16735 (N_16735,N_15271,N_16069);
xor U16736 (N_16736,N_15743,N_15889);
nand U16737 (N_16737,N_15744,N_16446);
or U16738 (N_16738,N_15097,N_15539);
xnor U16739 (N_16739,N_16416,N_15226);
or U16740 (N_16740,N_15687,N_16015);
xor U16741 (N_16741,N_16485,N_15876);
or U16742 (N_16742,N_16009,N_15377);
or U16743 (N_16743,N_15219,N_16078);
nor U16744 (N_16744,N_16002,N_15258);
or U16745 (N_16745,N_15553,N_15269);
and U16746 (N_16746,N_15434,N_16187);
nand U16747 (N_16747,N_15845,N_15039);
xnor U16748 (N_16748,N_15974,N_16247);
xnor U16749 (N_16749,N_16307,N_15941);
nand U16750 (N_16750,N_15666,N_15995);
and U16751 (N_16751,N_15644,N_15036);
nor U16752 (N_16752,N_16089,N_15952);
nand U16753 (N_16753,N_15211,N_16206);
nor U16754 (N_16754,N_16283,N_15528);
or U16755 (N_16755,N_15508,N_15869);
nand U16756 (N_16756,N_15704,N_15348);
xnor U16757 (N_16757,N_16098,N_15739);
xor U16758 (N_16758,N_15256,N_16161);
or U16759 (N_16759,N_16220,N_15166);
xor U16760 (N_16760,N_15297,N_16043);
or U16761 (N_16761,N_15499,N_16246);
and U16762 (N_16762,N_16385,N_15286);
and U16763 (N_16763,N_15988,N_16023);
or U16764 (N_16764,N_15622,N_15851);
or U16765 (N_16765,N_15458,N_15985);
nor U16766 (N_16766,N_16155,N_15780);
nand U16767 (N_16767,N_16088,N_15416);
nor U16768 (N_16768,N_15003,N_15886);
nor U16769 (N_16769,N_16014,N_16484);
or U16770 (N_16770,N_16243,N_15897);
or U16771 (N_16771,N_15173,N_15019);
and U16772 (N_16772,N_15817,N_15745);
nand U16773 (N_16773,N_15014,N_16175);
nand U16774 (N_16774,N_16186,N_15787);
xnor U16775 (N_16775,N_15327,N_15021);
nand U16776 (N_16776,N_15181,N_15657);
xnor U16777 (N_16777,N_15000,N_15705);
and U16778 (N_16778,N_16030,N_16488);
xor U16779 (N_16779,N_15629,N_15592);
nand U16780 (N_16780,N_16454,N_15915);
xor U16781 (N_16781,N_15872,N_15068);
or U16782 (N_16782,N_16152,N_16242);
or U16783 (N_16783,N_15954,N_15572);
nand U16784 (N_16784,N_16280,N_15688);
nor U16785 (N_16785,N_16334,N_16376);
nor U16786 (N_16786,N_15435,N_15141);
nor U16787 (N_16787,N_15963,N_15752);
nor U16788 (N_16788,N_16005,N_16189);
or U16789 (N_16789,N_15576,N_16346);
and U16790 (N_16790,N_15950,N_15848);
nor U16791 (N_16791,N_15762,N_16190);
nor U16792 (N_16792,N_15683,N_15852);
xor U16793 (N_16793,N_15673,N_15505);
and U16794 (N_16794,N_15301,N_16116);
or U16795 (N_16795,N_15101,N_16404);
or U16796 (N_16796,N_15463,N_15198);
nor U16797 (N_16797,N_16270,N_15066);
or U16798 (N_16798,N_15145,N_15051);
xnor U16799 (N_16799,N_15109,N_16011);
nor U16800 (N_16800,N_16185,N_16168);
nor U16801 (N_16801,N_15513,N_16383);
nand U16802 (N_16802,N_15077,N_15239);
nor U16803 (N_16803,N_16293,N_15502);
or U16804 (N_16804,N_16209,N_15496);
or U16805 (N_16805,N_15547,N_15969);
xnor U16806 (N_16806,N_16188,N_16066);
nor U16807 (N_16807,N_15682,N_15542);
xor U16808 (N_16808,N_15234,N_15796);
xnor U16809 (N_16809,N_15520,N_15679);
and U16810 (N_16810,N_15861,N_16128);
nor U16811 (N_16811,N_15004,N_15379);
xor U16812 (N_16812,N_15702,N_16305);
or U16813 (N_16813,N_15955,N_15769);
nor U16814 (N_16814,N_15923,N_15504);
and U16815 (N_16815,N_16431,N_15429);
xor U16816 (N_16816,N_16410,N_15052);
and U16817 (N_16817,N_16436,N_15372);
nand U16818 (N_16818,N_15625,N_15449);
nand U16819 (N_16819,N_15546,N_16028);
nand U16820 (N_16820,N_15918,N_16150);
or U16821 (N_16821,N_15027,N_15065);
nand U16822 (N_16822,N_16499,N_15841);
xor U16823 (N_16823,N_15959,N_16223);
or U16824 (N_16824,N_16164,N_15043);
nand U16825 (N_16825,N_16489,N_16438);
xor U16826 (N_16826,N_16425,N_15268);
or U16827 (N_16827,N_15797,N_16154);
nand U16828 (N_16828,N_15492,N_15050);
nand U16829 (N_16829,N_15346,N_16297);
nor U16830 (N_16830,N_15188,N_16211);
nand U16831 (N_16831,N_15510,N_16231);
or U16832 (N_16832,N_15111,N_15072);
nand U16833 (N_16833,N_15591,N_15038);
or U16834 (N_16834,N_16052,N_15760);
or U16835 (N_16835,N_15829,N_15531);
and U16836 (N_16836,N_16424,N_16369);
and U16837 (N_16837,N_15979,N_16387);
and U16838 (N_16838,N_15582,N_15989);
nand U16839 (N_16839,N_15380,N_15953);
and U16840 (N_16840,N_15484,N_15980);
and U16841 (N_16841,N_16146,N_15707);
or U16842 (N_16842,N_16085,N_16480);
nor U16843 (N_16843,N_15942,N_16456);
and U16844 (N_16844,N_15465,N_15208);
or U16845 (N_16845,N_15928,N_15423);
and U16846 (N_16846,N_16225,N_15500);
nor U16847 (N_16847,N_16309,N_16447);
xnor U16848 (N_16848,N_15814,N_15007);
and U16849 (N_16849,N_16160,N_15207);
or U16850 (N_16850,N_15824,N_15772);
or U16851 (N_16851,N_15961,N_15868);
nand U16852 (N_16852,N_15667,N_15471);
and U16853 (N_16853,N_16364,N_15321);
xnor U16854 (N_16854,N_15636,N_16020);
and U16855 (N_16855,N_15010,N_15803);
xor U16856 (N_16856,N_15873,N_16400);
nand U16857 (N_16857,N_15716,N_15560);
nand U16858 (N_16858,N_16406,N_15122);
nand U16859 (N_16859,N_16079,N_16255);
and U16860 (N_16860,N_15061,N_15709);
and U16861 (N_16861,N_15373,N_15457);
or U16862 (N_16862,N_16240,N_15891);
xor U16863 (N_16863,N_15503,N_16082);
and U16864 (N_16864,N_15445,N_16450);
xnor U16865 (N_16865,N_15024,N_16342);
nand U16866 (N_16866,N_15775,N_15501);
nor U16867 (N_16867,N_16421,N_15732);
nor U16868 (N_16868,N_15746,N_15722);
and U16869 (N_16869,N_15047,N_15229);
nor U16870 (N_16870,N_15907,N_15741);
xnor U16871 (N_16871,N_15108,N_15190);
xor U16872 (N_16872,N_16458,N_16166);
and U16873 (N_16873,N_16100,N_16452);
nor U16874 (N_16874,N_16019,N_15786);
and U16875 (N_16875,N_16121,N_15060);
xor U16876 (N_16876,N_15839,N_15919);
or U16877 (N_16877,N_15460,N_16322);
nor U16878 (N_16878,N_16372,N_16048);
and U16879 (N_16879,N_15535,N_16259);
nand U16880 (N_16880,N_16355,N_16013);
and U16881 (N_16881,N_15823,N_15064);
and U16882 (N_16882,N_15550,N_16256);
nand U16883 (N_16883,N_16165,N_16194);
nor U16884 (N_16884,N_15233,N_15761);
or U16885 (N_16885,N_16236,N_15074);
nand U16886 (N_16886,N_16235,N_16482);
nor U16887 (N_16887,N_15514,N_15300);
nand U16888 (N_16888,N_15202,N_16271);
or U16889 (N_16889,N_15696,N_15658);
and U16890 (N_16890,N_16481,N_15927);
xnor U16891 (N_16891,N_15192,N_15246);
or U16892 (N_16892,N_15124,N_15821);
xor U16893 (N_16893,N_15491,N_15844);
nand U16894 (N_16894,N_15882,N_15805);
or U16895 (N_16895,N_15526,N_15626);
nor U16896 (N_16896,N_16310,N_15247);
nand U16897 (N_16897,N_15731,N_15356);
xnor U16898 (N_16898,N_15225,N_15224);
nand U16899 (N_16899,N_16183,N_15395);
or U16900 (N_16900,N_16332,N_15571);
or U16901 (N_16901,N_15588,N_16024);
and U16902 (N_16902,N_15911,N_15903);
and U16903 (N_16903,N_16027,N_15476);
and U16904 (N_16904,N_15858,N_15424);
nand U16905 (N_16905,N_16101,N_15556);
and U16906 (N_16906,N_15978,N_15815);
xor U16907 (N_16907,N_15451,N_15645);
nor U16908 (N_16908,N_16279,N_15012);
and U16909 (N_16909,N_15337,N_16371);
xnor U16910 (N_16910,N_15619,N_15358);
xor U16911 (N_16911,N_15859,N_15660);
xnor U16912 (N_16912,N_15875,N_15639);
nand U16913 (N_16913,N_15326,N_16340);
xor U16914 (N_16914,N_16408,N_15098);
and U16915 (N_16915,N_16237,N_15776);
and U16916 (N_16916,N_16495,N_15818);
nor U16917 (N_16917,N_16197,N_16379);
and U16918 (N_16918,N_15235,N_15515);
xor U16919 (N_16919,N_15402,N_15511);
nand U16920 (N_16920,N_16050,N_16291);
and U16921 (N_16921,N_15866,N_16036);
and U16922 (N_16922,N_16304,N_16007);
nand U16923 (N_16923,N_15721,N_15983);
or U16924 (N_16924,N_16389,N_16106);
xor U16925 (N_16925,N_16151,N_16435);
or U16926 (N_16926,N_15338,N_16493);
xnor U16927 (N_16927,N_15446,N_16096);
nand U16928 (N_16928,N_15367,N_15374);
nand U16929 (N_16929,N_15042,N_16284);
and U16930 (N_16930,N_15750,N_15306);
and U16931 (N_16931,N_16388,N_15071);
nor U16932 (N_16932,N_15606,N_15857);
xor U16933 (N_16933,N_15399,N_15298);
nand U16934 (N_16934,N_15524,N_16017);
nand U16935 (N_16935,N_15922,N_16171);
xnor U16936 (N_16936,N_16316,N_15613);
or U16937 (N_16937,N_15648,N_16459);
or U16938 (N_16938,N_15581,N_16229);
xor U16939 (N_16939,N_16469,N_16357);
and U16940 (N_16940,N_16405,N_15396);
xor U16941 (N_16941,N_15128,N_15194);
or U16942 (N_16942,N_15257,N_15820);
or U16943 (N_16943,N_15630,N_15140);
or U16944 (N_16944,N_15703,N_15359);
or U16945 (N_16945,N_15037,N_16464);
nor U16946 (N_16946,N_15634,N_15662);
and U16947 (N_16947,N_16308,N_15360);
or U16948 (N_16948,N_15598,N_15250);
or U16949 (N_16949,N_15905,N_16059);
and U16950 (N_16950,N_15130,N_15620);
nor U16951 (N_16951,N_15984,N_15541);
and U16952 (N_16952,N_15125,N_15315);
nor U16953 (N_16953,N_15070,N_16118);
or U16954 (N_16954,N_15986,N_15411);
or U16955 (N_16955,N_15697,N_16001);
or U16956 (N_16956,N_16159,N_15439);
nor U16957 (N_16957,N_16207,N_16070);
nand U16958 (N_16958,N_15701,N_15148);
nor U16959 (N_16959,N_15783,N_16230);
or U16960 (N_16960,N_15264,N_15237);
xor U16961 (N_16961,N_15079,N_15669);
or U16962 (N_16962,N_15251,N_15023);
nor U16963 (N_16963,N_15864,N_15587);
xnor U16964 (N_16964,N_15512,N_15729);
nor U16965 (N_16965,N_15322,N_16016);
nand U16966 (N_16966,N_15585,N_15144);
or U16967 (N_16967,N_16093,N_15962);
or U16968 (N_16968,N_15405,N_15523);
xnor U16969 (N_16969,N_15227,N_15813);
nor U16970 (N_16970,N_15413,N_15084);
or U16971 (N_16971,N_15193,N_15162);
or U16972 (N_16972,N_15466,N_15908);
xnor U16973 (N_16973,N_15168,N_16184);
or U16974 (N_16974,N_16053,N_15187);
nor U16975 (N_16975,N_15779,N_15847);
nor U16976 (N_16976,N_16401,N_16466);
or U16977 (N_16977,N_16260,N_16345);
nand U16978 (N_16978,N_15715,N_15022);
xnor U16979 (N_16979,N_15191,N_16486);
nand U16980 (N_16980,N_15808,N_15375);
and U16981 (N_16981,N_15357,N_15933);
and U16982 (N_16982,N_15222,N_15419);
and U16983 (N_16983,N_15464,N_15121);
xor U16984 (N_16984,N_15165,N_15767);
nor U16985 (N_16985,N_16420,N_15452);
or U16986 (N_16986,N_16427,N_16338);
nand U16987 (N_16987,N_15305,N_15730);
xnor U16988 (N_16988,N_15624,N_15461);
nor U16989 (N_16989,N_15970,N_16081);
xnor U16990 (N_16990,N_15156,N_15310);
or U16991 (N_16991,N_15218,N_15473);
nand U16992 (N_16992,N_15252,N_15450);
nor U16993 (N_16993,N_15266,N_15407);
nor U16994 (N_16994,N_15368,N_16261);
nor U16995 (N_16995,N_15131,N_15621);
and U16996 (N_16996,N_15063,N_16344);
xnor U16997 (N_16997,N_16094,N_15519);
xnor U16998 (N_16998,N_15584,N_15672);
or U16999 (N_16999,N_15904,N_15663);
nand U17000 (N_17000,N_15863,N_15956);
xor U17001 (N_17001,N_15781,N_15966);
nor U17002 (N_17002,N_15112,N_16103);
nand U17003 (N_17003,N_15459,N_16149);
or U17004 (N_17004,N_15479,N_15353);
nand U17005 (N_17005,N_16465,N_15881);
or U17006 (N_17006,N_16462,N_15557);
nand U17007 (N_17007,N_16278,N_15478);
or U17008 (N_17008,N_16130,N_16470);
and U17009 (N_17009,N_16037,N_16313);
and U17010 (N_17010,N_15385,N_15265);
xnor U17011 (N_17011,N_15262,N_15811);
and U17012 (N_17012,N_15333,N_15714);
xor U17013 (N_17013,N_15307,N_15559);
or U17014 (N_17014,N_16269,N_16102);
xor U17015 (N_17015,N_15493,N_15167);
or U17016 (N_17016,N_15376,N_16041);
nor U17017 (N_17017,N_15160,N_15040);
or U17018 (N_17018,N_15299,N_16038);
nand U17019 (N_17019,N_15117,N_15944);
nand U17020 (N_17020,N_16108,N_15561);
or U17021 (N_17021,N_15147,N_15757);
nor U17022 (N_17022,N_15474,N_15602);
nand U17023 (N_17023,N_15275,N_15654);
and U17024 (N_17024,N_15751,N_15412);
xnor U17025 (N_17025,N_15389,N_15281);
or U17026 (N_17026,N_15604,N_16337);
or U17027 (N_17027,N_16492,N_16045);
or U17028 (N_17028,N_15341,N_15516);
nor U17029 (N_17029,N_15151,N_15993);
and U17030 (N_17030,N_16126,N_16478);
nand U17031 (N_17031,N_16418,N_15436);
nor U17032 (N_17032,N_16380,N_15331);
nand U17033 (N_17033,N_15795,N_15028);
and U17034 (N_17034,N_15344,N_15558);
nand U17035 (N_17035,N_15057,N_16330);
or U17036 (N_17036,N_15846,N_16006);
and U17037 (N_17037,N_16397,N_16244);
xnor U17038 (N_17038,N_15833,N_15390);
xnor U17039 (N_17039,N_15355,N_15653);
or U17040 (N_17040,N_16314,N_15045);
nor U17041 (N_17041,N_16250,N_15467);
or U17042 (N_17042,N_15155,N_15770);
nand U17043 (N_17043,N_15664,N_15579);
nand U17044 (N_17044,N_15916,N_15205);
nand U17045 (N_17045,N_15910,N_15822);
xnor U17046 (N_17046,N_16368,N_16145);
nand U17047 (N_17047,N_16413,N_15801);
or U17048 (N_17048,N_16142,N_15773);
and U17049 (N_17049,N_15293,N_15170);
and U17050 (N_17050,N_15318,N_15843);
or U17051 (N_17051,N_16326,N_15195);
and U17052 (N_17052,N_15771,N_15324);
xor U17053 (N_17053,N_15044,N_16430);
and U17054 (N_17054,N_15015,N_15486);
xor U17055 (N_17055,N_15462,N_15032);
xnor U17056 (N_17056,N_16074,N_15936);
nor U17057 (N_17057,N_16134,N_15537);
xor U17058 (N_17058,N_15755,N_16143);
and U17059 (N_17059,N_16412,N_15455);
xor U17060 (N_17060,N_15497,N_15490);
xor U17061 (N_17061,N_16140,N_15134);
nand U17062 (N_17062,N_15992,N_15865);
and U17063 (N_17063,N_15533,N_15228);
or U17064 (N_17064,N_15352,N_15006);
or U17065 (N_17065,N_15544,N_16054);
nand U17066 (N_17066,N_16177,N_15929);
nand U17067 (N_17067,N_15643,N_15548);
nand U17068 (N_17068,N_15943,N_16360);
xor U17069 (N_17069,N_15690,N_16381);
or U17070 (N_17070,N_16193,N_15831);
nand U17071 (N_17071,N_15827,N_16483);
or U17072 (N_17072,N_15563,N_15874);
or U17073 (N_17073,N_16268,N_15283);
nor U17074 (N_17074,N_15977,N_15578);
xor U17075 (N_17075,N_15480,N_15638);
and U17076 (N_17076,N_15734,N_15642);
nand U17077 (N_17077,N_15029,N_15958);
nand U17078 (N_17078,N_15738,N_15448);
or U17079 (N_17079,N_15614,N_16312);
nor U17080 (N_17080,N_16325,N_16403);
or U17081 (N_17081,N_16080,N_15913);
xnor U17082 (N_17082,N_15087,N_16252);
xor U17083 (N_17083,N_15589,N_15748);
nor U17084 (N_17084,N_16173,N_15255);
and U17085 (N_17085,N_16457,N_16443);
nor U17086 (N_17086,N_15999,N_16003);
xor U17087 (N_17087,N_16135,N_15336);
xnor U17088 (N_17088,N_16350,N_15174);
nor U17089 (N_17089,N_15651,N_16077);
nor U17090 (N_17090,N_15183,N_16051);
xor U17091 (N_17091,N_15319,N_16057);
and U17092 (N_17092,N_16373,N_15888);
and U17093 (N_17093,N_15253,N_16008);
and U17094 (N_17094,N_15611,N_15565);
nor U17095 (N_17095,N_16442,N_15890);
nor U17096 (N_17096,N_15899,N_15830);
nand U17097 (N_17097,N_16320,N_16351);
nand U17098 (N_17098,N_15349,N_15058);
or U17099 (N_17099,N_15804,N_15659);
xnor U17100 (N_17100,N_15694,N_15454);
xor U17101 (N_17101,N_15938,N_15917);
nand U17102 (N_17102,N_15498,N_15555);
xnor U17103 (N_17103,N_15947,N_16179);
and U17104 (N_17104,N_15132,N_15580);
nand U17105 (N_17105,N_15934,N_16333);
or U17106 (N_17106,N_16031,N_16455);
nand U17107 (N_17107,N_15835,N_16124);
and U17108 (N_17108,N_15671,N_15094);
and U17109 (N_17109,N_15199,N_16222);
nand U17110 (N_17110,N_15957,N_15453);
and U17111 (N_17111,N_15080,N_16022);
xnor U17112 (N_17112,N_15800,N_15317);
or U17113 (N_17113,N_15871,N_15756);
nand U17114 (N_17114,N_16044,N_15279);
xor U17115 (N_17115,N_15853,N_15856);
nor U17116 (N_17116,N_15627,N_15243);
and U17117 (N_17117,N_15422,N_15618);
nand U17118 (N_17118,N_15303,N_16107);
or U17119 (N_17119,N_15371,N_16203);
nor U17120 (N_17120,N_15427,N_15883);
nor U17121 (N_17121,N_16199,N_15213);
nor U17122 (N_17122,N_15313,N_15617);
and U17123 (N_17123,N_16282,N_15440);
or U17124 (N_17124,N_16331,N_16265);
xor U17125 (N_17125,N_15946,N_15388);
or U17126 (N_17126,N_15925,N_15401);
or U17127 (N_17127,N_16375,N_15896);
and U17128 (N_17128,N_15035,N_15798);
and U17129 (N_17129,N_16232,N_15534);
nand U17130 (N_17130,N_15517,N_15103);
and U17131 (N_17131,N_15048,N_15674);
nor U17132 (N_17132,N_16158,N_15836);
xnor U17133 (N_17133,N_15442,N_15073);
nand U17134 (N_17134,N_15116,N_15693);
or U17135 (N_17135,N_15632,N_15113);
nor U17136 (N_17136,N_15735,N_16277);
or U17137 (N_17137,N_15030,N_15607);
or U17138 (N_17138,N_16129,N_15009);
or U17139 (N_17139,N_16208,N_15393);
or U17140 (N_17140,N_15812,N_15059);
or U17141 (N_17141,N_15551,N_15067);
xor U17142 (N_17142,N_16075,N_15425);
nor U17143 (N_17143,N_15244,N_16294);
nor U17144 (N_17144,N_15996,N_16125);
or U17145 (N_17145,N_16099,N_16311);
nor U17146 (N_17146,N_15670,N_15180);
nor U17147 (N_17147,N_15718,N_15406);
nor U17148 (N_17148,N_15179,N_15139);
and U17149 (N_17149,N_16253,N_15184);
xnor U17150 (N_17150,N_15267,N_15033);
nor U17151 (N_17151,N_15740,N_15574);
and U17152 (N_17152,N_15325,N_15309);
nor U17153 (N_17153,N_15387,N_15417);
nor U17154 (N_17154,N_15178,N_15577);
nand U17155 (N_17155,N_15196,N_16274);
xnor U17156 (N_17156,N_15428,N_15834);
and U17157 (N_17157,N_15489,N_16092);
or U17158 (N_17158,N_15628,N_15221);
and U17159 (N_17159,N_16073,N_15991);
or U17160 (N_17160,N_15661,N_15135);
xor U17161 (N_17161,N_15034,N_15633);
xnor U17162 (N_17162,N_15906,N_16302);
xnor U17163 (N_17163,N_15940,N_16367);
or U17164 (N_17164,N_16398,N_15443);
xor U17165 (N_17165,N_15378,N_16473);
nand U17166 (N_17166,N_15867,N_15710);
or U17167 (N_17167,N_15075,N_15960);
and U17168 (N_17168,N_15487,N_15676);
and U17169 (N_17169,N_15737,N_15083);
nand U17170 (N_17170,N_15295,N_16285);
nand U17171 (N_17171,N_15594,N_15785);
xor U17172 (N_17172,N_16136,N_16300);
xnor U17173 (N_17173,N_16365,N_15736);
nor U17174 (N_17174,N_15093,N_15912);
or U17175 (N_17175,N_16228,N_16471);
nor U17176 (N_17176,N_15684,N_16390);
nand U17177 (N_17177,N_15647,N_15107);
or U17178 (N_17178,N_15431,N_15789);
nor U17179 (N_17179,N_15350,N_16363);
xor U17180 (N_17180,N_15878,N_16113);
and U17181 (N_17181,N_16241,N_15708);
nor U17182 (N_17182,N_16347,N_16463);
nor U17183 (N_17183,N_16095,N_16210);
and U17184 (N_17184,N_15880,N_15990);
xor U17185 (N_17185,N_15470,N_15713);
xnor U17186 (N_17186,N_15223,N_15261);
or U17187 (N_17187,N_16065,N_15282);
nor U17188 (N_17188,N_15096,N_15345);
or U17189 (N_17189,N_15114,N_15169);
or U17190 (N_17190,N_15287,N_15685);
nor U17191 (N_17191,N_16497,N_16286);
and U17192 (N_17192,N_15782,N_16214);
xnor U17193 (N_17193,N_15415,N_15926);
or U17194 (N_17194,N_15292,N_15110);
and U17195 (N_17195,N_15932,N_15656);
and U17196 (N_17196,N_15245,N_16174);
xnor U17197 (N_17197,N_15201,N_15711);
nand U17198 (N_17198,N_16224,N_15230);
or U17199 (N_17199,N_15725,N_15013);
nand U17200 (N_17200,N_15320,N_16288);
nand U17201 (N_17201,N_15182,N_16021);
or U17202 (N_17202,N_15433,N_15994);
nand U17203 (N_17203,N_15931,N_15409);
or U17204 (N_17204,N_16026,N_16025);
nand U17205 (N_17205,N_15157,N_15026);
or U17206 (N_17206,N_16040,N_15768);
or U17207 (N_17207,N_15884,N_16198);
or U17208 (N_17208,N_16004,N_15937);
nand U17209 (N_17209,N_15176,N_15469);
and U17210 (N_17210,N_15538,N_15005);
or U17211 (N_17211,N_16097,N_15171);
nand U17212 (N_17212,N_15695,N_16056);
nand U17213 (N_17213,N_16444,N_16029);
nor U17214 (N_17214,N_16083,N_15290);
xor U17215 (N_17215,N_15810,N_16234);
and U17216 (N_17216,N_15717,N_15403);
xor U17217 (N_17217,N_15900,N_15020);
nor U17218 (N_17218,N_15543,N_15971);
nor U17219 (N_17219,N_15583,N_15175);
nand U17220 (N_17220,N_16324,N_15383);
and U17221 (N_17221,N_16393,N_16382);
and U17222 (N_17222,N_15272,N_15284);
and U17223 (N_17223,N_15241,N_16180);
and U17224 (N_17224,N_15597,N_16144);
nand U17225 (N_17225,N_16167,N_15665);
nor U17226 (N_17226,N_15488,N_16328);
nand U17227 (N_17227,N_16391,N_16062);
nand U17228 (N_17228,N_16105,N_16437);
nor U17229 (N_17229,N_15031,N_15826);
xor U17230 (N_17230,N_16254,N_15152);
or U17231 (N_17231,N_15784,N_15475);
xor U17232 (N_17232,N_15220,N_16205);
nor U17233 (N_17233,N_15997,N_15323);
or U17234 (N_17234,N_15186,N_15605);
nand U17235 (N_17235,N_16318,N_15495);
nand U17236 (N_17236,N_15444,N_15430);
xnor U17237 (N_17237,N_16182,N_15753);
xnor U17238 (N_17238,N_16460,N_15329);
or U17239 (N_17239,N_15806,N_15363);
nand U17240 (N_17240,N_15091,N_15914);
nor U17241 (N_17241,N_15686,N_15016);
xnor U17242 (N_17242,N_16498,N_15163);
nand U17243 (N_17243,N_16414,N_16287);
nand U17244 (N_17244,N_16396,N_16127);
nand U17245 (N_17245,N_16423,N_15920);
xnor U17246 (N_17246,N_15468,N_15819);
nand U17247 (N_17247,N_15575,N_16215);
xnor U17248 (N_17248,N_15742,N_15689);
or U17249 (N_17249,N_15976,N_15285);
nor U17250 (N_17250,N_15081,N_16095);
and U17251 (N_17251,N_15395,N_16021);
or U17252 (N_17252,N_15921,N_15932);
and U17253 (N_17253,N_15954,N_16155);
nor U17254 (N_17254,N_16471,N_15667);
nor U17255 (N_17255,N_16209,N_15270);
or U17256 (N_17256,N_16166,N_15141);
nand U17257 (N_17257,N_15903,N_16007);
nand U17258 (N_17258,N_16126,N_15143);
nand U17259 (N_17259,N_16192,N_15699);
and U17260 (N_17260,N_16186,N_15884);
xor U17261 (N_17261,N_15087,N_15906);
or U17262 (N_17262,N_15513,N_15153);
and U17263 (N_17263,N_15132,N_15957);
xor U17264 (N_17264,N_15165,N_15111);
xor U17265 (N_17265,N_15052,N_16423);
and U17266 (N_17266,N_15148,N_15720);
or U17267 (N_17267,N_15776,N_15445);
nand U17268 (N_17268,N_15568,N_15755);
nor U17269 (N_17269,N_15274,N_15014);
nor U17270 (N_17270,N_16245,N_16124);
nor U17271 (N_17271,N_15056,N_15169);
nor U17272 (N_17272,N_16366,N_15737);
or U17273 (N_17273,N_15270,N_15048);
nor U17274 (N_17274,N_15088,N_15692);
xnor U17275 (N_17275,N_16148,N_15595);
nor U17276 (N_17276,N_16463,N_16046);
xnor U17277 (N_17277,N_15441,N_16156);
nor U17278 (N_17278,N_15828,N_15981);
or U17279 (N_17279,N_15879,N_15343);
or U17280 (N_17280,N_15588,N_15036);
and U17281 (N_17281,N_15729,N_16106);
xnor U17282 (N_17282,N_15056,N_15403);
or U17283 (N_17283,N_15952,N_15823);
nand U17284 (N_17284,N_16276,N_16238);
and U17285 (N_17285,N_15168,N_16055);
nor U17286 (N_17286,N_16127,N_15930);
nand U17287 (N_17287,N_16445,N_15681);
and U17288 (N_17288,N_16432,N_15753);
xnor U17289 (N_17289,N_15359,N_16434);
or U17290 (N_17290,N_15976,N_16106);
xor U17291 (N_17291,N_15146,N_16448);
xnor U17292 (N_17292,N_15648,N_15818);
xnor U17293 (N_17293,N_15214,N_16132);
and U17294 (N_17294,N_15213,N_15938);
xor U17295 (N_17295,N_15675,N_16448);
and U17296 (N_17296,N_15300,N_15107);
and U17297 (N_17297,N_15870,N_16394);
and U17298 (N_17298,N_15378,N_15077);
xor U17299 (N_17299,N_15268,N_15496);
and U17300 (N_17300,N_15817,N_15688);
nor U17301 (N_17301,N_15264,N_16437);
nand U17302 (N_17302,N_16207,N_15460);
or U17303 (N_17303,N_16195,N_16230);
nor U17304 (N_17304,N_15960,N_16425);
nand U17305 (N_17305,N_15064,N_16202);
xor U17306 (N_17306,N_15118,N_15161);
nor U17307 (N_17307,N_15794,N_16352);
nor U17308 (N_17308,N_16333,N_15485);
nor U17309 (N_17309,N_15266,N_16215);
xnor U17310 (N_17310,N_16191,N_16364);
xor U17311 (N_17311,N_15391,N_16279);
or U17312 (N_17312,N_16303,N_15831);
nor U17313 (N_17313,N_15147,N_16030);
or U17314 (N_17314,N_15811,N_16191);
nand U17315 (N_17315,N_15158,N_15847);
nor U17316 (N_17316,N_15481,N_15714);
nand U17317 (N_17317,N_16092,N_15095);
and U17318 (N_17318,N_15027,N_16007);
nand U17319 (N_17319,N_15104,N_16410);
or U17320 (N_17320,N_15887,N_15250);
nand U17321 (N_17321,N_15595,N_15189);
nand U17322 (N_17322,N_16405,N_15732);
xnor U17323 (N_17323,N_15851,N_15308);
nor U17324 (N_17324,N_15465,N_16011);
or U17325 (N_17325,N_15377,N_16053);
xnor U17326 (N_17326,N_15658,N_16117);
xor U17327 (N_17327,N_15580,N_16325);
nand U17328 (N_17328,N_16422,N_16488);
xnor U17329 (N_17329,N_16239,N_16282);
nor U17330 (N_17330,N_16449,N_15012);
and U17331 (N_17331,N_16309,N_15714);
and U17332 (N_17332,N_16426,N_16121);
or U17333 (N_17333,N_15809,N_16027);
nor U17334 (N_17334,N_15816,N_15705);
xnor U17335 (N_17335,N_15715,N_15946);
or U17336 (N_17336,N_15633,N_15446);
nand U17337 (N_17337,N_15834,N_16086);
nor U17338 (N_17338,N_16492,N_15304);
nand U17339 (N_17339,N_16345,N_15882);
or U17340 (N_17340,N_15582,N_16251);
nand U17341 (N_17341,N_15792,N_16311);
or U17342 (N_17342,N_15850,N_15986);
xor U17343 (N_17343,N_16202,N_15217);
or U17344 (N_17344,N_15205,N_16119);
xor U17345 (N_17345,N_15756,N_15651);
or U17346 (N_17346,N_15668,N_15650);
nand U17347 (N_17347,N_15036,N_15492);
xor U17348 (N_17348,N_15528,N_15851);
xnor U17349 (N_17349,N_15734,N_16172);
nor U17350 (N_17350,N_15925,N_15682);
or U17351 (N_17351,N_15450,N_15511);
nand U17352 (N_17352,N_15067,N_16443);
nand U17353 (N_17353,N_16175,N_15290);
nand U17354 (N_17354,N_15656,N_15571);
nor U17355 (N_17355,N_16256,N_15362);
or U17356 (N_17356,N_16290,N_15694);
nor U17357 (N_17357,N_15205,N_15643);
xor U17358 (N_17358,N_16483,N_15460);
xor U17359 (N_17359,N_15732,N_16148);
nand U17360 (N_17360,N_16394,N_16127);
nor U17361 (N_17361,N_16204,N_15342);
xnor U17362 (N_17362,N_16225,N_15892);
nand U17363 (N_17363,N_15863,N_15734);
nand U17364 (N_17364,N_15534,N_15140);
nor U17365 (N_17365,N_15240,N_16257);
nand U17366 (N_17366,N_15271,N_15074);
nor U17367 (N_17367,N_16086,N_15726);
nand U17368 (N_17368,N_15957,N_15938);
or U17369 (N_17369,N_16138,N_16261);
xnor U17370 (N_17370,N_15990,N_15833);
xnor U17371 (N_17371,N_15088,N_16031);
or U17372 (N_17372,N_15561,N_16188);
or U17373 (N_17373,N_15412,N_15569);
nor U17374 (N_17374,N_15620,N_16449);
or U17375 (N_17375,N_16193,N_15297);
nand U17376 (N_17376,N_15049,N_15249);
or U17377 (N_17377,N_16457,N_15706);
nor U17378 (N_17378,N_15789,N_15430);
and U17379 (N_17379,N_15939,N_15584);
xnor U17380 (N_17380,N_16356,N_16401);
nor U17381 (N_17381,N_16302,N_15960);
or U17382 (N_17382,N_16389,N_15556);
nor U17383 (N_17383,N_15718,N_15639);
nor U17384 (N_17384,N_16291,N_16425);
or U17385 (N_17385,N_15738,N_15869);
xor U17386 (N_17386,N_16424,N_15055);
and U17387 (N_17387,N_15074,N_15334);
xor U17388 (N_17388,N_15136,N_16040);
and U17389 (N_17389,N_15901,N_15014);
nand U17390 (N_17390,N_15894,N_15778);
and U17391 (N_17391,N_16208,N_15612);
nor U17392 (N_17392,N_16419,N_15632);
nor U17393 (N_17393,N_15229,N_16401);
xnor U17394 (N_17394,N_15690,N_15682);
nand U17395 (N_17395,N_16459,N_15367);
nor U17396 (N_17396,N_15796,N_16322);
nand U17397 (N_17397,N_15764,N_15668);
and U17398 (N_17398,N_15174,N_15826);
nand U17399 (N_17399,N_16240,N_16439);
nor U17400 (N_17400,N_15198,N_15076);
or U17401 (N_17401,N_16067,N_16319);
or U17402 (N_17402,N_15817,N_15890);
nand U17403 (N_17403,N_15782,N_15752);
nor U17404 (N_17404,N_16408,N_16483);
nand U17405 (N_17405,N_15166,N_15379);
xor U17406 (N_17406,N_15801,N_15609);
and U17407 (N_17407,N_15228,N_15089);
or U17408 (N_17408,N_15026,N_15643);
or U17409 (N_17409,N_16423,N_16489);
nand U17410 (N_17410,N_15096,N_15634);
or U17411 (N_17411,N_15804,N_15911);
or U17412 (N_17412,N_15595,N_16074);
nand U17413 (N_17413,N_16412,N_15004);
or U17414 (N_17414,N_15549,N_15894);
nand U17415 (N_17415,N_15157,N_15703);
nand U17416 (N_17416,N_15565,N_16147);
xnor U17417 (N_17417,N_16193,N_15549);
nor U17418 (N_17418,N_15879,N_15141);
or U17419 (N_17419,N_15394,N_16001);
or U17420 (N_17420,N_15302,N_16002);
or U17421 (N_17421,N_15984,N_15204);
nand U17422 (N_17422,N_15076,N_15392);
and U17423 (N_17423,N_15105,N_15551);
nor U17424 (N_17424,N_16101,N_15343);
and U17425 (N_17425,N_16106,N_15081);
nand U17426 (N_17426,N_15859,N_16489);
nor U17427 (N_17427,N_16296,N_15014);
nor U17428 (N_17428,N_15983,N_16364);
and U17429 (N_17429,N_16389,N_16034);
or U17430 (N_17430,N_15034,N_16420);
xnor U17431 (N_17431,N_15934,N_16455);
nand U17432 (N_17432,N_15777,N_15737);
and U17433 (N_17433,N_15735,N_15909);
or U17434 (N_17434,N_16470,N_15694);
nand U17435 (N_17435,N_15491,N_15403);
nor U17436 (N_17436,N_16045,N_15510);
xor U17437 (N_17437,N_16037,N_15380);
and U17438 (N_17438,N_15818,N_15862);
and U17439 (N_17439,N_16261,N_15256);
or U17440 (N_17440,N_15311,N_15740);
xnor U17441 (N_17441,N_16480,N_15562);
xor U17442 (N_17442,N_15911,N_15066);
nand U17443 (N_17443,N_16310,N_15590);
and U17444 (N_17444,N_16062,N_16407);
nand U17445 (N_17445,N_16455,N_16448);
or U17446 (N_17446,N_15996,N_15381);
or U17447 (N_17447,N_15173,N_16087);
or U17448 (N_17448,N_15061,N_15576);
or U17449 (N_17449,N_15162,N_16030);
nand U17450 (N_17450,N_15691,N_16311);
xor U17451 (N_17451,N_16170,N_15991);
nand U17452 (N_17452,N_16212,N_15738);
xor U17453 (N_17453,N_15400,N_15991);
xor U17454 (N_17454,N_15955,N_15147);
or U17455 (N_17455,N_16140,N_15337);
nand U17456 (N_17456,N_16498,N_15800);
nand U17457 (N_17457,N_15192,N_15961);
or U17458 (N_17458,N_15934,N_15216);
nor U17459 (N_17459,N_15121,N_15759);
nor U17460 (N_17460,N_15386,N_15783);
nor U17461 (N_17461,N_15985,N_15794);
or U17462 (N_17462,N_15127,N_15951);
nand U17463 (N_17463,N_16321,N_16041);
nor U17464 (N_17464,N_16374,N_15873);
nand U17465 (N_17465,N_16005,N_15609);
nor U17466 (N_17466,N_16261,N_15536);
nor U17467 (N_17467,N_15471,N_15359);
and U17468 (N_17468,N_15275,N_15964);
nand U17469 (N_17469,N_16377,N_15343);
nand U17470 (N_17470,N_15635,N_16468);
xor U17471 (N_17471,N_16226,N_15783);
and U17472 (N_17472,N_15955,N_16109);
and U17473 (N_17473,N_15488,N_16177);
or U17474 (N_17474,N_15564,N_15771);
nor U17475 (N_17475,N_15812,N_16428);
and U17476 (N_17476,N_16281,N_15630);
nor U17477 (N_17477,N_15696,N_15399);
xnor U17478 (N_17478,N_15991,N_16376);
nand U17479 (N_17479,N_16270,N_15702);
nor U17480 (N_17480,N_15036,N_16423);
xor U17481 (N_17481,N_15855,N_16262);
xor U17482 (N_17482,N_15891,N_15447);
nor U17483 (N_17483,N_15435,N_15978);
nand U17484 (N_17484,N_15085,N_16362);
nand U17485 (N_17485,N_15723,N_15126);
and U17486 (N_17486,N_16445,N_15651);
or U17487 (N_17487,N_15539,N_15283);
xnor U17488 (N_17488,N_16447,N_15199);
nor U17489 (N_17489,N_15897,N_15493);
xor U17490 (N_17490,N_15937,N_16167);
nor U17491 (N_17491,N_15243,N_15575);
nand U17492 (N_17492,N_15307,N_15469);
and U17493 (N_17493,N_15806,N_16119);
xnor U17494 (N_17494,N_15300,N_16179);
nor U17495 (N_17495,N_15962,N_16227);
and U17496 (N_17496,N_15935,N_15790);
nor U17497 (N_17497,N_16272,N_16088);
nand U17498 (N_17498,N_15656,N_16417);
and U17499 (N_17499,N_16455,N_15426);
or U17500 (N_17500,N_16134,N_15767);
nand U17501 (N_17501,N_15876,N_15514);
nand U17502 (N_17502,N_15295,N_16486);
and U17503 (N_17503,N_15733,N_15989);
or U17504 (N_17504,N_15489,N_15686);
or U17505 (N_17505,N_15269,N_15489);
and U17506 (N_17506,N_15160,N_15386);
xnor U17507 (N_17507,N_15104,N_15841);
xor U17508 (N_17508,N_16051,N_15787);
or U17509 (N_17509,N_16155,N_15830);
and U17510 (N_17510,N_15544,N_15764);
nor U17511 (N_17511,N_15897,N_16357);
nor U17512 (N_17512,N_16194,N_15202);
or U17513 (N_17513,N_16018,N_15994);
and U17514 (N_17514,N_15206,N_16368);
xnor U17515 (N_17515,N_16323,N_15836);
and U17516 (N_17516,N_15446,N_16081);
and U17517 (N_17517,N_15513,N_16374);
nand U17518 (N_17518,N_15686,N_15025);
xor U17519 (N_17519,N_16219,N_16088);
or U17520 (N_17520,N_15923,N_15666);
nor U17521 (N_17521,N_15642,N_15500);
nand U17522 (N_17522,N_15017,N_16185);
xor U17523 (N_17523,N_15209,N_15362);
nand U17524 (N_17524,N_15716,N_15224);
xor U17525 (N_17525,N_15974,N_15062);
xnor U17526 (N_17526,N_16450,N_16436);
or U17527 (N_17527,N_16019,N_15558);
xor U17528 (N_17528,N_15560,N_15505);
xor U17529 (N_17529,N_15412,N_16116);
nand U17530 (N_17530,N_16445,N_16435);
or U17531 (N_17531,N_16316,N_15869);
nor U17532 (N_17532,N_15051,N_15187);
nand U17533 (N_17533,N_16122,N_15159);
or U17534 (N_17534,N_16149,N_16413);
nand U17535 (N_17535,N_16268,N_16403);
xor U17536 (N_17536,N_15244,N_15171);
and U17537 (N_17537,N_16052,N_15432);
or U17538 (N_17538,N_15938,N_15187);
or U17539 (N_17539,N_16469,N_15452);
or U17540 (N_17540,N_15564,N_15728);
and U17541 (N_17541,N_16352,N_15228);
and U17542 (N_17542,N_15734,N_16047);
nor U17543 (N_17543,N_15171,N_15971);
or U17544 (N_17544,N_15371,N_16461);
and U17545 (N_17545,N_15367,N_15268);
nand U17546 (N_17546,N_15506,N_15223);
and U17547 (N_17547,N_16272,N_15685);
nor U17548 (N_17548,N_16420,N_16066);
and U17549 (N_17549,N_15739,N_15832);
and U17550 (N_17550,N_16122,N_15072);
xnor U17551 (N_17551,N_15950,N_15499);
nor U17552 (N_17552,N_15382,N_15001);
or U17553 (N_17553,N_15321,N_15240);
and U17554 (N_17554,N_16472,N_15133);
and U17555 (N_17555,N_16037,N_16212);
nor U17556 (N_17556,N_15967,N_15253);
nand U17557 (N_17557,N_16458,N_15605);
and U17558 (N_17558,N_15671,N_15894);
xnor U17559 (N_17559,N_15834,N_15139);
or U17560 (N_17560,N_15878,N_16362);
xnor U17561 (N_17561,N_16289,N_15099);
and U17562 (N_17562,N_15911,N_15552);
nor U17563 (N_17563,N_15068,N_15568);
or U17564 (N_17564,N_15496,N_15112);
and U17565 (N_17565,N_15376,N_15475);
and U17566 (N_17566,N_15749,N_16230);
or U17567 (N_17567,N_15360,N_15211);
or U17568 (N_17568,N_15499,N_15539);
nor U17569 (N_17569,N_15587,N_15010);
xor U17570 (N_17570,N_15998,N_15305);
or U17571 (N_17571,N_15171,N_16402);
nor U17572 (N_17572,N_15979,N_15744);
or U17573 (N_17573,N_15188,N_15763);
and U17574 (N_17574,N_15277,N_15074);
and U17575 (N_17575,N_16347,N_15220);
nand U17576 (N_17576,N_16176,N_15459);
and U17577 (N_17577,N_15669,N_15859);
xnor U17578 (N_17578,N_16048,N_15354);
xor U17579 (N_17579,N_16041,N_15125);
nand U17580 (N_17580,N_15798,N_15689);
xor U17581 (N_17581,N_15873,N_15955);
nand U17582 (N_17582,N_15398,N_15656);
nand U17583 (N_17583,N_15627,N_15475);
xor U17584 (N_17584,N_15021,N_16000);
xor U17585 (N_17585,N_15113,N_16167);
or U17586 (N_17586,N_15751,N_15048);
and U17587 (N_17587,N_15599,N_15592);
xor U17588 (N_17588,N_16290,N_15804);
xnor U17589 (N_17589,N_15175,N_16403);
nand U17590 (N_17590,N_15754,N_15117);
nand U17591 (N_17591,N_16351,N_15978);
or U17592 (N_17592,N_16432,N_16329);
or U17593 (N_17593,N_15994,N_15744);
or U17594 (N_17594,N_15875,N_16196);
or U17595 (N_17595,N_16230,N_15911);
or U17596 (N_17596,N_16284,N_15781);
or U17597 (N_17597,N_16021,N_15083);
nor U17598 (N_17598,N_15856,N_15734);
and U17599 (N_17599,N_15332,N_15412);
nor U17600 (N_17600,N_15428,N_15783);
nand U17601 (N_17601,N_16046,N_15971);
or U17602 (N_17602,N_15170,N_15689);
nand U17603 (N_17603,N_15371,N_15685);
nand U17604 (N_17604,N_15972,N_15085);
nor U17605 (N_17605,N_15912,N_15085);
xnor U17606 (N_17606,N_15711,N_15503);
nand U17607 (N_17607,N_15659,N_15576);
or U17608 (N_17608,N_15983,N_15346);
and U17609 (N_17609,N_15356,N_16049);
and U17610 (N_17610,N_15975,N_15902);
nor U17611 (N_17611,N_15165,N_15586);
and U17612 (N_17612,N_15035,N_15485);
and U17613 (N_17613,N_16094,N_15406);
or U17614 (N_17614,N_16339,N_15921);
nor U17615 (N_17615,N_15231,N_15808);
nand U17616 (N_17616,N_16464,N_15978);
nor U17617 (N_17617,N_16106,N_15908);
nor U17618 (N_17618,N_16406,N_16286);
xnor U17619 (N_17619,N_16399,N_15038);
nor U17620 (N_17620,N_15248,N_15656);
nor U17621 (N_17621,N_15669,N_16049);
and U17622 (N_17622,N_15728,N_16278);
nand U17623 (N_17623,N_15586,N_15621);
nand U17624 (N_17624,N_16223,N_15300);
nand U17625 (N_17625,N_15539,N_16320);
and U17626 (N_17626,N_16109,N_15806);
nor U17627 (N_17627,N_15724,N_15152);
nor U17628 (N_17628,N_15921,N_16368);
or U17629 (N_17629,N_16083,N_16093);
nand U17630 (N_17630,N_15562,N_15086);
xor U17631 (N_17631,N_15012,N_16023);
xor U17632 (N_17632,N_15667,N_15268);
nand U17633 (N_17633,N_15944,N_16263);
or U17634 (N_17634,N_16472,N_15324);
and U17635 (N_17635,N_15953,N_15397);
and U17636 (N_17636,N_15682,N_16432);
or U17637 (N_17637,N_15951,N_15066);
nor U17638 (N_17638,N_15814,N_16479);
nand U17639 (N_17639,N_15933,N_16212);
xnor U17640 (N_17640,N_15624,N_15726);
nor U17641 (N_17641,N_15897,N_15219);
and U17642 (N_17642,N_15490,N_16344);
nand U17643 (N_17643,N_15822,N_16057);
nand U17644 (N_17644,N_15344,N_15347);
xnor U17645 (N_17645,N_15618,N_16235);
or U17646 (N_17646,N_15164,N_15917);
nor U17647 (N_17647,N_15660,N_15919);
and U17648 (N_17648,N_15867,N_16488);
nor U17649 (N_17649,N_15711,N_15993);
xnor U17650 (N_17650,N_15004,N_15364);
xnor U17651 (N_17651,N_16110,N_16336);
nor U17652 (N_17652,N_16120,N_16367);
or U17653 (N_17653,N_15614,N_15101);
nand U17654 (N_17654,N_15799,N_15532);
and U17655 (N_17655,N_16360,N_15506);
nor U17656 (N_17656,N_16023,N_15931);
nand U17657 (N_17657,N_15650,N_16472);
or U17658 (N_17658,N_15428,N_16353);
nand U17659 (N_17659,N_15551,N_15463);
or U17660 (N_17660,N_15023,N_15947);
nor U17661 (N_17661,N_15992,N_16283);
nand U17662 (N_17662,N_16149,N_15695);
nor U17663 (N_17663,N_16115,N_15394);
xor U17664 (N_17664,N_15572,N_15034);
nor U17665 (N_17665,N_16248,N_16378);
nand U17666 (N_17666,N_15348,N_15920);
nor U17667 (N_17667,N_15916,N_15194);
nor U17668 (N_17668,N_16263,N_16414);
and U17669 (N_17669,N_16275,N_15381);
nand U17670 (N_17670,N_16319,N_16354);
nor U17671 (N_17671,N_16381,N_16180);
and U17672 (N_17672,N_15573,N_15825);
nor U17673 (N_17673,N_15487,N_15057);
xnor U17674 (N_17674,N_16337,N_16390);
xnor U17675 (N_17675,N_16353,N_16265);
nor U17676 (N_17676,N_15452,N_15346);
or U17677 (N_17677,N_16454,N_16115);
or U17678 (N_17678,N_15290,N_16251);
or U17679 (N_17679,N_16325,N_16263);
or U17680 (N_17680,N_15977,N_15505);
nand U17681 (N_17681,N_15921,N_16470);
xnor U17682 (N_17682,N_16039,N_16082);
nor U17683 (N_17683,N_16378,N_15728);
or U17684 (N_17684,N_16459,N_15909);
nand U17685 (N_17685,N_15117,N_15878);
nand U17686 (N_17686,N_16082,N_15915);
or U17687 (N_17687,N_15134,N_15663);
nor U17688 (N_17688,N_15828,N_15100);
xnor U17689 (N_17689,N_15826,N_15559);
nor U17690 (N_17690,N_15867,N_16217);
nand U17691 (N_17691,N_15889,N_16262);
nor U17692 (N_17692,N_15992,N_15233);
xnor U17693 (N_17693,N_16154,N_15072);
xor U17694 (N_17694,N_15007,N_15984);
or U17695 (N_17695,N_15213,N_15295);
or U17696 (N_17696,N_15682,N_15417);
and U17697 (N_17697,N_16468,N_15741);
xor U17698 (N_17698,N_15799,N_15679);
and U17699 (N_17699,N_16045,N_16315);
and U17700 (N_17700,N_16261,N_15095);
nand U17701 (N_17701,N_15107,N_16314);
nor U17702 (N_17702,N_16240,N_16218);
nand U17703 (N_17703,N_15059,N_15478);
nand U17704 (N_17704,N_15913,N_15777);
nor U17705 (N_17705,N_16412,N_15430);
nand U17706 (N_17706,N_16464,N_15820);
nor U17707 (N_17707,N_16429,N_15508);
and U17708 (N_17708,N_15482,N_16200);
nand U17709 (N_17709,N_16106,N_15436);
nand U17710 (N_17710,N_16410,N_16016);
xor U17711 (N_17711,N_15716,N_16044);
nand U17712 (N_17712,N_15132,N_15939);
nor U17713 (N_17713,N_15007,N_16284);
nand U17714 (N_17714,N_15039,N_16452);
nor U17715 (N_17715,N_16012,N_15360);
xor U17716 (N_17716,N_15414,N_16038);
xnor U17717 (N_17717,N_16261,N_15234);
or U17718 (N_17718,N_15764,N_16007);
or U17719 (N_17719,N_16146,N_15580);
nand U17720 (N_17720,N_15636,N_15808);
nor U17721 (N_17721,N_15586,N_16177);
xor U17722 (N_17722,N_15250,N_15024);
nand U17723 (N_17723,N_15303,N_15328);
or U17724 (N_17724,N_15668,N_16393);
and U17725 (N_17725,N_15016,N_16257);
or U17726 (N_17726,N_15302,N_15561);
nand U17727 (N_17727,N_15783,N_15262);
xnor U17728 (N_17728,N_15115,N_15810);
or U17729 (N_17729,N_15627,N_15352);
nor U17730 (N_17730,N_15696,N_15736);
and U17731 (N_17731,N_15078,N_16195);
xnor U17732 (N_17732,N_15095,N_16370);
or U17733 (N_17733,N_15698,N_16466);
nand U17734 (N_17734,N_16046,N_15044);
xor U17735 (N_17735,N_15458,N_16431);
xor U17736 (N_17736,N_16488,N_16386);
xor U17737 (N_17737,N_15750,N_16160);
nor U17738 (N_17738,N_16360,N_15780);
nor U17739 (N_17739,N_15124,N_15499);
nor U17740 (N_17740,N_16418,N_15424);
and U17741 (N_17741,N_15196,N_15487);
xor U17742 (N_17742,N_16487,N_15954);
nor U17743 (N_17743,N_15914,N_16269);
and U17744 (N_17744,N_15765,N_16406);
or U17745 (N_17745,N_15679,N_16103);
xnor U17746 (N_17746,N_16171,N_16016);
or U17747 (N_17747,N_16011,N_16426);
nand U17748 (N_17748,N_15460,N_16049);
and U17749 (N_17749,N_15292,N_15628);
or U17750 (N_17750,N_15193,N_15655);
nor U17751 (N_17751,N_15885,N_16249);
nand U17752 (N_17752,N_16045,N_16186);
and U17753 (N_17753,N_15698,N_16127);
and U17754 (N_17754,N_15036,N_16427);
nor U17755 (N_17755,N_15497,N_15738);
and U17756 (N_17756,N_15500,N_15656);
and U17757 (N_17757,N_16121,N_16392);
and U17758 (N_17758,N_15970,N_15964);
xnor U17759 (N_17759,N_15161,N_15773);
xnor U17760 (N_17760,N_16348,N_15917);
and U17761 (N_17761,N_15423,N_16353);
nor U17762 (N_17762,N_15318,N_15575);
nand U17763 (N_17763,N_15133,N_15213);
xnor U17764 (N_17764,N_15975,N_15186);
xor U17765 (N_17765,N_15111,N_16409);
or U17766 (N_17766,N_15823,N_15535);
nand U17767 (N_17767,N_15693,N_15801);
nor U17768 (N_17768,N_15581,N_15854);
xor U17769 (N_17769,N_15852,N_15842);
nand U17770 (N_17770,N_15564,N_15339);
nor U17771 (N_17771,N_15380,N_16465);
nand U17772 (N_17772,N_15767,N_15491);
or U17773 (N_17773,N_15646,N_16343);
nand U17774 (N_17774,N_16308,N_15365);
nor U17775 (N_17775,N_16118,N_15417);
xnor U17776 (N_17776,N_15994,N_15561);
nand U17777 (N_17777,N_15859,N_15555);
or U17778 (N_17778,N_16144,N_15721);
xnor U17779 (N_17779,N_15196,N_16145);
and U17780 (N_17780,N_16271,N_15702);
nor U17781 (N_17781,N_16115,N_15106);
or U17782 (N_17782,N_15776,N_15756);
nor U17783 (N_17783,N_15839,N_16329);
nor U17784 (N_17784,N_16434,N_15933);
and U17785 (N_17785,N_15778,N_15277);
nor U17786 (N_17786,N_15282,N_15464);
xor U17787 (N_17787,N_15251,N_15279);
xor U17788 (N_17788,N_16356,N_15327);
nand U17789 (N_17789,N_15188,N_15037);
nor U17790 (N_17790,N_15293,N_16278);
nor U17791 (N_17791,N_15866,N_15315);
nand U17792 (N_17792,N_16381,N_15477);
xor U17793 (N_17793,N_15750,N_15018);
nor U17794 (N_17794,N_15255,N_15773);
and U17795 (N_17795,N_15008,N_15174);
xnor U17796 (N_17796,N_16326,N_15841);
or U17797 (N_17797,N_16430,N_15588);
nand U17798 (N_17798,N_16168,N_15172);
and U17799 (N_17799,N_15879,N_15241);
nand U17800 (N_17800,N_15770,N_15776);
nand U17801 (N_17801,N_16220,N_15291);
xnor U17802 (N_17802,N_16263,N_15909);
or U17803 (N_17803,N_15071,N_16312);
or U17804 (N_17804,N_16146,N_15376);
xnor U17805 (N_17805,N_16352,N_15981);
xnor U17806 (N_17806,N_16075,N_15619);
xor U17807 (N_17807,N_15224,N_15250);
and U17808 (N_17808,N_16238,N_15344);
nand U17809 (N_17809,N_16374,N_15745);
nor U17810 (N_17810,N_15215,N_16413);
xnor U17811 (N_17811,N_15511,N_15217);
nor U17812 (N_17812,N_15216,N_16117);
or U17813 (N_17813,N_16034,N_16217);
xor U17814 (N_17814,N_15787,N_15029);
or U17815 (N_17815,N_15053,N_15590);
and U17816 (N_17816,N_15364,N_15946);
nor U17817 (N_17817,N_16464,N_15559);
nor U17818 (N_17818,N_16188,N_16388);
xor U17819 (N_17819,N_15087,N_15965);
or U17820 (N_17820,N_15661,N_15394);
nor U17821 (N_17821,N_15056,N_15537);
and U17822 (N_17822,N_15713,N_15428);
or U17823 (N_17823,N_16161,N_15704);
and U17824 (N_17824,N_16270,N_15497);
nand U17825 (N_17825,N_16165,N_15672);
nand U17826 (N_17826,N_15016,N_16489);
nor U17827 (N_17827,N_16387,N_15088);
nand U17828 (N_17828,N_15968,N_15605);
nor U17829 (N_17829,N_15151,N_15686);
or U17830 (N_17830,N_15712,N_15423);
or U17831 (N_17831,N_15993,N_16313);
xnor U17832 (N_17832,N_16140,N_15184);
and U17833 (N_17833,N_16177,N_15074);
xnor U17834 (N_17834,N_15429,N_15287);
nor U17835 (N_17835,N_15193,N_15155);
nand U17836 (N_17836,N_16413,N_15290);
and U17837 (N_17837,N_15822,N_16261);
nand U17838 (N_17838,N_16435,N_16239);
nor U17839 (N_17839,N_15188,N_15728);
and U17840 (N_17840,N_16406,N_15447);
xnor U17841 (N_17841,N_15619,N_15907);
nor U17842 (N_17842,N_15150,N_15973);
nor U17843 (N_17843,N_15166,N_16074);
xor U17844 (N_17844,N_15819,N_15573);
xnor U17845 (N_17845,N_15038,N_16290);
or U17846 (N_17846,N_16224,N_15234);
xnor U17847 (N_17847,N_16177,N_15025);
nor U17848 (N_17848,N_15140,N_16266);
nand U17849 (N_17849,N_15184,N_15433);
nor U17850 (N_17850,N_15142,N_15133);
nor U17851 (N_17851,N_15622,N_15465);
or U17852 (N_17852,N_15081,N_15253);
and U17853 (N_17853,N_15775,N_15232);
or U17854 (N_17854,N_15540,N_16318);
nor U17855 (N_17855,N_15784,N_15164);
and U17856 (N_17856,N_15275,N_15579);
xor U17857 (N_17857,N_16000,N_15978);
nand U17858 (N_17858,N_15292,N_15338);
nor U17859 (N_17859,N_15615,N_16469);
and U17860 (N_17860,N_15720,N_16253);
nand U17861 (N_17861,N_15965,N_15882);
and U17862 (N_17862,N_15681,N_15890);
and U17863 (N_17863,N_15346,N_15935);
xnor U17864 (N_17864,N_16474,N_15099);
and U17865 (N_17865,N_15865,N_15668);
or U17866 (N_17866,N_16425,N_16019);
nand U17867 (N_17867,N_15372,N_15174);
or U17868 (N_17868,N_16386,N_16325);
xnor U17869 (N_17869,N_16139,N_15845);
nand U17870 (N_17870,N_15173,N_15600);
xnor U17871 (N_17871,N_15979,N_16009);
xor U17872 (N_17872,N_15865,N_16312);
and U17873 (N_17873,N_15137,N_15739);
or U17874 (N_17874,N_15198,N_16496);
xnor U17875 (N_17875,N_15714,N_16001);
and U17876 (N_17876,N_16236,N_16075);
or U17877 (N_17877,N_16254,N_16265);
nand U17878 (N_17878,N_15598,N_15599);
nor U17879 (N_17879,N_15620,N_16386);
nor U17880 (N_17880,N_15989,N_15225);
xnor U17881 (N_17881,N_15444,N_16110);
or U17882 (N_17882,N_15340,N_15740);
nor U17883 (N_17883,N_15326,N_16369);
and U17884 (N_17884,N_15880,N_15220);
nor U17885 (N_17885,N_15295,N_16143);
xnor U17886 (N_17886,N_15766,N_15494);
nand U17887 (N_17887,N_16035,N_15222);
nand U17888 (N_17888,N_15566,N_15851);
xnor U17889 (N_17889,N_15534,N_15689);
and U17890 (N_17890,N_15246,N_15222);
nor U17891 (N_17891,N_15863,N_15523);
and U17892 (N_17892,N_15074,N_16340);
and U17893 (N_17893,N_16412,N_15533);
xnor U17894 (N_17894,N_16289,N_15692);
or U17895 (N_17895,N_16407,N_15377);
or U17896 (N_17896,N_15993,N_16421);
xnor U17897 (N_17897,N_15227,N_16458);
nand U17898 (N_17898,N_16409,N_16040);
xor U17899 (N_17899,N_16194,N_16193);
or U17900 (N_17900,N_15933,N_16318);
or U17901 (N_17901,N_15597,N_16282);
nor U17902 (N_17902,N_16273,N_16110);
and U17903 (N_17903,N_15898,N_15876);
and U17904 (N_17904,N_16040,N_16295);
xnor U17905 (N_17905,N_15194,N_16494);
xor U17906 (N_17906,N_16141,N_16387);
or U17907 (N_17907,N_15497,N_16052);
or U17908 (N_17908,N_16007,N_16300);
xnor U17909 (N_17909,N_15763,N_16017);
xnor U17910 (N_17910,N_15147,N_16196);
xor U17911 (N_17911,N_16189,N_16223);
or U17912 (N_17912,N_16468,N_15628);
and U17913 (N_17913,N_15185,N_15861);
nor U17914 (N_17914,N_16276,N_16487);
and U17915 (N_17915,N_15740,N_15446);
and U17916 (N_17916,N_16452,N_15276);
or U17917 (N_17917,N_15828,N_16279);
and U17918 (N_17918,N_16414,N_16192);
xor U17919 (N_17919,N_15720,N_16061);
nor U17920 (N_17920,N_15744,N_15379);
xor U17921 (N_17921,N_16282,N_16373);
xnor U17922 (N_17922,N_15656,N_15377);
or U17923 (N_17923,N_15161,N_16400);
xnor U17924 (N_17924,N_15845,N_16188);
and U17925 (N_17925,N_16335,N_15031);
nor U17926 (N_17926,N_16312,N_15239);
or U17927 (N_17927,N_15789,N_16107);
xnor U17928 (N_17928,N_15762,N_15904);
nor U17929 (N_17929,N_16047,N_16255);
xor U17930 (N_17930,N_15185,N_15903);
nor U17931 (N_17931,N_15791,N_15884);
nand U17932 (N_17932,N_16378,N_15141);
xnor U17933 (N_17933,N_15380,N_15034);
xor U17934 (N_17934,N_16365,N_15235);
or U17935 (N_17935,N_15991,N_15297);
nor U17936 (N_17936,N_15166,N_15106);
and U17937 (N_17937,N_15606,N_15622);
nand U17938 (N_17938,N_15964,N_16025);
and U17939 (N_17939,N_15913,N_15868);
nor U17940 (N_17940,N_15524,N_15402);
nor U17941 (N_17941,N_15528,N_16225);
xnor U17942 (N_17942,N_16020,N_15106);
nand U17943 (N_17943,N_15478,N_16464);
and U17944 (N_17944,N_16015,N_16271);
nor U17945 (N_17945,N_15328,N_16030);
nand U17946 (N_17946,N_15459,N_16298);
and U17947 (N_17947,N_15876,N_15395);
and U17948 (N_17948,N_15754,N_15829);
nand U17949 (N_17949,N_15199,N_15359);
or U17950 (N_17950,N_15764,N_15410);
or U17951 (N_17951,N_16119,N_15718);
or U17952 (N_17952,N_16461,N_16012);
and U17953 (N_17953,N_15783,N_16383);
nor U17954 (N_17954,N_15627,N_15848);
xnor U17955 (N_17955,N_16470,N_16268);
and U17956 (N_17956,N_15189,N_16228);
nor U17957 (N_17957,N_15238,N_15020);
or U17958 (N_17958,N_16078,N_15845);
nand U17959 (N_17959,N_15007,N_16127);
or U17960 (N_17960,N_16051,N_15030);
nor U17961 (N_17961,N_15254,N_15598);
or U17962 (N_17962,N_15570,N_15915);
nand U17963 (N_17963,N_15356,N_16162);
and U17964 (N_17964,N_15904,N_16187);
xor U17965 (N_17965,N_15532,N_16058);
nand U17966 (N_17966,N_15707,N_16399);
nand U17967 (N_17967,N_15102,N_15095);
nand U17968 (N_17968,N_16406,N_15509);
nand U17969 (N_17969,N_16161,N_15654);
xor U17970 (N_17970,N_15308,N_16483);
or U17971 (N_17971,N_16140,N_16496);
nand U17972 (N_17972,N_16302,N_16313);
nand U17973 (N_17973,N_15993,N_15844);
nor U17974 (N_17974,N_16188,N_15645);
nand U17975 (N_17975,N_16338,N_15759);
or U17976 (N_17976,N_15551,N_15157);
nor U17977 (N_17977,N_15723,N_15228);
nor U17978 (N_17978,N_15411,N_15115);
xnor U17979 (N_17979,N_15708,N_15205);
and U17980 (N_17980,N_15376,N_15058);
or U17981 (N_17981,N_15718,N_15053);
and U17982 (N_17982,N_16095,N_15025);
nor U17983 (N_17983,N_15155,N_15528);
nand U17984 (N_17984,N_16110,N_15922);
nor U17985 (N_17985,N_15463,N_16041);
nor U17986 (N_17986,N_16403,N_15977);
or U17987 (N_17987,N_15472,N_15159);
and U17988 (N_17988,N_15221,N_15945);
xor U17989 (N_17989,N_15015,N_15769);
and U17990 (N_17990,N_16055,N_15614);
nor U17991 (N_17991,N_16069,N_15368);
and U17992 (N_17992,N_15991,N_16024);
nand U17993 (N_17993,N_16495,N_16228);
and U17994 (N_17994,N_15540,N_15624);
xor U17995 (N_17995,N_15121,N_15519);
and U17996 (N_17996,N_15284,N_16025);
nand U17997 (N_17997,N_16355,N_15445);
nor U17998 (N_17998,N_15530,N_15475);
nor U17999 (N_17999,N_15326,N_15063);
and U18000 (N_18000,N_17123,N_16526);
nand U18001 (N_18001,N_16900,N_17440);
or U18002 (N_18002,N_16851,N_17978);
xnor U18003 (N_18003,N_17453,N_17035);
nor U18004 (N_18004,N_16812,N_16510);
or U18005 (N_18005,N_17677,N_17407);
xor U18006 (N_18006,N_16784,N_17504);
nand U18007 (N_18007,N_17061,N_17720);
xnor U18008 (N_18008,N_17853,N_17124);
xnor U18009 (N_18009,N_17591,N_17944);
nand U18010 (N_18010,N_17501,N_17881);
xnor U18011 (N_18011,N_17499,N_16745);
nand U18012 (N_18012,N_17638,N_16999);
nor U18013 (N_18013,N_17997,N_17816);
and U18014 (N_18014,N_16621,N_16930);
or U18015 (N_18015,N_17690,N_17454);
nor U18016 (N_18016,N_17423,N_16765);
nor U18017 (N_18017,N_16619,N_17420);
nor U18018 (N_18018,N_17526,N_17577);
and U18019 (N_18019,N_16558,N_16951);
xnor U18020 (N_18020,N_17076,N_17561);
xor U18021 (N_18021,N_17985,N_17915);
and U18022 (N_18022,N_17362,N_16569);
xnor U18023 (N_18023,N_17954,N_17968);
and U18024 (N_18024,N_16804,N_17823);
or U18025 (N_18025,N_16967,N_17898);
and U18026 (N_18026,N_17599,N_17660);
xor U18027 (N_18027,N_17410,N_17735);
and U18028 (N_18028,N_16799,N_17695);
nand U18029 (N_18029,N_17442,N_17405);
nor U18030 (N_18030,N_17525,N_17641);
nor U18031 (N_18031,N_17136,N_17221);
xor U18032 (N_18032,N_16743,N_17346);
xnor U18033 (N_18033,N_17073,N_17752);
nand U18034 (N_18034,N_17763,N_16889);
nand U18035 (N_18035,N_16964,N_16969);
nor U18036 (N_18036,N_16856,N_17108);
nor U18037 (N_18037,N_17810,N_17839);
or U18038 (N_18038,N_16956,N_16728);
nand U18039 (N_18039,N_16989,N_16600);
nand U18040 (N_18040,N_17072,N_16946);
xnor U18041 (N_18041,N_17884,N_17593);
or U18042 (N_18042,N_16533,N_17305);
nor U18043 (N_18043,N_17976,N_16673);
or U18044 (N_18044,N_16958,N_17357);
or U18045 (N_18045,N_16826,N_17329);
xnor U18046 (N_18046,N_17680,N_16845);
nor U18047 (N_18047,N_17862,N_16892);
or U18048 (N_18048,N_17077,N_16838);
xor U18049 (N_18049,N_16848,N_16737);
nor U18050 (N_18050,N_17718,N_17099);
or U18051 (N_18051,N_17046,N_17324);
or U18052 (N_18052,N_16603,N_16692);
xnor U18053 (N_18053,N_16731,N_16942);
or U18054 (N_18054,N_16780,N_17545);
xnor U18055 (N_18055,N_16870,N_17434);
nand U18056 (N_18056,N_17060,N_17254);
nand U18057 (N_18057,N_16786,N_16522);
or U18058 (N_18058,N_16565,N_17942);
and U18059 (N_18059,N_16920,N_17821);
and U18060 (N_18060,N_17737,N_17700);
nand U18061 (N_18061,N_17578,N_17066);
and U18062 (N_18062,N_17909,N_16871);
and U18063 (N_18063,N_16722,N_16516);
or U18064 (N_18064,N_16759,N_17387);
nor U18065 (N_18065,N_16719,N_16535);
nor U18066 (N_18066,N_17770,N_16730);
and U18067 (N_18067,N_16665,N_17714);
or U18068 (N_18068,N_17907,N_16595);
and U18069 (N_18069,N_16818,N_16664);
nor U18070 (N_18070,N_16615,N_17649);
nand U18071 (N_18071,N_16943,N_17286);
nand U18072 (N_18072,N_17102,N_16772);
nand U18073 (N_18073,N_17117,N_17993);
nand U18074 (N_18074,N_17247,N_17949);
and U18075 (N_18075,N_16977,N_17335);
and U18076 (N_18076,N_17438,N_17597);
nor U18077 (N_18077,N_17151,N_17250);
xnor U18078 (N_18078,N_17492,N_17157);
xnor U18079 (N_18079,N_17027,N_17918);
or U18080 (N_18080,N_17712,N_17041);
xnor U18081 (N_18081,N_17244,N_17683);
nand U18082 (N_18082,N_17604,N_17784);
and U18083 (N_18083,N_17082,N_16923);
nand U18084 (N_18084,N_17984,N_16701);
nand U18085 (N_18085,N_17461,N_16740);
nand U18086 (N_18086,N_17842,N_17302);
and U18087 (N_18087,N_17493,N_17894);
and U18088 (N_18088,N_17606,N_17478);
nor U18089 (N_18089,N_16631,N_17892);
or U18090 (N_18090,N_17512,N_16885);
nand U18091 (N_18091,N_16549,N_16931);
nor U18092 (N_18092,N_17462,N_17857);
or U18093 (N_18093,N_17541,N_16529);
nor U18094 (N_18094,N_17372,N_17742);
or U18095 (N_18095,N_17064,N_16911);
nor U18096 (N_18096,N_16577,N_17836);
nand U18097 (N_18097,N_17347,N_17276);
or U18098 (N_18098,N_16624,N_17464);
and U18099 (N_18099,N_16983,N_16864);
and U18100 (N_18100,N_17893,N_17473);
and U18101 (N_18101,N_16548,N_17111);
or U18102 (N_18102,N_17281,N_17678);
nor U18103 (N_18103,N_17125,N_17673);
nor U18104 (N_18104,N_17794,N_17234);
and U18105 (N_18105,N_16524,N_17001);
or U18106 (N_18106,N_16582,N_16584);
nor U18107 (N_18107,N_17260,N_16693);
nor U18108 (N_18108,N_16674,N_16869);
nand U18109 (N_18109,N_17208,N_16776);
nor U18110 (N_18110,N_17398,N_16820);
xnor U18111 (N_18111,N_16686,N_17910);
or U18112 (N_18112,N_17134,N_16854);
xor U18113 (N_18113,N_17105,N_17148);
xnor U18114 (N_18114,N_17343,N_17518);
nand U18115 (N_18115,N_16610,N_16552);
nor U18116 (N_18116,N_17452,N_17156);
xor U18117 (N_18117,N_17498,N_17081);
nand U18118 (N_18118,N_17052,N_17078);
xor U18119 (N_18119,N_17981,N_17284);
or U18120 (N_18120,N_16844,N_17919);
or U18121 (N_18121,N_17381,N_17962);
or U18122 (N_18122,N_17484,N_17091);
and U18123 (N_18123,N_17882,N_17211);
or U18124 (N_18124,N_16681,N_17249);
and U18125 (N_18125,N_16698,N_17280);
nand U18126 (N_18126,N_17846,N_17349);
and U18127 (N_18127,N_16816,N_16833);
and U18128 (N_18128,N_17559,N_16867);
nor U18129 (N_18129,N_17521,N_16978);
and U18130 (N_18130,N_17608,N_16771);
or U18131 (N_18131,N_17826,N_16625);
and U18132 (N_18132,N_17627,N_17131);
nor U18133 (N_18133,N_17671,N_17710);
nor U18134 (N_18134,N_17598,N_16908);
nand U18135 (N_18135,N_17992,N_16895);
and U18136 (N_18136,N_16909,N_17084);
nand U18137 (N_18137,N_16561,N_17845);
and U18138 (N_18138,N_17725,N_17554);
nand U18139 (N_18139,N_17380,N_17013);
nor U18140 (N_18140,N_17279,N_17093);
and U18141 (N_18141,N_17236,N_17886);
nand U18142 (N_18142,N_17419,N_17418);
and U18143 (N_18143,N_17971,N_17010);
or U18144 (N_18144,N_17797,N_17193);
nand U18145 (N_18145,N_16986,N_17307);
nand U18146 (N_18146,N_17580,N_16509);
or U18147 (N_18147,N_17607,N_16797);
nor U18148 (N_18148,N_16656,N_17414);
nand U18149 (N_18149,N_17549,N_16542);
nand U18150 (N_18150,N_17933,N_17092);
and U18151 (N_18151,N_17564,N_16960);
and U18152 (N_18152,N_17723,N_17183);
nand U18153 (N_18153,N_16865,N_17067);
nand U18154 (N_18154,N_16878,N_17195);
nand U18155 (N_18155,N_17016,N_16773);
or U18156 (N_18156,N_17594,N_17229);
xor U18157 (N_18157,N_17402,N_17864);
or U18158 (N_18158,N_16680,N_17689);
nor U18159 (N_18159,N_16988,N_16970);
or U18160 (N_18160,N_16781,N_16959);
nand U18161 (N_18161,N_17164,N_17548);
nor U18162 (N_18162,N_17255,N_16525);
nand U18163 (N_18163,N_16990,N_17068);
nor U18164 (N_18164,N_17761,N_16840);
or U18165 (N_18165,N_16517,N_17159);
nor U18166 (N_18166,N_17775,N_17474);
and U18167 (N_18167,N_17403,N_17334);
xor U18168 (N_18168,N_16606,N_17257);
xor U18169 (N_18169,N_17167,N_17514);
and U18170 (N_18170,N_16684,N_17535);
or U18171 (N_18171,N_17830,N_17458);
nor U18172 (N_18172,N_17177,N_17358);
xor U18173 (N_18173,N_17022,N_17282);
or U18174 (N_18174,N_16702,N_17270);
nor U18175 (N_18175,N_17231,N_16764);
xnor U18176 (N_18176,N_17391,N_17913);
xor U18177 (N_18177,N_17739,N_17706);
or U18178 (N_18178,N_17232,N_16763);
or U18179 (N_18179,N_17702,N_17506);
xnor U18180 (N_18180,N_17811,N_17767);
nor U18181 (N_18181,N_17018,N_17173);
and U18182 (N_18182,N_17336,N_17020);
nand U18183 (N_18183,N_17098,N_17443);
nand U18184 (N_18184,N_16783,N_16916);
nand U18185 (N_18185,N_17769,N_17668);
or U18186 (N_18186,N_17361,N_17003);
nand U18187 (N_18187,N_16585,N_17259);
and U18188 (N_18188,N_17872,N_16813);
xor U18189 (N_18189,N_16949,N_17153);
and U18190 (N_18190,N_16810,N_17070);
nor U18191 (N_18191,N_16766,N_16837);
and U18192 (N_18192,N_17552,N_17415);
nand U18193 (N_18193,N_16758,N_17116);
or U18194 (N_18194,N_17465,N_17646);
and U18195 (N_18195,N_16636,N_16753);
and U18196 (N_18196,N_16706,N_17180);
xor U18197 (N_18197,N_17294,N_16658);
xnor U18198 (N_18198,N_16563,N_17285);
xor U18199 (N_18199,N_17708,N_16592);
and U18200 (N_18200,N_17652,N_16891);
nand U18201 (N_18201,N_17112,N_17144);
and U18202 (N_18202,N_17531,N_17169);
and U18203 (N_18203,N_16917,N_17746);
xnor U18204 (N_18204,N_17792,N_17332);
nand U18205 (N_18205,N_17719,N_16748);
nor U18206 (N_18206,N_17736,N_16752);
nor U18207 (N_18207,N_16857,N_17146);
nor U18208 (N_18208,N_16770,N_17860);
and U18209 (N_18209,N_17048,N_17309);
nand U18210 (N_18210,N_17328,N_17870);
xor U18211 (N_18211,N_17669,N_16597);
or U18212 (N_18212,N_17914,N_17444);
and U18213 (N_18213,N_16667,N_17378);
or U18214 (N_18214,N_16550,N_17734);
and U18215 (N_18215,N_17936,N_17841);
and U18216 (N_18216,N_17047,N_17198);
xor U18217 (N_18217,N_17371,N_17867);
xor U18218 (N_18218,N_16849,N_17630);
nand U18219 (N_18219,N_17644,N_17687);
nand U18220 (N_18220,N_16630,N_16839);
and U18221 (N_18221,N_16963,N_17929);
or U18222 (N_18222,N_17912,N_16682);
xnor U18223 (N_18223,N_17691,N_17766);
nor U18224 (N_18224,N_17897,N_17982);
and U18225 (N_18225,N_16530,N_17953);
nand U18226 (N_18226,N_17701,N_17777);
nand U18227 (N_18227,N_17565,N_17196);
or U18228 (N_18228,N_17532,N_17296);
nand U18229 (N_18229,N_17460,N_17150);
nor U18230 (N_18230,N_16618,N_17631);
xnor U18231 (N_18231,N_17977,N_16858);
nand U18232 (N_18232,N_16703,N_16905);
xnor U18233 (N_18233,N_17029,N_17560);
nor U18234 (N_18234,N_17824,N_16641);
nor U18235 (N_18235,N_16629,N_17738);
nand U18236 (N_18236,N_17175,N_16705);
nand U18237 (N_18237,N_16755,N_16897);
nor U18238 (N_18238,N_17537,N_16863);
nand U18239 (N_18239,N_16587,N_16578);
and U18240 (N_18240,N_17654,N_17740);
nand U18241 (N_18241,N_16937,N_16623);
and U18242 (N_18242,N_17019,N_17456);
or U18243 (N_18243,N_16635,N_17868);
nand U18244 (N_18244,N_17904,N_16683);
nand U18245 (N_18245,N_16936,N_17017);
or U18246 (N_18246,N_17140,N_17413);
nor U18247 (N_18247,N_16950,N_17051);
nand U18248 (N_18248,N_16501,N_16711);
nand U18249 (N_18249,N_17058,N_17890);
nor U18250 (N_18250,N_17404,N_17980);
nor U18251 (N_18251,N_17203,N_17510);
nor U18252 (N_18252,N_17318,N_17692);
nor U18253 (N_18253,N_17728,N_17901);
nor U18254 (N_18254,N_16852,N_17426);
or U18255 (N_18255,N_17009,N_16880);
and U18256 (N_18256,N_17818,N_17764);
or U18257 (N_18257,N_16778,N_16998);
and U18258 (N_18258,N_16789,N_17130);
nand U18259 (N_18259,N_17781,N_17386);
nor U18260 (N_18260,N_17447,N_17483);
and U18261 (N_18261,N_17840,N_17163);
and U18262 (N_18262,N_16691,N_16769);
or U18263 (N_18263,N_17495,N_16940);
nor U18264 (N_18264,N_17004,N_17697);
xnor U18265 (N_18265,N_16735,N_17553);
nor U18266 (N_18266,N_17204,N_17439);
nand U18267 (N_18267,N_16596,N_17446);
nand U18268 (N_18268,N_17601,N_17288);
nor U18269 (N_18269,N_17972,N_17089);
xnor U18270 (N_18270,N_17471,N_16598);
xor U18271 (N_18271,N_17321,N_17351);
xor U18272 (N_18272,N_17103,N_16901);
or U18273 (N_18273,N_16997,N_17008);
xor U18274 (N_18274,N_17670,N_16634);
nand U18275 (N_18275,N_17433,N_16562);
xor U18276 (N_18276,N_17629,N_17304);
and U18277 (N_18277,N_16898,N_17273);
and U18278 (N_18278,N_17185,N_17875);
nor U18279 (N_18279,N_17620,N_17441);
nand U18280 (N_18280,N_16762,N_17158);
nand U18281 (N_18281,N_17905,N_16834);
nand U18282 (N_18282,N_16751,N_17315);
or U18283 (N_18283,N_17613,N_16828);
or U18284 (N_18284,N_17171,N_16579);
nand U18285 (N_18285,N_17828,N_17876);
or U18286 (N_18286,N_16756,N_17265);
nand U18287 (N_18287,N_17791,N_17724);
xnor U18288 (N_18288,N_17392,N_16645);
or U18289 (N_18289,N_17543,N_17104);
and U18290 (N_18290,N_16873,N_17617);
nor U18291 (N_18291,N_16742,N_17722);
nor U18292 (N_18292,N_17959,N_17119);
nand U18293 (N_18293,N_17705,N_17684);
nor U18294 (N_18294,N_17370,N_17323);
nand U18295 (N_18295,N_16543,N_16707);
and U18296 (N_18296,N_17256,N_16825);
nor U18297 (N_18297,N_17755,N_16754);
xor U18298 (N_18298,N_17534,N_17383);
nor U18299 (N_18299,N_16508,N_17584);
xor U18300 (N_18300,N_17186,N_17586);
nand U18301 (N_18301,N_17220,N_17717);
or U18302 (N_18302,N_17002,N_16609);
nand U18303 (N_18303,N_16557,N_17896);
and U18304 (N_18304,N_17359,N_17240);
nand U18305 (N_18305,N_16685,N_17576);
and U18306 (N_18306,N_17488,N_16503);
nor U18307 (N_18307,N_17160,N_17544);
and U18308 (N_18308,N_16935,N_17516);
and U18309 (N_18309,N_16594,N_17874);
and U18310 (N_18310,N_17348,N_17007);
nand U18311 (N_18311,N_17624,N_17448);
xor U18312 (N_18312,N_17128,N_17263);
xnor U18313 (N_18313,N_17055,N_17165);
or U18314 (N_18314,N_17658,N_17106);
xor U18315 (N_18315,N_17801,N_17952);
or U18316 (N_18316,N_16566,N_17772);
xnor U18317 (N_18317,N_17345,N_16973);
xor U18318 (N_18318,N_16775,N_17573);
nor U18319 (N_18319,N_17216,N_17765);
or U18320 (N_18320,N_16830,N_17809);
xor U18321 (N_18321,N_17437,N_17835);
or U18322 (N_18322,N_17341,N_17074);
or U18323 (N_18323,N_16984,N_17337);
nor U18324 (N_18324,N_17502,N_17973);
xor U18325 (N_18325,N_17485,N_16821);
and U18326 (N_18326,N_17685,N_17212);
nand U18327 (N_18327,N_17034,N_17790);
nand U18328 (N_18328,N_17562,N_17219);
xnor U18329 (N_18329,N_17612,N_17773);
xor U18330 (N_18330,N_17339,N_17353);
nor U18331 (N_18331,N_17648,N_17377);
and U18332 (N_18332,N_16955,N_17239);
and U18333 (N_18333,N_17056,N_17115);
xor U18334 (N_18334,N_16802,N_17109);
nand U18335 (N_18335,N_17258,N_17113);
nor U18336 (N_18336,N_17143,N_16941);
xor U18337 (N_18337,N_17486,N_17401);
nor U18338 (N_18338,N_17477,N_16952);
nand U18339 (N_18339,N_17551,N_17779);
or U18340 (N_18340,N_16532,N_17005);
nand U18341 (N_18341,N_17937,N_17045);
nor U18342 (N_18342,N_17923,N_17563);
nor U18343 (N_18343,N_16717,N_17194);
nand U18344 (N_18344,N_17431,N_17568);
xor U18345 (N_18345,N_16614,N_16612);
or U18346 (N_18346,N_17986,N_17831);
or U18347 (N_18347,N_17069,N_16991);
nor U18348 (N_18348,N_16690,N_17422);
and U18349 (N_18349,N_16734,N_16583);
or U18350 (N_18350,N_16945,N_17651);
nor U18351 (N_18351,N_17807,N_17623);
nand U18352 (N_18352,N_17289,N_17316);
xnor U18353 (N_18353,N_17214,N_17133);
and U18354 (N_18354,N_17364,N_17802);
nand U18355 (N_18355,N_16709,N_17891);
nand U18356 (N_18356,N_17399,N_16914);
or U18357 (N_18357,N_17319,N_16723);
xor U18358 (N_18358,N_16607,N_17911);
xor U18359 (N_18359,N_16500,N_17666);
and U18360 (N_18360,N_16678,N_16894);
nand U18361 (N_18361,N_16659,N_16912);
or U18362 (N_18362,N_17895,N_17928);
xnor U18363 (N_18363,N_17463,N_17955);
xor U18364 (N_18364,N_17759,N_16651);
xnor U18365 (N_18365,N_17015,N_17432);
or U18366 (N_18366,N_17957,N_17253);
nor U18367 (N_18367,N_17815,N_17916);
nor U18368 (N_18368,N_17595,N_16504);
xnor U18369 (N_18369,N_17201,N_17333);
nand U18370 (N_18370,N_17575,N_17813);
or U18371 (N_18371,N_17847,N_17268);
and U18372 (N_18372,N_17331,N_16640);
xnor U18373 (N_18373,N_16724,N_17470);
and U18374 (N_18374,N_17062,N_16853);
nor U18375 (N_18375,N_17344,N_16919);
xor U18376 (N_18376,N_17517,N_17054);
or U18377 (N_18377,N_17030,N_17455);
and U18378 (N_18378,N_17920,N_17162);
nand U18379 (N_18379,N_16729,N_17213);
nor U18380 (N_18380,N_17274,N_17887);
nor U18381 (N_18381,N_17025,N_17948);
nor U18382 (N_18382,N_17476,N_17650);
nand U18383 (N_18383,N_16616,N_17491);
nor U18384 (N_18384,N_17417,N_17472);
xnor U18385 (N_18385,N_17340,N_17667);
nor U18386 (N_18386,N_17118,N_16538);
or U18387 (N_18387,N_17466,N_17489);
and U18388 (N_18388,N_17819,N_17152);
nand U18389 (N_18389,N_17033,N_17057);
nand U18390 (N_18390,N_17424,N_17934);
nor U18391 (N_18391,N_17930,N_17950);
xor U18392 (N_18392,N_17547,N_16761);
and U18393 (N_18393,N_16660,N_17138);
nand U18394 (N_18394,N_17481,N_17833);
xor U18395 (N_18395,N_16666,N_17155);
and U18396 (N_18396,N_16805,N_17487);
and U18397 (N_18397,N_17969,N_17786);
nor U18398 (N_18398,N_17425,N_16980);
and U18399 (N_18399,N_17210,N_17075);
or U18400 (N_18400,N_16671,N_17771);
and U18401 (N_18401,N_17989,N_16886);
nor U18402 (N_18402,N_17961,N_16882);
xor U18403 (N_18403,N_16626,N_16622);
or U18404 (N_18404,N_17663,N_17524);
nor U18405 (N_18405,N_16687,N_16792);
xor U18406 (N_18406,N_16824,N_17379);
or U18407 (N_18407,N_17848,N_16801);
or U18408 (N_18408,N_17850,N_17854);
nand U18409 (N_18409,N_17745,N_17235);
or U18410 (N_18410,N_17696,N_16589);
and U18411 (N_18411,N_17271,N_17330);
nor U18412 (N_18412,N_17513,N_16732);
and U18413 (N_18413,N_16650,N_17127);
xor U18414 (N_18414,N_16588,N_17625);
and U18415 (N_18415,N_17511,N_17050);
nand U18416 (N_18416,N_17587,N_17360);
xor U18417 (N_18417,N_17843,N_16668);
nand U18418 (N_18418,N_16953,N_16974);
xor U18419 (N_18419,N_17400,N_17479);
and U18420 (N_18420,N_17042,N_17375);
nand U18421 (N_18421,N_17096,N_17181);
or U18422 (N_18422,N_16689,N_17311);
xor U18423 (N_18423,N_17983,N_17795);
or U18424 (N_18424,N_16646,N_17184);
and U18425 (N_18425,N_17190,N_16514);
xor U18426 (N_18426,N_17640,N_17979);
nand U18427 (N_18427,N_17793,N_16718);
nand U18428 (N_18428,N_17065,N_17012);
or U18429 (N_18429,N_17088,N_17110);
nor U18430 (N_18430,N_16803,N_17299);
nand U18431 (N_18431,N_17931,N_16720);
nand U18432 (N_18432,N_17783,N_17662);
nor U18433 (N_18433,N_17744,N_17283);
and U18434 (N_18434,N_17557,N_16904);
xnor U18435 (N_18435,N_16884,N_16938);
or U18436 (N_18436,N_17963,N_17246);
xnor U18437 (N_18437,N_16994,N_17664);
xor U18438 (N_18438,N_17675,N_17197);
nor U18439 (N_18439,N_16727,N_17788);
and U18440 (N_18440,N_17292,N_17806);
or U18441 (N_18441,N_17228,N_17086);
xor U18442 (N_18442,N_17393,N_17778);
xor U18443 (N_18443,N_17179,N_17226);
and U18444 (N_18444,N_17409,N_17233);
nand U18445 (N_18445,N_17428,N_17602);
or U18446 (N_18446,N_16918,N_17951);
xnor U18447 (N_18447,N_17605,N_17161);
or U18448 (N_18448,N_16648,N_17611);
or U18449 (N_18449,N_16899,N_17338);
nor U18450 (N_18450,N_17166,N_17411);
and U18451 (N_18451,N_16661,N_17202);
nor U18452 (N_18452,N_17326,N_17024);
and U18453 (N_18453,N_16921,N_17634);
xor U18454 (N_18454,N_17043,N_17805);
or U18455 (N_18455,N_16971,N_17320);
and U18456 (N_18456,N_16715,N_16750);
xnor U18457 (N_18457,N_17408,N_17827);
nor U18458 (N_18458,N_17590,N_17924);
nor U18459 (N_18459,N_16688,N_17178);
xnor U18460 (N_18460,N_17694,N_17698);
or U18461 (N_18461,N_17039,N_17053);
xnor U18462 (N_18462,N_17366,N_17275);
or U18463 (N_18463,N_17656,N_17509);
xnor U18464 (N_18464,N_16972,N_16846);
or U18465 (N_18465,N_17751,N_16511);
nand U18466 (N_18466,N_16637,N_16862);
or U18467 (N_18467,N_17938,N_16713);
nand U18468 (N_18468,N_17114,N_17031);
or U18469 (N_18469,N_16982,N_17365);
nor U18470 (N_18470,N_17312,N_16866);
nand U18471 (N_18471,N_17880,N_16591);
nand U18472 (N_18472,N_17369,N_17558);
nand U18473 (N_18473,N_17536,N_17291);
xor U18474 (N_18474,N_16992,N_16604);
and U18475 (N_18475,N_17796,N_16835);
xor U18476 (N_18476,N_17147,N_17715);
and U18477 (N_18477,N_17122,N_17374);
or U18478 (N_18478,N_16677,N_16655);
and U18479 (N_18479,N_17382,N_17036);
and U18480 (N_18480,N_17126,N_17154);
nand U18481 (N_18481,N_17237,N_17799);
xor U18482 (N_18482,N_17637,N_16893);
and U18483 (N_18483,N_17527,N_17429);
and U18484 (N_18484,N_17457,N_17500);
nor U18485 (N_18485,N_16617,N_16788);
nor U18486 (N_18486,N_16757,N_17610);
and U18487 (N_18487,N_17626,N_17191);
nand U18488 (N_18488,N_16652,N_16965);
xor U18489 (N_18489,N_16793,N_17303);
or U18490 (N_18490,N_17659,N_17095);
nand U18491 (N_18491,N_17657,N_16957);
nor U18492 (N_18492,N_16896,N_17800);
nand U18493 (N_18493,N_17879,N_16979);
nand U18494 (N_18494,N_16554,N_16791);
nor U18495 (N_18495,N_17248,N_16586);
or U18496 (N_18496,N_17217,N_17430);
and U18497 (N_18497,N_17956,N_17583);
xor U18498 (N_18498,N_17436,N_17990);
and U18499 (N_18499,N_17661,N_16795);
nor U18500 (N_18500,N_17932,N_17603);
and U18501 (N_18501,N_17206,N_16782);
and U18502 (N_18502,N_17427,N_16736);
or U18503 (N_18503,N_16574,N_17635);
and U18504 (N_18504,N_17988,N_16794);
nand U18505 (N_18505,N_16696,N_17100);
and U18506 (N_18506,N_17200,N_16739);
nor U18507 (N_18507,N_17519,N_16541);
xor U18508 (N_18508,N_16832,N_16874);
nor U18509 (N_18509,N_16842,N_16571);
nand U18510 (N_18510,N_17287,N_17459);
and U18511 (N_18511,N_17028,N_17699);
and U18512 (N_18512,N_17496,N_17592);
and U18513 (N_18513,N_16537,N_17182);
or U18514 (N_18514,N_17965,N_16877);
or U18515 (N_18515,N_16814,N_17925);
or U18516 (N_18516,N_16902,N_17782);
nand U18517 (N_18517,N_17906,N_17555);
nor U18518 (N_18518,N_17829,N_17676);
and U18519 (N_18519,N_17266,N_17885);
nand U18520 (N_18520,N_16527,N_17727);
nand U18521 (N_18521,N_17533,N_17747);
and U18522 (N_18522,N_17168,N_16890);
nor U18523 (N_18523,N_17482,N_17037);
and U18524 (N_18524,N_17014,N_16855);
nand U18525 (N_18525,N_17451,N_16590);
xor U18526 (N_18526,N_16551,N_17674);
nor U18527 (N_18527,N_16939,N_17899);
and U18528 (N_18528,N_17681,N_17633);
nand U18529 (N_18529,N_16547,N_16539);
and U18530 (N_18530,N_16553,N_16925);
or U18531 (N_18531,N_17803,N_17999);
xnor U18532 (N_18532,N_16746,N_16580);
nor U18533 (N_18533,N_17149,N_17528);
nand U18534 (N_18534,N_17903,N_17817);
nand U18535 (N_18535,N_17469,N_16887);
or U18536 (N_18536,N_17242,N_16695);
or U18537 (N_18537,N_16975,N_17515);
and U18538 (N_18538,N_16841,N_17542);
and U18539 (N_18539,N_17205,N_16639);
or U18540 (N_18540,N_17582,N_17679);
nand U18541 (N_18541,N_16861,N_17609);
nor U18542 (N_18542,N_17820,N_16714);
xnor U18543 (N_18543,N_16906,N_16774);
nor U18544 (N_18544,N_17926,N_17011);
nor U18545 (N_18545,N_16575,N_16534);
nand U18546 (N_18546,N_17958,N_17356);
and U18547 (N_18547,N_17390,N_17373);
xor U18548 (N_18548,N_17272,N_17585);
xor U18549 (N_18549,N_16747,N_16947);
and U18550 (N_18550,N_17450,N_17970);
nor U18551 (N_18551,N_17812,N_17137);
nand U18552 (N_18552,N_17269,N_16859);
xnor U18553 (N_18553,N_17588,N_17863);
and U18554 (N_18554,N_17888,N_16836);
and U18555 (N_18555,N_17352,N_17566);
and U18556 (N_18556,N_17021,N_16922);
nor U18557 (N_18557,N_17750,N_16515);
xor U18558 (N_18558,N_17449,N_16796);
or U18559 (N_18559,N_17300,N_16663);
nor U18560 (N_18560,N_16669,N_17943);
nand U18561 (N_18561,N_17861,N_16767);
or U18562 (N_18562,N_16850,N_17094);
or U18563 (N_18563,N_16829,N_16749);
nor U18564 (N_18564,N_17223,N_17416);
and U18565 (N_18565,N_17306,N_17176);
or U18566 (N_18566,N_16926,N_16638);
nand U18567 (N_18567,N_17384,N_17614);
or U18568 (N_18568,N_17768,N_16611);
or U18569 (N_18569,N_17480,N_17785);
and U18570 (N_18570,N_17000,N_16883);
nor U18571 (N_18571,N_17704,N_17278);
or U18572 (N_18572,N_16785,N_17855);
and U18573 (N_18573,N_16644,N_17688);
or U18574 (N_18574,N_17530,N_17758);
nand U18575 (N_18575,N_17902,N_16868);
xor U18576 (N_18576,N_17632,N_17224);
nand U18577 (N_18577,N_17787,N_16760);
nor U18578 (N_18578,N_16823,N_17974);
xor U18579 (N_18579,N_17574,N_16768);
nor U18580 (N_18580,N_16523,N_17693);
and U18581 (N_18581,N_16831,N_16995);
or U18582 (N_18582,N_16608,N_17798);
nor U18583 (N_18583,N_16996,N_16843);
nand U18584 (N_18584,N_17639,N_17686);
and U18585 (N_18585,N_16556,N_16576);
xor U18586 (N_18586,N_17743,N_16632);
nor U18587 (N_18587,N_17760,N_17729);
nand U18588 (N_18588,N_17825,N_17120);
nor U18589 (N_18589,N_17435,N_17227);
xnor U18590 (N_18590,N_17789,N_17310);
xor U18591 (N_18591,N_17085,N_17571);
and U18592 (N_18592,N_16540,N_16697);
and U18593 (N_18593,N_17188,N_16726);
and U18594 (N_18594,N_17350,N_16913);
and U18595 (N_18595,N_17921,N_17121);
xnor U18596 (N_18596,N_17367,N_17317);
or U18597 (N_18597,N_17245,N_16662);
or U18598 (N_18598,N_17927,N_17083);
nor U18599 (N_18599,N_17569,N_17642);
xor U18600 (N_18600,N_17129,N_17966);
and U18601 (N_18601,N_17878,N_17368);
and U18602 (N_18602,N_17187,N_17267);
and U18603 (N_18603,N_16976,N_17733);
nand U18604 (N_18604,N_17757,N_16822);
xor U18605 (N_18605,N_16777,N_16944);
nor U18606 (N_18606,N_17730,N_16654);
nor U18607 (N_18607,N_17445,N_17230);
and U18608 (N_18608,N_17189,N_17023);
xor U18609 (N_18609,N_16694,N_17837);
and U18610 (N_18610,N_16502,N_17858);
xor U18611 (N_18611,N_16672,N_17908);
nor U18612 (N_18612,N_16546,N_17780);
or U18613 (N_18613,N_16649,N_17505);
nor U18614 (N_18614,N_16601,N_16699);
and U18615 (N_18615,N_17941,N_17394);
or U18616 (N_18616,N_16910,N_17497);
xor U18617 (N_18617,N_17297,N_16741);
and U18618 (N_18618,N_17945,N_16744);
nor U18619 (N_18619,N_16555,N_17388);
nor U18620 (N_18620,N_17539,N_17600);
nand U18621 (N_18621,N_17540,N_17314);
and U18622 (N_18622,N_16948,N_17475);
nor U18623 (N_18623,N_17355,N_17922);
and U18624 (N_18624,N_17960,N_17529);
xnor U18625 (N_18625,N_17538,N_17238);
or U18626 (N_18626,N_16716,N_17762);
nand U18627 (N_18627,N_17354,N_16513);
nor U18628 (N_18628,N_16512,N_17709);
xor U18629 (N_18629,N_17753,N_17218);
and U18630 (N_18630,N_17917,N_17618);
nand U18631 (N_18631,N_16815,N_17856);
nand U18632 (N_18632,N_16643,N_17207);
nor U18633 (N_18633,N_17071,N_17508);
or U18634 (N_18634,N_16675,N_17814);
xnor U18635 (N_18635,N_17290,N_16581);
xor U18636 (N_18636,N_16653,N_16934);
and U18637 (N_18637,N_16819,N_16568);
nand U18638 (N_18638,N_17199,N_17040);
nor U18639 (N_18639,N_17090,N_16924);
and U18640 (N_18640,N_16875,N_16800);
xor U18641 (N_18641,N_16790,N_17038);
or U18642 (N_18642,N_17342,N_16993);
xor U18643 (N_18643,N_17834,N_16633);
or U18644 (N_18644,N_16700,N_16712);
or U18645 (N_18645,N_17832,N_17946);
nand U18646 (N_18646,N_17264,N_17101);
and U18647 (N_18647,N_17987,N_16721);
xor U18648 (N_18648,N_16506,N_17672);
nor U18649 (N_18649,N_17376,N_17277);
xnor U18650 (N_18650,N_16520,N_17215);
xor U18651 (N_18651,N_17859,N_16620);
or U18652 (N_18652,N_17774,N_16564);
nand U18653 (N_18653,N_17939,N_17741);
xor U18654 (N_18654,N_16738,N_17703);
or U18655 (N_18655,N_16670,N_17301);
or U18656 (N_18656,N_16966,N_16981);
nor U18657 (N_18657,N_17522,N_16879);
or U18658 (N_18658,N_17647,N_16572);
xnor U18659 (N_18659,N_17844,N_17252);
nand U18660 (N_18660,N_17822,N_17139);
nand U18661 (N_18661,N_16807,N_16605);
xor U18662 (N_18662,N_17589,N_17251);
or U18663 (N_18663,N_17995,N_16518);
xnor U18664 (N_18664,N_17883,N_17726);
nor U18665 (N_18665,N_17655,N_16808);
nor U18666 (N_18666,N_17412,N_17385);
and U18667 (N_18667,N_17998,N_17507);
nand U18668 (N_18668,N_17523,N_16657);
nor U18669 (N_18669,N_17241,N_17395);
xor U18670 (N_18670,N_17494,N_16531);
xor U18671 (N_18671,N_17996,N_16708);
nor U18672 (N_18672,N_17107,N_17327);
nor U18673 (N_18673,N_16733,N_17877);
and U18674 (N_18674,N_17621,N_17653);
nor U18675 (N_18675,N_17313,N_16903);
nor U18676 (N_18676,N_16505,N_16642);
nand U18677 (N_18677,N_16627,N_17994);
nor U18678 (N_18678,N_17940,N_16987);
nand U18679 (N_18679,N_17520,N_17225);
and U18680 (N_18680,N_16915,N_17293);
and U18681 (N_18681,N_17032,N_16599);
and U18682 (N_18682,N_17049,N_17581);
nand U18683 (N_18683,N_17776,N_16704);
and U18684 (N_18684,N_16570,N_16985);
or U18685 (N_18685,N_17873,N_17869);
nor U18686 (N_18686,N_17006,N_16560);
nand U18687 (N_18687,N_17141,N_17711);
and U18688 (N_18688,N_17947,N_16847);
nor U18689 (N_18689,N_17804,N_16559);
xnor U18690 (N_18690,N_17749,N_16932);
or U18691 (N_18691,N_17406,N_17636);
or U18692 (N_18692,N_16827,N_17967);
nand U18693 (N_18693,N_17087,N_16860);
and U18694 (N_18694,N_16519,N_17503);
xor U18695 (N_18695,N_16593,N_17026);
nand U18696 (N_18696,N_17209,N_17991);
and U18697 (N_18697,N_17871,N_16567);
xnor U18698 (N_18698,N_16881,N_17145);
nor U18699 (N_18699,N_16872,N_17059);
or U18700 (N_18700,N_17570,N_16962);
nand U18701 (N_18701,N_17322,N_16787);
nor U18702 (N_18702,N_16806,N_17754);
nor U18703 (N_18703,N_17325,N_17556);
nand U18704 (N_18704,N_17615,N_17389);
nor U18705 (N_18705,N_16961,N_16725);
or U18706 (N_18706,N_17261,N_17097);
and U18707 (N_18707,N_17866,N_17298);
xnor U18708 (N_18708,N_17132,N_17851);
and U18709 (N_18709,N_17616,N_17975);
nand U18710 (N_18710,N_16927,N_17308);
or U18711 (N_18711,N_17170,N_17865);
nand U18712 (N_18712,N_17808,N_17172);
or U18713 (N_18713,N_16809,N_17628);
nand U18714 (N_18714,N_16676,N_17080);
nor U18715 (N_18715,N_16817,N_16907);
nor U18716 (N_18716,N_17935,N_16545);
and U18717 (N_18717,N_17567,N_16798);
and U18718 (N_18718,N_17707,N_17964);
and U18719 (N_18719,N_16876,N_16602);
and U18720 (N_18720,N_16507,N_17622);
nand U18721 (N_18721,N_17748,N_17396);
nor U18722 (N_18722,N_17192,N_16628);
or U18723 (N_18723,N_17363,N_17262);
and U18724 (N_18724,N_16573,N_16888);
xor U18725 (N_18725,N_16521,N_16933);
and U18726 (N_18726,N_17619,N_17174);
and U18727 (N_18727,N_17243,N_17079);
nor U18728 (N_18728,N_17900,N_17838);
or U18729 (N_18729,N_17645,N_17682);
nand U18730 (N_18730,N_17572,N_17643);
nor U18731 (N_18731,N_17849,N_17142);
and U18732 (N_18732,N_16928,N_16647);
or U18733 (N_18733,N_16528,N_16954);
and U18734 (N_18734,N_17579,N_16968);
nand U18735 (N_18735,N_16613,N_17716);
or U18736 (N_18736,N_17889,N_17397);
or U18737 (N_18737,N_17731,N_17665);
or U18738 (N_18738,N_16779,N_17550);
xnor U18739 (N_18739,N_17490,N_16536);
nand U18740 (N_18740,N_16544,N_16811);
xor U18741 (N_18741,N_17852,N_17135);
nand U18742 (N_18742,N_17421,N_17721);
nor U18743 (N_18743,N_16679,N_17063);
or U18744 (N_18744,N_17295,N_17044);
or U18745 (N_18745,N_17596,N_17713);
and U18746 (N_18746,N_17756,N_17468);
nor U18747 (N_18747,N_16929,N_17467);
or U18748 (N_18748,N_17222,N_16710);
and U18749 (N_18749,N_17732,N_17546);
or U18750 (N_18750,N_16813,N_16657);
nand U18751 (N_18751,N_17520,N_17783);
nand U18752 (N_18752,N_17923,N_16784);
xor U18753 (N_18753,N_17388,N_17132);
nor U18754 (N_18754,N_17961,N_16914);
nor U18755 (N_18755,N_17426,N_17543);
and U18756 (N_18756,N_17671,N_17171);
xor U18757 (N_18757,N_17250,N_17141);
nor U18758 (N_18758,N_17254,N_16770);
or U18759 (N_18759,N_17902,N_16608);
and U18760 (N_18760,N_16759,N_17471);
or U18761 (N_18761,N_17628,N_17351);
xnor U18762 (N_18762,N_16890,N_17250);
or U18763 (N_18763,N_16512,N_17349);
nor U18764 (N_18764,N_17969,N_16526);
and U18765 (N_18765,N_17380,N_17552);
and U18766 (N_18766,N_16745,N_17390);
nand U18767 (N_18767,N_17515,N_17040);
xor U18768 (N_18768,N_17056,N_17107);
and U18769 (N_18769,N_16882,N_17380);
xor U18770 (N_18770,N_17879,N_16900);
or U18771 (N_18771,N_16712,N_17950);
nand U18772 (N_18772,N_16918,N_17658);
or U18773 (N_18773,N_17505,N_17761);
or U18774 (N_18774,N_17210,N_16577);
xor U18775 (N_18775,N_16744,N_16647);
and U18776 (N_18776,N_17008,N_17827);
and U18777 (N_18777,N_16757,N_17749);
nor U18778 (N_18778,N_17170,N_17917);
and U18779 (N_18779,N_16754,N_17514);
nand U18780 (N_18780,N_17879,N_17200);
or U18781 (N_18781,N_17068,N_17663);
or U18782 (N_18782,N_17989,N_17283);
xor U18783 (N_18783,N_17560,N_17748);
or U18784 (N_18784,N_17867,N_16662);
nand U18785 (N_18785,N_16675,N_17158);
or U18786 (N_18786,N_16536,N_16968);
or U18787 (N_18787,N_16988,N_16594);
or U18788 (N_18788,N_17991,N_17333);
nand U18789 (N_18789,N_17437,N_17847);
nor U18790 (N_18790,N_16916,N_17005);
xor U18791 (N_18791,N_16845,N_17067);
or U18792 (N_18792,N_17545,N_17297);
nand U18793 (N_18793,N_17584,N_17082);
nor U18794 (N_18794,N_16695,N_17202);
and U18795 (N_18795,N_17111,N_17040);
xnor U18796 (N_18796,N_17700,N_16582);
xor U18797 (N_18797,N_17695,N_17008);
nand U18798 (N_18798,N_17671,N_17057);
xnor U18799 (N_18799,N_17072,N_16845);
xor U18800 (N_18800,N_17749,N_16511);
or U18801 (N_18801,N_16517,N_16798);
xor U18802 (N_18802,N_17294,N_17751);
nor U18803 (N_18803,N_17861,N_17357);
or U18804 (N_18804,N_17978,N_17444);
xor U18805 (N_18805,N_17825,N_17136);
or U18806 (N_18806,N_16854,N_17583);
and U18807 (N_18807,N_17671,N_16914);
xor U18808 (N_18808,N_17229,N_17422);
or U18809 (N_18809,N_17819,N_16695);
and U18810 (N_18810,N_17594,N_16830);
xnor U18811 (N_18811,N_17570,N_17098);
nor U18812 (N_18812,N_16577,N_17986);
and U18813 (N_18813,N_17994,N_16650);
and U18814 (N_18814,N_17461,N_17381);
and U18815 (N_18815,N_17916,N_17074);
and U18816 (N_18816,N_17689,N_17962);
nand U18817 (N_18817,N_17220,N_16876);
nand U18818 (N_18818,N_17096,N_16875);
or U18819 (N_18819,N_17002,N_17781);
nand U18820 (N_18820,N_16982,N_17451);
and U18821 (N_18821,N_17860,N_16614);
and U18822 (N_18822,N_17606,N_17748);
xor U18823 (N_18823,N_17846,N_17234);
nor U18824 (N_18824,N_16827,N_16906);
nor U18825 (N_18825,N_16927,N_16729);
nor U18826 (N_18826,N_17947,N_17034);
or U18827 (N_18827,N_17078,N_16944);
xor U18828 (N_18828,N_17871,N_16613);
and U18829 (N_18829,N_17270,N_17985);
and U18830 (N_18830,N_16565,N_17979);
nor U18831 (N_18831,N_17168,N_17434);
nor U18832 (N_18832,N_16686,N_17070);
nand U18833 (N_18833,N_16956,N_17510);
or U18834 (N_18834,N_17052,N_17463);
xnor U18835 (N_18835,N_17429,N_17335);
and U18836 (N_18836,N_17908,N_16839);
nand U18837 (N_18837,N_17503,N_17802);
nor U18838 (N_18838,N_17163,N_17194);
nand U18839 (N_18839,N_16898,N_16547);
xnor U18840 (N_18840,N_16778,N_17138);
or U18841 (N_18841,N_17801,N_17854);
nand U18842 (N_18842,N_17867,N_16882);
or U18843 (N_18843,N_17106,N_17220);
or U18844 (N_18844,N_17873,N_17655);
nand U18845 (N_18845,N_16555,N_17268);
nor U18846 (N_18846,N_17630,N_16906);
and U18847 (N_18847,N_17332,N_17263);
nand U18848 (N_18848,N_17766,N_16568);
nor U18849 (N_18849,N_17297,N_17621);
nand U18850 (N_18850,N_17532,N_17000);
nor U18851 (N_18851,N_17199,N_17230);
nor U18852 (N_18852,N_17281,N_17888);
xor U18853 (N_18853,N_16538,N_17537);
and U18854 (N_18854,N_17504,N_16779);
nand U18855 (N_18855,N_17869,N_16956);
nor U18856 (N_18856,N_17408,N_17398);
xor U18857 (N_18857,N_17353,N_17006);
nor U18858 (N_18858,N_17861,N_17008);
nor U18859 (N_18859,N_16700,N_17094);
and U18860 (N_18860,N_16834,N_16742);
xnor U18861 (N_18861,N_17393,N_17366);
and U18862 (N_18862,N_17353,N_16595);
xnor U18863 (N_18863,N_16611,N_17307);
or U18864 (N_18864,N_17002,N_16861);
xor U18865 (N_18865,N_16749,N_17735);
nor U18866 (N_18866,N_16545,N_16606);
and U18867 (N_18867,N_17349,N_17229);
nand U18868 (N_18868,N_17857,N_17187);
nand U18869 (N_18869,N_16770,N_16990);
nand U18870 (N_18870,N_17520,N_16805);
or U18871 (N_18871,N_16836,N_16773);
xor U18872 (N_18872,N_16944,N_16636);
nand U18873 (N_18873,N_17712,N_17193);
and U18874 (N_18874,N_17212,N_17705);
nand U18875 (N_18875,N_17507,N_17798);
and U18876 (N_18876,N_17320,N_16757);
nor U18877 (N_18877,N_17069,N_17633);
and U18878 (N_18878,N_17353,N_17045);
nor U18879 (N_18879,N_17850,N_17205);
nand U18880 (N_18880,N_17235,N_16856);
xor U18881 (N_18881,N_17080,N_17433);
xor U18882 (N_18882,N_16804,N_16845);
xor U18883 (N_18883,N_17503,N_17153);
and U18884 (N_18884,N_16745,N_17264);
xor U18885 (N_18885,N_16636,N_16931);
xnor U18886 (N_18886,N_17867,N_17713);
or U18887 (N_18887,N_17825,N_17354);
or U18888 (N_18888,N_17282,N_17478);
xnor U18889 (N_18889,N_16651,N_17338);
or U18890 (N_18890,N_16681,N_16662);
xor U18891 (N_18891,N_16893,N_16933);
nand U18892 (N_18892,N_17941,N_17980);
or U18893 (N_18893,N_17545,N_17454);
and U18894 (N_18894,N_17502,N_17781);
or U18895 (N_18895,N_16564,N_17396);
xor U18896 (N_18896,N_17427,N_16822);
and U18897 (N_18897,N_17713,N_16764);
xnor U18898 (N_18898,N_16619,N_17882);
nor U18899 (N_18899,N_17549,N_16586);
xnor U18900 (N_18900,N_17261,N_17230);
nand U18901 (N_18901,N_16967,N_17253);
nand U18902 (N_18902,N_17390,N_17168);
and U18903 (N_18903,N_17598,N_17253);
or U18904 (N_18904,N_17150,N_16532);
xor U18905 (N_18905,N_17288,N_16618);
or U18906 (N_18906,N_16965,N_17759);
nor U18907 (N_18907,N_16506,N_16987);
and U18908 (N_18908,N_17823,N_17772);
or U18909 (N_18909,N_17016,N_17721);
or U18910 (N_18910,N_17057,N_17438);
nor U18911 (N_18911,N_16564,N_17505);
nor U18912 (N_18912,N_17090,N_16842);
or U18913 (N_18913,N_17201,N_17030);
and U18914 (N_18914,N_16634,N_17063);
xnor U18915 (N_18915,N_16649,N_17283);
or U18916 (N_18916,N_16822,N_17694);
and U18917 (N_18917,N_17382,N_16937);
nand U18918 (N_18918,N_17309,N_17907);
and U18919 (N_18919,N_16753,N_16511);
or U18920 (N_18920,N_17560,N_16820);
nand U18921 (N_18921,N_17142,N_17888);
nor U18922 (N_18922,N_17002,N_16906);
or U18923 (N_18923,N_17262,N_17253);
nand U18924 (N_18924,N_17848,N_17665);
nand U18925 (N_18925,N_17058,N_17545);
xnor U18926 (N_18926,N_17032,N_16885);
nand U18927 (N_18927,N_17157,N_17907);
and U18928 (N_18928,N_17369,N_17690);
xor U18929 (N_18929,N_17300,N_17341);
xnor U18930 (N_18930,N_17927,N_17949);
xnor U18931 (N_18931,N_17874,N_17115);
xor U18932 (N_18932,N_17884,N_17128);
nand U18933 (N_18933,N_16847,N_16957);
xor U18934 (N_18934,N_17403,N_17388);
nor U18935 (N_18935,N_16684,N_16627);
and U18936 (N_18936,N_16940,N_17551);
nor U18937 (N_18937,N_16985,N_17326);
and U18938 (N_18938,N_16519,N_17606);
xnor U18939 (N_18939,N_17168,N_17931);
nor U18940 (N_18940,N_17716,N_16869);
nand U18941 (N_18941,N_17227,N_17384);
nor U18942 (N_18942,N_16959,N_17256);
or U18943 (N_18943,N_17730,N_17594);
or U18944 (N_18944,N_17603,N_17586);
xnor U18945 (N_18945,N_17855,N_17369);
and U18946 (N_18946,N_17322,N_17241);
nand U18947 (N_18947,N_17114,N_17136);
and U18948 (N_18948,N_16636,N_17177);
nand U18949 (N_18949,N_17990,N_17896);
xnor U18950 (N_18950,N_17524,N_16849);
nor U18951 (N_18951,N_16870,N_16792);
nor U18952 (N_18952,N_16768,N_16818);
or U18953 (N_18953,N_17182,N_16518);
and U18954 (N_18954,N_16632,N_17859);
and U18955 (N_18955,N_17309,N_16955);
and U18956 (N_18956,N_17980,N_16829);
and U18957 (N_18957,N_16647,N_17456);
nor U18958 (N_18958,N_16611,N_17742);
and U18959 (N_18959,N_17362,N_17099);
nor U18960 (N_18960,N_16523,N_16546);
xor U18961 (N_18961,N_17285,N_17457);
and U18962 (N_18962,N_16990,N_17664);
and U18963 (N_18963,N_16572,N_17944);
nand U18964 (N_18964,N_17988,N_17500);
nand U18965 (N_18965,N_16770,N_17991);
and U18966 (N_18966,N_17646,N_17692);
xnor U18967 (N_18967,N_17092,N_16836);
nand U18968 (N_18968,N_17491,N_17433);
or U18969 (N_18969,N_17333,N_17035);
or U18970 (N_18970,N_16785,N_16580);
nand U18971 (N_18971,N_16922,N_16885);
and U18972 (N_18972,N_17730,N_17327);
xnor U18973 (N_18973,N_17981,N_16545);
and U18974 (N_18974,N_17192,N_17029);
and U18975 (N_18975,N_16944,N_16691);
nor U18976 (N_18976,N_17512,N_16840);
nand U18977 (N_18977,N_16679,N_16593);
or U18978 (N_18978,N_16796,N_17751);
or U18979 (N_18979,N_17912,N_17318);
xor U18980 (N_18980,N_16707,N_16573);
nor U18981 (N_18981,N_17557,N_17336);
and U18982 (N_18982,N_17886,N_17413);
nand U18983 (N_18983,N_16558,N_16900);
and U18984 (N_18984,N_16956,N_17198);
xnor U18985 (N_18985,N_16887,N_16939);
and U18986 (N_18986,N_17652,N_17545);
and U18987 (N_18987,N_16572,N_17903);
and U18988 (N_18988,N_16536,N_16783);
nor U18989 (N_18989,N_17556,N_17185);
xor U18990 (N_18990,N_17093,N_17824);
nand U18991 (N_18991,N_16722,N_16849);
nor U18992 (N_18992,N_17736,N_17772);
xnor U18993 (N_18993,N_17112,N_17389);
and U18994 (N_18994,N_17701,N_17823);
nand U18995 (N_18995,N_17977,N_17580);
or U18996 (N_18996,N_17649,N_17488);
xor U18997 (N_18997,N_16829,N_16880);
or U18998 (N_18998,N_17778,N_17293);
or U18999 (N_18999,N_16673,N_16603);
and U19000 (N_19000,N_17249,N_17389);
or U19001 (N_19001,N_17116,N_16978);
or U19002 (N_19002,N_16830,N_17715);
xnor U19003 (N_19003,N_17234,N_17070);
xor U19004 (N_19004,N_16694,N_17798);
or U19005 (N_19005,N_16779,N_16666);
and U19006 (N_19006,N_16603,N_17364);
nor U19007 (N_19007,N_17843,N_17356);
nand U19008 (N_19008,N_17593,N_17052);
nand U19009 (N_19009,N_16994,N_17994);
xnor U19010 (N_19010,N_16891,N_17589);
and U19011 (N_19011,N_17343,N_17395);
or U19012 (N_19012,N_17203,N_17613);
xnor U19013 (N_19013,N_17055,N_17641);
nand U19014 (N_19014,N_17446,N_17243);
nand U19015 (N_19015,N_16636,N_17173);
xor U19016 (N_19016,N_17804,N_17320);
nand U19017 (N_19017,N_17761,N_16923);
or U19018 (N_19018,N_17859,N_16896);
or U19019 (N_19019,N_17225,N_17466);
or U19020 (N_19020,N_17329,N_17173);
or U19021 (N_19021,N_17918,N_17902);
xnor U19022 (N_19022,N_16762,N_17047);
or U19023 (N_19023,N_17981,N_17051);
nand U19024 (N_19024,N_17548,N_17818);
or U19025 (N_19025,N_16950,N_16798);
nand U19026 (N_19026,N_17677,N_16699);
xor U19027 (N_19027,N_17271,N_16850);
nor U19028 (N_19028,N_17192,N_16849);
and U19029 (N_19029,N_17586,N_17051);
or U19030 (N_19030,N_17461,N_17067);
and U19031 (N_19031,N_17347,N_17252);
xor U19032 (N_19032,N_17682,N_16950);
nor U19033 (N_19033,N_17239,N_16901);
nor U19034 (N_19034,N_17295,N_17051);
and U19035 (N_19035,N_16783,N_17205);
nor U19036 (N_19036,N_17013,N_17191);
and U19037 (N_19037,N_17440,N_17997);
nor U19038 (N_19038,N_16675,N_16785);
and U19039 (N_19039,N_17686,N_16706);
and U19040 (N_19040,N_16992,N_16879);
nor U19041 (N_19041,N_17853,N_17762);
and U19042 (N_19042,N_17122,N_16989);
nor U19043 (N_19043,N_16863,N_16870);
xor U19044 (N_19044,N_17314,N_17425);
and U19045 (N_19045,N_16743,N_17021);
nand U19046 (N_19046,N_17059,N_16645);
or U19047 (N_19047,N_17182,N_16554);
and U19048 (N_19048,N_17193,N_16776);
xor U19049 (N_19049,N_17425,N_17116);
or U19050 (N_19050,N_16614,N_16604);
nand U19051 (N_19051,N_17975,N_16527);
or U19052 (N_19052,N_17917,N_17120);
xnor U19053 (N_19053,N_17682,N_17771);
nor U19054 (N_19054,N_17257,N_16945);
xor U19055 (N_19055,N_16838,N_17025);
xnor U19056 (N_19056,N_17749,N_17139);
or U19057 (N_19057,N_17916,N_17484);
xnor U19058 (N_19058,N_17592,N_16754);
nor U19059 (N_19059,N_17169,N_16566);
xnor U19060 (N_19060,N_16521,N_17074);
nor U19061 (N_19061,N_16934,N_16515);
xor U19062 (N_19062,N_16888,N_17538);
nand U19063 (N_19063,N_17569,N_17472);
or U19064 (N_19064,N_16573,N_16984);
xnor U19065 (N_19065,N_17761,N_17104);
nor U19066 (N_19066,N_16575,N_17982);
nand U19067 (N_19067,N_16855,N_16790);
xnor U19068 (N_19068,N_16866,N_16640);
xnor U19069 (N_19069,N_17972,N_17562);
or U19070 (N_19070,N_16673,N_17090);
nor U19071 (N_19071,N_17835,N_17075);
xnor U19072 (N_19072,N_17745,N_17625);
and U19073 (N_19073,N_16609,N_17921);
or U19074 (N_19074,N_17774,N_16536);
xnor U19075 (N_19075,N_17653,N_16866);
nor U19076 (N_19076,N_17844,N_16654);
nor U19077 (N_19077,N_17822,N_17088);
xnor U19078 (N_19078,N_17105,N_17668);
xnor U19079 (N_19079,N_16666,N_17499);
nor U19080 (N_19080,N_17891,N_17233);
or U19081 (N_19081,N_17149,N_17286);
or U19082 (N_19082,N_17175,N_17486);
and U19083 (N_19083,N_16510,N_17382);
nand U19084 (N_19084,N_16763,N_16687);
and U19085 (N_19085,N_17673,N_17523);
xor U19086 (N_19086,N_16942,N_17199);
xor U19087 (N_19087,N_17509,N_17219);
nand U19088 (N_19088,N_17330,N_16558);
or U19089 (N_19089,N_17344,N_17225);
and U19090 (N_19090,N_17308,N_17372);
nand U19091 (N_19091,N_17311,N_16695);
nand U19092 (N_19092,N_17371,N_17504);
and U19093 (N_19093,N_16849,N_16926);
xor U19094 (N_19094,N_17522,N_17068);
nand U19095 (N_19095,N_16967,N_16633);
nand U19096 (N_19096,N_17280,N_17697);
or U19097 (N_19097,N_17183,N_16661);
nor U19098 (N_19098,N_17743,N_16846);
or U19099 (N_19099,N_16894,N_17283);
nand U19100 (N_19100,N_17086,N_16695);
or U19101 (N_19101,N_17120,N_17257);
nand U19102 (N_19102,N_17883,N_17731);
xnor U19103 (N_19103,N_17483,N_17775);
nor U19104 (N_19104,N_17526,N_17676);
xnor U19105 (N_19105,N_17338,N_17243);
nor U19106 (N_19106,N_17001,N_16813);
and U19107 (N_19107,N_17306,N_17549);
xnor U19108 (N_19108,N_16542,N_17383);
and U19109 (N_19109,N_17020,N_16673);
nor U19110 (N_19110,N_17670,N_17171);
nand U19111 (N_19111,N_16913,N_17244);
nand U19112 (N_19112,N_17079,N_17119);
nand U19113 (N_19113,N_16571,N_17046);
nor U19114 (N_19114,N_17789,N_16668);
and U19115 (N_19115,N_16520,N_16636);
xnor U19116 (N_19116,N_16740,N_17899);
nor U19117 (N_19117,N_16577,N_17064);
or U19118 (N_19118,N_17737,N_17800);
and U19119 (N_19119,N_16642,N_16802);
or U19120 (N_19120,N_17968,N_16664);
and U19121 (N_19121,N_17234,N_17116);
nand U19122 (N_19122,N_16668,N_17955);
nand U19123 (N_19123,N_16653,N_16516);
and U19124 (N_19124,N_17262,N_16754);
nor U19125 (N_19125,N_17936,N_17159);
or U19126 (N_19126,N_17294,N_17217);
xnor U19127 (N_19127,N_17857,N_17505);
nor U19128 (N_19128,N_16607,N_17260);
nand U19129 (N_19129,N_17730,N_17586);
nand U19130 (N_19130,N_16534,N_17583);
nand U19131 (N_19131,N_17651,N_17232);
or U19132 (N_19132,N_17029,N_17853);
xor U19133 (N_19133,N_17844,N_16581);
nor U19134 (N_19134,N_17523,N_17869);
or U19135 (N_19135,N_17128,N_17962);
nor U19136 (N_19136,N_16899,N_17887);
or U19137 (N_19137,N_16810,N_17035);
nand U19138 (N_19138,N_17764,N_17136);
nor U19139 (N_19139,N_16705,N_16932);
xnor U19140 (N_19140,N_17835,N_17718);
nor U19141 (N_19141,N_17082,N_17640);
xnor U19142 (N_19142,N_17113,N_17091);
and U19143 (N_19143,N_17994,N_17436);
nand U19144 (N_19144,N_16919,N_17199);
nor U19145 (N_19145,N_17866,N_17635);
xor U19146 (N_19146,N_17282,N_17973);
or U19147 (N_19147,N_17112,N_17399);
or U19148 (N_19148,N_16694,N_17903);
and U19149 (N_19149,N_16541,N_17315);
xnor U19150 (N_19150,N_17712,N_17667);
or U19151 (N_19151,N_17740,N_17494);
and U19152 (N_19152,N_16771,N_16728);
xor U19153 (N_19153,N_16922,N_16526);
and U19154 (N_19154,N_17167,N_17693);
nand U19155 (N_19155,N_16831,N_16936);
xnor U19156 (N_19156,N_16898,N_16758);
nor U19157 (N_19157,N_16989,N_16565);
nand U19158 (N_19158,N_16869,N_16787);
nand U19159 (N_19159,N_16777,N_17159);
or U19160 (N_19160,N_17006,N_16588);
nand U19161 (N_19161,N_17038,N_16586);
or U19162 (N_19162,N_17335,N_16780);
nor U19163 (N_19163,N_17291,N_17754);
nand U19164 (N_19164,N_17634,N_17415);
and U19165 (N_19165,N_16621,N_17865);
nand U19166 (N_19166,N_16950,N_17411);
and U19167 (N_19167,N_16512,N_16617);
nor U19168 (N_19168,N_17481,N_17933);
xor U19169 (N_19169,N_16577,N_17784);
xor U19170 (N_19170,N_17672,N_17176);
xnor U19171 (N_19171,N_16811,N_17465);
nor U19172 (N_19172,N_17112,N_17756);
and U19173 (N_19173,N_16632,N_17620);
nand U19174 (N_19174,N_17839,N_16531);
xor U19175 (N_19175,N_16993,N_17706);
nor U19176 (N_19176,N_16798,N_16879);
nor U19177 (N_19177,N_16577,N_17538);
or U19178 (N_19178,N_16808,N_16886);
and U19179 (N_19179,N_16744,N_17156);
or U19180 (N_19180,N_16556,N_16623);
nor U19181 (N_19181,N_17200,N_17599);
or U19182 (N_19182,N_17186,N_17594);
nor U19183 (N_19183,N_16752,N_17158);
and U19184 (N_19184,N_17703,N_16606);
xnor U19185 (N_19185,N_16673,N_17813);
nand U19186 (N_19186,N_16733,N_17276);
or U19187 (N_19187,N_17624,N_16893);
nor U19188 (N_19188,N_17779,N_17366);
xor U19189 (N_19189,N_16514,N_16630);
nor U19190 (N_19190,N_16885,N_16835);
or U19191 (N_19191,N_17002,N_17918);
or U19192 (N_19192,N_17014,N_16625);
nor U19193 (N_19193,N_17701,N_17104);
nand U19194 (N_19194,N_17455,N_16985);
nor U19195 (N_19195,N_16833,N_17067);
nand U19196 (N_19196,N_16960,N_16616);
and U19197 (N_19197,N_16639,N_16683);
and U19198 (N_19198,N_16877,N_16887);
xor U19199 (N_19199,N_16733,N_16900);
xnor U19200 (N_19200,N_16899,N_17609);
or U19201 (N_19201,N_17874,N_16593);
and U19202 (N_19202,N_17763,N_17237);
xnor U19203 (N_19203,N_16861,N_17412);
nor U19204 (N_19204,N_17788,N_17326);
xor U19205 (N_19205,N_17093,N_17083);
or U19206 (N_19206,N_17329,N_17855);
nor U19207 (N_19207,N_17404,N_16822);
or U19208 (N_19208,N_17649,N_16964);
nand U19209 (N_19209,N_17250,N_17468);
xnor U19210 (N_19210,N_17591,N_17302);
nand U19211 (N_19211,N_16608,N_17467);
xor U19212 (N_19212,N_16839,N_17325);
nor U19213 (N_19213,N_17668,N_16879);
nand U19214 (N_19214,N_16567,N_17356);
nand U19215 (N_19215,N_17014,N_17857);
nand U19216 (N_19216,N_16805,N_17929);
and U19217 (N_19217,N_17852,N_16732);
and U19218 (N_19218,N_16878,N_16914);
or U19219 (N_19219,N_17779,N_17155);
nor U19220 (N_19220,N_16706,N_17962);
and U19221 (N_19221,N_17939,N_17710);
xnor U19222 (N_19222,N_17793,N_16716);
nand U19223 (N_19223,N_17721,N_16961);
or U19224 (N_19224,N_17779,N_17831);
xor U19225 (N_19225,N_16541,N_16994);
nand U19226 (N_19226,N_16964,N_17123);
nand U19227 (N_19227,N_17881,N_16945);
nor U19228 (N_19228,N_17543,N_17338);
or U19229 (N_19229,N_17748,N_16523);
nor U19230 (N_19230,N_17863,N_17717);
xor U19231 (N_19231,N_17875,N_17195);
and U19232 (N_19232,N_17780,N_16507);
xor U19233 (N_19233,N_17950,N_17902);
nor U19234 (N_19234,N_17893,N_17757);
xor U19235 (N_19235,N_17252,N_16626);
nand U19236 (N_19236,N_17777,N_16530);
nand U19237 (N_19237,N_17559,N_17952);
nor U19238 (N_19238,N_17584,N_17258);
nand U19239 (N_19239,N_16970,N_17466);
or U19240 (N_19240,N_16693,N_17204);
nor U19241 (N_19241,N_17094,N_16746);
and U19242 (N_19242,N_17815,N_17279);
or U19243 (N_19243,N_17778,N_16771);
or U19244 (N_19244,N_17098,N_17478);
or U19245 (N_19245,N_17715,N_17049);
xnor U19246 (N_19246,N_16994,N_17305);
or U19247 (N_19247,N_16638,N_17432);
xor U19248 (N_19248,N_16873,N_17573);
xnor U19249 (N_19249,N_17713,N_16847);
and U19250 (N_19250,N_16988,N_17644);
xor U19251 (N_19251,N_17238,N_16522);
nand U19252 (N_19252,N_16522,N_17754);
or U19253 (N_19253,N_17046,N_17885);
nor U19254 (N_19254,N_16849,N_16754);
or U19255 (N_19255,N_17240,N_17191);
nor U19256 (N_19256,N_17927,N_17180);
or U19257 (N_19257,N_16548,N_17834);
xor U19258 (N_19258,N_17915,N_17184);
nand U19259 (N_19259,N_17206,N_16999);
xor U19260 (N_19260,N_17797,N_16868);
xnor U19261 (N_19261,N_16653,N_16984);
xor U19262 (N_19262,N_17831,N_16800);
nand U19263 (N_19263,N_16690,N_16835);
nand U19264 (N_19264,N_17170,N_17868);
nand U19265 (N_19265,N_16937,N_16993);
nand U19266 (N_19266,N_17698,N_17856);
or U19267 (N_19267,N_16707,N_17859);
or U19268 (N_19268,N_17761,N_16739);
or U19269 (N_19269,N_17657,N_17935);
or U19270 (N_19270,N_17727,N_17538);
nor U19271 (N_19271,N_17838,N_17185);
xor U19272 (N_19272,N_16601,N_17003);
nand U19273 (N_19273,N_17652,N_17160);
nand U19274 (N_19274,N_16643,N_17432);
or U19275 (N_19275,N_16718,N_17629);
xor U19276 (N_19276,N_17077,N_17744);
nand U19277 (N_19277,N_17882,N_16652);
nand U19278 (N_19278,N_17544,N_17750);
nand U19279 (N_19279,N_17543,N_16817);
xor U19280 (N_19280,N_16894,N_17575);
or U19281 (N_19281,N_17306,N_17938);
and U19282 (N_19282,N_16710,N_17702);
nor U19283 (N_19283,N_16800,N_17814);
xor U19284 (N_19284,N_17833,N_16963);
nor U19285 (N_19285,N_17852,N_17876);
xor U19286 (N_19286,N_17644,N_17159);
or U19287 (N_19287,N_17348,N_17671);
nand U19288 (N_19288,N_17273,N_17092);
xnor U19289 (N_19289,N_16725,N_17113);
xor U19290 (N_19290,N_17779,N_17640);
nor U19291 (N_19291,N_16829,N_17728);
or U19292 (N_19292,N_17812,N_17670);
xnor U19293 (N_19293,N_17313,N_17204);
nor U19294 (N_19294,N_17164,N_17670);
nor U19295 (N_19295,N_17336,N_17346);
and U19296 (N_19296,N_17910,N_17715);
and U19297 (N_19297,N_17944,N_16801);
xor U19298 (N_19298,N_17194,N_17040);
and U19299 (N_19299,N_17277,N_17586);
xnor U19300 (N_19300,N_17139,N_17785);
nor U19301 (N_19301,N_17088,N_17174);
xor U19302 (N_19302,N_17052,N_16970);
nor U19303 (N_19303,N_16788,N_17020);
nand U19304 (N_19304,N_17746,N_17160);
or U19305 (N_19305,N_17143,N_17481);
or U19306 (N_19306,N_17218,N_16613);
and U19307 (N_19307,N_17622,N_17516);
nor U19308 (N_19308,N_17295,N_17024);
or U19309 (N_19309,N_17453,N_17471);
nand U19310 (N_19310,N_17892,N_17391);
nor U19311 (N_19311,N_17078,N_17699);
xor U19312 (N_19312,N_17403,N_17487);
or U19313 (N_19313,N_16761,N_17563);
nand U19314 (N_19314,N_17554,N_17806);
and U19315 (N_19315,N_16755,N_17180);
nor U19316 (N_19316,N_17467,N_16502);
nand U19317 (N_19317,N_17371,N_17563);
or U19318 (N_19318,N_17997,N_17877);
nor U19319 (N_19319,N_16672,N_16780);
and U19320 (N_19320,N_17744,N_16929);
and U19321 (N_19321,N_17544,N_16976);
nand U19322 (N_19322,N_17124,N_17020);
nor U19323 (N_19323,N_17061,N_17193);
nand U19324 (N_19324,N_16503,N_16730);
or U19325 (N_19325,N_17239,N_17404);
xor U19326 (N_19326,N_16938,N_17502);
or U19327 (N_19327,N_17409,N_16785);
nand U19328 (N_19328,N_17252,N_17796);
and U19329 (N_19329,N_17082,N_16798);
and U19330 (N_19330,N_16592,N_17093);
and U19331 (N_19331,N_16909,N_17157);
and U19332 (N_19332,N_17082,N_17660);
xor U19333 (N_19333,N_17980,N_16719);
and U19334 (N_19334,N_17259,N_16684);
or U19335 (N_19335,N_16530,N_17161);
nand U19336 (N_19336,N_16503,N_17283);
nor U19337 (N_19337,N_17167,N_17195);
nor U19338 (N_19338,N_17815,N_17660);
nand U19339 (N_19339,N_17448,N_17083);
nand U19340 (N_19340,N_17074,N_16933);
nor U19341 (N_19341,N_17406,N_17439);
nand U19342 (N_19342,N_16721,N_17794);
nand U19343 (N_19343,N_17869,N_17409);
nor U19344 (N_19344,N_16554,N_17290);
or U19345 (N_19345,N_17112,N_17373);
and U19346 (N_19346,N_16698,N_16672);
xnor U19347 (N_19347,N_17885,N_17569);
or U19348 (N_19348,N_17151,N_17271);
nand U19349 (N_19349,N_17998,N_17251);
nor U19350 (N_19350,N_16899,N_17592);
and U19351 (N_19351,N_17585,N_16924);
nor U19352 (N_19352,N_17567,N_17040);
nand U19353 (N_19353,N_17793,N_17683);
or U19354 (N_19354,N_17863,N_16545);
or U19355 (N_19355,N_16841,N_17911);
nor U19356 (N_19356,N_17974,N_16622);
and U19357 (N_19357,N_17534,N_16927);
nor U19358 (N_19358,N_17063,N_17754);
nand U19359 (N_19359,N_17725,N_17157);
nand U19360 (N_19360,N_17422,N_17740);
and U19361 (N_19361,N_17572,N_17855);
nor U19362 (N_19362,N_17550,N_16797);
or U19363 (N_19363,N_16885,N_17814);
nand U19364 (N_19364,N_17629,N_17441);
or U19365 (N_19365,N_17602,N_17455);
nand U19366 (N_19366,N_16726,N_16768);
and U19367 (N_19367,N_17780,N_16946);
or U19368 (N_19368,N_17675,N_17992);
xnor U19369 (N_19369,N_17159,N_17204);
and U19370 (N_19370,N_16919,N_17700);
and U19371 (N_19371,N_17842,N_16801);
xor U19372 (N_19372,N_16874,N_17650);
nand U19373 (N_19373,N_17327,N_17247);
xnor U19374 (N_19374,N_17985,N_17386);
or U19375 (N_19375,N_17969,N_17897);
nand U19376 (N_19376,N_17977,N_17671);
xor U19377 (N_19377,N_17473,N_17027);
or U19378 (N_19378,N_17153,N_16790);
and U19379 (N_19379,N_16503,N_17265);
nand U19380 (N_19380,N_16982,N_17260);
nor U19381 (N_19381,N_16807,N_17441);
or U19382 (N_19382,N_16973,N_17798);
nor U19383 (N_19383,N_17446,N_17786);
or U19384 (N_19384,N_17440,N_16862);
or U19385 (N_19385,N_17476,N_16886);
or U19386 (N_19386,N_17215,N_17793);
and U19387 (N_19387,N_16771,N_17370);
xor U19388 (N_19388,N_16884,N_17216);
nand U19389 (N_19389,N_16949,N_16802);
xor U19390 (N_19390,N_17949,N_16854);
nand U19391 (N_19391,N_16690,N_16541);
or U19392 (N_19392,N_16746,N_16620);
nand U19393 (N_19393,N_17865,N_17427);
xnor U19394 (N_19394,N_17691,N_17114);
and U19395 (N_19395,N_17872,N_17715);
or U19396 (N_19396,N_17208,N_17479);
or U19397 (N_19397,N_17158,N_16593);
and U19398 (N_19398,N_16590,N_16658);
xor U19399 (N_19399,N_17372,N_16695);
or U19400 (N_19400,N_17132,N_17372);
nor U19401 (N_19401,N_17858,N_17494);
and U19402 (N_19402,N_17434,N_17563);
xor U19403 (N_19403,N_17948,N_16887);
or U19404 (N_19404,N_16694,N_17528);
nand U19405 (N_19405,N_16846,N_17687);
or U19406 (N_19406,N_17458,N_16587);
or U19407 (N_19407,N_17385,N_17761);
nor U19408 (N_19408,N_17048,N_17872);
or U19409 (N_19409,N_17711,N_16974);
or U19410 (N_19410,N_17430,N_17059);
xor U19411 (N_19411,N_16915,N_16932);
xor U19412 (N_19412,N_17818,N_17135);
or U19413 (N_19413,N_17990,N_17449);
or U19414 (N_19414,N_17407,N_17729);
or U19415 (N_19415,N_17206,N_17364);
and U19416 (N_19416,N_17717,N_17024);
nand U19417 (N_19417,N_17910,N_17558);
nor U19418 (N_19418,N_17409,N_17221);
and U19419 (N_19419,N_16722,N_17726);
xor U19420 (N_19420,N_16604,N_16515);
and U19421 (N_19421,N_17108,N_17191);
xor U19422 (N_19422,N_16766,N_17961);
nand U19423 (N_19423,N_16623,N_17842);
and U19424 (N_19424,N_16842,N_16940);
nand U19425 (N_19425,N_17746,N_17667);
nor U19426 (N_19426,N_17797,N_16775);
and U19427 (N_19427,N_16592,N_16719);
nor U19428 (N_19428,N_17986,N_17441);
or U19429 (N_19429,N_17692,N_17267);
xnor U19430 (N_19430,N_17490,N_17947);
nor U19431 (N_19431,N_16999,N_17878);
nor U19432 (N_19432,N_16912,N_17306);
nand U19433 (N_19433,N_17259,N_17676);
xnor U19434 (N_19434,N_16882,N_17408);
xnor U19435 (N_19435,N_17836,N_17206);
xnor U19436 (N_19436,N_16860,N_17893);
xor U19437 (N_19437,N_16646,N_17453);
or U19438 (N_19438,N_17372,N_17819);
and U19439 (N_19439,N_17009,N_16876);
nand U19440 (N_19440,N_17956,N_16913);
and U19441 (N_19441,N_16763,N_17521);
nor U19442 (N_19442,N_17562,N_17687);
or U19443 (N_19443,N_17123,N_17013);
and U19444 (N_19444,N_17037,N_17312);
xor U19445 (N_19445,N_17816,N_17621);
nand U19446 (N_19446,N_16742,N_17755);
xor U19447 (N_19447,N_17192,N_17128);
or U19448 (N_19448,N_17082,N_17277);
nand U19449 (N_19449,N_16586,N_17515);
or U19450 (N_19450,N_17230,N_17126);
nor U19451 (N_19451,N_17773,N_17427);
xnor U19452 (N_19452,N_17848,N_17041);
nor U19453 (N_19453,N_17006,N_17819);
or U19454 (N_19454,N_17951,N_17922);
and U19455 (N_19455,N_17279,N_16738);
and U19456 (N_19456,N_17794,N_17603);
nor U19457 (N_19457,N_17469,N_17107);
or U19458 (N_19458,N_17366,N_17983);
and U19459 (N_19459,N_17258,N_17388);
or U19460 (N_19460,N_17967,N_17262);
or U19461 (N_19461,N_17382,N_17022);
and U19462 (N_19462,N_17734,N_17594);
and U19463 (N_19463,N_16975,N_17593);
and U19464 (N_19464,N_17477,N_16649);
xnor U19465 (N_19465,N_17979,N_17890);
or U19466 (N_19466,N_17607,N_16756);
and U19467 (N_19467,N_17484,N_17375);
nand U19468 (N_19468,N_16643,N_17684);
and U19469 (N_19469,N_17985,N_16967);
or U19470 (N_19470,N_16536,N_17326);
xor U19471 (N_19471,N_17485,N_17888);
and U19472 (N_19472,N_17541,N_17858);
and U19473 (N_19473,N_16578,N_17000);
nand U19474 (N_19474,N_16557,N_16809);
nor U19475 (N_19475,N_17884,N_17912);
xor U19476 (N_19476,N_17422,N_16888);
and U19477 (N_19477,N_17697,N_17801);
xor U19478 (N_19478,N_17491,N_16615);
nor U19479 (N_19479,N_16544,N_17902);
and U19480 (N_19480,N_17743,N_17469);
or U19481 (N_19481,N_17658,N_17363);
nand U19482 (N_19482,N_17300,N_17547);
nand U19483 (N_19483,N_17853,N_16840);
and U19484 (N_19484,N_16521,N_17268);
or U19485 (N_19485,N_17644,N_17065);
and U19486 (N_19486,N_17121,N_16838);
and U19487 (N_19487,N_17800,N_17282);
xnor U19488 (N_19488,N_17719,N_17796);
or U19489 (N_19489,N_16908,N_16800);
and U19490 (N_19490,N_16731,N_17738);
nand U19491 (N_19491,N_17769,N_17292);
or U19492 (N_19492,N_17043,N_17454);
or U19493 (N_19493,N_16539,N_17731);
xor U19494 (N_19494,N_17500,N_16653);
or U19495 (N_19495,N_17960,N_16562);
nor U19496 (N_19496,N_17404,N_17251);
nor U19497 (N_19497,N_16841,N_16626);
xor U19498 (N_19498,N_16816,N_16852);
xor U19499 (N_19499,N_17294,N_16812);
or U19500 (N_19500,N_18922,N_19383);
and U19501 (N_19501,N_19385,N_19189);
or U19502 (N_19502,N_18339,N_19138);
or U19503 (N_19503,N_19085,N_18522);
and U19504 (N_19504,N_18009,N_18533);
xor U19505 (N_19505,N_18890,N_18545);
nor U19506 (N_19506,N_19186,N_18470);
and U19507 (N_19507,N_18849,N_19192);
or U19508 (N_19508,N_19188,N_18923);
and U19509 (N_19509,N_18877,N_18137);
and U19510 (N_19510,N_18003,N_19087);
and U19511 (N_19511,N_18799,N_18175);
nand U19512 (N_19512,N_19113,N_19032);
and U19513 (N_19513,N_18089,N_18917);
or U19514 (N_19514,N_19246,N_18775);
and U19515 (N_19515,N_19309,N_18389);
nand U19516 (N_19516,N_18439,N_18631);
xnor U19517 (N_19517,N_18555,N_19447);
nand U19518 (N_19518,N_19218,N_18831);
or U19519 (N_19519,N_19417,N_19193);
and U19520 (N_19520,N_18664,N_18390);
or U19521 (N_19521,N_18220,N_19356);
xnor U19522 (N_19522,N_18094,N_18216);
nand U19523 (N_19523,N_18016,N_18876);
and U19524 (N_19524,N_19446,N_19004);
and U19525 (N_19525,N_19065,N_18237);
and U19526 (N_19526,N_18054,N_18346);
nor U19527 (N_19527,N_18403,N_18115);
or U19528 (N_19528,N_18297,N_18804);
nand U19529 (N_19529,N_18019,N_18540);
nor U19530 (N_19530,N_18402,N_19275);
xor U19531 (N_19531,N_18611,N_18709);
or U19532 (N_19532,N_19346,N_18875);
or U19533 (N_19533,N_19392,N_18000);
or U19534 (N_19534,N_19328,N_18474);
nor U19535 (N_19535,N_18110,N_18135);
xnor U19536 (N_19536,N_19498,N_18977);
or U19537 (N_19537,N_19190,N_18459);
and U19538 (N_19538,N_18340,N_18704);
nand U19539 (N_19539,N_19453,N_18935);
or U19540 (N_19540,N_18453,N_18226);
nor U19541 (N_19541,N_18008,N_19116);
nand U19542 (N_19542,N_19355,N_19177);
nand U19543 (N_19543,N_19072,N_18294);
and U19544 (N_19544,N_18868,N_19318);
nand U19545 (N_19545,N_19198,N_18651);
nor U19546 (N_19546,N_19341,N_18629);
nand U19547 (N_19547,N_19420,N_18599);
nor U19548 (N_19548,N_18145,N_19478);
xor U19549 (N_19549,N_18146,N_19155);
nand U19550 (N_19550,N_19001,N_19273);
or U19551 (N_19551,N_19289,N_18249);
nor U19552 (N_19552,N_18271,N_19093);
and U19553 (N_19553,N_18017,N_18218);
nor U19554 (N_19554,N_18335,N_19254);
nand U19555 (N_19555,N_18717,N_19316);
and U19556 (N_19556,N_18780,N_19130);
nor U19557 (N_19557,N_18621,N_18030);
xor U19558 (N_19558,N_18325,N_18375);
or U19559 (N_19559,N_19444,N_19399);
xor U19560 (N_19560,N_18743,N_19472);
and U19561 (N_19561,N_18666,N_19105);
nand U19562 (N_19562,N_18351,N_18131);
or U19563 (N_19563,N_18757,N_18910);
or U19564 (N_19564,N_18529,N_18207);
or U19565 (N_19565,N_19493,N_18685);
or U19566 (N_19566,N_19439,N_18268);
nor U19567 (N_19567,N_18612,N_18201);
and U19568 (N_19568,N_18803,N_18984);
nor U19569 (N_19569,N_18365,N_19062);
nor U19570 (N_19570,N_19243,N_18998);
xnor U19571 (N_19571,N_18515,N_18819);
and U19572 (N_19572,N_19495,N_18475);
and U19573 (N_19573,N_18916,N_18565);
xor U19574 (N_19574,N_18858,N_18253);
nand U19575 (N_19575,N_19252,N_18992);
xnor U19576 (N_19576,N_19121,N_18034);
or U19577 (N_19577,N_19018,N_19250);
nand U19578 (N_19578,N_18681,N_19055);
nor U19579 (N_19579,N_19384,N_19357);
and U19580 (N_19580,N_19184,N_18193);
and U19581 (N_19581,N_18307,N_18878);
xnor U19582 (N_19582,N_18314,N_18993);
and U19583 (N_19583,N_19408,N_18396);
nand U19584 (N_19584,N_18020,N_18200);
xnor U19585 (N_19585,N_18760,N_18980);
nand U19586 (N_19586,N_18236,N_18885);
or U19587 (N_19587,N_18357,N_19460);
xor U19588 (N_19588,N_19479,N_18842);
nor U19589 (N_19589,N_18978,N_18443);
or U19590 (N_19590,N_18063,N_18418);
and U19591 (N_19591,N_18416,N_19031);
nor U19592 (N_19592,N_18726,N_19148);
or U19593 (N_19593,N_19078,N_19156);
nand U19594 (N_19594,N_18245,N_18300);
nor U19595 (N_19595,N_18288,N_18759);
and U19596 (N_19596,N_18598,N_18729);
or U19597 (N_19597,N_19211,N_18927);
nor U19598 (N_19598,N_18290,N_18725);
xor U19599 (N_19599,N_19152,N_19313);
nor U19600 (N_19600,N_19069,N_18446);
nand U19601 (N_19601,N_18506,N_18329);
and U19602 (N_19602,N_19304,N_18635);
nand U19603 (N_19603,N_18058,N_18574);
or U19604 (N_19604,N_18251,N_19435);
and U19605 (N_19605,N_18082,N_18051);
or U19606 (N_19606,N_19285,N_19061);
xor U19607 (N_19607,N_18005,N_18167);
nor U19608 (N_19608,N_19373,N_18667);
nand U19609 (N_19609,N_18940,N_19083);
xor U19610 (N_19610,N_18953,N_18974);
xnor U19611 (N_19611,N_19253,N_18445);
xor U19612 (N_19612,N_18733,N_19306);
or U19613 (N_19613,N_19416,N_18383);
and U19614 (N_19614,N_19100,N_18693);
nand U19615 (N_19615,N_18069,N_18045);
xnor U19616 (N_19616,N_18101,N_19003);
and U19617 (N_19617,N_18258,N_19277);
xor U19618 (N_19618,N_18350,N_18333);
and U19619 (N_19619,N_19168,N_18208);
and U19620 (N_19620,N_18289,N_18263);
nor U19621 (N_19621,N_18705,N_19164);
nor U19622 (N_19622,N_18711,N_18093);
nor U19623 (N_19623,N_19034,N_18720);
nor U19624 (N_19624,N_19238,N_18280);
nand U19625 (N_19625,N_19452,N_18634);
or U19626 (N_19626,N_18581,N_18739);
or U19627 (N_19627,N_18646,N_19333);
or U19628 (N_19628,N_18809,N_18961);
xor U19629 (N_19629,N_18792,N_18904);
nor U19630 (N_19630,N_18941,N_18802);
nor U19631 (N_19631,N_19009,N_18412);
nand U19632 (N_19632,N_18433,N_19450);
xor U19633 (N_19633,N_18838,N_18751);
and U19634 (N_19634,N_19262,N_19268);
and U19635 (N_19635,N_18811,N_18587);
nand U19636 (N_19636,N_18343,N_19215);
or U19637 (N_19637,N_18963,N_18500);
or U19638 (N_19638,N_19287,N_18192);
nand U19639 (N_19639,N_18186,N_19220);
or U19640 (N_19640,N_19013,N_18815);
nand U19641 (N_19641,N_18930,N_19411);
nor U19642 (N_19642,N_18795,N_19282);
nand U19643 (N_19643,N_18643,N_18088);
nand U19644 (N_19644,N_18912,N_18728);
and U19645 (N_19645,N_18584,N_18462);
xnor U19646 (N_19646,N_18550,N_19213);
and U19647 (N_19647,N_18805,N_18310);
or U19648 (N_19648,N_19343,N_18098);
xnor U19649 (N_19649,N_19387,N_18590);
or U19650 (N_19650,N_18936,N_18524);
or U19651 (N_19651,N_18542,N_18388);
or U19652 (N_19652,N_19425,N_19021);
or U19653 (N_19653,N_19162,N_19281);
nand U19654 (N_19654,N_18369,N_18668);
nand U19655 (N_19655,N_18287,N_18790);
nor U19656 (N_19656,N_18764,N_18066);
or U19657 (N_19657,N_19465,N_18971);
or U19658 (N_19658,N_19086,N_18495);
or U19659 (N_19659,N_18523,N_19326);
nand U19660 (N_19660,N_18356,N_19437);
nor U19661 (N_19661,N_18274,N_18719);
nand U19662 (N_19662,N_19308,N_18492);
xnor U19663 (N_19663,N_19167,N_19020);
and U19664 (N_19664,N_19187,N_18257);
xor U19665 (N_19665,N_18223,N_18042);
xnor U19666 (N_19666,N_19299,N_18173);
nor U19667 (N_19667,N_19208,N_18671);
or U19668 (N_19668,N_18102,N_19056);
xnor U19669 (N_19669,N_19362,N_18426);
nand U19670 (N_19670,N_19456,N_19183);
xor U19671 (N_19671,N_19048,N_18494);
nand U19672 (N_19672,N_18514,N_18750);
and U19673 (N_19673,N_18091,N_18076);
or U19674 (N_19674,N_18139,N_19487);
or U19675 (N_19675,N_18376,N_19063);
and U19676 (N_19676,N_18723,N_19217);
xor U19677 (N_19677,N_19301,N_19106);
or U19678 (N_19678,N_19266,N_18129);
and U19679 (N_19679,N_19006,N_19467);
and U19680 (N_19680,N_18434,N_18969);
or U19681 (N_19681,N_18559,N_18684);
nand U19682 (N_19682,N_18296,N_18832);
or U19683 (N_19683,N_18421,N_18588);
xor U19684 (N_19684,N_18182,N_18266);
nor U19685 (N_19685,N_19388,N_18517);
or U19686 (N_19686,N_19348,N_19209);
and U19687 (N_19687,N_19418,N_19283);
xor U19688 (N_19688,N_19461,N_19426);
nand U19689 (N_19689,N_19127,N_19036);
nor U19690 (N_19690,N_18820,N_18901);
nand U19691 (N_19691,N_19323,N_18558);
nor U19692 (N_19692,N_18456,N_18417);
and U19693 (N_19693,N_18577,N_18222);
or U19694 (N_19694,N_19429,N_18084);
or U19695 (N_19695,N_18564,N_19321);
xor U19696 (N_19696,N_18883,N_18487);
nor U19697 (N_19697,N_19248,N_19485);
nand U19698 (N_19698,N_18055,N_19117);
nand U19699 (N_19699,N_18349,N_18441);
and U19700 (N_19700,N_18013,N_18585);
or U19701 (N_19701,N_19149,N_18537);
and U19702 (N_19702,N_18853,N_18707);
and U19703 (N_19703,N_18670,N_18463);
and U19704 (N_19704,N_18413,N_19463);
xor U19705 (N_19705,N_18583,N_18230);
nand U19706 (N_19706,N_18505,N_19258);
or U19707 (N_19707,N_18464,N_18718);
nor U19708 (N_19708,N_18015,N_18848);
nand U19709 (N_19709,N_18779,N_19310);
xor U19710 (N_19710,N_18136,N_19494);
nor U19711 (N_19711,N_18948,N_18282);
and U19712 (N_19712,N_19067,N_18269);
and U19713 (N_19713,N_19368,N_18428);
nor U19714 (N_19714,N_18722,N_19363);
and U19715 (N_19715,N_18852,N_18489);
or U19716 (N_19716,N_18669,N_18509);
nor U19717 (N_19717,N_18945,N_18014);
nor U19718 (N_19718,N_18080,N_18399);
nand U19719 (N_19719,N_19475,N_18106);
xnor U19720 (N_19720,N_18732,N_18767);
xor U19721 (N_19721,N_18111,N_18814);
and U19722 (N_19722,N_18960,N_18158);
nor U19723 (N_19723,N_18188,N_18074);
nand U19724 (N_19724,N_18293,N_19372);
nand U19725 (N_19725,N_19071,N_18304);
nand U19726 (N_19726,N_18658,N_19389);
or U19727 (N_19727,N_18233,N_18516);
xor U19728 (N_19728,N_18143,N_19102);
nand U19729 (N_19729,N_19174,N_18839);
xor U19730 (N_19730,N_19015,N_18401);
or U19731 (N_19731,N_18202,N_18580);
xnor U19732 (N_19732,N_18538,N_19204);
nand U19733 (N_19733,N_18273,N_18863);
nor U19734 (N_19734,N_18007,N_18036);
or U19735 (N_19735,N_19410,N_18134);
or U19736 (N_19736,N_19471,N_18606);
or U19737 (N_19737,N_19140,N_19235);
or U19738 (N_19738,N_19210,N_18845);
nor U19739 (N_19739,N_18278,N_18968);
and U19740 (N_19740,N_18122,N_18393);
and U19741 (N_19741,N_19421,N_18452);
xnor U19742 (N_19742,N_19312,N_19074);
nor U19743 (N_19743,N_18121,N_19068);
or U19744 (N_19744,N_19349,N_18437);
xnor U19745 (N_19745,N_19137,N_19286);
xor U19746 (N_19746,N_19172,N_18800);
xor U19747 (N_19747,N_18267,N_19000);
nand U19748 (N_19748,N_19377,N_18797);
xnor U19749 (N_19749,N_18962,N_18114);
or U19750 (N_19750,N_18873,N_18661);
xnor U19751 (N_19751,N_18057,N_18353);
and U19752 (N_19752,N_18386,N_18241);
nand U19753 (N_19753,N_18699,N_18752);
or U19754 (N_19754,N_18286,N_19375);
or U19755 (N_19755,N_19352,N_19237);
and U19756 (N_19756,N_19202,N_19432);
xnor U19757 (N_19757,N_18126,N_19104);
or U19758 (N_19758,N_19497,N_19300);
or U19759 (N_19759,N_18373,N_18265);
and U19760 (N_19760,N_18663,N_18133);
nand U19761 (N_19761,N_19111,N_18461);
and U19762 (N_19762,N_18778,N_18985);
nand U19763 (N_19763,N_18065,N_18438);
and U19764 (N_19764,N_18525,N_18050);
xor U19765 (N_19765,N_18486,N_18213);
and U19766 (N_19766,N_18181,N_19334);
nor U19767 (N_19767,N_18191,N_19434);
nand U19768 (N_19768,N_18116,N_18784);
and U19769 (N_19769,N_18690,N_18336);
xnor U19770 (N_19770,N_18731,N_18568);
nor U19771 (N_19771,N_18482,N_18543);
and U19772 (N_19772,N_18561,N_18614);
nor U19773 (N_19773,N_18377,N_18306);
and U19774 (N_19774,N_18119,N_19199);
and U19775 (N_19775,N_18604,N_18983);
nor U19776 (N_19776,N_19403,N_18469);
xor U19777 (N_19777,N_18323,N_19280);
or U19778 (N_19778,N_18113,N_18090);
xor U19779 (N_19779,N_19180,N_18465);
nor U19780 (N_19780,N_18712,N_19366);
nand U19781 (N_19781,N_18378,N_18630);
and U19782 (N_19782,N_19331,N_18988);
nor U19783 (N_19783,N_19492,N_18370);
nor U19784 (N_19784,N_18232,N_19466);
nand U19785 (N_19785,N_18806,N_18163);
or U19786 (N_19786,N_18672,N_19491);
nand U19787 (N_19787,N_18761,N_18594);
nand U19788 (N_19788,N_19200,N_18198);
nor U19789 (N_19789,N_19260,N_18311);
and U19790 (N_19790,N_18716,N_19438);
nor U19791 (N_19791,N_18322,N_18640);
xor U19792 (N_19792,N_19226,N_19119);
nor U19793 (N_19793,N_19097,N_18768);
or U19794 (N_19794,N_19296,N_19405);
and U19795 (N_19795,N_19081,N_19241);
nand U19796 (N_19796,N_18737,N_19436);
and U19797 (N_19797,N_18148,N_19043);
nor U19798 (N_19798,N_18501,N_18841);
nand U19799 (N_19799,N_18449,N_18773);
or U19800 (N_19800,N_19358,N_19222);
nor U19801 (N_19801,N_18504,N_18225);
xnor U19802 (N_19802,N_18075,N_19454);
or U19803 (N_19803,N_19263,N_18099);
nand U19804 (N_19804,N_19109,N_18881);
nor U19805 (N_19805,N_19040,N_19115);
nor U19806 (N_19806,N_18644,N_19090);
or U19807 (N_19807,N_19096,N_19367);
or U19808 (N_19808,N_18818,N_18560);
nand U19809 (N_19809,N_18966,N_18478);
and U19810 (N_19810,N_18214,N_19007);
xnor U19811 (N_19811,N_18822,N_18721);
nor U19812 (N_19812,N_18476,N_19247);
nor U19813 (N_19813,N_18925,N_18603);
or U19814 (N_19814,N_18552,N_19413);
nand U19815 (N_19815,N_19473,N_19047);
nor U19816 (N_19816,N_19279,N_18676);
nor U19817 (N_19817,N_18578,N_19158);
or U19818 (N_19818,N_18851,N_18184);
or U19819 (N_19819,N_18813,N_18107);
xor U19820 (N_19820,N_18793,N_18535);
nor U19821 (N_19821,N_19276,N_19054);
xnor U19822 (N_19822,N_18547,N_18682);
and U19823 (N_19823,N_18331,N_18586);
and U19824 (N_19824,N_18123,N_19433);
nand U19825 (N_19825,N_18435,N_18391);
nor U19826 (N_19826,N_18947,N_19256);
nor U19827 (N_19827,N_18632,N_19342);
nor U19828 (N_19828,N_18837,N_18490);
and U19829 (N_19829,N_18865,N_18301);
xnor U19830 (N_19830,N_18758,N_18738);
or U19831 (N_19831,N_18924,N_18234);
or U19832 (N_19832,N_18355,N_18755);
and U19833 (N_19833,N_18384,N_18965);
or U19834 (N_19834,N_18913,N_18899);
and U19835 (N_19835,N_18688,N_18468);
xnor U19836 (N_19836,N_18344,N_19374);
xnor U19837 (N_19837,N_18436,N_18746);
nand U19838 (N_19838,N_18451,N_18763);
nand U19839 (N_19839,N_19404,N_18637);
nand U19840 (N_19840,N_18411,N_18601);
or U19841 (N_19841,N_18534,N_18382);
xnor U19842 (N_19842,N_18695,N_18109);
nand U19843 (N_19843,N_18964,N_18169);
nor U19844 (N_19844,N_18518,N_18931);
xor U19845 (N_19845,N_19207,N_19236);
nor U19846 (N_19846,N_18785,N_18556);
xor U19847 (N_19847,N_18613,N_18367);
nand U19848 (N_19848,N_19302,N_18911);
nor U19849 (N_19849,N_19365,N_18150);
nor U19850 (N_19850,N_18703,N_19203);
nor U19851 (N_19851,N_18056,N_19371);
nand U19852 (N_19852,N_18209,N_19060);
nand U19853 (N_19853,N_19094,N_18649);
xnor U19854 (N_19854,N_18986,N_18946);
or U19855 (N_19855,N_18829,N_19415);
or U19856 (N_19856,N_19298,N_19288);
nor U19857 (N_19857,N_19039,N_19407);
or U19858 (N_19858,N_19151,N_18168);
and U19859 (N_19859,N_18165,N_18155);
and U19860 (N_19860,N_19242,N_19011);
xnor U19861 (N_19861,N_18281,N_19058);
nand U19862 (N_19862,N_18582,N_18740);
and U19863 (N_19863,N_18400,N_19332);
nor U19864 (N_19864,N_18954,N_18149);
xor U19865 (N_19865,N_18179,N_19319);
nand U19866 (N_19866,N_19153,N_18077);
or U19867 (N_19867,N_19025,N_19139);
nor U19868 (N_19868,N_19143,N_19245);
or U19869 (N_19869,N_18609,N_18364);
nand U19870 (N_19870,N_18420,N_18921);
nor U19871 (N_19871,N_18526,N_18995);
xnor U19872 (N_19872,N_18031,N_18835);
or U19873 (N_19873,N_19154,N_18843);
or U19874 (N_19874,N_18432,N_18745);
xnor U19875 (N_19875,N_19161,N_19422);
nor U19876 (N_19876,N_19294,N_19354);
xnor U19877 (N_19877,N_18347,N_18907);
and U19878 (N_19878,N_18154,N_18850);
nand U19879 (N_19879,N_18153,N_19108);
nor U19880 (N_19880,N_19041,N_18087);
nand U19881 (N_19881,N_18053,N_18352);
and U19882 (N_19882,N_18252,N_18826);
and U19883 (N_19883,N_18410,N_18513);
nand U19884 (N_19884,N_18419,N_18937);
or U19885 (N_19885,N_18519,N_18976);
nand U19886 (N_19886,N_18319,N_19027);
xnor U19887 (N_19887,N_18029,N_19214);
nor U19888 (N_19888,N_19259,N_19128);
xnor U19889 (N_19889,N_18284,N_18934);
and U19890 (N_19890,N_18942,N_18562);
or U19891 (N_19891,N_19486,N_18104);
or U19892 (N_19892,N_18250,N_19396);
xor U19893 (N_19893,N_18205,N_18888);
nand U19894 (N_19894,N_19066,N_18210);
or U19895 (N_19895,N_19219,N_19150);
and U19896 (N_19896,N_19181,N_18591);
and U19897 (N_19897,N_19076,N_18011);
and U19898 (N_19898,N_18337,N_18302);
xor U19899 (N_19899,N_18787,N_18455);
xnor U19900 (N_19900,N_18283,N_19325);
xnor U19901 (N_19901,N_19244,N_18554);
or U19902 (N_19902,N_18683,N_19176);
nor U19903 (N_19903,N_18987,N_19216);
and U19904 (N_19904,N_18164,N_19114);
xor U19905 (N_19905,N_19095,N_18387);
and U19906 (N_19906,N_18955,N_18100);
xor U19907 (N_19907,N_19175,N_18747);
and U19908 (N_19908,N_18212,N_18328);
nor U19909 (N_19909,N_19488,N_18033);
xnor U19910 (N_19910,N_18855,N_19134);
or U19911 (N_19911,N_19477,N_18471);
nor U19912 (N_19912,N_18915,N_18821);
xor U19913 (N_19913,N_18275,N_19295);
and U19914 (N_19914,N_18847,N_18472);
or U19915 (N_19915,N_19118,N_19147);
and U19916 (N_19916,N_19091,N_19171);
and U19917 (N_19917,N_19430,N_18157);
and U19918 (N_19918,N_19376,N_18359);
nand U19919 (N_19919,N_19132,N_18914);
and U19920 (N_19920,N_18424,N_18654);
nand U19921 (N_19921,N_18046,N_19489);
nor U19922 (N_19922,N_19293,N_18407);
nand U19923 (N_19923,N_19324,N_19322);
or U19924 (N_19924,N_18141,N_18096);
nand U19925 (N_19925,N_19073,N_18639);
or U19926 (N_19926,N_18010,N_18317);
nor U19927 (N_19927,N_18025,N_18762);
or U19928 (N_19928,N_18052,N_18361);
or U19929 (N_19929,N_18769,N_18366);
or U19930 (N_19930,N_18197,N_18548);
or U19931 (N_19931,N_19035,N_18497);
nand U19932 (N_19932,N_18589,N_18862);
and U19933 (N_19933,N_19320,N_18744);
and U19934 (N_19934,N_19394,N_18162);
xnor U19935 (N_19935,N_18140,N_18348);
xnor U19936 (N_19936,N_18686,N_19391);
and U19937 (N_19937,N_19157,N_18772);
nor U19938 (N_19938,N_19469,N_18532);
and U19939 (N_19939,N_19379,N_18636);
or U19940 (N_19940,N_18484,N_19103);
and U19941 (N_19941,N_18394,N_18950);
nand U19942 (N_19942,N_19476,N_19307);
xnor U19943 (N_19943,N_18004,N_19225);
nand U19944 (N_19944,N_19206,N_18512);
xnor U19945 (N_19945,N_19344,N_18291);
or U19946 (N_19946,N_18520,N_18624);
xor U19947 (N_19947,N_18919,N_18483);
or U19948 (N_19948,N_19290,N_18130);
nand U19949 (N_19949,N_18576,N_19353);
xor U19950 (N_19950,N_18891,N_18457);
or U19951 (N_19951,N_18678,N_18423);
nor U19952 (N_19952,N_19125,N_18753);
nor U19953 (N_19953,N_18674,N_18617);
nand U19954 (N_19954,N_18037,N_18180);
or U19955 (N_19955,N_19329,N_19194);
nand U19956 (N_19956,N_18929,N_19030);
nand U19957 (N_19957,N_19084,N_19080);
or U19958 (N_19958,N_18622,N_18546);
xor U19959 (N_19959,N_18810,N_18623);
nand U19960 (N_19960,N_18238,N_19023);
nor U19961 (N_19961,N_19327,N_19445);
or U19962 (N_19962,N_19272,N_19464);
or U19963 (N_19963,N_19033,N_18754);
or U19964 (N_19964,N_18272,N_18170);
and U19965 (N_19965,N_18765,N_19017);
nor U19966 (N_19966,N_18264,N_19008);
nor U19967 (N_19967,N_19338,N_19005);
or U19968 (N_19968,N_19046,N_18616);
or U19969 (N_19969,N_19441,N_18259);
and U19970 (N_19970,N_19024,N_19449);
nor U19971 (N_19971,N_18006,N_18896);
and U19972 (N_19972,N_18303,N_19112);
xnor U19973 (N_19973,N_18493,N_18648);
nand U19974 (N_19974,N_18127,N_18228);
and U19975 (N_19975,N_18068,N_19233);
or U19976 (N_19976,N_18724,N_18766);
nor U19977 (N_19977,N_18566,N_18982);
and U19978 (N_19978,N_18156,N_18909);
nand U19979 (N_19979,N_19197,N_18177);
xnor U19980 (N_19980,N_18567,N_19099);
and U19981 (N_19981,N_19378,N_18206);
nor U19982 (N_19982,N_18933,N_18477);
nor U19983 (N_19983,N_18144,N_19160);
or U19984 (N_19984,N_18970,N_18596);
nand U19985 (N_19985,N_18900,N_19428);
nand U19986 (N_19986,N_18001,N_18926);
xnor U19987 (N_19987,N_18659,N_19077);
nor U19988 (N_19988,N_19468,N_18072);
and U19989 (N_19989,N_18638,N_18330);
nor U19990 (N_19990,N_19201,N_18893);
nor U19991 (N_19991,N_18103,N_18081);
nand U19992 (N_19992,N_19381,N_18794);
xnor U19993 (N_19993,N_19165,N_18125);
nand U19994 (N_19994,N_19496,N_18879);
or U19995 (N_19995,N_18480,N_18159);
xnor U19996 (N_19996,N_18444,N_18860);
and U19997 (N_19997,N_18508,N_19443);
nor U19998 (N_19998,N_18415,N_18215);
or U19999 (N_19999,N_18801,N_19278);
and U20000 (N_20000,N_18427,N_19480);
and U20001 (N_20001,N_18642,N_18834);
and U20002 (N_20002,N_18048,N_18748);
nor U20003 (N_20003,N_18026,N_18756);
xor U20004 (N_20004,N_18939,N_18895);
xnor U20005 (N_20005,N_18187,N_18991);
or U20006 (N_20006,N_18142,N_18903);
nor U20007 (N_20007,N_19265,N_18118);
nor U20008 (N_20008,N_18138,N_19053);
or U20009 (N_20009,N_18830,N_18521);
nand U20010 (N_20010,N_18360,N_18864);
and U20011 (N_20011,N_18447,N_19402);
xnor U20012 (N_20012,N_18246,N_18405);
or U20013 (N_20013,N_18626,N_18791);
nand U20014 (N_20014,N_18183,N_19234);
or U20015 (N_20015,N_18078,N_19136);
or U20016 (N_20016,N_19110,N_18828);
xnor U20017 (N_20017,N_18247,N_18700);
nand U20018 (N_20018,N_18327,N_18527);
nor U20019 (N_20019,N_18292,N_18467);
or U20020 (N_20020,N_19261,N_19038);
nor U20021 (N_20021,N_19330,N_18796);
nor U20022 (N_20022,N_19409,N_18836);
nor U20023 (N_20023,N_18615,N_18032);
nor U20024 (N_20024,N_19382,N_18067);
xor U20025 (N_20025,N_19231,N_18431);
xor U20026 (N_20026,N_19284,N_19251);
xnor U20027 (N_20027,N_18996,N_18918);
nor U20028 (N_20028,N_18256,N_18990);
nand U20029 (N_20029,N_18872,N_19386);
xor U20030 (N_20030,N_19098,N_18244);
nor U20031 (N_20031,N_18221,N_18172);
nand U20032 (N_20032,N_18812,N_18060);
xor U20033 (N_20033,N_18354,N_19166);
or U20034 (N_20034,N_18650,N_18023);
xor U20035 (N_20035,N_18833,N_18619);
or U20036 (N_20036,N_18318,N_18044);
or U20037 (N_20037,N_18741,N_18656);
xnor U20038 (N_20038,N_19145,N_18952);
nor U20039 (N_20039,N_18285,N_18880);
nand U20040 (N_20040,N_18697,N_18908);
and U20041 (N_20041,N_18362,N_18313);
or U20042 (N_20042,N_18511,N_18660);
xnor U20043 (N_20043,N_18299,N_18777);
xor U20044 (N_20044,N_19141,N_18315);
nand U20045 (N_20045,N_19303,N_19019);
or U20046 (N_20046,N_18742,N_19305);
or U20047 (N_20047,N_18610,N_19014);
xnor U20048 (N_20048,N_18645,N_18124);
nor U20049 (N_20049,N_18458,N_18694);
xnor U20050 (N_20050,N_18481,N_18312);
xor U20051 (N_20051,N_18092,N_19457);
xor U20052 (N_20052,N_18840,N_18673);
and U20053 (N_20053,N_19131,N_18536);
nand U20054 (N_20054,N_19462,N_18385);
or U20055 (N_20055,N_18049,N_19317);
or U20056 (N_20056,N_18341,N_18530);
or U20057 (N_20057,N_19022,N_19400);
xnor U20058 (N_20058,N_18132,N_18979);
or U20059 (N_20059,N_18043,N_18117);
xor U20060 (N_20060,N_18363,N_19107);
xor U20061 (N_20061,N_18392,N_18038);
xnor U20062 (N_20062,N_19345,N_18569);
xnor U20063 (N_20063,N_18372,N_19412);
nor U20064 (N_20064,N_18570,N_18662);
nor U20065 (N_20065,N_18696,N_18321);
xnor U20066 (N_20066,N_19051,N_19037);
and U20067 (N_20067,N_19224,N_18808);
or U20068 (N_20068,N_19028,N_18827);
and U20069 (N_20069,N_18166,N_19490);
and U20070 (N_20070,N_18295,N_18507);
nor U20071 (N_20071,N_19481,N_18789);
or U20072 (N_20072,N_19424,N_19340);
and U20073 (N_20073,N_18380,N_18414);
nand U20074 (N_20074,N_18368,N_19390);
nor U20075 (N_20075,N_18665,N_19124);
nand U20076 (N_20076,N_18227,N_19135);
nand U20077 (N_20077,N_19227,N_18553);
or U20078 (N_20078,N_19380,N_18846);
nand U20079 (N_20079,N_18095,N_19364);
or U20080 (N_20080,N_18714,N_19499);
or U20081 (N_20081,N_19442,N_19010);
and U20082 (N_20082,N_18279,N_19239);
nand U20083 (N_20083,N_18605,N_18194);
or U20084 (N_20084,N_18204,N_19458);
and U20085 (N_20085,N_18749,N_18374);
and U20086 (N_20086,N_18894,N_18774);
nor U20087 (N_20087,N_18240,N_18857);
or U20088 (N_20088,N_18071,N_19240);
xor U20089 (N_20089,N_18625,N_18086);
nor U20090 (N_20090,N_19339,N_19070);
nand U20091 (N_20091,N_18185,N_18406);
nand U20092 (N_20092,N_18866,N_18975);
and U20093 (N_20093,N_18231,N_18309);
and U20094 (N_20094,N_19257,N_18687);
nand U20095 (N_20095,N_18932,N_18059);
or U20096 (N_20096,N_19016,N_18844);
nor U20097 (N_20097,N_18047,N_18442);
nand U20098 (N_20098,N_18677,N_18981);
and U20099 (N_20099,N_19350,N_18499);
nand U20100 (N_20100,N_18854,N_18943);
xor U20101 (N_20101,N_18905,N_19101);
or U20102 (N_20102,N_18460,N_19052);
xnor U20103 (N_20103,N_18571,N_19212);
or U20104 (N_20104,N_18680,N_18781);
nand U20105 (N_20105,N_18706,N_18152);
and U20106 (N_20106,N_19274,N_18859);
nor U20107 (N_20107,N_19232,N_19002);
nand U20108 (N_20108,N_18199,N_18422);
and U20109 (N_20109,N_18999,N_18260);
xor U20110 (N_20110,N_18920,N_18620);
or U20111 (N_20111,N_19029,N_18211);
and U20112 (N_20112,N_18973,N_18120);
and U20113 (N_20113,N_18628,N_19044);
nor U20114 (N_20114,N_19144,N_18647);
or U20115 (N_20115,N_19178,N_18572);
nand U20116 (N_20116,N_19269,N_18174);
or U20117 (N_20117,N_18938,N_18097);
and U20118 (N_20118,N_19335,N_19360);
nor U20119 (N_20119,N_19205,N_18338);
xor U20120 (N_20120,N_18870,N_19026);
and U20121 (N_20121,N_18105,N_18024);
and U20122 (N_20122,N_18381,N_19146);
nand U20123 (N_20123,N_19483,N_18408);
nand U20124 (N_20124,N_18219,N_18771);
and U20125 (N_20125,N_19195,N_18064);
xnor U20126 (N_20126,N_18679,N_18994);
xnor U20127 (N_20127,N_18735,N_18786);
or U20128 (N_20128,N_18397,N_18128);
and U20129 (N_20129,N_18783,N_19123);
nor U20130 (N_20130,N_19045,N_18958);
or U20131 (N_20131,N_19297,N_18479);
nand U20132 (N_20132,N_18178,N_18592);
xnor U20133 (N_20133,N_18972,N_18653);
and U20134 (N_20134,N_18886,N_18021);
and U20135 (N_20135,N_19482,N_18702);
and U20136 (N_20136,N_18404,N_18358);
xor U20137 (N_20137,N_19361,N_18022);
nor U20138 (N_20138,N_19182,N_19314);
nor U20139 (N_20139,N_18430,N_18607);
nor U20140 (N_20140,N_18817,N_18882);
xnor U20141 (N_20141,N_19455,N_18887);
nor U20142 (N_20142,N_18262,N_19075);
and U20143 (N_20143,N_18736,N_18466);
nor U20144 (N_20144,N_18502,N_19291);
or U20145 (N_20145,N_18203,N_18503);
nor U20146 (N_20146,N_19470,N_18398);
or U20147 (N_20147,N_19401,N_18597);
and U20148 (N_20148,N_18957,N_18967);
xnor U20149 (N_20149,N_18147,N_19270);
xnor U20150 (N_20150,N_18255,N_19474);
nand U20151 (N_20151,N_18689,N_19397);
nor U20152 (N_20152,N_18041,N_19347);
and U20153 (N_20153,N_19370,N_18316);
nor U20154 (N_20154,N_18324,N_18701);
and U20155 (N_20155,N_19271,N_18254);
or U20156 (N_20156,N_19142,N_18491);
nor U20157 (N_20157,N_18788,N_18691);
xnor U20158 (N_20158,N_19336,N_18320);
xnor U20159 (N_20159,N_18593,N_19255);
xnor U20160 (N_20160,N_18675,N_18528);
nand U20161 (N_20161,N_18473,N_19398);
and U20162 (N_20162,N_18652,N_18730);
xnor U20163 (N_20163,N_18235,N_19431);
or U20164 (N_20164,N_18326,N_18450);
xnor U20165 (N_20165,N_18884,N_18345);
nand U20166 (N_20166,N_19351,N_18782);
and U20167 (N_20167,N_18070,N_19133);
nand U20168 (N_20168,N_18083,N_18298);
and U20169 (N_20169,N_19170,N_18575);
or U20170 (N_20170,N_19089,N_18035);
nand U20171 (N_20171,N_18770,N_18488);
nor U20172 (N_20172,N_18549,N_18002);
and U20173 (N_20173,N_18869,N_18485);
nor U20174 (N_20174,N_19230,N_19264);
or U20175 (N_20175,N_18608,N_18734);
or U20176 (N_20176,N_18959,N_18541);
xor U20177 (N_20177,N_19092,N_18334);
nand U20178 (N_20178,N_18627,N_19315);
nand U20179 (N_20179,N_19173,N_18028);
nor U20180 (N_20180,N_18816,N_18708);
nor U20181 (N_20181,N_18305,N_18261);
xnor U20182 (N_20182,N_19369,N_19292);
nor U20183 (N_20183,N_18498,N_18573);
nand U20184 (N_20184,N_18600,N_19059);
nand U20185 (N_20185,N_18897,N_19440);
nor U20186 (N_20186,N_18332,N_18713);
xor U20187 (N_20187,N_18425,N_18557);
xnor U20188 (N_20188,N_19311,N_18190);
xor U20189 (N_20189,N_18715,N_18039);
or U20190 (N_20190,N_18108,N_18902);
or U20191 (N_20191,N_18928,N_19042);
and U20192 (N_20192,N_18061,N_18727);
nand U20193 (N_20193,N_19221,N_18012);
xor U20194 (N_20194,N_18633,N_19448);
or U20195 (N_20195,N_19169,N_18563);
and U20196 (N_20196,N_18448,N_19406);
nand U20197 (N_20197,N_18151,N_18161);
and U20198 (N_20198,N_19082,N_19451);
xor U20199 (N_20199,N_19120,N_18956);
nor U20200 (N_20200,N_19163,N_19423);
xor U20201 (N_20201,N_19079,N_18308);
or U20202 (N_20202,N_18807,N_19223);
and U20203 (N_20203,N_19191,N_18825);
nor U20204 (N_20204,N_19427,N_18224);
nand U20205 (N_20205,N_18602,N_18409);
xor U20206 (N_20206,N_18898,N_18270);
nand U20207 (N_20207,N_18189,N_19459);
nand U20208 (N_20208,N_18657,N_19395);
nor U20209 (N_20209,N_18544,N_19129);
and U20210 (N_20210,N_18618,N_18579);
xnor U20211 (N_20211,N_18595,N_18944);
nand U20212 (N_20212,N_19088,N_18989);
nor U20213 (N_20213,N_18242,N_19122);
nand U20214 (N_20214,N_18371,N_18276);
xnor U20215 (N_20215,N_18510,N_18160);
and U20216 (N_20216,N_18874,N_18856);
and U20217 (N_20217,N_18824,N_18823);
nand U20218 (N_20218,N_19267,N_18027);
or U20219 (N_20219,N_19337,N_19196);
nor U20220 (N_20220,N_18171,N_19249);
nand U20221 (N_20221,N_18892,N_18889);
nor U20222 (N_20222,N_19057,N_19228);
xnor U20223 (N_20223,N_18641,N_18949);
or U20224 (N_20224,N_18018,N_19064);
nor U20225 (N_20225,N_18217,N_18229);
and U20226 (N_20226,N_19126,N_18539);
nor U20227 (N_20227,N_18906,N_18531);
and U20228 (N_20228,N_18079,N_19484);
and U20229 (N_20229,N_19359,N_18867);
xor U20230 (N_20230,N_18861,N_19012);
nand U20231 (N_20231,N_18176,N_19159);
and U20232 (N_20232,N_18798,N_19414);
nor U20233 (N_20233,N_19229,N_18112);
nor U20234 (N_20234,N_18496,N_18655);
nand U20235 (N_20235,N_18040,N_18073);
xnor U20236 (N_20236,N_18551,N_18454);
and U20237 (N_20237,N_18379,N_18196);
xor U20238 (N_20238,N_19050,N_18085);
nor U20239 (N_20239,N_19179,N_18239);
or U20240 (N_20240,N_18062,N_18195);
nand U20241 (N_20241,N_19185,N_18871);
nand U20242 (N_20242,N_18951,N_19393);
xor U20243 (N_20243,N_18243,N_18429);
nand U20244 (N_20244,N_18698,N_19419);
nand U20245 (N_20245,N_18395,N_18776);
nand U20246 (N_20246,N_19049,N_18342);
nor U20247 (N_20247,N_18277,N_18248);
or U20248 (N_20248,N_18710,N_18440);
or U20249 (N_20249,N_18692,N_18997);
and U20250 (N_20250,N_18106,N_18250);
nor U20251 (N_20251,N_18547,N_18894);
or U20252 (N_20252,N_19364,N_18903);
xnor U20253 (N_20253,N_18932,N_18539);
xor U20254 (N_20254,N_19444,N_18377);
or U20255 (N_20255,N_18435,N_18096);
or U20256 (N_20256,N_19029,N_18162);
or U20257 (N_20257,N_18670,N_18613);
nor U20258 (N_20258,N_18768,N_19209);
xor U20259 (N_20259,N_19262,N_19330);
nor U20260 (N_20260,N_19171,N_18313);
nand U20261 (N_20261,N_18858,N_19292);
nand U20262 (N_20262,N_18926,N_19318);
and U20263 (N_20263,N_19457,N_18975);
or U20264 (N_20264,N_18875,N_18826);
or U20265 (N_20265,N_19016,N_18446);
and U20266 (N_20266,N_18328,N_18530);
xor U20267 (N_20267,N_18727,N_19066);
or U20268 (N_20268,N_18084,N_18492);
or U20269 (N_20269,N_18767,N_19010);
and U20270 (N_20270,N_18656,N_19036);
or U20271 (N_20271,N_18087,N_18270);
xnor U20272 (N_20272,N_18376,N_18638);
xor U20273 (N_20273,N_18315,N_18104);
xor U20274 (N_20274,N_18946,N_18175);
xnor U20275 (N_20275,N_18333,N_18538);
nor U20276 (N_20276,N_18114,N_18392);
or U20277 (N_20277,N_19154,N_18823);
nor U20278 (N_20278,N_18776,N_19118);
or U20279 (N_20279,N_19294,N_18670);
and U20280 (N_20280,N_18413,N_18673);
xor U20281 (N_20281,N_18978,N_18509);
nand U20282 (N_20282,N_19372,N_19329);
nor U20283 (N_20283,N_18149,N_18186);
xnor U20284 (N_20284,N_19477,N_18400);
nor U20285 (N_20285,N_18831,N_18024);
and U20286 (N_20286,N_19239,N_19176);
or U20287 (N_20287,N_18472,N_18560);
or U20288 (N_20288,N_18102,N_18713);
nor U20289 (N_20289,N_18259,N_18239);
nand U20290 (N_20290,N_18492,N_18601);
xnor U20291 (N_20291,N_19444,N_18091);
and U20292 (N_20292,N_18521,N_18295);
nand U20293 (N_20293,N_18895,N_19179);
nand U20294 (N_20294,N_19447,N_19443);
xor U20295 (N_20295,N_18714,N_18266);
xnor U20296 (N_20296,N_18153,N_19480);
nor U20297 (N_20297,N_19308,N_18282);
nor U20298 (N_20298,N_19220,N_19042);
and U20299 (N_20299,N_18064,N_18315);
nor U20300 (N_20300,N_18519,N_19108);
nor U20301 (N_20301,N_19379,N_18664);
and U20302 (N_20302,N_18834,N_18911);
xor U20303 (N_20303,N_18868,N_19359);
or U20304 (N_20304,N_18899,N_18264);
and U20305 (N_20305,N_18953,N_18972);
nand U20306 (N_20306,N_18775,N_18844);
xnor U20307 (N_20307,N_18900,N_18636);
nand U20308 (N_20308,N_18690,N_19012);
nor U20309 (N_20309,N_18717,N_19040);
xor U20310 (N_20310,N_18286,N_18121);
nor U20311 (N_20311,N_18594,N_19344);
nor U20312 (N_20312,N_19121,N_19341);
nor U20313 (N_20313,N_18314,N_18306);
xor U20314 (N_20314,N_19137,N_18457);
nand U20315 (N_20315,N_18302,N_19433);
nand U20316 (N_20316,N_18073,N_18929);
nand U20317 (N_20317,N_19179,N_19461);
xor U20318 (N_20318,N_19448,N_19485);
nand U20319 (N_20319,N_18006,N_19382);
nand U20320 (N_20320,N_18196,N_18370);
xor U20321 (N_20321,N_18554,N_19187);
nand U20322 (N_20322,N_19424,N_18770);
and U20323 (N_20323,N_19285,N_19433);
or U20324 (N_20324,N_18100,N_18259);
or U20325 (N_20325,N_19354,N_18612);
xor U20326 (N_20326,N_18471,N_19008);
nand U20327 (N_20327,N_19322,N_18773);
or U20328 (N_20328,N_18150,N_18936);
xor U20329 (N_20329,N_18319,N_18815);
nor U20330 (N_20330,N_18489,N_19095);
xor U20331 (N_20331,N_18031,N_19025);
xor U20332 (N_20332,N_18035,N_18091);
or U20333 (N_20333,N_18887,N_19175);
nand U20334 (N_20334,N_19109,N_18095);
nor U20335 (N_20335,N_19375,N_18283);
or U20336 (N_20336,N_19053,N_18666);
xnor U20337 (N_20337,N_18035,N_18895);
xor U20338 (N_20338,N_19064,N_18472);
nand U20339 (N_20339,N_18186,N_19377);
xor U20340 (N_20340,N_19480,N_18766);
nand U20341 (N_20341,N_18796,N_18176);
nor U20342 (N_20342,N_18954,N_19283);
nand U20343 (N_20343,N_18776,N_18405);
nor U20344 (N_20344,N_18579,N_19334);
or U20345 (N_20345,N_19322,N_18746);
or U20346 (N_20346,N_19240,N_19160);
nor U20347 (N_20347,N_18075,N_18269);
nor U20348 (N_20348,N_19323,N_18346);
nor U20349 (N_20349,N_18110,N_18389);
xnor U20350 (N_20350,N_18476,N_18721);
or U20351 (N_20351,N_18148,N_19110);
or U20352 (N_20352,N_18440,N_19432);
or U20353 (N_20353,N_18283,N_19128);
nand U20354 (N_20354,N_18225,N_18754);
or U20355 (N_20355,N_18117,N_18973);
and U20356 (N_20356,N_19323,N_18276);
xnor U20357 (N_20357,N_19439,N_19081);
nand U20358 (N_20358,N_18192,N_19149);
nor U20359 (N_20359,N_18084,N_18520);
nand U20360 (N_20360,N_18841,N_19082);
nor U20361 (N_20361,N_18270,N_18839);
xor U20362 (N_20362,N_18636,N_19066);
nand U20363 (N_20363,N_18609,N_18921);
or U20364 (N_20364,N_19036,N_18509);
nand U20365 (N_20365,N_19466,N_18305);
or U20366 (N_20366,N_19309,N_19399);
xnor U20367 (N_20367,N_18631,N_19436);
or U20368 (N_20368,N_18370,N_18811);
xnor U20369 (N_20369,N_18277,N_18044);
or U20370 (N_20370,N_18906,N_18374);
and U20371 (N_20371,N_18309,N_19146);
nand U20372 (N_20372,N_18367,N_18297);
and U20373 (N_20373,N_19109,N_18628);
xnor U20374 (N_20374,N_18547,N_18262);
and U20375 (N_20375,N_18340,N_18706);
nand U20376 (N_20376,N_18413,N_18705);
or U20377 (N_20377,N_18418,N_18801);
xor U20378 (N_20378,N_18348,N_19397);
or U20379 (N_20379,N_18613,N_19369);
xor U20380 (N_20380,N_18941,N_18587);
xnor U20381 (N_20381,N_18923,N_19126);
nor U20382 (N_20382,N_18839,N_18784);
and U20383 (N_20383,N_19477,N_18445);
or U20384 (N_20384,N_19305,N_18334);
or U20385 (N_20385,N_18062,N_19006);
and U20386 (N_20386,N_19325,N_19331);
and U20387 (N_20387,N_19215,N_18325);
and U20388 (N_20388,N_18285,N_19424);
or U20389 (N_20389,N_18572,N_18832);
nand U20390 (N_20390,N_18163,N_19397);
and U20391 (N_20391,N_18849,N_18734);
and U20392 (N_20392,N_19047,N_19075);
and U20393 (N_20393,N_19215,N_19421);
or U20394 (N_20394,N_18102,N_18055);
and U20395 (N_20395,N_18200,N_18032);
xnor U20396 (N_20396,N_18925,N_18725);
and U20397 (N_20397,N_18050,N_19461);
nand U20398 (N_20398,N_19202,N_18987);
nor U20399 (N_20399,N_18042,N_18906);
or U20400 (N_20400,N_18281,N_18761);
and U20401 (N_20401,N_19231,N_18116);
nand U20402 (N_20402,N_19086,N_19277);
xnor U20403 (N_20403,N_18685,N_19271);
nor U20404 (N_20404,N_18994,N_18306);
and U20405 (N_20405,N_18427,N_18799);
nor U20406 (N_20406,N_18579,N_18774);
or U20407 (N_20407,N_18198,N_18663);
nand U20408 (N_20408,N_18796,N_18913);
nor U20409 (N_20409,N_19183,N_19372);
nand U20410 (N_20410,N_18391,N_19444);
nor U20411 (N_20411,N_18812,N_19119);
xor U20412 (N_20412,N_18357,N_19479);
nor U20413 (N_20413,N_18232,N_19293);
or U20414 (N_20414,N_18225,N_18876);
and U20415 (N_20415,N_19278,N_18915);
and U20416 (N_20416,N_19104,N_18556);
nor U20417 (N_20417,N_19013,N_19008);
and U20418 (N_20418,N_19383,N_19210);
nand U20419 (N_20419,N_19329,N_18580);
nor U20420 (N_20420,N_19394,N_18605);
nor U20421 (N_20421,N_18469,N_18501);
nor U20422 (N_20422,N_18497,N_18345);
nand U20423 (N_20423,N_18096,N_18315);
nor U20424 (N_20424,N_19346,N_19311);
nor U20425 (N_20425,N_18099,N_19296);
or U20426 (N_20426,N_18884,N_18150);
xor U20427 (N_20427,N_18354,N_18839);
xor U20428 (N_20428,N_18584,N_18258);
nand U20429 (N_20429,N_18780,N_19059);
nand U20430 (N_20430,N_18436,N_19032);
nor U20431 (N_20431,N_19148,N_18343);
xor U20432 (N_20432,N_18815,N_18068);
xnor U20433 (N_20433,N_18394,N_19451);
and U20434 (N_20434,N_18010,N_18756);
or U20435 (N_20435,N_18659,N_18970);
xnor U20436 (N_20436,N_18522,N_18443);
nand U20437 (N_20437,N_18642,N_18675);
nand U20438 (N_20438,N_19202,N_19201);
xnor U20439 (N_20439,N_18021,N_18765);
and U20440 (N_20440,N_19310,N_19233);
or U20441 (N_20441,N_18120,N_18047);
and U20442 (N_20442,N_19336,N_19012);
and U20443 (N_20443,N_18816,N_19472);
or U20444 (N_20444,N_19212,N_19114);
xor U20445 (N_20445,N_18433,N_19341);
xor U20446 (N_20446,N_18036,N_19101);
nor U20447 (N_20447,N_18186,N_18299);
nor U20448 (N_20448,N_18745,N_18830);
or U20449 (N_20449,N_18515,N_18854);
and U20450 (N_20450,N_18141,N_18465);
nor U20451 (N_20451,N_19027,N_18669);
and U20452 (N_20452,N_19376,N_18161);
xnor U20453 (N_20453,N_19368,N_19340);
and U20454 (N_20454,N_18706,N_18564);
nor U20455 (N_20455,N_18698,N_19411);
or U20456 (N_20456,N_19364,N_19389);
nand U20457 (N_20457,N_19325,N_19476);
xnor U20458 (N_20458,N_18099,N_18026);
and U20459 (N_20459,N_18346,N_18006);
or U20460 (N_20460,N_19200,N_18103);
xnor U20461 (N_20461,N_18834,N_19434);
and U20462 (N_20462,N_19223,N_19045);
and U20463 (N_20463,N_18422,N_18498);
or U20464 (N_20464,N_18738,N_18537);
xnor U20465 (N_20465,N_18086,N_18667);
and U20466 (N_20466,N_18709,N_18148);
nand U20467 (N_20467,N_18792,N_18756);
or U20468 (N_20468,N_18857,N_18787);
xnor U20469 (N_20469,N_18880,N_19422);
nand U20470 (N_20470,N_18825,N_18798);
nand U20471 (N_20471,N_18011,N_18430);
or U20472 (N_20472,N_18480,N_18696);
or U20473 (N_20473,N_19281,N_19317);
nor U20474 (N_20474,N_18820,N_18361);
xor U20475 (N_20475,N_19351,N_18377);
nor U20476 (N_20476,N_18478,N_19193);
nor U20477 (N_20477,N_19134,N_18267);
nor U20478 (N_20478,N_19263,N_19028);
and U20479 (N_20479,N_19071,N_18862);
xnor U20480 (N_20480,N_18709,N_18458);
or U20481 (N_20481,N_19259,N_19425);
and U20482 (N_20482,N_18193,N_19179);
and U20483 (N_20483,N_18501,N_18034);
nor U20484 (N_20484,N_19094,N_19418);
and U20485 (N_20485,N_18421,N_19416);
nand U20486 (N_20486,N_19114,N_18835);
nor U20487 (N_20487,N_18339,N_18908);
nor U20488 (N_20488,N_18869,N_18044);
or U20489 (N_20489,N_18566,N_18323);
xnor U20490 (N_20490,N_18208,N_18994);
or U20491 (N_20491,N_18166,N_18772);
and U20492 (N_20492,N_18895,N_18611);
nor U20493 (N_20493,N_18750,N_19473);
or U20494 (N_20494,N_19232,N_18795);
and U20495 (N_20495,N_18058,N_19093);
nand U20496 (N_20496,N_19065,N_19001);
and U20497 (N_20497,N_18178,N_18980);
or U20498 (N_20498,N_18284,N_18876);
and U20499 (N_20499,N_19495,N_18288);
nand U20500 (N_20500,N_19222,N_18372);
nor U20501 (N_20501,N_19284,N_18514);
nand U20502 (N_20502,N_18265,N_18649);
and U20503 (N_20503,N_19458,N_18626);
nor U20504 (N_20504,N_18996,N_19357);
nor U20505 (N_20505,N_18157,N_19343);
or U20506 (N_20506,N_19446,N_19103);
nand U20507 (N_20507,N_19040,N_19131);
nor U20508 (N_20508,N_18430,N_19404);
or U20509 (N_20509,N_18496,N_18523);
xnor U20510 (N_20510,N_19277,N_19438);
nor U20511 (N_20511,N_19108,N_18502);
or U20512 (N_20512,N_18095,N_18870);
nand U20513 (N_20513,N_18310,N_19363);
nor U20514 (N_20514,N_18734,N_19103);
or U20515 (N_20515,N_18427,N_19067);
nand U20516 (N_20516,N_19325,N_18303);
or U20517 (N_20517,N_18625,N_19272);
and U20518 (N_20518,N_18535,N_19240);
xnor U20519 (N_20519,N_18105,N_18604);
or U20520 (N_20520,N_19197,N_18399);
or U20521 (N_20521,N_19159,N_19162);
nand U20522 (N_20522,N_18475,N_19363);
nand U20523 (N_20523,N_18087,N_18899);
or U20524 (N_20524,N_19489,N_19452);
nand U20525 (N_20525,N_18655,N_18857);
xor U20526 (N_20526,N_18810,N_18514);
and U20527 (N_20527,N_18864,N_18888);
and U20528 (N_20528,N_19133,N_18675);
nand U20529 (N_20529,N_18035,N_18489);
xor U20530 (N_20530,N_18155,N_18272);
and U20531 (N_20531,N_19490,N_18172);
nand U20532 (N_20532,N_18233,N_19275);
xor U20533 (N_20533,N_18246,N_18930);
nand U20534 (N_20534,N_18353,N_18487);
xor U20535 (N_20535,N_19191,N_18880);
or U20536 (N_20536,N_19080,N_18770);
and U20537 (N_20537,N_19298,N_18242);
xor U20538 (N_20538,N_19253,N_18909);
xnor U20539 (N_20539,N_18649,N_18627);
nand U20540 (N_20540,N_18155,N_18383);
nand U20541 (N_20541,N_18558,N_18000);
xor U20542 (N_20542,N_19082,N_19275);
nand U20543 (N_20543,N_19488,N_19119);
nand U20544 (N_20544,N_19389,N_18189);
or U20545 (N_20545,N_18310,N_18908);
and U20546 (N_20546,N_19283,N_19061);
nor U20547 (N_20547,N_18403,N_18110);
and U20548 (N_20548,N_18153,N_19025);
nor U20549 (N_20549,N_18849,N_19092);
or U20550 (N_20550,N_19402,N_18030);
or U20551 (N_20551,N_18655,N_18817);
or U20552 (N_20552,N_18524,N_19110);
nand U20553 (N_20553,N_19386,N_18369);
and U20554 (N_20554,N_18679,N_18307);
xnor U20555 (N_20555,N_18121,N_18993);
or U20556 (N_20556,N_18543,N_18824);
or U20557 (N_20557,N_18661,N_18833);
and U20558 (N_20558,N_18898,N_19006);
and U20559 (N_20559,N_19207,N_18338);
or U20560 (N_20560,N_18220,N_18072);
and U20561 (N_20561,N_18162,N_18800);
or U20562 (N_20562,N_19265,N_18252);
nor U20563 (N_20563,N_18624,N_19098);
nor U20564 (N_20564,N_18860,N_18005);
nor U20565 (N_20565,N_19279,N_19478);
nand U20566 (N_20566,N_18762,N_19260);
and U20567 (N_20567,N_19004,N_18474);
or U20568 (N_20568,N_18866,N_18534);
or U20569 (N_20569,N_19243,N_18643);
nand U20570 (N_20570,N_18128,N_19203);
or U20571 (N_20571,N_19199,N_18263);
nand U20572 (N_20572,N_18515,N_19392);
nor U20573 (N_20573,N_19132,N_18424);
nor U20574 (N_20574,N_19400,N_18322);
and U20575 (N_20575,N_18574,N_18609);
nand U20576 (N_20576,N_18645,N_18714);
or U20577 (N_20577,N_18414,N_18521);
nor U20578 (N_20578,N_18455,N_18351);
xor U20579 (N_20579,N_18033,N_18043);
nand U20580 (N_20580,N_18352,N_18800);
and U20581 (N_20581,N_18943,N_18765);
and U20582 (N_20582,N_18077,N_18469);
xor U20583 (N_20583,N_18089,N_19279);
xnor U20584 (N_20584,N_18986,N_19167);
nand U20585 (N_20585,N_18832,N_18413);
and U20586 (N_20586,N_19159,N_18458);
nand U20587 (N_20587,N_18674,N_18412);
nor U20588 (N_20588,N_18375,N_19089);
or U20589 (N_20589,N_19297,N_19380);
or U20590 (N_20590,N_18998,N_19126);
xor U20591 (N_20591,N_18560,N_18891);
and U20592 (N_20592,N_18422,N_18593);
or U20593 (N_20593,N_18872,N_19373);
nor U20594 (N_20594,N_18738,N_18321);
or U20595 (N_20595,N_19424,N_18258);
nor U20596 (N_20596,N_18956,N_19418);
and U20597 (N_20597,N_18500,N_18747);
or U20598 (N_20598,N_18808,N_18448);
nor U20599 (N_20599,N_18855,N_19436);
and U20600 (N_20600,N_19017,N_18990);
and U20601 (N_20601,N_18762,N_18818);
and U20602 (N_20602,N_19383,N_19186);
nand U20603 (N_20603,N_19175,N_18755);
xnor U20604 (N_20604,N_19434,N_18572);
or U20605 (N_20605,N_18233,N_19401);
nand U20606 (N_20606,N_19464,N_18917);
and U20607 (N_20607,N_18231,N_18673);
nand U20608 (N_20608,N_18313,N_18027);
and U20609 (N_20609,N_19025,N_18488);
nor U20610 (N_20610,N_19181,N_18123);
or U20611 (N_20611,N_19040,N_18183);
nor U20612 (N_20612,N_18457,N_18129);
nor U20613 (N_20613,N_18581,N_18885);
nor U20614 (N_20614,N_18027,N_19078);
nand U20615 (N_20615,N_19033,N_19391);
xor U20616 (N_20616,N_18271,N_18510);
nor U20617 (N_20617,N_18072,N_18203);
xor U20618 (N_20618,N_18508,N_18008);
and U20619 (N_20619,N_18924,N_18152);
nor U20620 (N_20620,N_19444,N_18564);
nor U20621 (N_20621,N_18590,N_18363);
nand U20622 (N_20622,N_19063,N_18794);
nor U20623 (N_20623,N_18011,N_18708);
and U20624 (N_20624,N_18865,N_18803);
and U20625 (N_20625,N_19093,N_19282);
or U20626 (N_20626,N_18641,N_19375);
or U20627 (N_20627,N_19496,N_19008);
or U20628 (N_20628,N_19292,N_18296);
nand U20629 (N_20629,N_18429,N_19348);
xnor U20630 (N_20630,N_18161,N_18236);
and U20631 (N_20631,N_18372,N_18462);
and U20632 (N_20632,N_19378,N_19037);
nor U20633 (N_20633,N_18789,N_18250);
nand U20634 (N_20634,N_18101,N_18694);
and U20635 (N_20635,N_19352,N_18993);
nor U20636 (N_20636,N_19484,N_18988);
or U20637 (N_20637,N_19246,N_19426);
xor U20638 (N_20638,N_18049,N_18146);
or U20639 (N_20639,N_18442,N_19398);
or U20640 (N_20640,N_18640,N_18226);
xnor U20641 (N_20641,N_18066,N_19040);
xnor U20642 (N_20642,N_18897,N_18735);
nor U20643 (N_20643,N_18298,N_19210);
nor U20644 (N_20644,N_18551,N_18285);
or U20645 (N_20645,N_19281,N_18990);
or U20646 (N_20646,N_18659,N_18404);
nor U20647 (N_20647,N_18650,N_18181);
nand U20648 (N_20648,N_18783,N_19072);
xnor U20649 (N_20649,N_19254,N_18626);
and U20650 (N_20650,N_18502,N_18119);
nor U20651 (N_20651,N_19458,N_18003);
and U20652 (N_20652,N_19423,N_19022);
nor U20653 (N_20653,N_18305,N_18008);
xor U20654 (N_20654,N_19133,N_18386);
nor U20655 (N_20655,N_19053,N_18144);
xor U20656 (N_20656,N_18712,N_19404);
and U20657 (N_20657,N_18985,N_19227);
or U20658 (N_20658,N_18004,N_18844);
or U20659 (N_20659,N_18442,N_18043);
and U20660 (N_20660,N_19033,N_18738);
nand U20661 (N_20661,N_19366,N_19252);
nand U20662 (N_20662,N_18964,N_19324);
nor U20663 (N_20663,N_19078,N_19237);
or U20664 (N_20664,N_18719,N_18670);
nor U20665 (N_20665,N_18579,N_18524);
xnor U20666 (N_20666,N_19471,N_19205);
nand U20667 (N_20667,N_18402,N_18017);
xnor U20668 (N_20668,N_18370,N_18855);
xnor U20669 (N_20669,N_18506,N_19481);
or U20670 (N_20670,N_18195,N_19233);
and U20671 (N_20671,N_18873,N_19058);
and U20672 (N_20672,N_18347,N_18089);
and U20673 (N_20673,N_18089,N_18745);
nand U20674 (N_20674,N_19148,N_18513);
nand U20675 (N_20675,N_19463,N_18402);
or U20676 (N_20676,N_19259,N_18157);
nor U20677 (N_20677,N_18552,N_18080);
or U20678 (N_20678,N_18498,N_18181);
and U20679 (N_20679,N_19038,N_18705);
xnor U20680 (N_20680,N_19265,N_19102);
nand U20681 (N_20681,N_18919,N_19420);
and U20682 (N_20682,N_18578,N_18704);
nor U20683 (N_20683,N_18344,N_19378);
and U20684 (N_20684,N_18868,N_18135);
or U20685 (N_20685,N_18353,N_19068);
nand U20686 (N_20686,N_18035,N_18169);
nor U20687 (N_20687,N_18382,N_19383);
and U20688 (N_20688,N_18498,N_18228);
or U20689 (N_20689,N_19151,N_19010);
nand U20690 (N_20690,N_19335,N_19426);
nand U20691 (N_20691,N_18326,N_18273);
xor U20692 (N_20692,N_18224,N_18626);
nand U20693 (N_20693,N_18507,N_18004);
and U20694 (N_20694,N_19155,N_18894);
or U20695 (N_20695,N_18550,N_19395);
or U20696 (N_20696,N_18254,N_19107);
or U20697 (N_20697,N_19080,N_18992);
or U20698 (N_20698,N_18132,N_18569);
xnor U20699 (N_20699,N_18503,N_19305);
or U20700 (N_20700,N_18524,N_19129);
nor U20701 (N_20701,N_19262,N_19102);
or U20702 (N_20702,N_19221,N_18208);
nand U20703 (N_20703,N_19173,N_18955);
and U20704 (N_20704,N_18292,N_19417);
xor U20705 (N_20705,N_18180,N_18421);
or U20706 (N_20706,N_18376,N_18048);
nor U20707 (N_20707,N_19105,N_19153);
xor U20708 (N_20708,N_18500,N_19394);
or U20709 (N_20709,N_19294,N_18572);
nand U20710 (N_20710,N_19296,N_18017);
nor U20711 (N_20711,N_19485,N_18202);
nand U20712 (N_20712,N_19064,N_18550);
xor U20713 (N_20713,N_19263,N_18286);
xnor U20714 (N_20714,N_19178,N_19038);
and U20715 (N_20715,N_18019,N_18022);
or U20716 (N_20716,N_18349,N_18296);
nor U20717 (N_20717,N_18634,N_18812);
nand U20718 (N_20718,N_18044,N_19281);
or U20719 (N_20719,N_19411,N_18205);
nand U20720 (N_20720,N_19449,N_18065);
xor U20721 (N_20721,N_18750,N_19367);
and U20722 (N_20722,N_19282,N_19207);
nor U20723 (N_20723,N_19232,N_18318);
or U20724 (N_20724,N_18724,N_18382);
nand U20725 (N_20725,N_18822,N_18952);
and U20726 (N_20726,N_18015,N_19416);
or U20727 (N_20727,N_18742,N_18643);
nor U20728 (N_20728,N_18536,N_18496);
nand U20729 (N_20729,N_19363,N_18391);
and U20730 (N_20730,N_18472,N_18166);
nor U20731 (N_20731,N_18526,N_19250);
nor U20732 (N_20732,N_19362,N_18916);
nand U20733 (N_20733,N_18562,N_19231);
nand U20734 (N_20734,N_18707,N_18788);
nand U20735 (N_20735,N_18553,N_18237);
nor U20736 (N_20736,N_18605,N_19277);
xnor U20737 (N_20737,N_19133,N_18912);
or U20738 (N_20738,N_18119,N_19298);
xor U20739 (N_20739,N_18763,N_19368);
xor U20740 (N_20740,N_19428,N_19294);
and U20741 (N_20741,N_18697,N_19151);
nor U20742 (N_20742,N_19317,N_18974);
and U20743 (N_20743,N_18516,N_19046);
nand U20744 (N_20744,N_18514,N_19217);
xor U20745 (N_20745,N_18974,N_18123);
xnor U20746 (N_20746,N_18484,N_18948);
nand U20747 (N_20747,N_19416,N_18133);
xnor U20748 (N_20748,N_18643,N_18446);
nand U20749 (N_20749,N_18767,N_18390);
nor U20750 (N_20750,N_19387,N_18401);
and U20751 (N_20751,N_18074,N_19357);
nand U20752 (N_20752,N_19483,N_18115);
nand U20753 (N_20753,N_19114,N_18925);
nand U20754 (N_20754,N_18181,N_18015);
and U20755 (N_20755,N_18282,N_18428);
xor U20756 (N_20756,N_19366,N_18479);
or U20757 (N_20757,N_18723,N_18968);
xor U20758 (N_20758,N_18763,N_19003);
and U20759 (N_20759,N_19158,N_18148);
and U20760 (N_20760,N_18690,N_19353);
xnor U20761 (N_20761,N_18765,N_18110);
nand U20762 (N_20762,N_19079,N_18012);
xnor U20763 (N_20763,N_18948,N_18927);
xor U20764 (N_20764,N_19351,N_18937);
nor U20765 (N_20765,N_19044,N_19275);
and U20766 (N_20766,N_18047,N_19359);
nor U20767 (N_20767,N_19177,N_18735);
xor U20768 (N_20768,N_18278,N_18618);
and U20769 (N_20769,N_18801,N_18368);
xnor U20770 (N_20770,N_19313,N_18748);
or U20771 (N_20771,N_18530,N_19322);
nand U20772 (N_20772,N_18858,N_18139);
nor U20773 (N_20773,N_19070,N_18285);
nand U20774 (N_20774,N_18347,N_18930);
xor U20775 (N_20775,N_18418,N_19486);
or U20776 (N_20776,N_18414,N_19168);
and U20777 (N_20777,N_19292,N_19363);
nor U20778 (N_20778,N_18254,N_19082);
xor U20779 (N_20779,N_18651,N_18464);
nand U20780 (N_20780,N_18821,N_18207);
nor U20781 (N_20781,N_18885,N_18476);
xor U20782 (N_20782,N_18722,N_18923);
xor U20783 (N_20783,N_19325,N_19195);
nor U20784 (N_20784,N_18391,N_18702);
nor U20785 (N_20785,N_18918,N_19397);
nor U20786 (N_20786,N_18269,N_19365);
nand U20787 (N_20787,N_18440,N_19323);
nor U20788 (N_20788,N_19094,N_18271);
and U20789 (N_20789,N_19084,N_18207);
and U20790 (N_20790,N_18251,N_19204);
nor U20791 (N_20791,N_18559,N_19045);
or U20792 (N_20792,N_19321,N_19016);
nand U20793 (N_20793,N_19131,N_19217);
nand U20794 (N_20794,N_19136,N_18964);
nand U20795 (N_20795,N_19334,N_19141);
nor U20796 (N_20796,N_18691,N_18538);
xnor U20797 (N_20797,N_19014,N_18159);
and U20798 (N_20798,N_18064,N_19217);
xnor U20799 (N_20799,N_19371,N_19050);
and U20800 (N_20800,N_18828,N_18290);
xnor U20801 (N_20801,N_18788,N_18513);
and U20802 (N_20802,N_18858,N_18726);
nor U20803 (N_20803,N_18002,N_19108);
xor U20804 (N_20804,N_18604,N_18241);
or U20805 (N_20805,N_18495,N_18757);
xnor U20806 (N_20806,N_18871,N_18710);
nor U20807 (N_20807,N_18292,N_18096);
xor U20808 (N_20808,N_19160,N_19414);
nor U20809 (N_20809,N_18520,N_18328);
or U20810 (N_20810,N_19133,N_18637);
nor U20811 (N_20811,N_19416,N_18494);
nor U20812 (N_20812,N_18236,N_18540);
and U20813 (N_20813,N_18657,N_18600);
nor U20814 (N_20814,N_18975,N_18269);
nand U20815 (N_20815,N_19338,N_19390);
xor U20816 (N_20816,N_18553,N_19016);
and U20817 (N_20817,N_18845,N_19099);
nor U20818 (N_20818,N_19275,N_18846);
or U20819 (N_20819,N_18295,N_18666);
xnor U20820 (N_20820,N_18577,N_19397);
nand U20821 (N_20821,N_18525,N_19369);
xor U20822 (N_20822,N_19051,N_18433);
nand U20823 (N_20823,N_18903,N_19322);
nand U20824 (N_20824,N_18546,N_18552);
xnor U20825 (N_20825,N_19092,N_19147);
xor U20826 (N_20826,N_18505,N_18578);
or U20827 (N_20827,N_18115,N_19404);
or U20828 (N_20828,N_19431,N_18725);
or U20829 (N_20829,N_19152,N_18557);
or U20830 (N_20830,N_19087,N_18650);
nand U20831 (N_20831,N_18783,N_18480);
xnor U20832 (N_20832,N_18556,N_19280);
nand U20833 (N_20833,N_19377,N_18850);
or U20834 (N_20834,N_18460,N_18408);
nand U20835 (N_20835,N_19199,N_19333);
or U20836 (N_20836,N_18367,N_18667);
xnor U20837 (N_20837,N_19019,N_18348);
nand U20838 (N_20838,N_18115,N_19149);
nor U20839 (N_20839,N_18622,N_19469);
and U20840 (N_20840,N_18881,N_18061);
nor U20841 (N_20841,N_18156,N_18231);
nor U20842 (N_20842,N_18305,N_18074);
or U20843 (N_20843,N_18446,N_18752);
nor U20844 (N_20844,N_19457,N_19384);
or U20845 (N_20845,N_19338,N_18810);
and U20846 (N_20846,N_19421,N_19441);
nand U20847 (N_20847,N_18207,N_18391);
and U20848 (N_20848,N_19252,N_18119);
nor U20849 (N_20849,N_18255,N_18423);
or U20850 (N_20850,N_18323,N_18641);
xor U20851 (N_20851,N_19341,N_18888);
nand U20852 (N_20852,N_18454,N_18641);
or U20853 (N_20853,N_19166,N_18893);
xor U20854 (N_20854,N_18398,N_18206);
or U20855 (N_20855,N_19093,N_18447);
nand U20856 (N_20856,N_18952,N_19090);
nand U20857 (N_20857,N_18040,N_18711);
nand U20858 (N_20858,N_18308,N_18437);
nor U20859 (N_20859,N_18762,N_19087);
xnor U20860 (N_20860,N_19400,N_18170);
nand U20861 (N_20861,N_18215,N_18691);
xor U20862 (N_20862,N_18555,N_18032);
or U20863 (N_20863,N_18512,N_18910);
xor U20864 (N_20864,N_18103,N_18016);
and U20865 (N_20865,N_19071,N_19153);
or U20866 (N_20866,N_18863,N_18049);
and U20867 (N_20867,N_18284,N_18760);
nor U20868 (N_20868,N_18864,N_19321);
xor U20869 (N_20869,N_18636,N_18155);
xor U20870 (N_20870,N_19487,N_18992);
xnor U20871 (N_20871,N_18798,N_19096);
xor U20872 (N_20872,N_19307,N_18261);
xnor U20873 (N_20873,N_18809,N_18325);
nor U20874 (N_20874,N_18643,N_18725);
nand U20875 (N_20875,N_18174,N_18567);
or U20876 (N_20876,N_19171,N_19041);
or U20877 (N_20877,N_18386,N_19356);
nor U20878 (N_20878,N_18899,N_19102);
xor U20879 (N_20879,N_19068,N_18064);
or U20880 (N_20880,N_18642,N_19363);
or U20881 (N_20881,N_18322,N_18507);
xnor U20882 (N_20882,N_18317,N_18265);
xnor U20883 (N_20883,N_18638,N_19464);
and U20884 (N_20884,N_19269,N_18699);
nand U20885 (N_20885,N_19079,N_19105);
or U20886 (N_20886,N_18204,N_19168);
or U20887 (N_20887,N_18757,N_18827);
and U20888 (N_20888,N_18008,N_18718);
xnor U20889 (N_20889,N_19141,N_19048);
nand U20890 (N_20890,N_18214,N_18237);
nor U20891 (N_20891,N_19251,N_19494);
xor U20892 (N_20892,N_18020,N_18776);
nor U20893 (N_20893,N_19275,N_18352);
and U20894 (N_20894,N_18266,N_19146);
xor U20895 (N_20895,N_18308,N_19090);
or U20896 (N_20896,N_19174,N_19498);
nor U20897 (N_20897,N_18735,N_18285);
xor U20898 (N_20898,N_19184,N_18021);
or U20899 (N_20899,N_18772,N_19420);
and U20900 (N_20900,N_19294,N_19218);
nor U20901 (N_20901,N_18336,N_18320);
xnor U20902 (N_20902,N_18507,N_19460);
and U20903 (N_20903,N_19292,N_18084);
nand U20904 (N_20904,N_19102,N_18572);
and U20905 (N_20905,N_18968,N_19010);
or U20906 (N_20906,N_19417,N_19077);
or U20907 (N_20907,N_18152,N_18316);
and U20908 (N_20908,N_18500,N_19329);
or U20909 (N_20909,N_18415,N_18653);
nand U20910 (N_20910,N_18129,N_18765);
nor U20911 (N_20911,N_19140,N_19233);
or U20912 (N_20912,N_18878,N_18731);
and U20913 (N_20913,N_19447,N_18752);
xnor U20914 (N_20914,N_18369,N_19302);
or U20915 (N_20915,N_18509,N_18081);
nand U20916 (N_20916,N_18942,N_18239);
or U20917 (N_20917,N_18117,N_19018);
and U20918 (N_20918,N_18717,N_18988);
or U20919 (N_20919,N_18185,N_18113);
xor U20920 (N_20920,N_18124,N_18131);
nand U20921 (N_20921,N_18673,N_18400);
nor U20922 (N_20922,N_18631,N_18709);
nand U20923 (N_20923,N_18904,N_18768);
nor U20924 (N_20924,N_18148,N_18115);
xor U20925 (N_20925,N_18271,N_19423);
and U20926 (N_20926,N_18523,N_18526);
and U20927 (N_20927,N_19034,N_18238);
xnor U20928 (N_20928,N_18966,N_19023);
nor U20929 (N_20929,N_18182,N_19128);
or U20930 (N_20930,N_18900,N_18464);
nor U20931 (N_20931,N_18570,N_18385);
or U20932 (N_20932,N_18563,N_19010);
or U20933 (N_20933,N_18747,N_18844);
nand U20934 (N_20934,N_18060,N_19469);
or U20935 (N_20935,N_18780,N_19119);
or U20936 (N_20936,N_18954,N_19347);
xnor U20937 (N_20937,N_18306,N_18635);
or U20938 (N_20938,N_19385,N_18621);
xor U20939 (N_20939,N_19443,N_18197);
and U20940 (N_20940,N_18423,N_18577);
or U20941 (N_20941,N_19457,N_18816);
and U20942 (N_20942,N_19120,N_19421);
and U20943 (N_20943,N_18526,N_19008);
and U20944 (N_20944,N_19467,N_18753);
and U20945 (N_20945,N_18959,N_18642);
nand U20946 (N_20946,N_18618,N_19125);
xnor U20947 (N_20947,N_18935,N_19007);
xor U20948 (N_20948,N_18094,N_18793);
nand U20949 (N_20949,N_18928,N_19155);
or U20950 (N_20950,N_19494,N_18956);
or U20951 (N_20951,N_18489,N_18261);
or U20952 (N_20952,N_19353,N_19249);
nor U20953 (N_20953,N_18405,N_18946);
nand U20954 (N_20954,N_19182,N_18718);
xor U20955 (N_20955,N_18256,N_18860);
and U20956 (N_20956,N_19012,N_19237);
or U20957 (N_20957,N_18601,N_18326);
xor U20958 (N_20958,N_19164,N_18985);
and U20959 (N_20959,N_19433,N_19076);
xor U20960 (N_20960,N_18547,N_18180);
and U20961 (N_20961,N_19402,N_19051);
nor U20962 (N_20962,N_18837,N_18041);
nor U20963 (N_20963,N_19369,N_19268);
nand U20964 (N_20964,N_18887,N_18929);
nand U20965 (N_20965,N_18214,N_18244);
nand U20966 (N_20966,N_19042,N_18830);
and U20967 (N_20967,N_18249,N_18242);
or U20968 (N_20968,N_19312,N_18108);
nor U20969 (N_20969,N_19360,N_18160);
or U20970 (N_20970,N_18331,N_18281);
nand U20971 (N_20971,N_19122,N_18422);
and U20972 (N_20972,N_19014,N_18533);
and U20973 (N_20973,N_19405,N_19441);
or U20974 (N_20974,N_19353,N_19473);
nor U20975 (N_20975,N_18750,N_18959);
nor U20976 (N_20976,N_18696,N_18179);
and U20977 (N_20977,N_19031,N_19102);
and U20978 (N_20978,N_18657,N_18461);
xor U20979 (N_20979,N_18610,N_18954);
and U20980 (N_20980,N_19098,N_18957);
xnor U20981 (N_20981,N_18848,N_18100);
and U20982 (N_20982,N_19340,N_18392);
xor U20983 (N_20983,N_18423,N_19133);
nor U20984 (N_20984,N_18290,N_19092);
xnor U20985 (N_20985,N_19078,N_19198);
and U20986 (N_20986,N_18301,N_18607);
and U20987 (N_20987,N_18771,N_18021);
xor U20988 (N_20988,N_18317,N_18852);
nand U20989 (N_20989,N_18090,N_19481);
and U20990 (N_20990,N_18025,N_18749);
or U20991 (N_20991,N_18902,N_18504);
nor U20992 (N_20992,N_19452,N_19398);
and U20993 (N_20993,N_19259,N_18799);
nand U20994 (N_20994,N_19223,N_18878);
nor U20995 (N_20995,N_18790,N_19373);
xnor U20996 (N_20996,N_18371,N_19301);
nand U20997 (N_20997,N_19093,N_18689);
nand U20998 (N_20998,N_18801,N_18750);
nand U20999 (N_20999,N_18387,N_18237);
nor U21000 (N_21000,N_20301,N_19614);
and U21001 (N_21001,N_20684,N_19855);
or U21002 (N_21002,N_20814,N_20618);
and U21003 (N_21003,N_20158,N_20332);
nor U21004 (N_21004,N_20037,N_19937);
and U21005 (N_21005,N_20006,N_20792);
nand U21006 (N_21006,N_19655,N_20511);
nand U21007 (N_21007,N_20045,N_20808);
nand U21008 (N_21008,N_20778,N_20348);
and U21009 (N_21009,N_20421,N_20382);
nor U21010 (N_21010,N_19945,N_20193);
xor U21011 (N_21011,N_20950,N_19668);
nand U21012 (N_21012,N_19892,N_20420);
or U21013 (N_21013,N_20172,N_20296);
nor U21014 (N_21014,N_20940,N_19504);
or U21015 (N_21015,N_20634,N_20327);
or U21016 (N_21016,N_20241,N_20031);
xor U21017 (N_21017,N_20957,N_20072);
xnor U21018 (N_21018,N_20519,N_19547);
and U21019 (N_21019,N_20265,N_20608);
and U21020 (N_21020,N_20110,N_20208);
nor U21021 (N_21021,N_19871,N_20611);
xor U21022 (N_21022,N_20998,N_20777);
nand U21023 (N_21023,N_20169,N_20850);
nor U21024 (N_21024,N_20727,N_20503);
or U21025 (N_21025,N_20047,N_20779);
xnor U21026 (N_21026,N_19631,N_20381);
nor U21027 (N_21027,N_19864,N_20932);
and U21028 (N_21028,N_19827,N_19860);
or U21029 (N_21029,N_20641,N_20055);
or U21030 (N_21030,N_20350,N_20418);
nor U21031 (N_21031,N_20996,N_20472);
nor U21032 (N_21032,N_20165,N_19604);
xnor U21033 (N_21033,N_19581,N_20823);
nand U21034 (N_21034,N_20685,N_19633);
xnor U21035 (N_21035,N_20657,N_20754);
nor U21036 (N_21036,N_19874,N_20580);
nand U21037 (N_21037,N_20951,N_19663);
xor U21038 (N_21038,N_20293,N_20275);
or U21039 (N_21039,N_19769,N_20197);
or U21040 (N_21040,N_20590,N_19993);
or U21041 (N_21041,N_19500,N_19972);
and U21042 (N_21042,N_20459,N_19763);
and U21043 (N_21043,N_20105,N_20461);
and U21044 (N_21044,N_20475,N_20123);
nor U21045 (N_21045,N_19841,N_19988);
nand U21046 (N_21046,N_20783,N_19897);
nand U21047 (N_21047,N_20261,N_20786);
nor U21048 (N_21048,N_19930,N_20152);
nand U21049 (N_21049,N_20127,N_19902);
and U21050 (N_21050,N_20153,N_20274);
or U21051 (N_21051,N_19625,N_19856);
xnor U21052 (N_21052,N_20336,N_20976);
nand U21053 (N_21053,N_20672,N_19576);
nor U21054 (N_21054,N_20946,N_20021);
nor U21055 (N_21055,N_19552,N_20411);
xnor U21056 (N_21056,N_19743,N_20030);
xor U21057 (N_21057,N_19608,N_19679);
nand U21058 (N_21058,N_19698,N_20116);
nand U21059 (N_21059,N_19861,N_20943);
and U21060 (N_21060,N_20745,N_19825);
nand U21061 (N_21061,N_20060,N_20582);
xnor U21062 (N_21062,N_19738,N_20528);
or U21063 (N_21063,N_19671,N_20321);
xor U21064 (N_21064,N_19853,N_20358);
nor U21065 (N_21065,N_19796,N_20191);
nand U21066 (N_21066,N_20505,N_20357);
and U21067 (N_21067,N_20266,N_20020);
or U21068 (N_21068,N_20470,N_19899);
nand U21069 (N_21069,N_20442,N_20170);
nor U21070 (N_21070,N_20757,N_20283);
and U21071 (N_21071,N_20906,N_20465);
and U21072 (N_21072,N_20662,N_20385);
or U21073 (N_21073,N_20439,N_20595);
xnor U21074 (N_21074,N_20225,N_19715);
nor U21075 (N_21075,N_20562,N_20180);
nand U21076 (N_21076,N_20676,N_19792);
nor U21077 (N_21077,N_20803,N_19741);
and U21078 (N_21078,N_19685,N_20949);
nand U21079 (N_21079,N_19757,N_20794);
nand U21080 (N_21080,N_20359,N_20237);
nor U21081 (N_21081,N_20686,N_19705);
xnor U21082 (N_21082,N_19620,N_20877);
xor U21083 (N_21083,N_19506,N_20203);
xnor U21084 (N_21084,N_19677,N_19977);
or U21085 (N_21085,N_20510,N_19508);
xor U21086 (N_21086,N_20986,N_20973);
nand U21087 (N_21087,N_20181,N_19777);
nand U21088 (N_21088,N_19915,N_20065);
and U21089 (N_21089,N_19645,N_19987);
and U21090 (N_21090,N_20196,N_20583);
nor U21091 (N_21091,N_19744,N_20092);
nor U21092 (N_21092,N_20379,N_19755);
nor U21093 (N_21093,N_20100,N_20244);
xnor U21094 (N_21094,N_19695,N_19816);
nor U21095 (N_21095,N_20854,N_19661);
or U21096 (N_21096,N_19578,N_19805);
nand U21097 (N_21097,N_19650,N_20124);
nor U21098 (N_21098,N_20085,N_20542);
and U21099 (N_21099,N_20547,N_19691);
nand U21100 (N_21100,N_20206,N_20842);
xor U21101 (N_21101,N_19501,N_20372);
xor U21102 (N_21102,N_19593,N_20975);
nor U21103 (N_21103,N_20145,N_19660);
nor U21104 (N_21104,N_19801,N_20066);
xnor U21105 (N_21105,N_20469,N_20128);
nand U21106 (N_21106,N_20650,N_20329);
xor U21107 (N_21107,N_20330,N_19727);
and U21108 (N_21108,N_20767,N_19797);
and U21109 (N_21109,N_20787,N_20003);
nor U21110 (N_21110,N_19720,N_20617);
xor U21111 (N_21111,N_20768,N_19847);
and U21112 (N_21112,N_20772,N_20119);
and U21113 (N_21113,N_20610,N_20015);
and U21114 (N_21114,N_20781,N_20924);
nand U21115 (N_21115,N_20102,N_20551);
xnor U21116 (N_21116,N_19824,N_20023);
xnor U21117 (N_21117,N_20619,N_20167);
or U21118 (N_21118,N_19959,N_19725);
xnor U21119 (N_21119,N_19640,N_19814);
or U21120 (N_21120,N_20520,N_19692);
nand U21121 (N_21121,N_20228,N_20432);
xor U21122 (N_21122,N_20623,N_20163);
xor U21123 (N_21123,N_19617,N_20680);
or U21124 (N_21124,N_20373,N_20605);
xor U21125 (N_21125,N_20424,N_19599);
nor U21126 (N_21126,N_20488,N_20088);
nand U21127 (N_21127,N_19833,N_19719);
nor U21128 (N_21128,N_20915,N_19703);
xor U21129 (N_21129,N_19817,N_19551);
xnor U21130 (N_21130,N_19994,N_19809);
nor U21131 (N_21131,N_20649,N_20199);
nand U21132 (N_21132,N_20438,N_20326);
nor U21133 (N_21133,N_19819,N_20160);
nor U21134 (N_21134,N_19564,N_20639);
nand U21135 (N_21135,N_19942,N_20426);
xor U21136 (N_21136,N_20095,N_20454);
and U21137 (N_21137,N_20747,N_20916);
and U21138 (N_21138,N_19866,N_20829);
nand U21139 (N_21139,N_20449,N_19838);
nand U21140 (N_21140,N_20937,N_20134);
xor U21141 (N_21141,N_20972,N_19546);
and U21142 (N_21142,N_20215,N_19531);
nor U21143 (N_21143,N_20004,N_19654);
nor U21144 (N_21144,N_20168,N_20809);
or U21145 (N_21145,N_20417,N_19976);
nand U21146 (N_21146,N_19549,N_20371);
nor U21147 (N_21147,N_20213,N_20585);
or U21148 (N_21148,N_20981,N_19784);
and U21149 (N_21149,N_20064,N_20271);
nand U21150 (N_21150,N_20435,N_20082);
and U21151 (N_21151,N_19764,N_19658);
nor U21152 (N_21152,N_20890,N_19693);
and U21153 (N_21153,N_20462,N_20310);
nand U21154 (N_21154,N_19510,N_20240);
or U21155 (N_21155,N_19590,N_20891);
xor U21156 (N_21156,N_20069,N_19895);
or U21157 (N_21157,N_20554,N_20759);
nand U21158 (N_21158,N_19932,N_20679);
nor U21159 (N_21159,N_20930,N_20252);
xnor U21160 (N_21160,N_19525,N_19718);
nor U21161 (N_21161,N_20603,N_19516);
xnor U21162 (N_21162,N_19828,N_19558);
nor U21163 (N_21163,N_19785,N_20750);
or U21164 (N_21164,N_20337,N_20784);
nor U21165 (N_21165,N_20892,N_20239);
xnor U21166 (N_21166,N_20405,N_19731);
nor U21167 (N_21167,N_20356,N_20481);
or U21168 (N_21168,N_20540,N_19935);
and U21169 (N_21169,N_19543,N_20247);
xor U21170 (N_21170,N_19779,N_20107);
nand U21171 (N_21171,N_19971,N_20224);
or U21172 (N_21172,N_20207,N_20818);
nor U21173 (N_21173,N_20433,N_20307);
or U21174 (N_21174,N_20028,N_20304);
nand U21175 (N_21175,N_19835,N_20303);
nor U21176 (N_21176,N_20306,N_20625);
nand U21177 (N_21177,N_20075,N_20393);
nor U21178 (N_21178,N_19647,N_20067);
nor U21179 (N_21179,N_20230,N_19623);
nor U21180 (N_21180,N_19951,N_20502);
nor U21181 (N_21181,N_20368,N_20987);
nor U21182 (N_21182,N_19539,N_19808);
nand U21183 (N_21183,N_20340,N_20250);
or U21184 (N_21184,N_19821,N_20183);
nor U21185 (N_21185,N_20185,N_20796);
xor U21186 (N_21186,N_19707,N_20458);
nor U21187 (N_21187,N_20501,N_19813);
nand U21188 (N_21188,N_20315,N_20353);
nor U21189 (N_21189,N_20844,N_20837);
xor U21190 (N_21190,N_20366,N_20232);
nor U21191 (N_21191,N_20059,N_20367);
nand U21192 (N_21192,N_19820,N_20791);
nor U21193 (N_21193,N_20493,N_19591);
nand U21194 (N_21194,N_20399,N_19798);
nor U21195 (N_21195,N_20576,N_20712);
nor U21196 (N_21196,N_20632,N_20961);
and U21197 (N_21197,N_20612,N_20647);
and U21198 (N_21198,N_20968,N_20828);
or U21199 (N_21199,N_19873,N_20925);
nand U21200 (N_21200,N_20309,N_19709);
and U21201 (N_21201,N_20601,N_20833);
nand U21202 (N_21202,N_20299,N_19862);
xor U21203 (N_21203,N_19653,N_20113);
xnor U21204 (N_21204,N_19610,N_20707);
xnor U21205 (N_21205,N_20383,N_20851);
xnor U21206 (N_21206,N_20575,N_20947);
xor U21207 (N_21207,N_20194,N_19664);
xor U21208 (N_21208,N_20245,N_19753);
nand U21209 (N_21209,N_20855,N_19529);
and U21210 (N_21210,N_20954,N_20220);
and U21211 (N_21211,N_20847,N_20734);
nand U21212 (N_21212,N_20347,N_19950);
nand U21213 (N_21213,N_19519,N_19553);
and U21214 (N_21214,N_19834,N_20944);
nand U21215 (N_21215,N_19849,N_19925);
and U21216 (N_21216,N_20962,N_19712);
nor U21217 (N_21217,N_20428,N_20600);
xor U21218 (N_21218,N_19982,N_20670);
and U21219 (N_21219,N_20678,N_19583);
or U21220 (N_21220,N_20517,N_20518);
nor U21221 (N_21221,N_19986,N_20209);
xor U21222 (N_21222,N_20074,N_20663);
nor U21223 (N_21223,N_20606,N_20345);
xor U21224 (N_21224,N_19635,N_20121);
nor U21225 (N_21225,N_20885,N_19766);
nand U21226 (N_21226,N_20485,N_20553);
nand U21227 (N_21227,N_20538,N_20441);
or U21228 (N_21228,N_20051,N_19587);
and U21229 (N_21229,N_20893,N_20574);
xnor U21230 (N_21230,N_20083,N_19944);
xor U21231 (N_21231,N_20084,N_20819);
nor U21232 (N_21232,N_20572,N_20635);
and U21233 (N_21233,N_19966,N_19722);
and U21234 (N_21234,N_20443,N_19742);
nand U21235 (N_21235,N_19960,N_19615);
and U21236 (N_21236,N_19975,N_19839);
and U21237 (N_21237,N_20188,N_20229);
or U21238 (N_21238,N_19845,N_20038);
xnor U21239 (N_21239,N_19515,N_20970);
nor U21240 (N_21240,N_19939,N_19810);
and U21241 (N_21241,N_20886,N_19804);
and U21242 (N_21242,N_20744,N_19984);
or U21243 (N_21243,N_20776,N_20835);
nand U21244 (N_21244,N_20888,N_20236);
and U21245 (N_21245,N_20997,N_20911);
and U21246 (N_21246,N_20813,N_20314);
nand U21247 (N_21247,N_20151,N_20008);
or U21248 (N_21248,N_20969,N_20450);
xor U21249 (N_21249,N_20523,N_19990);
and U21250 (N_21250,N_19511,N_20544);
and U21251 (N_21251,N_19687,N_19783);
and U21252 (N_21252,N_20564,N_20821);
xor U21253 (N_21253,N_19673,N_20039);
nor U21254 (N_21254,N_19759,N_20009);
and U21255 (N_21255,N_20966,N_20764);
and U21256 (N_21256,N_20322,N_19884);
nor U21257 (N_21257,N_19887,N_19585);
xnor U21258 (N_21258,N_20834,N_20016);
nand U21259 (N_21259,N_20751,N_20217);
xnor U21260 (N_21260,N_20187,N_20810);
and U21261 (N_21261,N_19793,N_20471);
nor U21262 (N_21262,N_19566,N_20507);
nor U21263 (N_21263,N_20651,N_20466);
and U21264 (N_21264,N_19606,N_20876);
nor U21265 (N_21265,N_20269,N_20222);
nand U21266 (N_21266,N_20254,N_19642);
nand U21267 (N_21267,N_19621,N_20482);
xnor U21268 (N_21268,N_19848,N_20588);
xor U21269 (N_21269,N_20256,N_19961);
nor U21270 (N_21270,N_20104,N_19688);
nand U21271 (N_21271,N_20335,N_19927);
xor U21272 (N_21272,N_19710,N_20741);
xnor U21273 (N_21273,N_20831,N_20896);
or U21274 (N_21274,N_20057,N_20688);
and U21275 (N_21275,N_19605,N_19559);
xnor U21276 (N_21276,N_20827,N_19596);
nor U21277 (N_21277,N_20774,N_20945);
xor U21278 (N_21278,N_19791,N_20934);
and U21279 (N_21279,N_20728,N_19563);
nand U21280 (N_21280,N_20040,N_20097);
or U21281 (N_21281,N_19619,N_20483);
or U21282 (N_21282,N_19851,N_20742);
or U21283 (N_21283,N_20171,N_19686);
or U21284 (N_21284,N_20248,N_20980);
nor U21285 (N_21285,N_20198,N_19865);
and U21286 (N_21286,N_20044,N_19962);
and U21287 (N_21287,N_19842,N_19600);
nand U21288 (N_21288,N_19729,N_20607);
and U21289 (N_21289,N_19928,N_20111);
nand U21290 (N_21290,N_20011,N_20636);
and U21291 (N_21291,N_20598,N_19646);
or U21292 (N_21292,N_20354,N_19748);
and U21293 (N_21293,N_20740,N_20691);
nor U21294 (N_21294,N_20820,N_20677);
or U21295 (N_21295,N_20627,N_19973);
or U21296 (N_21296,N_20723,N_20905);
or U21297 (N_21297,N_20628,N_20917);
or U21298 (N_21298,N_20956,N_20012);
and U21299 (N_21299,N_20845,N_20630);
nand U21300 (N_21300,N_20017,N_19750);
nand U21301 (N_21301,N_19906,N_20141);
xnor U21302 (N_21302,N_19918,N_19948);
xnor U21303 (N_21303,N_19891,N_20762);
xor U21304 (N_21304,N_20077,N_20249);
nand U21305 (N_21305,N_20866,N_20577);
nor U21306 (N_21306,N_20025,N_19876);
nor U21307 (N_21307,N_20509,N_19917);
xnor U21308 (N_21308,N_20593,N_19978);
xnor U21309 (N_21309,N_20887,N_20579);
xnor U21310 (N_21310,N_20150,N_19542);
nand U21311 (N_21311,N_20597,N_20931);
or U21312 (N_21312,N_19936,N_19674);
and U21313 (N_21313,N_20156,N_19974);
nor U21314 (N_21314,N_19683,N_20451);
or U21315 (N_21315,N_20868,N_19924);
or U21316 (N_21316,N_19812,N_19586);
nand U21317 (N_21317,N_20964,N_20312);
xor U21318 (N_21318,N_20115,N_20880);
or U21319 (N_21319,N_20161,N_19518);
xor U21320 (N_21320,N_19562,N_19634);
or U21321 (N_21321,N_20062,N_20656);
or U21322 (N_21322,N_19611,N_19811);
and U21323 (N_21323,N_20913,N_20255);
nand U21324 (N_21324,N_20640,N_19595);
or U21325 (N_21325,N_19776,N_20709);
xor U21326 (N_21326,N_20173,N_20898);
xnor U21327 (N_21327,N_20638,N_20305);
nor U21328 (N_21328,N_20497,N_20070);
xor U21329 (N_21329,N_20280,N_20653);
nand U21330 (N_21330,N_20260,N_20392);
nor U21331 (N_21331,N_20027,N_20720);
and U21332 (N_21332,N_20408,N_19644);
and U21333 (N_21333,N_20109,N_20515);
xnor U21334 (N_21334,N_20955,N_19980);
nand U21335 (N_21335,N_20690,N_20713);
nand U21336 (N_21336,N_20994,N_19863);
and U21337 (N_21337,N_19622,N_20174);
xnor U21338 (N_21338,N_19636,N_20807);
xor U21339 (N_21339,N_20360,N_20089);
xor U21340 (N_21340,N_20278,N_20537);
and U21341 (N_21341,N_19609,N_20702);
xor U21342 (N_21342,N_20013,N_19706);
or U21343 (N_21343,N_20375,N_20463);
nand U21344 (N_21344,N_20971,N_19868);
and U21345 (N_21345,N_20920,N_20046);
xnor U21346 (N_21346,N_19770,N_19616);
nand U21347 (N_21347,N_19965,N_20131);
or U21348 (N_21348,N_19740,N_20129);
nand U21349 (N_21349,N_19538,N_20568);
and U21350 (N_21350,N_19822,N_20952);
nor U21351 (N_21351,N_20730,N_20334);
nor U21352 (N_21352,N_19735,N_20512);
nor U21353 (N_21353,N_19765,N_19916);
nand U21354 (N_21354,N_20234,N_20189);
nor U21355 (N_21355,N_20508,N_20394);
or U21356 (N_21356,N_20374,N_20071);
nor U21357 (N_21357,N_20253,N_19667);
or U21358 (N_21358,N_19905,N_20853);
xnor U21359 (N_21359,N_19567,N_20561);
nand U21360 (N_21360,N_20226,N_19775);
and U21361 (N_21361,N_20883,N_19732);
or U21362 (N_21362,N_20346,N_20711);
nor U21363 (N_21363,N_19565,N_19794);
nand U21364 (N_21364,N_19837,N_20860);
xor U21365 (N_21365,N_20212,N_20144);
nor U21366 (N_21366,N_20655,N_20534);
xor U21367 (N_21367,N_20802,N_20789);
or U21368 (N_21368,N_20725,N_19953);
nor U21369 (N_21369,N_19657,N_20233);
or U21370 (N_21370,N_20719,N_20029);
and U21371 (N_21371,N_20755,N_19651);
xor U21372 (N_21372,N_20316,N_20793);
nor U21373 (N_21373,N_19739,N_19528);
nor U21374 (N_21374,N_20861,N_20870);
nor U21375 (N_21375,N_19522,N_20532);
nand U21376 (N_21376,N_20795,N_20546);
xor U21377 (N_21377,N_19734,N_20313);
nand U21378 (N_21378,N_20164,N_20324);
nand U21379 (N_21379,N_20277,N_19662);
or U21380 (N_21380,N_20864,N_20846);
and U21381 (N_21381,N_20096,N_20959);
and U21382 (N_21382,N_20895,N_19666);
nand U21383 (N_21383,N_20642,N_19681);
and U21384 (N_21384,N_20661,N_20763);
xnor U21385 (N_21385,N_19726,N_20291);
nand U21386 (N_21386,N_20705,N_20993);
and U21387 (N_21387,N_20136,N_20349);
nor U21388 (N_21388,N_20902,N_20524);
nor U21389 (N_21389,N_20182,N_20231);
xnor U21390 (N_21390,N_20130,N_20543);
nor U21391 (N_21391,N_20178,N_19846);
or U21392 (N_21392,N_20756,N_19530);
xor U21393 (N_21393,N_19570,N_20448);
and U21394 (N_21394,N_19630,N_20406);
nand U21395 (N_21395,N_20571,N_20325);
nand U21396 (N_21396,N_19882,N_20122);
or U21397 (N_21397,N_20380,N_19985);
and U21398 (N_21398,N_19721,N_19632);
or U21399 (N_21399,N_19886,N_20881);
nand U21400 (N_21400,N_19665,N_20377);
xnor U21401 (N_21401,N_19893,N_20473);
nor U21402 (N_21402,N_19826,N_20942);
nor U21403 (N_21403,N_19878,N_20566);
or U21404 (N_21404,N_19992,N_20753);
xnor U21405 (N_21405,N_19676,N_19730);
xor U21406 (N_21406,N_20871,N_20991);
and U21407 (N_21407,N_20024,N_19774);
xor U21408 (N_21408,N_19507,N_20484);
and U21409 (N_21409,N_20863,N_20616);
xnor U21410 (N_21410,N_20660,N_20106);
xnor U21411 (N_21411,N_20716,N_20053);
nand U21412 (N_21412,N_19762,N_20862);
and U21413 (N_21413,N_20729,N_20531);
or U21414 (N_21414,N_20637,N_19883);
and U21415 (N_21415,N_20186,N_20290);
nor U21416 (N_21416,N_19818,N_20749);
or U21417 (N_21417,N_19602,N_20557);
nor U21418 (N_21418,N_20223,N_20276);
or U21419 (N_21419,N_20192,N_19780);
and U21420 (N_21420,N_20726,N_19588);
nand U21421 (N_21421,N_20586,N_19699);
nand U21422 (N_21422,N_19885,N_19761);
xnor U21423 (N_21423,N_19955,N_19575);
nor U21424 (N_21424,N_19524,N_20281);
or U21425 (N_21425,N_20801,N_20648);
and U21426 (N_21426,N_19523,N_20257);
nor U21427 (N_21427,N_20320,N_20822);
and U21428 (N_21428,N_20370,N_20043);
nand U21429 (N_21429,N_19535,N_20056);
and U21430 (N_21430,N_19675,N_19795);
xnor U21431 (N_21431,N_20514,N_20548);
or U21432 (N_21432,N_20401,N_19789);
nand U21433 (N_21433,N_19624,N_19901);
xnor U21434 (N_21434,N_20592,N_19781);
or U21435 (N_21435,N_20694,N_19749);
nand U21436 (N_21436,N_20963,N_20118);
and U21437 (N_21437,N_20423,N_19670);
nor U21438 (N_21438,N_20879,N_20396);
or U21439 (N_21439,N_20782,N_20721);
nand U21440 (N_21440,N_19858,N_20633);
or U21441 (N_21441,N_20919,N_19696);
nand U21442 (N_21442,N_20935,N_20545);
or U21443 (N_21443,N_19713,N_20369);
and U21444 (N_21444,N_20434,N_19997);
nor U21445 (N_21445,N_20328,N_20960);
nand U21446 (N_21446,N_20995,N_20843);
and U21447 (N_21447,N_20609,N_19717);
xor U21448 (N_21448,N_19970,N_20621);
and U21449 (N_21449,N_20733,N_20687);
xor U21450 (N_21450,N_20440,N_20022);
nor U21451 (N_21451,N_19708,N_20268);
nand U21452 (N_21452,N_20142,N_20133);
xnor U21453 (N_21453,N_19637,N_20457);
xor U21454 (N_21454,N_20455,N_20695);
or U21455 (N_21455,N_19626,N_20416);
or U21456 (N_21456,N_19723,N_19571);
or U21457 (N_21457,N_20175,N_20965);
nand U21458 (N_21458,N_20839,N_20317);
nor U21459 (N_21459,N_20108,N_20570);
or U21460 (N_21460,N_19823,N_20549);
nor U21461 (N_21461,N_19513,N_20806);
nand U21462 (N_21462,N_20500,N_20589);
and U21463 (N_21463,N_20875,N_19648);
xnor U21464 (N_21464,N_20032,N_20388);
and U21465 (N_21465,N_20927,N_19716);
or U21466 (N_21466,N_20780,N_19520);
nand U21467 (N_21467,N_20526,N_20041);
nor U21468 (N_21468,N_19584,N_20700);
xnor U21469 (N_21469,N_20298,N_20273);
or U21470 (N_21470,N_20387,N_19701);
and U21471 (N_21471,N_20613,N_20696);
xor U21472 (N_21472,N_19733,N_19758);
nor U21473 (N_21473,N_19704,N_20235);
nand U21474 (N_21474,N_20149,N_19700);
and U21475 (N_21475,N_19556,N_20536);
or U21476 (N_21476,N_19772,N_20732);
xnor U21477 (N_21477,N_19931,N_20923);
nor U21478 (N_21478,N_20897,N_20114);
and U21479 (N_21479,N_20785,N_19947);
or U21480 (N_21480,N_20599,N_20456);
nor U21481 (N_21481,N_19618,N_20221);
xor U21482 (N_21482,N_20147,N_20157);
or U21483 (N_21483,N_20362,N_19888);
or U21484 (N_21484,N_19968,N_20529);
or U21485 (N_21485,N_20659,N_20413);
and U21486 (N_21486,N_20626,N_20901);
and U21487 (N_21487,N_20771,N_19641);
or U21488 (N_21488,N_19983,N_20311);
or U21489 (N_21489,N_20527,N_20513);
xor U21490 (N_21490,N_20091,N_20550);
and U21491 (N_21491,N_19958,N_20427);
or U21492 (N_21492,N_19502,N_19881);
nor U21493 (N_21493,N_20120,N_20714);
and U21494 (N_21494,N_19728,N_20992);
or U21495 (N_21495,N_20743,N_19767);
nand U21496 (N_21496,N_20323,N_19714);
or U21497 (N_21497,N_19840,N_20094);
xnor U21498 (N_21498,N_19752,N_20019);
or U21499 (N_21499,N_20594,N_20722);
nor U21500 (N_21500,N_20918,N_20140);
xnor U21501 (N_21501,N_20263,N_19573);
and U21502 (N_21502,N_19607,N_19852);
or U21503 (N_21503,N_20251,N_20737);
and U21504 (N_21504,N_20431,N_19680);
nor U21505 (N_21505,N_19746,N_20495);
and U21506 (N_21506,N_19908,N_20643);
nor U21507 (N_21507,N_19702,N_20126);
nand U21508 (N_21508,N_20146,N_20176);
xor U21509 (N_21509,N_20715,N_20953);
xnor U21510 (N_21510,N_20629,N_20302);
and U21511 (N_21511,N_19904,N_19697);
nand U21512 (N_21512,N_19669,N_19934);
nand U21513 (N_21513,N_19806,N_19786);
or U21514 (N_21514,N_20364,N_20058);
nand U21515 (N_21515,N_20735,N_20272);
or U21516 (N_21516,N_20101,N_20474);
and U21517 (N_21517,N_20219,N_20139);
or U21518 (N_21518,N_19612,N_19579);
xor U21519 (N_21519,N_19509,N_19536);
nand U21520 (N_21520,N_20338,N_20922);
or U21521 (N_21521,N_19568,N_20389);
and U21522 (N_21522,N_20018,N_20202);
nor U21523 (N_21523,N_20631,N_19690);
nand U21524 (N_21524,N_19979,N_19582);
xnor U21525 (N_21525,N_20453,N_19870);
and U21526 (N_21526,N_20800,N_20479);
and U21527 (N_21527,N_20867,N_20098);
nor U21528 (N_21528,N_20376,N_20099);
or U21529 (N_21529,N_20179,N_19545);
and U21530 (N_21530,N_20429,N_20666);
and U21531 (N_21531,N_20758,N_20068);
nand U21532 (N_21532,N_19598,N_20425);
nor U21533 (N_21533,N_19773,N_20415);
nor U21534 (N_21534,N_20658,N_19949);
nor U21535 (N_21535,N_19537,N_19991);
and U21536 (N_21536,N_20926,N_20218);
nor U21537 (N_21537,N_20525,N_20909);
nor U21538 (N_21538,N_20352,N_20587);
xnor U21539 (N_21539,N_20262,N_20007);
and U21540 (N_21540,N_20050,N_20731);
xnor U21541 (N_21541,N_20002,N_20988);
or U21542 (N_21542,N_19514,N_20766);
or U21543 (N_21543,N_20087,N_20560);
nand U21544 (N_21544,N_20565,N_19920);
or U21545 (N_21545,N_19954,N_20125);
xor U21546 (N_21546,N_20578,N_19603);
and U21547 (N_21547,N_20386,N_20410);
nor U21548 (N_21548,N_19843,N_19555);
nor U21549 (N_21549,N_20668,N_20010);
xor U21550 (N_21550,N_20914,N_20869);
or U21551 (N_21551,N_20177,N_19903);
nor U21552 (N_21552,N_20216,N_19832);
nor U21553 (N_21553,N_19957,N_20765);
nand U21554 (N_21554,N_20884,N_19649);
or U21555 (N_21555,N_20076,N_20644);
and U21556 (N_21556,N_20210,N_19643);
or U21557 (N_21557,N_19768,N_20259);
nand U21558 (N_21558,N_20817,N_19922);
xor U21559 (N_21559,N_20584,N_20409);
nand U21560 (N_21560,N_20135,N_20339);
or U21561 (N_21561,N_19678,N_20155);
xnor U21562 (N_21562,N_19532,N_20936);
and U21563 (N_21563,N_19574,N_19802);
or U21564 (N_21564,N_20446,N_20805);
xnor U21565 (N_21565,N_20614,N_19527);
nand U21566 (N_21566,N_20026,N_20447);
and U21567 (N_21567,N_20402,N_20788);
and U21568 (N_21568,N_19938,N_19517);
and U21569 (N_21569,N_20541,N_20499);
nor U21570 (N_21570,N_20344,N_20361);
nor U21571 (N_21571,N_20422,N_20319);
or U21572 (N_21572,N_20138,N_20333);
nand U21573 (N_21573,N_20243,N_19580);
xnor U21574 (N_21574,N_19877,N_20974);
or U21575 (N_21575,N_20005,N_20282);
or U21576 (N_21576,N_20491,N_20667);
and U21577 (N_21577,N_20397,N_19613);
nor U21578 (N_21578,N_20848,N_19998);
nor U21579 (N_21579,N_20073,N_19747);
or U21580 (N_21580,N_19778,N_20738);
and U21581 (N_21581,N_20824,N_20445);
nor U21582 (N_21582,N_20984,N_19969);
and U21583 (N_21583,N_20214,N_20227);
nand U21584 (N_21584,N_19787,N_19995);
nor U21585 (N_21585,N_20132,N_19736);
nor U21586 (N_21586,N_20899,N_20103);
nor U21587 (N_21587,N_20555,N_20498);
and U21588 (N_21588,N_19859,N_19503);
xor U21589 (N_21589,N_20929,N_19964);
nor U21590 (N_21590,N_19940,N_20063);
xnor U21591 (N_21591,N_20830,N_20490);
nor U21592 (N_21592,N_20289,N_19900);
or U21593 (N_21593,N_20878,N_19541);
xor U21594 (N_21594,N_20036,N_20812);
or U21595 (N_21595,N_20211,N_19771);
or U21596 (N_21596,N_20400,N_20849);
and U21597 (N_21597,N_20355,N_20398);
and U21598 (N_21598,N_19912,N_20799);
nor U21599 (N_21599,N_20378,N_19745);
nor U21600 (N_21600,N_20581,N_20404);
xnor U21601 (N_21601,N_20014,N_20790);
nor U21602 (N_21602,N_19941,N_19869);
and U21603 (N_21603,N_20693,N_20468);
nor U21604 (N_21604,N_19548,N_20948);
and U21605 (N_21605,N_20928,N_19577);
nor U21606 (N_21606,N_20204,N_20363);
xnor U21607 (N_21607,N_20033,N_19919);
and U21608 (N_21608,N_20112,N_20989);
xor U21609 (N_21609,N_20436,N_19572);
xor U21610 (N_21610,N_19754,N_20137);
nand U21611 (N_21611,N_20894,N_19996);
nand U21612 (N_21612,N_20889,N_20288);
xor U21613 (N_21613,N_20798,N_19724);
nor U21614 (N_21614,N_20983,N_19836);
nand U21615 (N_21615,N_19629,N_20910);
nand U21616 (N_21616,N_20384,N_20804);
xor U21617 (N_21617,N_20000,N_20706);
nand U21618 (N_21618,N_20669,N_19933);
nor U21619 (N_21619,N_20300,N_20591);
nand U21620 (N_21620,N_20035,N_19815);
and U21621 (N_21621,N_20620,N_20117);
or U21622 (N_21622,N_20391,N_19909);
and U21623 (N_21623,N_20452,N_20090);
nand U21624 (N_21624,N_20859,N_20294);
and U21625 (N_21625,N_20078,N_20052);
or U21626 (N_21626,N_19534,N_19557);
xnor U21627 (N_21627,N_20285,N_20318);
nor U21628 (N_21628,N_19540,N_19533);
xnor U21629 (N_21629,N_20437,N_20292);
xnor U21630 (N_21630,N_20717,N_19526);
xnor U21631 (N_21631,N_19896,N_19989);
and U21632 (N_21632,N_20912,N_20205);
nor U21633 (N_21633,N_19601,N_20826);
or U21634 (N_21634,N_20086,N_20365);
nor U21635 (N_21635,N_20414,N_19656);
xor U21636 (N_21636,N_19689,N_20904);
nor U21637 (N_21637,N_20708,N_19597);
xor U21638 (N_21638,N_20907,N_20724);
or U21639 (N_21639,N_20351,N_20516);
xor U21640 (N_21640,N_20675,N_20521);
or U21641 (N_21641,N_20710,N_19999);
xnor U21642 (N_21642,N_20815,N_20419);
or U21643 (N_21643,N_20563,N_20903);
nand U21644 (N_21644,N_20154,N_19929);
and U21645 (N_21645,N_19910,N_19592);
nor U21646 (N_21646,N_20978,N_20238);
nor U21647 (N_21647,N_20748,N_20622);
and U21648 (N_21648,N_19807,N_20166);
nand U21649 (N_21649,N_20034,N_20143);
xnor U21650 (N_21650,N_19890,N_19694);
nand U21651 (N_21651,N_19682,N_20985);
xnor U21652 (N_21652,N_20760,N_20395);
nand U21653 (N_21653,N_20042,N_20048);
nor U21654 (N_21654,N_20933,N_19652);
xnor U21655 (N_21655,N_20761,N_20080);
or U21656 (N_21656,N_20697,N_20287);
nand U21657 (N_21657,N_20856,N_20836);
nor U21658 (N_21658,N_19638,N_19639);
nand U21659 (N_21659,N_20444,N_19914);
or U21660 (N_21660,N_20939,N_19512);
or U21661 (N_21661,N_20486,N_20874);
nor U21662 (N_21662,N_20873,N_19751);
or U21663 (N_21663,N_20703,N_19867);
xor U21664 (N_21664,N_19790,N_20770);
nand U21665 (N_21665,N_20797,N_19911);
xnor U21666 (N_21666,N_19857,N_20773);
nor U21667 (N_21667,N_20492,N_20900);
and U21668 (N_21668,N_20682,N_20407);
or U21669 (N_21669,N_19956,N_19875);
and U21670 (N_21670,N_20559,N_20195);
or U21671 (N_21671,N_19963,N_20496);
xor U21672 (N_21672,N_19907,N_20201);
or U21673 (N_21673,N_20504,N_20701);
nor U21674 (N_21674,N_20739,N_19854);
xor U21675 (N_21675,N_19628,N_19505);
and U21676 (N_21676,N_20811,N_19829);
xnor U21677 (N_21677,N_20487,N_20673);
nor U21678 (N_21678,N_20692,N_20342);
or U21679 (N_21679,N_19894,N_20539);
and U21680 (N_21680,N_19659,N_19554);
nand U21681 (N_21681,N_20390,N_19921);
nor U21682 (N_21682,N_20494,N_20552);
or U21683 (N_21683,N_19560,N_20664);
xor U21684 (N_21684,N_19561,N_19788);
nand U21685 (N_21685,N_20752,N_20746);
and U21686 (N_21686,N_20522,N_20840);
and U21687 (N_21687,N_20530,N_20683);
and U21688 (N_21688,N_20489,N_20478);
nand U21689 (N_21689,N_19952,N_20646);
xnor U21690 (N_21690,N_20941,N_19799);
or U21691 (N_21691,N_20689,N_20148);
and U21692 (N_21692,N_20624,N_19684);
and U21693 (N_21693,N_20184,N_19913);
xnor U21694 (N_21694,N_20343,N_20769);
nand U21695 (N_21695,N_19803,N_19889);
and U21696 (N_21696,N_20460,N_20506);
or U21697 (N_21697,N_20412,N_20297);
xnor U21698 (N_21698,N_20736,N_20982);
xor U21699 (N_21699,N_20556,N_20558);
nor U21700 (N_21700,N_20569,N_19967);
xor U21701 (N_21701,N_20999,N_19981);
or U21702 (N_21702,N_20242,N_20967);
and U21703 (N_21703,N_20464,N_20775);
xnor U21704 (N_21704,N_20841,N_19672);
xor U21705 (N_21705,N_20865,N_20190);
xnor U21706 (N_21706,N_20279,N_20681);
nor U21707 (N_21707,N_20246,N_20093);
nor U21708 (N_21708,N_19946,N_20477);
nor U21709 (N_21709,N_20908,N_20654);
and U21710 (N_21710,N_20665,N_20858);
nor U21711 (N_21711,N_20295,N_20480);
or U21712 (N_21712,N_19589,N_19800);
or U21713 (N_21713,N_20162,N_20001);
nand U21714 (N_21714,N_20284,N_20857);
nor U21715 (N_21715,N_19737,N_19898);
and U21716 (N_21716,N_20264,N_20615);
xor U21717 (N_21717,N_20308,N_20200);
xnor U21718 (N_21718,N_20403,N_20430);
and U21719 (N_21719,N_20872,N_20467);
xor U21720 (N_21720,N_19831,N_20533);
or U21721 (N_21721,N_20671,N_20270);
or U21722 (N_21722,N_20832,N_20267);
and U21723 (N_21723,N_20699,N_20604);
and U21724 (N_21724,N_19844,N_20258);
or U21725 (N_21725,N_20286,N_19850);
nor U21726 (N_21726,N_20674,N_20838);
and U21727 (N_21727,N_19923,N_20958);
nand U21728 (N_21728,N_20535,N_20977);
or U21729 (N_21729,N_20341,N_20079);
xor U21730 (N_21730,N_19926,N_19521);
xnor U21731 (N_21731,N_20698,N_19711);
and U21732 (N_21732,N_20652,N_19879);
nor U21733 (N_21733,N_20704,N_19569);
or U21734 (N_21734,N_20852,N_19594);
or U21735 (N_21735,N_20049,N_20331);
and U21736 (N_21736,N_19830,N_20921);
xor U21737 (N_21737,N_19627,N_20990);
xor U21738 (N_21738,N_20816,N_19544);
nor U21739 (N_21739,N_20882,N_20645);
nand U21740 (N_21740,N_20602,N_19756);
xnor U21741 (N_21741,N_19872,N_20476);
nor U21742 (N_21742,N_19782,N_19943);
and U21743 (N_21743,N_20979,N_20159);
nand U21744 (N_21744,N_20938,N_20596);
or U21745 (N_21745,N_20825,N_20718);
xor U21746 (N_21746,N_19550,N_20567);
xor U21747 (N_21747,N_19760,N_20081);
or U21748 (N_21748,N_20054,N_20573);
nand U21749 (N_21749,N_19880,N_20061);
or U21750 (N_21750,N_20991,N_19616);
or U21751 (N_21751,N_20611,N_20937);
xor U21752 (N_21752,N_20336,N_19564);
xnor U21753 (N_21753,N_19639,N_19865);
or U21754 (N_21754,N_19721,N_20651);
nor U21755 (N_21755,N_20869,N_19592);
or U21756 (N_21756,N_20921,N_19825);
nor U21757 (N_21757,N_19923,N_20795);
nand U21758 (N_21758,N_20421,N_20749);
nand U21759 (N_21759,N_20064,N_20611);
xnor U21760 (N_21760,N_20583,N_19645);
and U21761 (N_21761,N_20277,N_20187);
and U21762 (N_21762,N_20030,N_20129);
xor U21763 (N_21763,N_19834,N_20067);
nand U21764 (N_21764,N_20545,N_20383);
nor U21765 (N_21765,N_19793,N_20510);
xor U21766 (N_21766,N_20255,N_20095);
or U21767 (N_21767,N_20242,N_20396);
and U21768 (N_21768,N_20521,N_20827);
nor U21769 (N_21769,N_20559,N_20865);
nor U21770 (N_21770,N_20013,N_20206);
xnor U21771 (N_21771,N_20986,N_19500);
nand U21772 (N_21772,N_20333,N_20672);
nand U21773 (N_21773,N_20358,N_20370);
or U21774 (N_21774,N_20506,N_20486);
nand U21775 (N_21775,N_20170,N_20847);
nor U21776 (N_21776,N_20897,N_19879);
and U21777 (N_21777,N_19722,N_20416);
and U21778 (N_21778,N_20604,N_19735);
nor U21779 (N_21779,N_19958,N_19914);
and U21780 (N_21780,N_20024,N_19911);
nand U21781 (N_21781,N_20233,N_20841);
nand U21782 (N_21782,N_19668,N_19748);
xnor U21783 (N_21783,N_19866,N_20105);
nor U21784 (N_21784,N_20257,N_20352);
and U21785 (N_21785,N_19925,N_19768);
nand U21786 (N_21786,N_19676,N_20548);
xnor U21787 (N_21787,N_20928,N_20804);
nor U21788 (N_21788,N_19930,N_20854);
xnor U21789 (N_21789,N_20569,N_20224);
xor U21790 (N_21790,N_20309,N_19763);
nor U21791 (N_21791,N_20297,N_20133);
xor U21792 (N_21792,N_20414,N_20265);
nand U21793 (N_21793,N_19901,N_19655);
nand U21794 (N_21794,N_19508,N_20996);
nand U21795 (N_21795,N_20015,N_20260);
and U21796 (N_21796,N_20353,N_19580);
or U21797 (N_21797,N_20766,N_20303);
or U21798 (N_21798,N_20715,N_20650);
xor U21799 (N_21799,N_20237,N_20570);
xor U21800 (N_21800,N_20564,N_19938);
nor U21801 (N_21801,N_19697,N_20497);
and U21802 (N_21802,N_20438,N_20658);
nand U21803 (N_21803,N_20576,N_20446);
xnor U21804 (N_21804,N_20179,N_19592);
and U21805 (N_21805,N_19660,N_20198);
nand U21806 (N_21806,N_20693,N_19537);
or U21807 (N_21807,N_20503,N_19884);
nor U21808 (N_21808,N_20622,N_20273);
or U21809 (N_21809,N_20589,N_20792);
xor U21810 (N_21810,N_20679,N_20768);
nor U21811 (N_21811,N_19771,N_20136);
nand U21812 (N_21812,N_20889,N_19596);
nand U21813 (N_21813,N_20829,N_19623);
nor U21814 (N_21814,N_20730,N_19872);
or U21815 (N_21815,N_20609,N_20503);
or U21816 (N_21816,N_19724,N_20792);
xor U21817 (N_21817,N_19903,N_19749);
xor U21818 (N_21818,N_20992,N_19720);
or U21819 (N_21819,N_19933,N_20261);
nor U21820 (N_21820,N_20788,N_20891);
nor U21821 (N_21821,N_20903,N_20353);
nor U21822 (N_21822,N_20892,N_20098);
nor U21823 (N_21823,N_20592,N_20779);
and U21824 (N_21824,N_20958,N_20680);
nand U21825 (N_21825,N_20523,N_20564);
nand U21826 (N_21826,N_20641,N_19544);
nor U21827 (N_21827,N_20233,N_20124);
nand U21828 (N_21828,N_20557,N_20969);
nor U21829 (N_21829,N_20828,N_20911);
nand U21830 (N_21830,N_19553,N_20528);
nand U21831 (N_21831,N_20677,N_20667);
and U21832 (N_21832,N_20708,N_19831);
nor U21833 (N_21833,N_20018,N_20955);
nand U21834 (N_21834,N_20085,N_20945);
nand U21835 (N_21835,N_19568,N_19632);
nor U21836 (N_21836,N_19812,N_20492);
nand U21837 (N_21837,N_20664,N_20338);
or U21838 (N_21838,N_19657,N_20909);
nor U21839 (N_21839,N_20475,N_19533);
and U21840 (N_21840,N_20970,N_20839);
xor U21841 (N_21841,N_20262,N_19730);
or U21842 (N_21842,N_20357,N_19610);
and U21843 (N_21843,N_20835,N_19732);
and U21844 (N_21844,N_20222,N_20823);
or U21845 (N_21845,N_19597,N_20713);
xnor U21846 (N_21846,N_20385,N_20767);
nor U21847 (N_21847,N_20858,N_19885);
nand U21848 (N_21848,N_19630,N_20641);
xor U21849 (N_21849,N_20983,N_20136);
or U21850 (N_21850,N_20710,N_20940);
xnor U21851 (N_21851,N_20316,N_19729);
xor U21852 (N_21852,N_20232,N_20474);
xnor U21853 (N_21853,N_19846,N_20874);
nand U21854 (N_21854,N_19911,N_20502);
nand U21855 (N_21855,N_19570,N_19608);
nand U21856 (N_21856,N_20494,N_19565);
or U21857 (N_21857,N_20971,N_19510);
nor U21858 (N_21858,N_20173,N_20946);
or U21859 (N_21859,N_20758,N_19722);
and U21860 (N_21860,N_20616,N_20093);
and U21861 (N_21861,N_20425,N_19845);
nor U21862 (N_21862,N_20088,N_20439);
nand U21863 (N_21863,N_19992,N_20765);
or U21864 (N_21864,N_20456,N_19859);
nand U21865 (N_21865,N_19716,N_20746);
nand U21866 (N_21866,N_19924,N_20973);
or U21867 (N_21867,N_20470,N_20060);
nor U21868 (N_21868,N_20974,N_19827);
xor U21869 (N_21869,N_19584,N_20315);
or U21870 (N_21870,N_20522,N_20520);
nor U21871 (N_21871,N_20190,N_19955);
or U21872 (N_21872,N_20218,N_20757);
nor U21873 (N_21873,N_20714,N_20308);
or U21874 (N_21874,N_20458,N_20334);
or U21875 (N_21875,N_20406,N_19505);
and U21876 (N_21876,N_19634,N_20723);
nand U21877 (N_21877,N_20671,N_19635);
nand U21878 (N_21878,N_20210,N_20169);
nand U21879 (N_21879,N_19587,N_19743);
or U21880 (N_21880,N_19776,N_20392);
nor U21881 (N_21881,N_20929,N_19751);
nand U21882 (N_21882,N_19669,N_19579);
or U21883 (N_21883,N_19804,N_20096);
nand U21884 (N_21884,N_20579,N_19725);
or U21885 (N_21885,N_19985,N_19740);
nand U21886 (N_21886,N_20282,N_19946);
nand U21887 (N_21887,N_20157,N_19995);
and U21888 (N_21888,N_20292,N_19802);
nand U21889 (N_21889,N_20024,N_19964);
nor U21890 (N_21890,N_20433,N_20634);
and U21891 (N_21891,N_19550,N_20974);
and U21892 (N_21892,N_19655,N_19796);
or U21893 (N_21893,N_20576,N_20987);
nor U21894 (N_21894,N_20259,N_20417);
or U21895 (N_21895,N_20193,N_19796);
nor U21896 (N_21896,N_20370,N_19652);
and U21897 (N_21897,N_20413,N_20591);
xor U21898 (N_21898,N_20408,N_20065);
xnor U21899 (N_21899,N_20379,N_19904);
nand U21900 (N_21900,N_20733,N_19792);
xnor U21901 (N_21901,N_20528,N_20182);
nand U21902 (N_21902,N_20914,N_19553);
nor U21903 (N_21903,N_20120,N_20821);
or U21904 (N_21904,N_20136,N_20340);
nand U21905 (N_21905,N_20317,N_19500);
nor U21906 (N_21906,N_20898,N_20096);
nor U21907 (N_21907,N_19623,N_19750);
nand U21908 (N_21908,N_19736,N_20230);
nor U21909 (N_21909,N_19629,N_19842);
nand U21910 (N_21910,N_20033,N_19695);
or U21911 (N_21911,N_20892,N_20589);
and U21912 (N_21912,N_20377,N_20228);
or U21913 (N_21913,N_20107,N_20785);
and U21914 (N_21914,N_20945,N_20663);
xnor U21915 (N_21915,N_19594,N_20035);
nor U21916 (N_21916,N_20544,N_20242);
nor U21917 (N_21917,N_20383,N_20816);
or U21918 (N_21918,N_20789,N_20858);
nor U21919 (N_21919,N_20826,N_20937);
and U21920 (N_21920,N_20297,N_20719);
nor U21921 (N_21921,N_20718,N_20666);
nor U21922 (N_21922,N_20239,N_19545);
and U21923 (N_21923,N_19506,N_20431);
and U21924 (N_21924,N_20145,N_20379);
and U21925 (N_21925,N_20809,N_20903);
nor U21926 (N_21926,N_19886,N_20193);
and U21927 (N_21927,N_19859,N_20286);
xnor U21928 (N_21928,N_19779,N_19802);
nor U21929 (N_21929,N_20187,N_20252);
xnor U21930 (N_21930,N_20171,N_20781);
nor U21931 (N_21931,N_20045,N_20208);
or U21932 (N_21932,N_20913,N_20661);
xor U21933 (N_21933,N_19850,N_20813);
nand U21934 (N_21934,N_20439,N_20043);
and U21935 (N_21935,N_20160,N_19628);
or U21936 (N_21936,N_20674,N_20048);
nand U21937 (N_21937,N_19852,N_19906);
nand U21938 (N_21938,N_19983,N_20714);
and U21939 (N_21939,N_20271,N_19922);
nor U21940 (N_21940,N_20300,N_20481);
nand U21941 (N_21941,N_20464,N_19678);
nand U21942 (N_21942,N_20098,N_19729);
or U21943 (N_21943,N_20504,N_20412);
nand U21944 (N_21944,N_20980,N_20047);
xor U21945 (N_21945,N_20503,N_20946);
or U21946 (N_21946,N_19791,N_20123);
and U21947 (N_21947,N_19825,N_20020);
nor U21948 (N_21948,N_20976,N_19595);
xor U21949 (N_21949,N_20019,N_20078);
nor U21950 (N_21950,N_19748,N_20922);
xor U21951 (N_21951,N_20332,N_19507);
nor U21952 (N_21952,N_19643,N_19888);
or U21953 (N_21953,N_20715,N_19850);
nor U21954 (N_21954,N_19973,N_19753);
and U21955 (N_21955,N_20263,N_20449);
nand U21956 (N_21956,N_20283,N_20935);
nand U21957 (N_21957,N_19755,N_19836);
and U21958 (N_21958,N_19726,N_20305);
nor U21959 (N_21959,N_19972,N_19693);
or U21960 (N_21960,N_20132,N_20779);
nor U21961 (N_21961,N_19728,N_19750);
nor U21962 (N_21962,N_19976,N_19542);
nor U21963 (N_21963,N_20801,N_20905);
nand U21964 (N_21964,N_20860,N_20150);
nand U21965 (N_21965,N_20396,N_20496);
and U21966 (N_21966,N_20285,N_20995);
or U21967 (N_21967,N_20810,N_19913);
xor U21968 (N_21968,N_20461,N_20555);
nor U21969 (N_21969,N_20970,N_20930);
and U21970 (N_21970,N_19999,N_20579);
and U21971 (N_21971,N_19845,N_20517);
or U21972 (N_21972,N_20545,N_19571);
nor U21973 (N_21973,N_20908,N_19813);
or U21974 (N_21974,N_20178,N_20452);
or U21975 (N_21975,N_20407,N_19982);
and U21976 (N_21976,N_19734,N_20419);
nor U21977 (N_21977,N_20823,N_20068);
xor U21978 (N_21978,N_19906,N_20800);
nand U21979 (N_21979,N_19600,N_20779);
xnor U21980 (N_21980,N_20160,N_20590);
nand U21981 (N_21981,N_20247,N_19779);
nor U21982 (N_21982,N_19742,N_20252);
nor U21983 (N_21983,N_19898,N_20189);
nor U21984 (N_21984,N_19879,N_20421);
xor U21985 (N_21985,N_19993,N_20095);
nor U21986 (N_21986,N_20055,N_19669);
nand U21987 (N_21987,N_20965,N_19651);
or U21988 (N_21988,N_19788,N_20892);
xor U21989 (N_21989,N_20490,N_20232);
nor U21990 (N_21990,N_20208,N_20719);
or U21991 (N_21991,N_20412,N_20714);
nor U21992 (N_21992,N_19556,N_20560);
xor U21993 (N_21993,N_20505,N_19637);
nor U21994 (N_21994,N_20466,N_20073);
nand U21995 (N_21995,N_20802,N_19850);
nand U21996 (N_21996,N_20045,N_19766);
nand U21997 (N_21997,N_20319,N_20207);
nand U21998 (N_21998,N_20987,N_20152);
or U21999 (N_21999,N_19701,N_20692);
nand U22000 (N_22000,N_20034,N_20339);
xor U22001 (N_22001,N_20742,N_19647);
xor U22002 (N_22002,N_20710,N_20671);
and U22003 (N_22003,N_19699,N_20435);
and U22004 (N_22004,N_20511,N_20167);
or U22005 (N_22005,N_20634,N_20466);
and U22006 (N_22006,N_20627,N_20339);
nand U22007 (N_22007,N_20340,N_20130);
or U22008 (N_22008,N_20644,N_19807);
and U22009 (N_22009,N_20979,N_20029);
and U22010 (N_22010,N_19555,N_20561);
nor U22011 (N_22011,N_19761,N_19577);
nand U22012 (N_22012,N_20128,N_20918);
and U22013 (N_22013,N_20538,N_19755);
nand U22014 (N_22014,N_19575,N_20004);
nand U22015 (N_22015,N_19885,N_19813);
nand U22016 (N_22016,N_19669,N_19596);
nor U22017 (N_22017,N_20521,N_20559);
nor U22018 (N_22018,N_19556,N_20411);
and U22019 (N_22019,N_20470,N_20946);
xor U22020 (N_22020,N_20572,N_20996);
nor U22021 (N_22021,N_19972,N_20139);
nor U22022 (N_22022,N_19752,N_20756);
nor U22023 (N_22023,N_20677,N_20334);
nor U22024 (N_22024,N_20767,N_20261);
nor U22025 (N_22025,N_20779,N_20492);
nand U22026 (N_22026,N_19539,N_20607);
xor U22027 (N_22027,N_20383,N_20427);
xor U22028 (N_22028,N_20274,N_19771);
and U22029 (N_22029,N_20196,N_19533);
or U22030 (N_22030,N_20321,N_19958);
or U22031 (N_22031,N_19543,N_20765);
nor U22032 (N_22032,N_19824,N_20192);
nand U22033 (N_22033,N_20668,N_20480);
nor U22034 (N_22034,N_19571,N_19532);
nor U22035 (N_22035,N_20145,N_20821);
nor U22036 (N_22036,N_19829,N_19576);
nor U22037 (N_22037,N_20818,N_19836);
or U22038 (N_22038,N_20666,N_20694);
and U22039 (N_22039,N_20054,N_20754);
or U22040 (N_22040,N_20946,N_20413);
or U22041 (N_22041,N_20269,N_20348);
nand U22042 (N_22042,N_19519,N_20934);
nand U22043 (N_22043,N_19574,N_20164);
nor U22044 (N_22044,N_19781,N_19696);
nor U22045 (N_22045,N_20917,N_20089);
nor U22046 (N_22046,N_19516,N_20463);
or U22047 (N_22047,N_20326,N_20581);
nand U22048 (N_22048,N_20033,N_20325);
and U22049 (N_22049,N_20241,N_20426);
and U22050 (N_22050,N_20709,N_19874);
nand U22051 (N_22051,N_20638,N_20525);
or U22052 (N_22052,N_20332,N_20141);
or U22053 (N_22053,N_20980,N_20172);
and U22054 (N_22054,N_20632,N_20834);
xnor U22055 (N_22055,N_19538,N_20203);
and U22056 (N_22056,N_20770,N_19718);
nand U22057 (N_22057,N_20344,N_19950);
or U22058 (N_22058,N_20768,N_20137);
and U22059 (N_22059,N_20564,N_20092);
nand U22060 (N_22060,N_19960,N_19766);
xor U22061 (N_22061,N_20206,N_20779);
or U22062 (N_22062,N_20932,N_19612);
nor U22063 (N_22063,N_20674,N_19867);
and U22064 (N_22064,N_19530,N_20110);
nand U22065 (N_22065,N_20776,N_19661);
nor U22066 (N_22066,N_20106,N_19763);
and U22067 (N_22067,N_19771,N_20754);
or U22068 (N_22068,N_20755,N_20106);
or U22069 (N_22069,N_20312,N_20283);
and U22070 (N_22070,N_20640,N_20418);
nor U22071 (N_22071,N_20351,N_19899);
xnor U22072 (N_22072,N_19590,N_19579);
nand U22073 (N_22073,N_20668,N_20700);
xor U22074 (N_22074,N_20756,N_20153);
nand U22075 (N_22075,N_20372,N_19962);
xor U22076 (N_22076,N_20460,N_20331);
nand U22077 (N_22077,N_20745,N_20839);
and U22078 (N_22078,N_19550,N_20435);
nor U22079 (N_22079,N_19566,N_20277);
nand U22080 (N_22080,N_19611,N_20820);
xnor U22081 (N_22081,N_20549,N_19608);
nand U22082 (N_22082,N_19848,N_20579);
xnor U22083 (N_22083,N_20755,N_20561);
nand U22084 (N_22084,N_20252,N_20462);
nand U22085 (N_22085,N_20452,N_20607);
nor U22086 (N_22086,N_19929,N_20735);
or U22087 (N_22087,N_20219,N_20483);
xor U22088 (N_22088,N_19835,N_20044);
and U22089 (N_22089,N_20681,N_20820);
nor U22090 (N_22090,N_19525,N_20268);
and U22091 (N_22091,N_19611,N_20921);
xor U22092 (N_22092,N_19949,N_19968);
and U22093 (N_22093,N_20094,N_20443);
xnor U22094 (N_22094,N_19715,N_19975);
nor U22095 (N_22095,N_20450,N_19589);
and U22096 (N_22096,N_20925,N_20125);
and U22097 (N_22097,N_20845,N_20962);
and U22098 (N_22098,N_20420,N_20203);
nand U22099 (N_22099,N_20005,N_19694);
nand U22100 (N_22100,N_19838,N_19950);
nor U22101 (N_22101,N_20892,N_20148);
and U22102 (N_22102,N_20881,N_19859);
xnor U22103 (N_22103,N_20578,N_20541);
and U22104 (N_22104,N_20073,N_20557);
or U22105 (N_22105,N_19662,N_19915);
nor U22106 (N_22106,N_19948,N_19987);
or U22107 (N_22107,N_19973,N_20686);
nand U22108 (N_22108,N_19652,N_20456);
nand U22109 (N_22109,N_20363,N_19666);
or U22110 (N_22110,N_19519,N_19775);
xor U22111 (N_22111,N_20304,N_20331);
and U22112 (N_22112,N_19648,N_20572);
nor U22113 (N_22113,N_20207,N_20820);
or U22114 (N_22114,N_20674,N_19531);
and U22115 (N_22115,N_19550,N_20036);
xnor U22116 (N_22116,N_19659,N_20499);
or U22117 (N_22117,N_20763,N_20171);
and U22118 (N_22118,N_19957,N_19872);
xor U22119 (N_22119,N_19844,N_20367);
xor U22120 (N_22120,N_20595,N_19944);
or U22121 (N_22121,N_20421,N_19687);
and U22122 (N_22122,N_20282,N_20866);
nand U22123 (N_22123,N_20000,N_20586);
or U22124 (N_22124,N_20226,N_19935);
and U22125 (N_22125,N_20260,N_20926);
nor U22126 (N_22126,N_20778,N_19776);
nor U22127 (N_22127,N_20642,N_19711);
or U22128 (N_22128,N_20330,N_20826);
or U22129 (N_22129,N_19905,N_20772);
and U22130 (N_22130,N_20743,N_20154);
or U22131 (N_22131,N_19655,N_20326);
nor U22132 (N_22132,N_19727,N_20729);
nor U22133 (N_22133,N_20284,N_20520);
and U22134 (N_22134,N_20944,N_19708);
or U22135 (N_22135,N_20531,N_20709);
nand U22136 (N_22136,N_20473,N_19852);
and U22137 (N_22137,N_20224,N_19783);
and U22138 (N_22138,N_20489,N_20006);
or U22139 (N_22139,N_20965,N_20555);
xnor U22140 (N_22140,N_20556,N_19922);
or U22141 (N_22141,N_20587,N_20379);
and U22142 (N_22142,N_20311,N_20351);
nand U22143 (N_22143,N_20528,N_20228);
or U22144 (N_22144,N_20769,N_20674);
xor U22145 (N_22145,N_19902,N_20121);
or U22146 (N_22146,N_20477,N_20485);
nand U22147 (N_22147,N_20865,N_19533);
nor U22148 (N_22148,N_20399,N_20885);
and U22149 (N_22149,N_20645,N_20377);
xor U22150 (N_22150,N_20654,N_20968);
or U22151 (N_22151,N_20053,N_19823);
and U22152 (N_22152,N_20566,N_19675);
xnor U22153 (N_22153,N_19920,N_19530);
xor U22154 (N_22154,N_20265,N_20357);
xor U22155 (N_22155,N_20773,N_19681);
xnor U22156 (N_22156,N_19713,N_20281);
and U22157 (N_22157,N_19616,N_19655);
and U22158 (N_22158,N_20987,N_19602);
xnor U22159 (N_22159,N_20152,N_20712);
xnor U22160 (N_22160,N_20157,N_19664);
xor U22161 (N_22161,N_19617,N_20272);
xnor U22162 (N_22162,N_20924,N_20180);
nand U22163 (N_22163,N_20805,N_19978);
xnor U22164 (N_22164,N_20779,N_20709);
nor U22165 (N_22165,N_20738,N_20100);
nand U22166 (N_22166,N_20326,N_20194);
or U22167 (N_22167,N_20909,N_20108);
xnor U22168 (N_22168,N_19737,N_20906);
xor U22169 (N_22169,N_19551,N_20489);
and U22170 (N_22170,N_20498,N_20049);
nor U22171 (N_22171,N_20079,N_19939);
nor U22172 (N_22172,N_19763,N_20722);
nand U22173 (N_22173,N_20841,N_20581);
and U22174 (N_22174,N_19693,N_19584);
and U22175 (N_22175,N_20421,N_19922);
nand U22176 (N_22176,N_20599,N_20040);
or U22177 (N_22177,N_20832,N_19950);
and U22178 (N_22178,N_20853,N_19623);
xnor U22179 (N_22179,N_19627,N_20197);
nand U22180 (N_22180,N_20204,N_19919);
xor U22181 (N_22181,N_19809,N_19592);
xor U22182 (N_22182,N_19546,N_20833);
or U22183 (N_22183,N_19722,N_20573);
xor U22184 (N_22184,N_20707,N_19586);
or U22185 (N_22185,N_20889,N_19530);
or U22186 (N_22186,N_20992,N_20121);
nand U22187 (N_22187,N_19509,N_20543);
xnor U22188 (N_22188,N_20160,N_20913);
nand U22189 (N_22189,N_20030,N_20696);
or U22190 (N_22190,N_19650,N_20991);
xor U22191 (N_22191,N_20222,N_20903);
and U22192 (N_22192,N_19517,N_19585);
nor U22193 (N_22193,N_20958,N_20923);
xor U22194 (N_22194,N_19831,N_20421);
or U22195 (N_22195,N_19526,N_20566);
and U22196 (N_22196,N_19987,N_19582);
nor U22197 (N_22197,N_20160,N_19720);
or U22198 (N_22198,N_19681,N_20168);
xnor U22199 (N_22199,N_20026,N_19501);
and U22200 (N_22200,N_20048,N_19694);
and U22201 (N_22201,N_19945,N_19861);
and U22202 (N_22202,N_19988,N_19615);
nor U22203 (N_22203,N_20540,N_19705);
nand U22204 (N_22204,N_20522,N_20366);
nor U22205 (N_22205,N_20332,N_20986);
nand U22206 (N_22206,N_20212,N_19734);
nor U22207 (N_22207,N_19961,N_19791);
or U22208 (N_22208,N_20034,N_20896);
nor U22209 (N_22209,N_20008,N_20378);
or U22210 (N_22210,N_19594,N_20635);
and U22211 (N_22211,N_20666,N_19659);
nor U22212 (N_22212,N_19885,N_19523);
nand U22213 (N_22213,N_20619,N_19736);
nor U22214 (N_22214,N_20598,N_19818);
xor U22215 (N_22215,N_19524,N_19906);
nor U22216 (N_22216,N_20812,N_19530);
xor U22217 (N_22217,N_19960,N_20277);
or U22218 (N_22218,N_20760,N_20574);
or U22219 (N_22219,N_20025,N_19895);
and U22220 (N_22220,N_20587,N_20234);
xnor U22221 (N_22221,N_19500,N_19790);
or U22222 (N_22222,N_20009,N_20534);
and U22223 (N_22223,N_20191,N_20939);
nor U22224 (N_22224,N_20119,N_19548);
nor U22225 (N_22225,N_20847,N_20228);
nand U22226 (N_22226,N_20030,N_20886);
nand U22227 (N_22227,N_20981,N_20200);
xnor U22228 (N_22228,N_19641,N_19887);
and U22229 (N_22229,N_20826,N_19560);
or U22230 (N_22230,N_19747,N_20605);
or U22231 (N_22231,N_19747,N_19976);
and U22232 (N_22232,N_20979,N_20503);
nand U22233 (N_22233,N_20471,N_20289);
and U22234 (N_22234,N_20609,N_20275);
xor U22235 (N_22235,N_20022,N_19686);
xnor U22236 (N_22236,N_20779,N_20470);
and U22237 (N_22237,N_20082,N_19543);
xnor U22238 (N_22238,N_19807,N_20398);
xor U22239 (N_22239,N_20455,N_20042);
nor U22240 (N_22240,N_20506,N_20815);
xor U22241 (N_22241,N_20297,N_19518);
xnor U22242 (N_22242,N_19828,N_20260);
and U22243 (N_22243,N_20944,N_20831);
nor U22244 (N_22244,N_19763,N_20754);
or U22245 (N_22245,N_20736,N_20437);
and U22246 (N_22246,N_20285,N_20138);
nor U22247 (N_22247,N_19777,N_20529);
and U22248 (N_22248,N_19527,N_20872);
nand U22249 (N_22249,N_20387,N_19842);
or U22250 (N_22250,N_20229,N_19517);
and U22251 (N_22251,N_20930,N_20542);
and U22252 (N_22252,N_20734,N_20348);
xnor U22253 (N_22253,N_20523,N_20790);
or U22254 (N_22254,N_19795,N_20949);
or U22255 (N_22255,N_19962,N_20961);
or U22256 (N_22256,N_20745,N_20318);
or U22257 (N_22257,N_20405,N_20119);
and U22258 (N_22258,N_19685,N_19896);
nand U22259 (N_22259,N_20847,N_20739);
xnor U22260 (N_22260,N_19799,N_20865);
or U22261 (N_22261,N_19997,N_20648);
and U22262 (N_22262,N_20705,N_20501);
or U22263 (N_22263,N_19616,N_19521);
nand U22264 (N_22264,N_19929,N_20731);
xnor U22265 (N_22265,N_20359,N_19925);
nor U22266 (N_22266,N_20956,N_19579);
xnor U22267 (N_22267,N_20179,N_20802);
nand U22268 (N_22268,N_19721,N_20317);
and U22269 (N_22269,N_20963,N_19597);
and U22270 (N_22270,N_20430,N_19688);
xnor U22271 (N_22271,N_20163,N_19875);
xnor U22272 (N_22272,N_20200,N_20198);
nor U22273 (N_22273,N_20079,N_20173);
nor U22274 (N_22274,N_20523,N_19751);
nand U22275 (N_22275,N_20613,N_19947);
and U22276 (N_22276,N_19909,N_19538);
xor U22277 (N_22277,N_20343,N_20717);
xnor U22278 (N_22278,N_19513,N_19904);
nor U22279 (N_22279,N_20261,N_19944);
xnor U22280 (N_22280,N_20889,N_19681);
nor U22281 (N_22281,N_19511,N_19627);
and U22282 (N_22282,N_20587,N_20561);
xnor U22283 (N_22283,N_20849,N_20990);
nand U22284 (N_22284,N_20588,N_20307);
nand U22285 (N_22285,N_20755,N_19962);
and U22286 (N_22286,N_20432,N_20174);
nor U22287 (N_22287,N_19939,N_20251);
nand U22288 (N_22288,N_20842,N_20762);
or U22289 (N_22289,N_20527,N_19752);
xor U22290 (N_22290,N_19697,N_20915);
xnor U22291 (N_22291,N_19578,N_19745);
nor U22292 (N_22292,N_20401,N_20251);
nor U22293 (N_22293,N_19746,N_20679);
and U22294 (N_22294,N_20181,N_20687);
and U22295 (N_22295,N_20372,N_20842);
nor U22296 (N_22296,N_20421,N_19553);
nor U22297 (N_22297,N_20983,N_19647);
nand U22298 (N_22298,N_19719,N_20981);
nor U22299 (N_22299,N_20813,N_19683);
nand U22300 (N_22300,N_20607,N_19601);
nor U22301 (N_22301,N_20205,N_20298);
xnor U22302 (N_22302,N_19941,N_20370);
nand U22303 (N_22303,N_20645,N_20526);
xnor U22304 (N_22304,N_20441,N_20036);
or U22305 (N_22305,N_19978,N_19651);
nand U22306 (N_22306,N_19689,N_20664);
or U22307 (N_22307,N_19862,N_19836);
nand U22308 (N_22308,N_19674,N_20299);
nor U22309 (N_22309,N_20692,N_20439);
and U22310 (N_22310,N_19879,N_20686);
nand U22311 (N_22311,N_20162,N_20425);
nor U22312 (N_22312,N_20478,N_19778);
xor U22313 (N_22313,N_20971,N_20599);
nor U22314 (N_22314,N_20971,N_20436);
and U22315 (N_22315,N_19732,N_20695);
xor U22316 (N_22316,N_20851,N_19796);
nor U22317 (N_22317,N_19705,N_20505);
and U22318 (N_22318,N_20382,N_20301);
and U22319 (N_22319,N_19533,N_19722);
and U22320 (N_22320,N_20584,N_19722);
nand U22321 (N_22321,N_20637,N_19985);
nor U22322 (N_22322,N_20573,N_20177);
nor U22323 (N_22323,N_20075,N_20994);
nand U22324 (N_22324,N_20778,N_20990);
xor U22325 (N_22325,N_20430,N_20462);
nand U22326 (N_22326,N_19872,N_19826);
nand U22327 (N_22327,N_19966,N_19713);
nor U22328 (N_22328,N_20901,N_20620);
nor U22329 (N_22329,N_19913,N_20067);
xnor U22330 (N_22330,N_20474,N_20458);
nor U22331 (N_22331,N_20465,N_20601);
nand U22332 (N_22332,N_20351,N_20775);
xnor U22333 (N_22333,N_20967,N_20979);
nand U22334 (N_22334,N_20749,N_20836);
nor U22335 (N_22335,N_19849,N_19869);
xor U22336 (N_22336,N_20394,N_20171);
nor U22337 (N_22337,N_19543,N_19822);
nor U22338 (N_22338,N_19837,N_19625);
xor U22339 (N_22339,N_19622,N_20682);
or U22340 (N_22340,N_19720,N_20538);
nand U22341 (N_22341,N_19814,N_20905);
and U22342 (N_22342,N_19747,N_20108);
xor U22343 (N_22343,N_20715,N_19687);
nand U22344 (N_22344,N_20819,N_20996);
nand U22345 (N_22345,N_20989,N_19859);
or U22346 (N_22346,N_20894,N_20020);
or U22347 (N_22347,N_19761,N_19797);
nand U22348 (N_22348,N_19595,N_20494);
xnor U22349 (N_22349,N_20988,N_20959);
nor U22350 (N_22350,N_20592,N_19941);
nor U22351 (N_22351,N_20270,N_20844);
or U22352 (N_22352,N_20433,N_20442);
and U22353 (N_22353,N_19668,N_20621);
nor U22354 (N_22354,N_19828,N_20591);
nand U22355 (N_22355,N_20953,N_20415);
xnor U22356 (N_22356,N_20007,N_19640);
xor U22357 (N_22357,N_20434,N_20075);
nand U22358 (N_22358,N_20349,N_20082);
nor U22359 (N_22359,N_20271,N_20159);
or U22360 (N_22360,N_20020,N_19517);
nand U22361 (N_22361,N_20101,N_19501);
or U22362 (N_22362,N_19997,N_19909);
and U22363 (N_22363,N_19835,N_19531);
nand U22364 (N_22364,N_20196,N_20328);
nand U22365 (N_22365,N_20307,N_20533);
or U22366 (N_22366,N_19666,N_19855);
nor U22367 (N_22367,N_20155,N_20364);
nor U22368 (N_22368,N_20883,N_20291);
nor U22369 (N_22369,N_20516,N_20117);
nor U22370 (N_22370,N_20103,N_19598);
nor U22371 (N_22371,N_20876,N_19846);
nor U22372 (N_22372,N_20148,N_20747);
and U22373 (N_22373,N_19814,N_20146);
and U22374 (N_22374,N_20712,N_20346);
xor U22375 (N_22375,N_20096,N_19783);
xnor U22376 (N_22376,N_20461,N_20339);
nand U22377 (N_22377,N_20599,N_19515);
xnor U22378 (N_22378,N_20552,N_20691);
or U22379 (N_22379,N_19621,N_20119);
xnor U22380 (N_22380,N_20259,N_20048);
nand U22381 (N_22381,N_20293,N_20962);
and U22382 (N_22382,N_20736,N_20610);
xor U22383 (N_22383,N_20702,N_19849);
nor U22384 (N_22384,N_20942,N_20450);
or U22385 (N_22385,N_19612,N_20347);
or U22386 (N_22386,N_20704,N_20423);
and U22387 (N_22387,N_19512,N_20115);
nand U22388 (N_22388,N_20875,N_20553);
and U22389 (N_22389,N_20174,N_20169);
nand U22390 (N_22390,N_20997,N_20545);
xor U22391 (N_22391,N_20545,N_19560);
xnor U22392 (N_22392,N_19651,N_19705);
nor U22393 (N_22393,N_20780,N_20031);
nand U22394 (N_22394,N_20331,N_19780);
or U22395 (N_22395,N_19722,N_19578);
nand U22396 (N_22396,N_20819,N_20954);
nor U22397 (N_22397,N_19982,N_20079);
or U22398 (N_22398,N_19998,N_20233);
and U22399 (N_22399,N_20408,N_20438);
xor U22400 (N_22400,N_20362,N_19508);
xor U22401 (N_22401,N_19658,N_20747);
xor U22402 (N_22402,N_20025,N_20329);
and U22403 (N_22403,N_20975,N_20784);
and U22404 (N_22404,N_20913,N_19874);
xnor U22405 (N_22405,N_19680,N_19774);
nand U22406 (N_22406,N_20563,N_20841);
nand U22407 (N_22407,N_20489,N_19522);
or U22408 (N_22408,N_20747,N_19578);
nor U22409 (N_22409,N_20197,N_20917);
nor U22410 (N_22410,N_19671,N_19575);
or U22411 (N_22411,N_19989,N_20139);
nor U22412 (N_22412,N_19950,N_20885);
nand U22413 (N_22413,N_20372,N_19977);
or U22414 (N_22414,N_20033,N_20370);
xnor U22415 (N_22415,N_20825,N_19519);
or U22416 (N_22416,N_19899,N_20839);
or U22417 (N_22417,N_19931,N_19891);
nand U22418 (N_22418,N_20919,N_20616);
nand U22419 (N_22419,N_20692,N_20104);
and U22420 (N_22420,N_20513,N_20633);
or U22421 (N_22421,N_20082,N_20818);
nand U22422 (N_22422,N_20886,N_20278);
nor U22423 (N_22423,N_19834,N_19900);
nor U22424 (N_22424,N_20586,N_20151);
or U22425 (N_22425,N_20739,N_20887);
or U22426 (N_22426,N_20690,N_19873);
xor U22427 (N_22427,N_19978,N_20260);
nor U22428 (N_22428,N_19599,N_19814);
xor U22429 (N_22429,N_20562,N_20229);
xor U22430 (N_22430,N_20562,N_19535);
or U22431 (N_22431,N_19683,N_20852);
nand U22432 (N_22432,N_19828,N_20453);
nand U22433 (N_22433,N_19766,N_20244);
xnor U22434 (N_22434,N_19862,N_20703);
and U22435 (N_22435,N_20496,N_20692);
nor U22436 (N_22436,N_19941,N_20457);
xnor U22437 (N_22437,N_20828,N_20311);
nor U22438 (N_22438,N_20684,N_20033);
nor U22439 (N_22439,N_20374,N_19912);
xor U22440 (N_22440,N_20708,N_20074);
nand U22441 (N_22441,N_19895,N_19845);
xnor U22442 (N_22442,N_20872,N_20065);
or U22443 (N_22443,N_19614,N_19964);
nand U22444 (N_22444,N_19611,N_20699);
xnor U22445 (N_22445,N_20159,N_19631);
or U22446 (N_22446,N_20383,N_19511);
and U22447 (N_22447,N_20579,N_20194);
or U22448 (N_22448,N_20707,N_19890);
and U22449 (N_22449,N_20061,N_20024);
nor U22450 (N_22450,N_19649,N_20640);
or U22451 (N_22451,N_20081,N_19523);
nor U22452 (N_22452,N_20467,N_20448);
xnor U22453 (N_22453,N_20148,N_20766);
nand U22454 (N_22454,N_20034,N_19786);
xnor U22455 (N_22455,N_19681,N_19821);
or U22456 (N_22456,N_20718,N_20604);
or U22457 (N_22457,N_20857,N_20983);
nor U22458 (N_22458,N_20221,N_19581);
or U22459 (N_22459,N_20435,N_20167);
nor U22460 (N_22460,N_20991,N_20477);
or U22461 (N_22461,N_20729,N_19793);
nor U22462 (N_22462,N_20656,N_19627);
and U22463 (N_22463,N_20503,N_19779);
nand U22464 (N_22464,N_20668,N_20420);
xor U22465 (N_22465,N_19833,N_20966);
nor U22466 (N_22466,N_20768,N_20897);
and U22467 (N_22467,N_19703,N_20656);
nand U22468 (N_22468,N_20526,N_20546);
or U22469 (N_22469,N_20032,N_20250);
nand U22470 (N_22470,N_19792,N_20764);
xor U22471 (N_22471,N_20487,N_20942);
nand U22472 (N_22472,N_19801,N_19866);
nand U22473 (N_22473,N_20766,N_19988);
xor U22474 (N_22474,N_20382,N_20900);
nor U22475 (N_22475,N_19709,N_20959);
or U22476 (N_22476,N_20852,N_20621);
nand U22477 (N_22477,N_19604,N_20501);
nand U22478 (N_22478,N_19921,N_19710);
or U22479 (N_22479,N_19890,N_20291);
and U22480 (N_22480,N_19553,N_19752);
and U22481 (N_22481,N_20360,N_20569);
nand U22482 (N_22482,N_19855,N_20014);
or U22483 (N_22483,N_20464,N_19915);
nand U22484 (N_22484,N_20488,N_20816);
or U22485 (N_22485,N_20130,N_20306);
nor U22486 (N_22486,N_19537,N_20079);
or U22487 (N_22487,N_19747,N_19916);
nor U22488 (N_22488,N_20477,N_19999);
nand U22489 (N_22489,N_20232,N_20148);
xor U22490 (N_22490,N_20639,N_20119);
and U22491 (N_22491,N_20194,N_20121);
and U22492 (N_22492,N_20561,N_20010);
nand U22493 (N_22493,N_20397,N_20236);
and U22494 (N_22494,N_19640,N_20798);
nor U22495 (N_22495,N_19652,N_19662);
xnor U22496 (N_22496,N_19773,N_20844);
and U22497 (N_22497,N_20503,N_20514);
xor U22498 (N_22498,N_20840,N_20195);
xnor U22499 (N_22499,N_20559,N_20673);
nand U22500 (N_22500,N_21484,N_21413);
nand U22501 (N_22501,N_22170,N_21086);
xor U22502 (N_22502,N_22121,N_21813);
nand U22503 (N_22503,N_22471,N_22235);
xnor U22504 (N_22504,N_21850,N_22130);
or U22505 (N_22505,N_21639,N_21949);
nor U22506 (N_22506,N_21960,N_21728);
nand U22507 (N_22507,N_21750,N_22340);
and U22508 (N_22508,N_21723,N_21306);
xor U22509 (N_22509,N_21556,N_21001);
and U22510 (N_22510,N_21385,N_21738);
or U22511 (N_22511,N_21171,N_22279);
and U22512 (N_22512,N_21580,N_21319);
nand U22513 (N_22513,N_21979,N_21276);
nor U22514 (N_22514,N_22006,N_22023);
nor U22515 (N_22515,N_21336,N_21618);
and U22516 (N_22516,N_22445,N_22193);
or U22517 (N_22517,N_21403,N_22200);
nor U22518 (N_22518,N_21449,N_21169);
xnor U22519 (N_22519,N_22073,N_22368);
nor U22520 (N_22520,N_21012,N_21654);
nor U22521 (N_22521,N_22143,N_21679);
or U22522 (N_22522,N_22428,N_21454);
and U22523 (N_22523,N_21530,N_21234);
nand U22524 (N_22524,N_21715,N_22353);
nand U22525 (N_22525,N_22302,N_21225);
or U22526 (N_22526,N_21831,N_22350);
nor U22527 (N_22527,N_21082,N_21840);
nand U22528 (N_22528,N_22425,N_21818);
nand U22529 (N_22529,N_21571,N_22265);
or U22530 (N_22530,N_21548,N_21295);
nand U22531 (N_22531,N_21474,N_21810);
and U22532 (N_22532,N_21933,N_22267);
and U22533 (N_22533,N_21724,N_21190);
nor U22534 (N_22534,N_21433,N_21322);
or U22535 (N_22535,N_21749,N_21861);
xnor U22536 (N_22536,N_21983,N_22079);
or U22537 (N_22537,N_22015,N_22082);
xor U22538 (N_22538,N_21896,N_21281);
or U22539 (N_22539,N_22002,N_21343);
nor U22540 (N_22540,N_21809,N_21976);
nand U22541 (N_22541,N_21819,N_21080);
nor U22542 (N_22542,N_21758,N_21998);
nor U22543 (N_22543,N_22278,N_22078);
nand U22544 (N_22544,N_21874,N_22145);
nor U22545 (N_22545,N_21131,N_22258);
and U22546 (N_22546,N_21664,N_21019);
nor U22547 (N_22547,N_21047,N_22323);
xnor U22548 (N_22548,N_21858,N_21803);
nor U22549 (N_22549,N_22198,N_21994);
xnor U22550 (N_22550,N_21613,N_21946);
and U22551 (N_22551,N_21686,N_22185);
nand U22552 (N_22552,N_21305,N_22228);
and U22553 (N_22553,N_21666,N_22106);
xnor U22554 (N_22554,N_21699,N_21646);
nand U22555 (N_22555,N_21718,N_21529);
nand U22556 (N_22556,N_21538,N_22105);
nand U22557 (N_22557,N_21505,N_21263);
xnor U22558 (N_22558,N_21521,N_22150);
and U22559 (N_22559,N_21923,N_21503);
nor U22560 (N_22560,N_21212,N_21962);
or U22561 (N_22561,N_21910,N_22245);
nor U22562 (N_22562,N_21106,N_21761);
or U22563 (N_22563,N_22019,N_22036);
or U22564 (N_22564,N_22196,N_22379);
and U22565 (N_22565,N_22155,N_22303);
or U22566 (N_22566,N_22022,N_22418);
nor U22567 (N_22567,N_21161,N_21844);
xor U22568 (N_22568,N_21648,N_21703);
xor U22569 (N_22569,N_21271,N_21692);
or U22570 (N_22570,N_21149,N_21203);
nor U22571 (N_22571,N_21342,N_21873);
xnor U22572 (N_22572,N_21172,N_22383);
or U22573 (N_22573,N_21720,N_22238);
or U22574 (N_22574,N_21637,N_22210);
xnor U22575 (N_22575,N_21845,N_21722);
or U22576 (N_22576,N_21359,N_21997);
nand U22577 (N_22577,N_21045,N_21361);
nand U22578 (N_22578,N_21440,N_21763);
or U22579 (N_22579,N_21445,N_21003);
xor U22580 (N_22580,N_21489,N_21768);
nor U22581 (N_22581,N_21655,N_21292);
nor U22582 (N_22582,N_21783,N_21363);
nor U22583 (N_22583,N_21888,N_21643);
and U22584 (N_22584,N_21901,N_21553);
nor U22585 (N_22585,N_22049,N_22342);
or U22586 (N_22586,N_22024,N_21132);
nor U22587 (N_22587,N_21074,N_21140);
nand U22588 (N_22588,N_21255,N_22415);
and U22589 (N_22589,N_21407,N_21875);
nor U22590 (N_22590,N_21437,N_21789);
or U22591 (N_22591,N_22239,N_21536);
or U22592 (N_22592,N_21100,N_21855);
xnor U22593 (N_22593,N_21352,N_22213);
nand U22594 (N_22594,N_21682,N_21614);
nand U22595 (N_22595,N_21137,N_21830);
nor U22596 (N_22596,N_21220,N_21545);
xnor U22597 (N_22597,N_22014,N_21041);
or U22598 (N_22598,N_21675,N_22395);
nor U22599 (N_22599,N_21727,N_21817);
and U22600 (N_22600,N_21714,N_21439);
and U22601 (N_22601,N_22467,N_22042);
or U22602 (N_22602,N_21911,N_22160);
or U22603 (N_22603,N_22183,N_21357);
or U22604 (N_22604,N_21611,N_22236);
nand U22605 (N_22605,N_21173,N_21154);
nor U22606 (N_22606,N_22360,N_22206);
and U22607 (N_22607,N_21434,N_21564);
and U22608 (N_22608,N_21381,N_21573);
xnor U22609 (N_22609,N_22435,N_21869);
nor U22610 (N_22610,N_22404,N_21460);
nor U22611 (N_22611,N_22133,N_21656);
nor U22612 (N_22612,N_21448,N_21967);
nand U22613 (N_22613,N_21044,N_21288);
xor U22614 (N_22614,N_22362,N_21522);
nor U22615 (N_22615,N_22240,N_22306);
or U22616 (N_22616,N_22068,N_21591);
or U22617 (N_22617,N_21891,N_22051);
nand U22618 (N_22618,N_21287,N_21630);
nand U22619 (N_22619,N_21252,N_21547);
xor U22620 (N_22620,N_21283,N_22461);
or U22621 (N_22621,N_22394,N_21067);
nand U22622 (N_22622,N_21502,N_21755);
nor U22623 (N_22623,N_21954,N_22232);
or U22624 (N_22624,N_22046,N_21272);
and U22625 (N_22625,N_21736,N_22005);
and U22626 (N_22626,N_21575,N_22347);
nor U22627 (N_22627,N_22080,N_22016);
or U22628 (N_22628,N_21739,N_22473);
xor U22629 (N_22629,N_21446,N_22411);
xor U22630 (N_22630,N_21774,N_22289);
or U22631 (N_22631,N_21133,N_21752);
or U22632 (N_22632,N_21174,N_22187);
and U22633 (N_22633,N_21216,N_21313);
and U22634 (N_22634,N_21661,N_21631);
nand U22635 (N_22635,N_21790,N_21531);
or U22636 (N_22636,N_21370,N_22189);
or U22637 (N_22637,N_21918,N_21237);
or U22638 (N_22638,N_22367,N_22077);
xor U22639 (N_22639,N_21912,N_21982);
xor U22640 (N_22640,N_21092,N_22241);
and U22641 (N_22641,N_21827,N_22431);
or U22642 (N_22642,N_22484,N_21590);
xnor U22643 (N_22643,N_21680,N_22021);
nor U22644 (N_22644,N_22216,N_21985);
and U22645 (N_22645,N_21146,N_21649);
nor U22646 (N_22646,N_22380,N_22389);
nand U22647 (N_22647,N_22297,N_21138);
xor U22648 (N_22648,N_22172,N_21963);
or U22649 (N_22649,N_21898,N_21170);
nor U22650 (N_22650,N_21984,N_21841);
nor U22651 (N_22651,N_22357,N_21640);
or U22652 (N_22652,N_22136,N_21353);
xnor U22653 (N_22653,N_21696,N_21026);
and U22654 (N_22654,N_22163,N_22139);
or U22655 (N_22655,N_21641,N_22178);
nor U22656 (N_22656,N_22407,N_21540);
and U22657 (N_22657,N_21043,N_21475);
and U22658 (N_22658,N_21593,N_21602);
nand U22659 (N_22659,N_21002,N_22045);
nand U22660 (N_22660,N_21953,N_21355);
nand U22661 (N_22661,N_21064,N_21402);
and U22662 (N_22662,N_22413,N_21691);
and U22663 (N_22663,N_21205,N_21859);
xnor U22664 (N_22664,N_21491,N_21596);
or U22665 (N_22665,N_22094,N_21307);
or U22666 (N_22666,N_21990,N_22040);
or U22667 (N_22667,N_21156,N_21846);
or U22668 (N_22668,N_21384,N_21430);
nand U22669 (N_22669,N_21835,N_21121);
or U22670 (N_22670,N_21629,N_21122);
nor U22671 (N_22671,N_21606,N_21419);
xor U22672 (N_22672,N_22218,N_22260);
nor U22673 (N_22673,N_21551,N_21392);
xnor U22674 (N_22674,N_21552,N_22287);
nor U22675 (N_22675,N_22332,N_21730);
nand U22676 (N_22676,N_21334,N_21936);
nand U22677 (N_22677,N_21158,N_21317);
and U22678 (N_22678,N_21472,N_21777);
and U22679 (N_22679,N_21023,N_21324);
nand U22680 (N_22680,N_21500,N_22304);
and U22681 (N_22681,N_22345,N_22424);
nand U22682 (N_22682,N_21337,N_21128);
xnor U22683 (N_22683,N_22153,N_21127);
or U22684 (N_22684,N_21470,N_21110);
or U22685 (N_22685,N_21671,N_21525);
xor U22686 (N_22686,N_21665,N_21151);
and U22687 (N_22687,N_21136,N_22305);
and U22688 (N_22688,N_21259,N_21235);
nor U22689 (N_22689,N_22157,N_21424);
nand U22690 (N_22690,N_22169,N_21969);
or U22691 (N_22691,N_22086,N_22122);
xnor U22692 (N_22692,N_21612,N_22038);
or U22693 (N_22693,N_22430,N_21134);
nor U22694 (N_22694,N_22039,N_21988);
or U22695 (N_22695,N_21729,N_21488);
nand U22696 (N_22696,N_21465,N_22470);
nor U22697 (N_22697,N_21479,N_22041);
and U22698 (N_22698,N_21285,N_21678);
xor U22699 (N_22699,N_21247,N_21050);
or U22700 (N_22700,N_21597,N_21093);
or U22701 (N_22701,N_22207,N_21016);
or U22702 (N_22702,N_21458,N_21964);
and U22703 (N_22703,N_21579,N_21406);
and U22704 (N_22704,N_22284,N_21404);
nor U22705 (N_22705,N_21076,N_22351);
nand U22706 (N_22706,N_22165,N_22377);
xnor U22707 (N_22707,N_21717,N_22399);
nand U22708 (N_22708,N_21296,N_21327);
xor U22709 (N_22709,N_22453,N_21786);
and U22710 (N_22710,N_22468,N_22254);
and U22711 (N_22711,N_21583,N_21609);
and U22712 (N_22712,N_22075,N_21248);
nor U22713 (N_22713,N_22249,N_22203);
and U22714 (N_22714,N_22017,N_21557);
xnor U22715 (N_22715,N_22371,N_22375);
and U22716 (N_22716,N_21528,N_21354);
nor U22717 (N_22717,N_21084,N_21759);
nor U22718 (N_22718,N_21632,N_22147);
nor U22719 (N_22719,N_21034,N_21395);
nand U22720 (N_22720,N_21326,N_21516);
nand U22721 (N_22721,N_21834,N_21226);
or U22722 (N_22722,N_22188,N_21107);
nand U22723 (N_22723,N_21401,N_22363);
nor U22724 (N_22724,N_21275,N_22293);
nor U22725 (N_22725,N_21396,N_21518);
or U22726 (N_22726,N_21892,N_21941);
nand U22727 (N_22727,N_22124,N_22382);
nand U22728 (N_22728,N_22137,N_22223);
or U22729 (N_22729,N_22234,N_21471);
or U22730 (N_22730,N_21356,N_22171);
nand U22731 (N_22731,N_21496,N_21367);
nand U22732 (N_22732,N_22104,N_21265);
nand U22733 (N_22733,N_22199,N_21509);
or U22734 (N_22734,N_21523,N_21822);
xor U22735 (N_22735,N_21622,N_22409);
or U22736 (N_22736,N_21344,N_22361);
nand U22737 (N_22737,N_21376,N_21927);
xor U22738 (N_22738,N_21013,N_22119);
nand U22739 (N_22739,N_21719,N_21456);
or U22740 (N_22740,N_21186,N_22149);
xnor U22741 (N_22741,N_21436,N_21996);
nor U22742 (N_22742,N_22099,N_21812);
or U22743 (N_22743,N_22277,N_21486);
nor U22744 (N_22744,N_21077,N_22202);
or U22745 (N_22745,N_21558,N_21742);
or U22746 (N_22746,N_21346,N_21358);
nor U22747 (N_22747,N_21669,N_22091);
and U22748 (N_22748,N_21196,N_21181);
and U22749 (N_22749,N_21708,N_21599);
xnor U22750 (N_22750,N_21115,N_22455);
xnor U22751 (N_22751,N_22312,N_22176);
nor U22752 (N_22752,N_21857,N_21210);
or U22753 (N_22753,N_21177,N_21040);
and U22754 (N_22754,N_22055,N_21239);
and U22755 (N_22755,N_22346,N_21435);
or U22756 (N_22756,N_21236,N_21464);
nand U22757 (N_22757,N_21139,N_22285);
nand U22758 (N_22758,N_21231,N_22369);
or U22759 (N_22759,N_21821,N_21610);
nor U22760 (N_22760,N_21792,N_21908);
xor U22761 (N_22761,N_22333,N_21560);
nor U22762 (N_22762,N_22283,N_21520);
or U22763 (N_22763,N_22372,N_22412);
nor U22764 (N_22764,N_22164,N_21483);
or U22765 (N_22765,N_21124,N_21194);
and U22766 (N_22766,N_21673,N_21219);
xor U22767 (N_22767,N_22443,N_22292);
xnor U22768 (N_22768,N_21847,N_21498);
or U22769 (N_22769,N_22403,N_21224);
nand U22770 (N_22770,N_21069,N_22489);
or U22771 (N_22771,N_21088,N_21141);
or U22772 (N_22772,N_22324,N_21517);
and U22773 (N_22773,N_22151,N_21785);
nand U22774 (N_22774,N_22182,N_22250);
nor U22775 (N_22775,N_22309,N_21201);
xnor U22776 (N_22776,N_21348,N_21974);
nand U22777 (N_22777,N_21762,N_21278);
or U22778 (N_22778,N_21005,N_21431);
nor U22779 (N_22779,N_21290,N_21147);
and U22780 (N_22780,N_22269,N_22112);
and U22781 (N_22781,N_22209,N_22387);
and U22782 (N_22782,N_21716,N_22261);
or U22783 (N_22783,N_22111,N_21427);
and U22784 (N_22784,N_21198,N_21565);
nand U22785 (N_22785,N_21094,N_21603);
nor U22786 (N_22786,N_21162,N_21339);
nor U22787 (N_22787,N_21549,N_21176);
nor U22788 (N_22788,N_21600,N_21024);
or U22789 (N_22789,N_22220,N_21684);
nor U22790 (N_22790,N_21906,N_22328);
nand U22791 (N_22791,N_21709,N_21090);
and U22792 (N_22792,N_22339,N_21737);
xnor U22793 (N_22793,N_21770,N_22414);
nand U22794 (N_22794,N_21808,N_21443);
xnor U22795 (N_22795,N_21331,N_22444);
nand U22796 (N_22796,N_21797,N_21350);
or U22797 (N_22797,N_22081,N_21939);
nand U22798 (N_22798,N_21119,N_22497);
nor U22799 (N_22799,N_21644,N_21543);
xnor U22800 (N_22800,N_22156,N_21950);
nand U22801 (N_22801,N_21900,N_22201);
nor U22802 (N_22802,N_21102,N_21633);
and U22803 (N_22803,N_22276,N_21153);
and U22804 (N_22804,N_22483,N_22442);
and U22805 (N_22805,N_22295,N_22364);
nand U22806 (N_22806,N_21227,N_22402);
or U22807 (N_22807,N_21981,N_21452);
nor U22808 (N_22808,N_21754,N_21061);
or U22809 (N_22809,N_21148,N_21405);
and U22810 (N_22810,N_22013,N_21389);
and U22811 (N_22811,N_22233,N_21364);
nand U22812 (N_22812,N_21189,N_21380);
nand U22813 (N_22813,N_21662,N_21320);
or U22814 (N_22814,N_21214,N_21200);
xnor U22815 (N_22815,N_21929,N_21282);
or U22816 (N_22816,N_21550,N_21059);
xor U22817 (N_22817,N_22034,N_21126);
nand U22818 (N_22818,N_22438,N_21347);
or U22819 (N_22819,N_21109,N_21078);
and U22820 (N_22820,N_22001,N_21542);
xor U22821 (N_22821,N_21721,N_22102);
or U22822 (N_22822,N_21638,N_21693);
or U22823 (N_22823,N_21453,N_21928);
xnor U22824 (N_22824,N_22307,N_21595);
or U22825 (N_22825,N_21025,N_21297);
xnor U22826 (N_22826,N_21607,N_22381);
and U22827 (N_22827,N_21302,N_21561);
or U22828 (N_22828,N_21624,N_21152);
nand U22829 (N_22829,N_21410,N_21877);
or U22830 (N_22830,N_21804,N_21280);
and U22831 (N_22831,N_21300,N_22495);
and U22832 (N_22832,N_21568,N_21702);
nand U22833 (N_22833,N_21011,N_21065);
or U22834 (N_22834,N_21805,N_21033);
and U22835 (N_22835,N_22370,N_22141);
or U22836 (N_22836,N_21240,N_21164);
nor U22837 (N_22837,N_21291,N_22230);
xnor U22838 (N_22838,N_22474,N_22158);
or U22839 (N_22839,N_22074,N_21249);
xnor U22840 (N_22840,N_21885,N_21418);
or U22841 (N_22841,N_21921,N_22067);
or U22842 (N_22842,N_21112,N_21698);
and U22843 (N_22843,N_21099,N_22162);
nor U22844 (N_22844,N_21793,N_22174);
or U22845 (N_22845,N_21802,N_21965);
and U22846 (N_22846,N_21746,N_21031);
nand U22847 (N_22847,N_22101,N_22486);
nand U22848 (N_22848,N_21052,N_21992);
or U22849 (N_22849,N_21987,N_22492);
nand U22850 (N_22850,N_22208,N_21116);
and U22851 (N_22851,N_22215,N_21743);
xor U22852 (N_22852,N_21938,N_21944);
xnor U22853 (N_22853,N_21837,N_21986);
or U22854 (N_22854,N_22173,N_21261);
nand U22855 (N_22855,N_21254,N_22427);
nor U22856 (N_22856,N_21039,N_22439);
or U22857 (N_22857,N_21940,N_21694);
or U22858 (N_22858,N_21771,N_22134);
nor U22859 (N_22859,N_21318,N_21676);
and U22860 (N_22860,N_22028,N_22008);
nand U22861 (N_22861,N_22088,N_21499);
or U22862 (N_22862,N_22222,N_22378);
or U22863 (N_22863,N_21245,N_22392);
or U22864 (N_22864,N_21586,N_22098);
or U22865 (N_22865,N_21206,N_22450);
and U22866 (N_22866,N_21776,N_22437);
nor U22867 (N_22867,N_21178,N_21241);
and U22868 (N_22868,N_22298,N_22263);
nor U22869 (N_22869,N_22408,N_21461);
nand U22870 (N_22870,N_21796,N_21250);
and U22871 (N_22871,N_22114,N_22063);
xnor U22872 (N_22872,N_22460,N_22491);
nand U22873 (N_22873,N_22469,N_22354);
nor U22874 (N_22874,N_22374,N_21879);
or U22875 (N_22875,N_21087,N_21180);
nor U22876 (N_22876,N_22376,N_22103);
or U22877 (N_22877,N_21183,N_22396);
and U22878 (N_22878,N_21316,N_22142);
xnor U22879 (N_22879,N_22211,N_21604);
or U22880 (N_22880,N_22499,N_21242);
nand U22881 (N_22881,N_21924,N_22476);
nand U22882 (N_22882,N_21398,N_21130);
xor U22883 (N_22883,N_21243,N_21379);
or U22884 (N_22884,N_21815,N_22388);
xor U22885 (N_22885,N_21883,N_21978);
or U22886 (N_22886,N_21199,N_21021);
nand U22887 (N_22887,N_21386,N_22494);
nor U22888 (N_22888,N_22115,N_21187);
or U22889 (N_22889,N_22186,N_21876);
nor U22890 (N_22890,N_21415,N_21592);
xnor U22891 (N_22891,N_21791,N_22047);
and U22892 (N_22892,N_22320,N_21991);
or U22893 (N_22893,N_21626,N_22026);
and U22894 (N_22894,N_22288,N_21753);
or U22895 (N_22895,N_21351,N_21382);
nor U22896 (N_22896,N_21289,N_21383);
nor U22897 (N_22897,N_21251,N_21325);
xor U22898 (N_22898,N_21215,N_21469);
nand U22899 (N_22899,N_22004,N_21208);
nor U22900 (N_22900,N_21362,N_21029);
nand U22901 (N_22901,N_22107,N_22027);
nand U22902 (N_22902,N_21046,N_22059);
and U22903 (N_22903,N_21301,N_22062);
xor U22904 (N_22904,N_22144,N_21393);
xnor U22905 (N_22905,N_21537,N_22480);
or U22906 (N_22906,N_22432,N_22048);
or U22907 (N_22907,N_21416,N_21233);
or U22908 (N_22908,N_21444,N_21782);
and U22909 (N_22909,N_22393,N_21497);
nor U22910 (N_22910,N_21833,N_21634);
nor U22911 (N_22911,N_22448,N_21204);
nand U22912 (N_22912,N_21507,N_21478);
nor U22913 (N_22913,N_21066,N_22066);
nand U22914 (N_22914,N_22031,N_21732);
nor U22915 (N_22915,N_21970,N_21056);
nor U22916 (N_22916,N_21660,N_21482);
nand U22917 (N_22917,N_21349,N_22251);
or U22918 (N_22918,N_22069,N_21333);
nor U22919 (N_22919,N_21922,N_21390);
nand U22920 (N_22920,N_21309,N_22128);
xor U22921 (N_22921,N_21995,N_21651);
nor U22922 (N_22922,N_21246,N_21764);
nor U22923 (N_22923,N_22154,N_22282);
and U22924 (N_22924,N_21269,N_21935);
nor U22925 (N_22925,N_21956,N_22253);
nor U22926 (N_22926,N_21806,N_21798);
xor U22927 (N_22927,N_21951,N_22029);
or U22928 (N_22928,N_21229,N_22168);
nor U22929 (N_22929,N_21925,N_21903);
and U22930 (N_22930,N_21527,N_21495);
and U22931 (N_22931,N_21756,N_22030);
and U22932 (N_22932,N_22053,N_22058);
nor U22933 (N_22933,N_21218,N_22365);
or U22934 (N_22934,N_21142,N_22390);
nand U22935 (N_22935,N_21778,N_21563);
nor U22936 (N_22936,N_22300,N_22272);
nor U22937 (N_22937,N_21711,N_21476);
and U22938 (N_22938,N_22205,N_21731);
nand U22939 (N_22939,N_21532,N_21658);
and U22940 (N_22940,N_21501,N_21620);
nor U22941 (N_22941,N_22226,N_21773);
and U22942 (N_22942,N_21878,N_21823);
or U22943 (N_22943,N_22366,N_21519);
xnor U22944 (N_22944,N_21865,N_22336);
nand U22945 (N_22945,N_21825,N_21411);
nor U22946 (N_22946,N_22127,N_21057);
nor U22947 (N_22947,N_22341,N_22330);
and U22948 (N_22948,N_22264,N_22132);
nor U22949 (N_22949,N_21304,N_22018);
or U22950 (N_22950,N_22123,N_21615);
or U22951 (N_22951,N_22299,N_22237);
nor U22952 (N_22952,N_21747,N_21569);
nand U22953 (N_22953,N_21868,N_21089);
nand U22954 (N_22954,N_21657,N_21387);
or U22955 (N_22955,N_21480,N_22093);
xnor U22956 (N_22956,N_22070,N_21957);
nor U22957 (N_22957,N_22025,N_21168);
nand U22958 (N_22958,N_21725,N_21635);
and U22959 (N_22959,N_22487,N_21972);
nand U22960 (N_22960,N_22152,N_21293);
nor U22961 (N_22961,N_21959,N_21980);
nor U22962 (N_22962,N_22225,N_22227);
nand U22963 (N_22963,N_22020,N_21150);
and U22964 (N_22964,N_22076,N_21576);
and U22965 (N_22965,N_21735,N_21018);
or U22966 (N_22966,N_22419,N_22310);
and U22967 (N_22967,N_21884,N_21438);
and U22968 (N_22968,N_22175,N_21188);
nand U22969 (N_22969,N_21706,N_22064);
and U22970 (N_22970,N_21726,N_21075);
nor U22971 (N_22971,N_21417,N_21185);
nand U22972 (N_22972,N_22440,N_21695);
xnor U22973 (N_22973,N_22212,N_21765);
nor U22974 (N_22974,N_21866,N_21704);
or U22975 (N_22975,N_22057,N_21705);
nand U22976 (N_22976,N_22311,N_22397);
nor U22977 (N_22977,N_21211,N_21191);
and U22978 (N_22978,N_21388,N_21374);
or U22979 (N_22979,N_21849,N_21504);
xnor U22980 (N_22980,N_21429,N_22246);
xor U22981 (N_22981,N_22257,N_21232);
and U22982 (N_22982,N_22325,N_21572);
nor U22983 (N_22983,N_22286,N_21030);
nand U22984 (N_22984,N_22252,N_21085);
nand U22985 (N_22985,N_22481,N_21298);
or U22986 (N_22986,N_22011,N_21989);
and U22987 (N_22987,N_21934,N_21467);
and U22988 (N_22988,N_21584,N_22477);
xnor U22989 (N_22989,N_21890,N_22319);
nor U22990 (N_22990,N_22457,N_22458);
nor U22991 (N_22991,N_21973,N_22090);
and U22992 (N_22992,N_21104,N_21862);
or U22993 (N_22993,N_22243,N_21312);
nor U22994 (N_22994,N_21485,N_21993);
and U22995 (N_22995,N_21952,N_22033);
and U22996 (N_22996,N_21103,N_22056);
xor U22997 (N_22997,N_22385,N_22335);
nor U22998 (N_22998,N_21566,N_21165);
and U22999 (N_22999,N_22337,N_22485);
and U23000 (N_23000,N_21455,N_22177);
nand U23001 (N_23001,N_21787,N_22358);
or U23002 (N_23002,N_21468,N_21083);
nand U23003 (N_23003,N_22420,N_21853);
and U23004 (N_23004,N_22398,N_21340);
nand U23005 (N_23005,N_21256,N_21451);
or U23006 (N_23006,N_22129,N_21035);
nor U23007 (N_23007,N_21931,N_21447);
xnor U23008 (N_23008,N_22113,N_21687);
xor U23009 (N_23009,N_21017,N_21854);
and U23010 (N_23010,N_21423,N_21555);
nand U23011 (N_23011,N_22433,N_21966);
xnor U23012 (N_23012,N_21882,N_21734);
nor U23013 (N_23013,N_22092,N_21073);
nor U23014 (N_23014,N_21314,N_21111);
or U23015 (N_23015,N_21378,N_22463);
nand U23016 (N_23016,N_21038,N_21114);
nand U23017 (N_23017,N_21535,N_21627);
nand U23018 (N_23018,N_21621,N_22426);
xnor U23019 (N_23019,N_21477,N_21070);
or U23020 (N_23020,N_21713,N_22054);
or U23021 (N_23021,N_22343,N_21917);
or U23022 (N_23022,N_21769,N_21000);
xor U23023 (N_23023,N_22356,N_22052);
xnor U23024 (N_23024,N_21788,N_21570);
and U23025 (N_23025,N_22010,N_22296);
or U23026 (N_23026,N_21608,N_21009);
xor U23027 (N_23027,N_22043,N_22096);
nor U23028 (N_23028,N_21048,N_21541);
xnor U23029 (N_23029,N_22308,N_21578);
and U23030 (N_23030,N_22181,N_22231);
xnor U23031 (N_23031,N_21027,N_21155);
xor U23032 (N_23032,N_21697,N_21668);
nor U23033 (N_23033,N_21072,N_21975);
nand U23034 (N_23034,N_22032,N_21807);
nor U23035 (N_23035,N_21377,N_21864);
xor U23036 (N_23036,N_22221,N_22479);
nor U23037 (N_23037,N_21659,N_21311);
nor U23038 (N_23038,N_21838,N_22416);
nor U23039 (N_23039,N_21744,N_22214);
xor U23040 (N_23040,N_22349,N_21328);
and U23041 (N_23041,N_21870,N_21015);
xor U23042 (N_23042,N_22274,N_21167);
and U23043 (N_23043,N_22498,N_21179);
xnor U23044 (N_23044,N_21867,N_21457);
nand U23045 (N_23045,N_21667,N_21303);
or U23046 (N_23046,N_22259,N_22301);
nand U23047 (N_23047,N_21968,N_21372);
or U23048 (N_23048,N_21459,N_21897);
and U23049 (N_23049,N_21049,N_21587);
nor U23050 (N_23050,N_22291,N_22184);
nand U23051 (N_23051,N_22195,N_21412);
nand U23052 (N_23052,N_22410,N_21712);
nand U23053 (N_23053,N_21270,N_21098);
nand U23054 (N_23054,N_21829,N_22247);
nand U23055 (N_23055,N_21617,N_21894);
nor U23056 (N_23056,N_22044,N_22120);
and U23057 (N_23057,N_21733,N_22204);
xnor U23058 (N_23058,N_21526,N_21828);
nor U23059 (N_23059,N_22244,N_22421);
nor U23060 (N_23060,N_22192,N_21871);
nand U23061 (N_23061,N_21144,N_22400);
xnor U23062 (N_23062,N_22447,N_21286);
xor U23063 (N_23063,N_21588,N_21195);
nand U23064 (N_23064,N_21800,N_21157);
nand U23065 (N_23065,N_21071,N_21096);
nor U23066 (N_23066,N_21253,N_21268);
and U23067 (N_23067,N_22109,N_21345);
nand U23068 (N_23068,N_21581,N_22466);
xnor U23069 (N_23069,N_22138,N_21909);
or U23070 (N_23070,N_22190,N_22217);
and U23071 (N_23071,N_22327,N_21399);
xnor U23072 (N_23072,N_21097,N_22472);
nand U23073 (N_23073,N_21492,N_21244);
xor U23074 (N_23074,N_22454,N_21330);
nor U23075 (N_23075,N_21811,N_21125);
and U23076 (N_23076,N_21945,N_22035);
or U23077 (N_23077,N_21081,N_21801);
nand U23078 (N_23078,N_21284,N_21707);
nand U23079 (N_23079,N_21262,N_21450);
and U23080 (N_23080,N_22060,N_21848);
nor U23081 (N_23081,N_21701,N_22315);
nor U23082 (N_23082,N_21619,N_21863);
or U23083 (N_23083,N_22087,N_21279);
and U23084 (N_23084,N_21683,N_22313);
or U23085 (N_23085,N_22161,N_21487);
or U23086 (N_23086,N_21123,N_21799);
or U23087 (N_23087,N_21192,N_21163);
nor U23088 (N_23088,N_21108,N_21533);
nor U23089 (N_23089,N_21310,N_22423);
nor U23090 (N_23090,N_22050,N_21741);
and U23091 (N_23091,N_22334,N_21221);
nand U23092 (N_23092,N_21913,N_21915);
or U23093 (N_23093,N_21397,N_21400);
xnor U23094 (N_23094,N_22290,N_21751);
and U23095 (N_23095,N_22117,N_21510);
nand U23096 (N_23096,N_21338,N_21032);
nor U23097 (N_23097,N_21308,N_21118);
or U23098 (N_23098,N_22148,N_22100);
nand U23099 (N_23099,N_21422,N_21902);
nand U23100 (N_23100,N_21539,N_22179);
and U23101 (N_23101,N_21512,N_21645);
nand U23102 (N_23102,N_21795,N_21274);
nand U23103 (N_23103,N_22434,N_22003);
xor U23104 (N_23104,N_21315,N_21961);
nor U23105 (N_23105,N_21230,N_21373);
nor U23106 (N_23106,N_21880,N_21091);
nand U23107 (N_23107,N_21843,N_21832);
xnor U23108 (N_23108,N_21554,N_21095);
nand U23109 (N_23109,N_21159,N_21166);
nand U23110 (N_23110,N_21062,N_21856);
nor U23111 (N_23111,N_21893,N_21582);
xnor U23112 (N_23112,N_21574,N_21760);
nand U23113 (N_23113,N_21914,N_22326);
or U23114 (N_23114,N_22271,N_21685);
nor U23115 (N_23115,N_22314,N_21365);
or U23116 (N_23116,N_22373,N_21567);
xnor U23117 (N_23117,N_21420,N_22478);
nor U23118 (N_23118,N_22266,N_22449);
nand U23119 (N_23119,N_22012,N_21905);
and U23120 (N_23120,N_22095,N_22131);
or U23121 (N_23121,N_21663,N_21534);
nor U23122 (N_23122,N_22462,N_21129);
nor U23123 (N_23123,N_21544,N_21916);
nor U23124 (N_23124,N_21160,N_21625);
nand U23125 (N_23125,N_21036,N_21616);
nand U23126 (N_23126,N_22242,N_22359);
xor U23127 (N_23127,N_21428,N_22280);
nand U23128 (N_23128,N_22490,N_21779);
nor U23129 (N_23129,N_21299,N_21101);
nand U23130 (N_23130,N_21394,N_21442);
nor U23131 (N_23131,N_21636,N_21546);
nand U23132 (N_23132,N_21184,N_22496);
nand U23133 (N_23133,N_21264,N_21852);
and U23134 (N_23134,N_21466,N_21942);
and U23135 (N_23135,N_21820,N_21368);
nand U23136 (N_23136,N_22167,N_21238);
and U23137 (N_23137,N_21217,N_22270);
and U23138 (N_23138,N_22255,N_22256);
xnor U23139 (N_23139,N_21135,N_21068);
nor U23140 (N_23140,N_22180,N_21055);
nor U23141 (N_23141,N_21182,N_21999);
nor U23142 (N_23142,N_21202,N_21511);
or U23143 (N_23143,N_21674,N_21947);
xor U23144 (N_23144,N_21601,N_21197);
xnor U23145 (N_23145,N_21513,N_22118);
nand U23146 (N_23146,N_21335,N_22331);
or U23147 (N_23147,N_21872,N_21010);
or U23148 (N_23148,N_21710,N_21672);
nand U23149 (N_23149,N_21958,N_22275);
nand U23150 (N_23150,N_21409,N_21932);
nor U23151 (N_23151,N_21079,N_21767);
nor U23152 (N_23152,N_21360,N_22197);
nand U23153 (N_23153,N_21004,N_21260);
and U23154 (N_23154,N_22436,N_21473);
or U23155 (N_23155,N_22007,N_21775);
nand U23156 (N_23156,N_21514,N_22316);
and U23157 (N_23157,N_22321,N_21926);
or U23158 (N_23158,N_21824,N_21977);
nand U23159 (N_23159,N_21781,N_21559);
or U23160 (N_23160,N_21899,N_21042);
and U23161 (N_23161,N_21481,N_21508);
xor U23162 (N_23162,N_22452,N_21425);
and U23163 (N_23163,N_21213,N_22352);
nor U23164 (N_23164,N_21277,N_22401);
nand U23165 (N_23165,N_22248,N_21022);
nand U23166 (N_23166,N_21594,N_21919);
nand U23167 (N_23167,N_21294,N_21839);
nand U23168 (N_23168,N_21490,N_21677);
xor U23169 (N_23169,N_21426,N_22085);
nor U23170 (N_23170,N_21369,N_22089);
xor U23171 (N_23171,N_22108,N_22262);
or U23172 (N_23172,N_21653,N_21836);
and U23173 (N_23173,N_21740,N_22406);
xnor U23174 (N_23174,N_21223,N_21700);
nor U23175 (N_23175,N_22441,N_21391);
nand U23176 (N_23176,N_21816,N_21889);
xor U23177 (N_23177,N_22322,N_21757);
and U23178 (N_23178,N_22061,N_21037);
xor U23179 (N_23179,N_21881,N_21745);
nor U23180 (N_23180,N_21652,N_21895);
and U23181 (N_23181,N_22146,N_21826);
and U23182 (N_23182,N_21054,N_21670);
and U23183 (N_23183,N_21907,N_21943);
or U23184 (N_23184,N_22429,N_22348);
nor U23185 (N_23185,N_21060,N_22135);
nand U23186 (N_23186,N_21222,N_22459);
nor U23187 (N_23187,N_21266,N_22126);
and U23188 (N_23188,N_22405,N_22391);
or U23189 (N_23189,N_21814,N_22009);
or U23190 (N_23190,N_21784,N_21628);
nor U23191 (N_23191,N_21766,N_21332);
xor U23192 (N_23192,N_21053,N_21058);
nand U23193 (N_23193,N_21690,N_21937);
nand U23194 (N_23194,N_22116,N_21366);
xor U23195 (N_23195,N_21051,N_21008);
and U23196 (N_23196,N_21494,N_21441);
nor U23197 (N_23197,N_21273,N_21780);
nand U23198 (N_23198,N_22488,N_22166);
nand U23199 (N_23199,N_21971,N_21257);
nor U23200 (N_23200,N_21228,N_21207);
or U23201 (N_23201,N_22386,N_22084);
xnor U23202 (N_23202,N_21598,N_22125);
nand U23203 (N_23203,N_22417,N_21113);
or U23204 (N_23204,N_21028,N_21143);
nor U23205 (N_23205,N_21642,N_21329);
and U23206 (N_23206,N_21562,N_22329);
and U23207 (N_23207,N_21887,N_22273);
nand U23208 (N_23208,N_21267,N_21421);
and U23209 (N_23209,N_22229,N_22037);
or U23210 (N_23210,N_21515,N_22065);
nor U23211 (N_23211,N_22493,N_21145);
or U23212 (N_23212,N_21577,N_22464);
or U23213 (N_23213,N_21323,N_21920);
nor U23214 (N_23214,N_21506,N_22456);
and U23215 (N_23215,N_22384,N_21689);
nor U23216 (N_23216,N_21321,N_21851);
nand U23217 (N_23217,N_21105,N_21063);
nor U23218 (N_23218,N_22194,N_21605);
nor U23219 (N_23219,N_22159,N_21886);
or U23220 (N_23220,N_21408,N_21120);
xnor U23221 (N_23221,N_21794,N_22071);
xnor U23222 (N_23222,N_21341,N_22355);
nand U23223 (N_23223,N_21524,N_21688);
xnor U23224 (N_23224,N_21493,N_21007);
nand U23225 (N_23225,N_22465,N_22317);
nor U23226 (N_23226,N_22422,N_21955);
and U23227 (N_23227,N_21585,N_21175);
or U23228 (N_23228,N_22224,N_21463);
nand U23229 (N_23229,N_21014,N_22446);
or U23230 (N_23230,N_22268,N_21209);
xnor U23231 (N_23231,N_21006,N_21258);
nand U23232 (N_23232,N_22000,N_21860);
or U23233 (N_23233,N_21772,N_21930);
nand U23234 (N_23234,N_22083,N_21842);
or U23235 (N_23235,N_22191,N_22318);
xnor U23236 (N_23236,N_21647,N_21589);
nor U23237 (N_23237,N_22072,N_22475);
nor U23238 (N_23238,N_21375,N_21371);
or U23239 (N_23239,N_21432,N_21904);
nor U23240 (N_23240,N_22219,N_21948);
nand U23241 (N_23241,N_22482,N_22281);
and U23242 (N_23242,N_21193,N_22294);
nand U23243 (N_23243,N_22338,N_22344);
nand U23244 (N_23244,N_22451,N_21462);
nor U23245 (N_23245,N_22097,N_21117);
and U23246 (N_23246,N_22110,N_21650);
and U23247 (N_23247,N_21414,N_21623);
nand U23248 (N_23248,N_22140,N_21748);
or U23249 (N_23249,N_21681,N_21020);
xnor U23250 (N_23250,N_21518,N_22166);
or U23251 (N_23251,N_21424,N_21118);
and U23252 (N_23252,N_21059,N_21849);
nand U23253 (N_23253,N_21157,N_21281);
or U23254 (N_23254,N_21836,N_21991);
nor U23255 (N_23255,N_21292,N_22078);
nor U23256 (N_23256,N_21458,N_21108);
nand U23257 (N_23257,N_21985,N_22234);
nand U23258 (N_23258,N_21482,N_21858);
nand U23259 (N_23259,N_21733,N_22338);
nor U23260 (N_23260,N_21907,N_22393);
nand U23261 (N_23261,N_22151,N_21272);
and U23262 (N_23262,N_21770,N_21681);
or U23263 (N_23263,N_21751,N_21362);
nand U23264 (N_23264,N_22110,N_21450);
nand U23265 (N_23265,N_22242,N_21791);
nor U23266 (N_23266,N_21544,N_21238);
or U23267 (N_23267,N_22482,N_22315);
xnor U23268 (N_23268,N_22289,N_22231);
nor U23269 (N_23269,N_21768,N_21684);
xor U23270 (N_23270,N_21710,N_21590);
nand U23271 (N_23271,N_22265,N_21407);
and U23272 (N_23272,N_21679,N_21270);
nor U23273 (N_23273,N_22416,N_21611);
and U23274 (N_23274,N_22092,N_22285);
nand U23275 (N_23275,N_21122,N_22337);
nor U23276 (N_23276,N_22132,N_22236);
xnor U23277 (N_23277,N_22207,N_21551);
nand U23278 (N_23278,N_21670,N_21888);
nor U23279 (N_23279,N_22167,N_21420);
or U23280 (N_23280,N_22028,N_22086);
xor U23281 (N_23281,N_21410,N_22328);
xnor U23282 (N_23282,N_21288,N_21681);
xnor U23283 (N_23283,N_21592,N_21972);
xnor U23284 (N_23284,N_21628,N_21227);
nand U23285 (N_23285,N_21264,N_21909);
nand U23286 (N_23286,N_22074,N_22363);
xnor U23287 (N_23287,N_21944,N_21906);
nor U23288 (N_23288,N_21050,N_21600);
xnor U23289 (N_23289,N_21505,N_22325);
nor U23290 (N_23290,N_22088,N_21856);
and U23291 (N_23291,N_21537,N_22342);
nor U23292 (N_23292,N_21941,N_21658);
nor U23293 (N_23293,N_21897,N_22420);
nor U23294 (N_23294,N_22132,N_21618);
and U23295 (N_23295,N_22195,N_22454);
and U23296 (N_23296,N_21619,N_21180);
xnor U23297 (N_23297,N_22415,N_21792);
nand U23298 (N_23298,N_21688,N_22199);
xor U23299 (N_23299,N_21464,N_21376);
nor U23300 (N_23300,N_22237,N_21801);
nand U23301 (N_23301,N_22280,N_22128);
or U23302 (N_23302,N_22214,N_21145);
and U23303 (N_23303,N_22225,N_21548);
and U23304 (N_23304,N_21561,N_21012);
or U23305 (N_23305,N_22111,N_22316);
nand U23306 (N_23306,N_21223,N_21407);
nand U23307 (N_23307,N_22127,N_21433);
xnor U23308 (N_23308,N_21280,N_21106);
or U23309 (N_23309,N_22425,N_21251);
nor U23310 (N_23310,N_21629,N_21377);
nor U23311 (N_23311,N_21537,N_22353);
nor U23312 (N_23312,N_21832,N_21597);
and U23313 (N_23313,N_22279,N_22118);
xor U23314 (N_23314,N_21830,N_21226);
xnor U23315 (N_23315,N_21330,N_21283);
nand U23316 (N_23316,N_21118,N_21946);
or U23317 (N_23317,N_21103,N_21737);
and U23318 (N_23318,N_21234,N_21005);
nor U23319 (N_23319,N_22499,N_21270);
nor U23320 (N_23320,N_21192,N_21984);
nor U23321 (N_23321,N_21027,N_21467);
nor U23322 (N_23322,N_21488,N_22251);
and U23323 (N_23323,N_21637,N_21144);
nor U23324 (N_23324,N_21953,N_21851);
and U23325 (N_23325,N_22337,N_22089);
and U23326 (N_23326,N_22449,N_22312);
or U23327 (N_23327,N_22281,N_21535);
and U23328 (N_23328,N_22460,N_22117);
nor U23329 (N_23329,N_22478,N_21303);
xnor U23330 (N_23330,N_22453,N_21895);
xor U23331 (N_23331,N_21491,N_22036);
nand U23332 (N_23332,N_21500,N_21248);
xnor U23333 (N_23333,N_22028,N_21540);
xnor U23334 (N_23334,N_22157,N_21030);
and U23335 (N_23335,N_22413,N_21198);
nand U23336 (N_23336,N_21105,N_21908);
or U23337 (N_23337,N_21275,N_22416);
nand U23338 (N_23338,N_22247,N_21182);
nor U23339 (N_23339,N_22006,N_22250);
nor U23340 (N_23340,N_21589,N_22472);
nor U23341 (N_23341,N_21358,N_21459);
xnor U23342 (N_23342,N_21593,N_22375);
nand U23343 (N_23343,N_22168,N_22260);
and U23344 (N_23344,N_21762,N_21196);
nor U23345 (N_23345,N_22248,N_21046);
nor U23346 (N_23346,N_21555,N_21290);
nand U23347 (N_23347,N_21723,N_22224);
or U23348 (N_23348,N_21235,N_21635);
xnor U23349 (N_23349,N_21492,N_21084);
and U23350 (N_23350,N_21499,N_22281);
nand U23351 (N_23351,N_22000,N_21293);
and U23352 (N_23352,N_21337,N_21200);
and U23353 (N_23353,N_21542,N_22418);
nand U23354 (N_23354,N_21049,N_22369);
or U23355 (N_23355,N_22248,N_21023);
xnor U23356 (N_23356,N_21352,N_21651);
xnor U23357 (N_23357,N_21165,N_22293);
and U23358 (N_23358,N_22047,N_21827);
and U23359 (N_23359,N_21416,N_21061);
nand U23360 (N_23360,N_21775,N_21143);
xnor U23361 (N_23361,N_21821,N_21776);
xnor U23362 (N_23362,N_22053,N_21090);
nand U23363 (N_23363,N_22347,N_22434);
and U23364 (N_23364,N_22407,N_21314);
xor U23365 (N_23365,N_21791,N_21404);
or U23366 (N_23366,N_21929,N_21130);
and U23367 (N_23367,N_21450,N_21045);
nand U23368 (N_23368,N_21281,N_22369);
nand U23369 (N_23369,N_21686,N_21882);
or U23370 (N_23370,N_21804,N_21164);
nand U23371 (N_23371,N_21578,N_21932);
nor U23372 (N_23372,N_21272,N_21250);
and U23373 (N_23373,N_21715,N_22255);
and U23374 (N_23374,N_22057,N_21272);
nand U23375 (N_23375,N_22263,N_22092);
or U23376 (N_23376,N_21690,N_22442);
nand U23377 (N_23377,N_21758,N_21757);
xnor U23378 (N_23378,N_22483,N_22344);
nor U23379 (N_23379,N_22217,N_21812);
nand U23380 (N_23380,N_21553,N_22237);
nor U23381 (N_23381,N_21536,N_21114);
nor U23382 (N_23382,N_22436,N_21432);
and U23383 (N_23383,N_21536,N_21977);
nor U23384 (N_23384,N_21399,N_21229);
or U23385 (N_23385,N_21664,N_21322);
xor U23386 (N_23386,N_21248,N_22154);
nand U23387 (N_23387,N_21599,N_22242);
or U23388 (N_23388,N_21247,N_22457);
or U23389 (N_23389,N_22248,N_21747);
and U23390 (N_23390,N_22313,N_22334);
or U23391 (N_23391,N_21220,N_22483);
and U23392 (N_23392,N_22301,N_22076);
and U23393 (N_23393,N_22220,N_22077);
xor U23394 (N_23394,N_22014,N_22078);
nand U23395 (N_23395,N_21505,N_21391);
nor U23396 (N_23396,N_21757,N_22327);
nand U23397 (N_23397,N_21975,N_22453);
nand U23398 (N_23398,N_22441,N_21427);
or U23399 (N_23399,N_21297,N_21047);
xor U23400 (N_23400,N_22406,N_22295);
or U23401 (N_23401,N_21964,N_22257);
xor U23402 (N_23402,N_21891,N_21308);
nand U23403 (N_23403,N_21893,N_22357);
or U23404 (N_23404,N_22161,N_21961);
or U23405 (N_23405,N_22341,N_21549);
xor U23406 (N_23406,N_21821,N_21229);
nor U23407 (N_23407,N_21221,N_21978);
xor U23408 (N_23408,N_22478,N_22369);
xnor U23409 (N_23409,N_22143,N_21860);
nand U23410 (N_23410,N_22340,N_22073);
and U23411 (N_23411,N_21368,N_22221);
nand U23412 (N_23412,N_21124,N_22434);
and U23413 (N_23413,N_21811,N_21824);
or U23414 (N_23414,N_22193,N_21588);
nor U23415 (N_23415,N_22390,N_22101);
or U23416 (N_23416,N_21077,N_22448);
and U23417 (N_23417,N_21481,N_21473);
nand U23418 (N_23418,N_21741,N_21474);
nand U23419 (N_23419,N_22295,N_22009);
and U23420 (N_23420,N_21377,N_22149);
or U23421 (N_23421,N_22488,N_21377);
nor U23422 (N_23422,N_21585,N_21947);
nand U23423 (N_23423,N_21978,N_21517);
nor U23424 (N_23424,N_21320,N_21948);
nand U23425 (N_23425,N_22479,N_22185);
nor U23426 (N_23426,N_22177,N_21389);
nor U23427 (N_23427,N_21586,N_22148);
xnor U23428 (N_23428,N_22469,N_21665);
xnor U23429 (N_23429,N_21479,N_21477);
and U23430 (N_23430,N_21004,N_21441);
or U23431 (N_23431,N_21284,N_21779);
nand U23432 (N_23432,N_21070,N_22255);
or U23433 (N_23433,N_21632,N_22140);
nor U23434 (N_23434,N_21029,N_21255);
nand U23435 (N_23435,N_22017,N_21657);
and U23436 (N_23436,N_21517,N_21401);
nand U23437 (N_23437,N_21203,N_21594);
nor U23438 (N_23438,N_21750,N_22450);
nor U23439 (N_23439,N_21122,N_22195);
nand U23440 (N_23440,N_21650,N_22467);
and U23441 (N_23441,N_21291,N_21829);
xnor U23442 (N_23442,N_21559,N_22276);
or U23443 (N_23443,N_21094,N_21318);
and U23444 (N_23444,N_22194,N_21438);
or U23445 (N_23445,N_22328,N_21134);
and U23446 (N_23446,N_22090,N_21025);
or U23447 (N_23447,N_21558,N_22417);
and U23448 (N_23448,N_21467,N_22172);
nand U23449 (N_23449,N_21028,N_21800);
or U23450 (N_23450,N_21490,N_21634);
or U23451 (N_23451,N_22136,N_21675);
nor U23452 (N_23452,N_21670,N_21826);
nand U23453 (N_23453,N_21375,N_22411);
or U23454 (N_23454,N_21398,N_21272);
nand U23455 (N_23455,N_21065,N_22351);
or U23456 (N_23456,N_21963,N_21396);
xnor U23457 (N_23457,N_21046,N_21538);
or U23458 (N_23458,N_21362,N_22190);
or U23459 (N_23459,N_21199,N_22474);
or U23460 (N_23460,N_21486,N_22455);
xnor U23461 (N_23461,N_21935,N_21430);
xor U23462 (N_23462,N_22118,N_21024);
xor U23463 (N_23463,N_21522,N_21618);
xnor U23464 (N_23464,N_21523,N_21276);
or U23465 (N_23465,N_21624,N_21568);
and U23466 (N_23466,N_21097,N_21576);
xnor U23467 (N_23467,N_21994,N_21357);
and U23468 (N_23468,N_21059,N_22495);
nor U23469 (N_23469,N_22324,N_21977);
xor U23470 (N_23470,N_21293,N_22060);
nor U23471 (N_23471,N_22009,N_21551);
xor U23472 (N_23472,N_22417,N_21781);
or U23473 (N_23473,N_21505,N_21991);
or U23474 (N_23474,N_21628,N_22301);
nor U23475 (N_23475,N_21928,N_22235);
and U23476 (N_23476,N_22496,N_21226);
xor U23477 (N_23477,N_21924,N_22127);
nand U23478 (N_23478,N_22102,N_21858);
or U23479 (N_23479,N_21106,N_22183);
or U23480 (N_23480,N_21521,N_21507);
and U23481 (N_23481,N_21758,N_21802);
xnor U23482 (N_23482,N_21068,N_22202);
nor U23483 (N_23483,N_21571,N_21392);
xnor U23484 (N_23484,N_21809,N_21890);
nor U23485 (N_23485,N_22233,N_21628);
nor U23486 (N_23486,N_21749,N_22024);
xnor U23487 (N_23487,N_21820,N_21971);
and U23488 (N_23488,N_21791,N_21675);
and U23489 (N_23489,N_22411,N_22263);
and U23490 (N_23490,N_21505,N_22170);
nor U23491 (N_23491,N_22335,N_21778);
xnor U23492 (N_23492,N_21262,N_21673);
and U23493 (N_23493,N_21915,N_22415);
xnor U23494 (N_23494,N_21886,N_21008);
nor U23495 (N_23495,N_22025,N_22327);
nand U23496 (N_23496,N_22035,N_21563);
xnor U23497 (N_23497,N_21896,N_21943);
xnor U23498 (N_23498,N_21266,N_22139);
nand U23499 (N_23499,N_21201,N_22223);
and U23500 (N_23500,N_22086,N_22050);
xnor U23501 (N_23501,N_22360,N_21554);
nand U23502 (N_23502,N_21741,N_21650);
and U23503 (N_23503,N_21445,N_21684);
and U23504 (N_23504,N_21304,N_21405);
and U23505 (N_23505,N_21531,N_21487);
or U23506 (N_23506,N_21435,N_22233);
and U23507 (N_23507,N_21257,N_21827);
xnor U23508 (N_23508,N_22483,N_21412);
or U23509 (N_23509,N_21340,N_22424);
nor U23510 (N_23510,N_22161,N_22340);
nand U23511 (N_23511,N_21235,N_21865);
and U23512 (N_23512,N_22499,N_21621);
and U23513 (N_23513,N_22157,N_22414);
nor U23514 (N_23514,N_21235,N_21315);
xor U23515 (N_23515,N_22037,N_21949);
or U23516 (N_23516,N_21968,N_21005);
nand U23517 (N_23517,N_22421,N_22314);
and U23518 (N_23518,N_22096,N_21296);
nand U23519 (N_23519,N_21232,N_22492);
xor U23520 (N_23520,N_21859,N_21796);
and U23521 (N_23521,N_22244,N_21492);
nand U23522 (N_23522,N_21628,N_21497);
xnor U23523 (N_23523,N_22073,N_22488);
nor U23524 (N_23524,N_21454,N_21385);
nor U23525 (N_23525,N_21325,N_22291);
nand U23526 (N_23526,N_21244,N_21473);
and U23527 (N_23527,N_22025,N_21394);
and U23528 (N_23528,N_21787,N_21588);
xor U23529 (N_23529,N_22213,N_21779);
nor U23530 (N_23530,N_21127,N_21572);
nand U23531 (N_23531,N_21490,N_21132);
xnor U23532 (N_23532,N_21113,N_21332);
xor U23533 (N_23533,N_21835,N_22238);
or U23534 (N_23534,N_21242,N_22193);
or U23535 (N_23535,N_21414,N_21037);
xnor U23536 (N_23536,N_21490,N_22323);
nand U23537 (N_23537,N_22445,N_21997);
or U23538 (N_23538,N_22224,N_21376);
or U23539 (N_23539,N_22487,N_21476);
or U23540 (N_23540,N_21323,N_21315);
and U23541 (N_23541,N_21472,N_21465);
xnor U23542 (N_23542,N_21128,N_22472);
and U23543 (N_23543,N_21096,N_21607);
and U23544 (N_23544,N_21121,N_22056);
nand U23545 (N_23545,N_21992,N_21207);
xor U23546 (N_23546,N_22397,N_21244);
xnor U23547 (N_23547,N_21468,N_22059);
or U23548 (N_23548,N_21140,N_22242);
xor U23549 (N_23549,N_21962,N_22194);
nor U23550 (N_23550,N_21836,N_21671);
or U23551 (N_23551,N_21181,N_22319);
and U23552 (N_23552,N_22428,N_22321);
nand U23553 (N_23553,N_21750,N_21252);
or U23554 (N_23554,N_21930,N_21173);
or U23555 (N_23555,N_22438,N_21851);
and U23556 (N_23556,N_21490,N_21570);
xnor U23557 (N_23557,N_21873,N_21427);
or U23558 (N_23558,N_21653,N_22268);
and U23559 (N_23559,N_21778,N_21359);
or U23560 (N_23560,N_22271,N_21106);
nand U23561 (N_23561,N_22172,N_21815);
nor U23562 (N_23562,N_21798,N_22228);
nand U23563 (N_23563,N_22479,N_21619);
or U23564 (N_23564,N_21710,N_22403);
nor U23565 (N_23565,N_22249,N_21323);
xnor U23566 (N_23566,N_21650,N_21807);
nand U23567 (N_23567,N_22287,N_21105);
nor U23568 (N_23568,N_21855,N_21501);
and U23569 (N_23569,N_22083,N_21764);
nand U23570 (N_23570,N_22455,N_21577);
nor U23571 (N_23571,N_22438,N_21335);
or U23572 (N_23572,N_21129,N_21874);
xnor U23573 (N_23573,N_21123,N_22361);
nand U23574 (N_23574,N_22489,N_22174);
nor U23575 (N_23575,N_22105,N_22443);
or U23576 (N_23576,N_21546,N_21198);
nand U23577 (N_23577,N_21391,N_21372);
or U23578 (N_23578,N_21223,N_21404);
nand U23579 (N_23579,N_21217,N_22377);
and U23580 (N_23580,N_21904,N_21654);
or U23581 (N_23581,N_21448,N_22444);
and U23582 (N_23582,N_21321,N_22216);
and U23583 (N_23583,N_21434,N_22057);
or U23584 (N_23584,N_22002,N_21404);
or U23585 (N_23585,N_21887,N_22402);
nor U23586 (N_23586,N_21500,N_21001);
or U23587 (N_23587,N_22032,N_21658);
xor U23588 (N_23588,N_21507,N_21398);
and U23589 (N_23589,N_21626,N_21679);
nor U23590 (N_23590,N_21104,N_21643);
xor U23591 (N_23591,N_22222,N_21910);
or U23592 (N_23592,N_21939,N_21959);
nor U23593 (N_23593,N_22403,N_22038);
nor U23594 (N_23594,N_22016,N_22006);
or U23595 (N_23595,N_21314,N_21517);
and U23596 (N_23596,N_21856,N_21369);
and U23597 (N_23597,N_22415,N_22482);
or U23598 (N_23598,N_22475,N_21871);
nor U23599 (N_23599,N_21380,N_21042);
nor U23600 (N_23600,N_21833,N_21467);
or U23601 (N_23601,N_21690,N_21435);
or U23602 (N_23602,N_21577,N_21597);
and U23603 (N_23603,N_21287,N_21623);
and U23604 (N_23604,N_21665,N_22385);
nand U23605 (N_23605,N_22016,N_21560);
and U23606 (N_23606,N_21251,N_21283);
nand U23607 (N_23607,N_21793,N_21890);
nor U23608 (N_23608,N_21271,N_21741);
or U23609 (N_23609,N_22022,N_21633);
xnor U23610 (N_23610,N_21567,N_21282);
and U23611 (N_23611,N_21598,N_21375);
nor U23612 (N_23612,N_21340,N_22089);
or U23613 (N_23613,N_21513,N_21905);
nand U23614 (N_23614,N_21527,N_22215);
nor U23615 (N_23615,N_22360,N_21852);
or U23616 (N_23616,N_21336,N_21360);
or U23617 (N_23617,N_22429,N_21467);
nor U23618 (N_23618,N_22228,N_21196);
xnor U23619 (N_23619,N_22306,N_21211);
or U23620 (N_23620,N_22336,N_22203);
and U23621 (N_23621,N_22265,N_21640);
and U23622 (N_23622,N_22430,N_22424);
nor U23623 (N_23623,N_21843,N_22184);
nand U23624 (N_23624,N_21623,N_21884);
and U23625 (N_23625,N_21220,N_21279);
or U23626 (N_23626,N_22436,N_21652);
xor U23627 (N_23627,N_21903,N_22215);
or U23628 (N_23628,N_21203,N_21592);
xnor U23629 (N_23629,N_22205,N_22112);
xor U23630 (N_23630,N_22071,N_22076);
or U23631 (N_23631,N_21190,N_21845);
xor U23632 (N_23632,N_22425,N_21126);
or U23633 (N_23633,N_22092,N_22247);
and U23634 (N_23634,N_21786,N_21991);
and U23635 (N_23635,N_22019,N_21364);
and U23636 (N_23636,N_21680,N_22120);
nor U23637 (N_23637,N_21167,N_22334);
nand U23638 (N_23638,N_22258,N_21115);
nand U23639 (N_23639,N_22009,N_21598);
xor U23640 (N_23640,N_21048,N_21062);
nor U23641 (N_23641,N_21814,N_22116);
or U23642 (N_23642,N_21252,N_21768);
nor U23643 (N_23643,N_21804,N_21060);
and U23644 (N_23644,N_22185,N_21548);
nor U23645 (N_23645,N_21972,N_22110);
nor U23646 (N_23646,N_22478,N_21605);
xnor U23647 (N_23647,N_22332,N_21986);
nand U23648 (N_23648,N_21054,N_21400);
nor U23649 (N_23649,N_21763,N_22180);
nor U23650 (N_23650,N_21253,N_22337);
nand U23651 (N_23651,N_21152,N_22090);
and U23652 (N_23652,N_21406,N_22313);
nand U23653 (N_23653,N_21698,N_22136);
and U23654 (N_23654,N_21359,N_21664);
nor U23655 (N_23655,N_21573,N_22398);
and U23656 (N_23656,N_21681,N_22218);
or U23657 (N_23657,N_21310,N_21164);
nand U23658 (N_23658,N_21196,N_22439);
and U23659 (N_23659,N_21589,N_21705);
nor U23660 (N_23660,N_22244,N_22268);
nor U23661 (N_23661,N_21030,N_22384);
nor U23662 (N_23662,N_21932,N_22353);
nor U23663 (N_23663,N_21450,N_22091);
or U23664 (N_23664,N_21150,N_21214);
xnor U23665 (N_23665,N_22447,N_21275);
xnor U23666 (N_23666,N_22092,N_21386);
xor U23667 (N_23667,N_21873,N_22156);
nor U23668 (N_23668,N_21201,N_22062);
and U23669 (N_23669,N_21468,N_21169);
or U23670 (N_23670,N_22368,N_21432);
xnor U23671 (N_23671,N_21887,N_22433);
nor U23672 (N_23672,N_21960,N_21890);
or U23673 (N_23673,N_21043,N_21784);
and U23674 (N_23674,N_22487,N_22388);
and U23675 (N_23675,N_22002,N_22463);
nor U23676 (N_23676,N_22283,N_21440);
xor U23677 (N_23677,N_21908,N_22001);
and U23678 (N_23678,N_21668,N_21552);
nand U23679 (N_23679,N_21422,N_22200);
nand U23680 (N_23680,N_21216,N_22188);
and U23681 (N_23681,N_21822,N_21723);
nand U23682 (N_23682,N_21979,N_21286);
nand U23683 (N_23683,N_22463,N_21349);
nand U23684 (N_23684,N_22195,N_21885);
or U23685 (N_23685,N_21555,N_22240);
and U23686 (N_23686,N_22446,N_21409);
and U23687 (N_23687,N_21781,N_21990);
xor U23688 (N_23688,N_21481,N_22254);
and U23689 (N_23689,N_21528,N_21406);
xor U23690 (N_23690,N_22128,N_21783);
xor U23691 (N_23691,N_21247,N_21098);
nor U23692 (N_23692,N_22196,N_22210);
and U23693 (N_23693,N_22395,N_22078);
nor U23694 (N_23694,N_21929,N_21063);
and U23695 (N_23695,N_21495,N_21437);
nand U23696 (N_23696,N_21393,N_21633);
and U23697 (N_23697,N_21825,N_22462);
and U23698 (N_23698,N_21094,N_21331);
or U23699 (N_23699,N_21557,N_22360);
xnor U23700 (N_23700,N_22453,N_21766);
xnor U23701 (N_23701,N_22040,N_21824);
nand U23702 (N_23702,N_22013,N_21337);
and U23703 (N_23703,N_21656,N_21260);
xnor U23704 (N_23704,N_22157,N_21261);
or U23705 (N_23705,N_22364,N_21333);
or U23706 (N_23706,N_21584,N_21613);
xnor U23707 (N_23707,N_21586,N_22424);
or U23708 (N_23708,N_22496,N_22146);
nor U23709 (N_23709,N_22335,N_21472);
xnor U23710 (N_23710,N_22074,N_22448);
xnor U23711 (N_23711,N_22292,N_22228);
or U23712 (N_23712,N_21001,N_21098);
nand U23713 (N_23713,N_22253,N_21627);
and U23714 (N_23714,N_21938,N_22066);
xor U23715 (N_23715,N_21411,N_22280);
nor U23716 (N_23716,N_22117,N_21425);
and U23717 (N_23717,N_21851,N_21057);
xnor U23718 (N_23718,N_21558,N_21253);
nand U23719 (N_23719,N_21233,N_21799);
or U23720 (N_23720,N_21600,N_22077);
nand U23721 (N_23721,N_21595,N_21071);
nand U23722 (N_23722,N_21184,N_21875);
and U23723 (N_23723,N_21299,N_21714);
nor U23724 (N_23724,N_22366,N_21653);
xor U23725 (N_23725,N_22286,N_22478);
or U23726 (N_23726,N_21121,N_22259);
xnor U23727 (N_23727,N_21380,N_21653);
nor U23728 (N_23728,N_22005,N_21582);
xnor U23729 (N_23729,N_21088,N_21940);
nor U23730 (N_23730,N_21585,N_22175);
xor U23731 (N_23731,N_21017,N_22340);
nor U23732 (N_23732,N_22290,N_21603);
or U23733 (N_23733,N_22441,N_21778);
and U23734 (N_23734,N_21318,N_22162);
or U23735 (N_23735,N_22133,N_22170);
and U23736 (N_23736,N_21183,N_21639);
nand U23737 (N_23737,N_21122,N_21983);
or U23738 (N_23738,N_22378,N_22316);
or U23739 (N_23739,N_22139,N_22080);
nand U23740 (N_23740,N_21556,N_21864);
xor U23741 (N_23741,N_22220,N_21807);
nand U23742 (N_23742,N_21044,N_21107);
nor U23743 (N_23743,N_22114,N_21186);
xor U23744 (N_23744,N_21505,N_21611);
nor U23745 (N_23745,N_21588,N_22269);
and U23746 (N_23746,N_21455,N_22096);
and U23747 (N_23747,N_21077,N_21591);
nor U23748 (N_23748,N_22020,N_21464);
xor U23749 (N_23749,N_21767,N_21666);
nand U23750 (N_23750,N_22308,N_21281);
nand U23751 (N_23751,N_21622,N_22155);
or U23752 (N_23752,N_21895,N_22413);
nor U23753 (N_23753,N_22134,N_21121);
and U23754 (N_23754,N_21205,N_22455);
and U23755 (N_23755,N_21250,N_21411);
or U23756 (N_23756,N_21204,N_21639);
xnor U23757 (N_23757,N_21740,N_21068);
or U23758 (N_23758,N_21847,N_22442);
xnor U23759 (N_23759,N_22464,N_21574);
xor U23760 (N_23760,N_22200,N_21925);
xnor U23761 (N_23761,N_21335,N_22237);
nand U23762 (N_23762,N_21739,N_22225);
xnor U23763 (N_23763,N_21417,N_22491);
nor U23764 (N_23764,N_21315,N_21151);
nor U23765 (N_23765,N_21037,N_22196);
xor U23766 (N_23766,N_21837,N_21076);
xnor U23767 (N_23767,N_21761,N_21697);
and U23768 (N_23768,N_21303,N_21776);
xnor U23769 (N_23769,N_21273,N_21494);
nand U23770 (N_23770,N_21525,N_22325);
or U23771 (N_23771,N_21891,N_21497);
nand U23772 (N_23772,N_22454,N_21234);
nand U23773 (N_23773,N_22112,N_22251);
nor U23774 (N_23774,N_22173,N_21437);
and U23775 (N_23775,N_21974,N_22314);
xnor U23776 (N_23776,N_21562,N_22180);
xor U23777 (N_23777,N_21026,N_21422);
nand U23778 (N_23778,N_22425,N_21045);
and U23779 (N_23779,N_21333,N_22459);
nand U23780 (N_23780,N_22498,N_22066);
xnor U23781 (N_23781,N_22376,N_21348);
nor U23782 (N_23782,N_21892,N_22453);
nand U23783 (N_23783,N_21161,N_21504);
xnor U23784 (N_23784,N_21433,N_21494);
or U23785 (N_23785,N_22247,N_21347);
xor U23786 (N_23786,N_21295,N_21561);
xor U23787 (N_23787,N_22292,N_22208);
or U23788 (N_23788,N_21408,N_22490);
nand U23789 (N_23789,N_21628,N_21464);
and U23790 (N_23790,N_21300,N_21345);
xnor U23791 (N_23791,N_22123,N_21856);
or U23792 (N_23792,N_21858,N_21891);
and U23793 (N_23793,N_21339,N_22405);
xor U23794 (N_23794,N_21167,N_22065);
and U23795 (N_23795,N_22385,N_21874);
or U23796 (N_23796,N_21321,N_21405);
and U23797 (N_23797,N_21590,N_21841);
nand U23798 (N_23798,N_21333,N_21024);
and U23799 (N_23799,N_22089,N_21750);
or U23800 (N_23800,N_21033,N_22300);
and U23801 (N_23801,N_22317,N_21782);
xnor U23802 (N_23802,N_21055,N_21775);
nand U23803 (N_23803,N_22045,N_21257);
nand U23804 (N_23804,N_21664,N_21469);
or U23805 (N_23805,N_22341,N_21215);
nand U23806 (N_23806,N_22157,N_22330);
nor U23807 (N_23807,N_21479,N_21470);
or U23808 (N_23808,N_21396,N_21925);
and U23809 (N_23809,N_22266,N_21419);
nor U23810 (N_23810,N_22191,N_22082);
xor U23811 (N_23811,N_21963,N_21329);
nand U23812 (N_23812,N_21602,N_22277);
nor U23813 (N_23813,N_21816,N_21210);
nor U23814 (N_23814,N_21862,N_21957);
nor U23815 (N_23815,N_22298,N_22412);
or U23816 (N_23816,N_22244,N_22241);
nand U23817 (N_23817,N_22343,N_22359);
nand U23818 (N_23818,N_21304,N_21513);
xor U23819 (N_23819,N_21866,N_21993);
or U23820 (N_23820,N_21504,N_22368);
xor U23821 (N_23821,N_21698,N_21402);
and U23822 (N_23822,N_21314,N_21788);
and U23823 (N_23823,N_21533,N_21226);
nand U23824 (N_23824,N_21608,N_21432);
nand U23825 (N_23825,N_22333,N_22436);
nand U23826 (N_23826,N_22133,N_22141);
xor U23827 (N_23827,N_22031,N_22232);
nor U23828 (N_23828,N_21731,N_21253);
and U23829 (N_23829,N_21402,N_21796);
nand U23830 (N_23830,N_22416,N_22264);
or U23831 (N_23831,N_21946,N_21253);
xnor U23832 (N_23832,N_21700,N_21758);
nand U23833 (N_23833,N_21967,N_21171);
and U23834 (N_23834,N_22043,N_21802);
nor U23835 (N_23835,N_21922,N_22462);
nand U23836 (N_23836,N_22277,N_21202);
xnor U23837 (N_23837,N_22070,N_21243);
or U23838 (N_23838,N_21152,N_22071);
nor U23839 (N_23839,N_21781,N_21709);
or U23840 (N_23840,N_21288,N_21766);
and U23841 (N_23841,N_22085,N_22355);
nor U23842 (N_23842,N_21182,N_22414);
or U23843 (N_23843,N_21803,N_21433);
nand U23844 (N_23844,N_21142,N_21927);
or U23845 (N_23845,N_21676,N_22497);
or U23846 (N_23846,N_21167,N_21713);
or U23847 (N_23847,N_21700,N_21295);
xnor U23848 (N_23848,N_21295,N_21285);
or U23849 (N_23849,N_21258,N_22485);
nor U23850 (N_23850,N_21925,N_21002);
or U23851 (N_23851,N_21693,N_22359);
xnor U23852 (N_23852,N_21897,N_22405);
or U23853 (N_23853,N_21298,N_21200);
and U23854 (N_23854,N_21954,N_21825);
nor U23855 (N_23855,N_21213,N_21591);
nand U23856 (N_23856,N_22330,N_22176);
xor U23857 (N_23857,N_21699,N_21840);
and U23858 (N_23858,N_21734,N_21707);
xnor U23859 (N_23859,N_22314,N_22195);
xor U23860 (N_23860,N_21031,N_21638);
xor U23861 (N_23861,N_22302,N_22191);
or U23862 (N_23862,N_21793,N_21873);
nor U23863 (N_23863,N_21564,N_21771);
or U23864 (N_23864,N_22182,N_21221);
or U23865 (N_23865,N_21437,N_21717);
and U23866 (N_23866,N_21734,N_21685);
or U23867 (N_23867,N_21769,N_22248);
xor U23868 (N_23868,N_21832,N_21613);
nand U23869 (N_23869,N_21105,N_21304);
xor U23870 (N_23870,N_21976,N_22255);
or U23871 (N_23871,N_21839,N_21679);
and U23872 (N_23872,N_21550,N_21288);
nor U23873 (N_23873,N_22236,N_21986);
nand U23874 (N_23874,N_22165,N_22142);
or U23875 (N_23875,N_21526,N_21082);
nand U23876 (N_23876,N_21108,N_22453);
nand U23877 (N_23877,N_21890,N_21990);
and U23878 (N_23878,N_21950,N_21514);
nor U23879 (N_23879,N_21003,N_21994);
xor U23880 (N_23880,N_21383,N_21221);
and U23881 (N_23881,N_22081,N_22226);
or U23882 (N_23882,N_21592,N_21216);
or U23883 (N_23883,N_22081,N_22027);
nand U23884 (N_23884,N_21148,N_21783);
xor U23885 (N_23885,N_21632,N_21319);
nor U23886 (N_23886,N_22199,N_21725);
nand U23887 (N_23887,N_21328,N_21474);
xor U23888 (N_23888,N_21782,N_21120);
or U23889 (N_23889,N_21673,N_22239);
and U23890 (N_23890,N_21259,N_21823);
and U23891 (N_23891,N_21545,N_21961);
xor U23892 (N_23892,N_21674,N_21843);
or U23893 (N_23893,N_21501,N_22472);
xor U23894 (N_23894,N_22335,N_21375);
and U23895 (N_23895,N_21829,N_22417);
nand U23896 (N_23896,N_21806,N_22185);
and U23897 (N_23897,N_21590,N_22367);
nor U23898 (N_23898,N_22310,N_21796);
nand U23899 (N_23899,N_21534,N_21978);
xor U23900 (N_23900,N_21939,N_21592);
nor U23901 (N_23901,N_22023,N_21645);
nor U23902 (N_23902,N_21331,N_21672);
and U23903 (N_23903,N_22239,N_21183);
nand U23904 (N_23904,N_21769,N_21690);
nor U23905 (N_23905,N_21775,N_22062);
xnor U23906 (N_23906,N_21176,N_21499);
or U23907 (N_23907,N_22223,N_21190);
and U23908 (N_23908,N_21902,N_21382);
nand U23909 (N_23909,N_21728,N_21475);
and U23910 (N_23910,N_22280,N_22462);
and U23911 (N_23911,N_21059,N_21595);
and U23912 (N_23912,N_21928,N_21782);
xnor U23913 (N_23913,N_21682,N_21089);
or U23914 (N_23914,N_21278,N_21633);
xor U23915 (N_23915,N_22439,N_21713);
xnor U23916 (N_23916,N_21892,N_22074);
or U23917 (N_23917,N_22353,N_21364);
nor U23918 (N_23918,N_22430,N_21077);
xnor U23919 (N_23919,N_22490,N_22401);
xor U23920 (N_23920,N_21183,N_21423);
or U23921 (N_23921,N_21655,N_21537);
xor U23922 (N_23922,N_21819,N_22083);
and U23923 (N_23923,N_21554,N_21050);
nor U23924 (N_23924,N_22046,N_21988);
or U23925 (N_23925,N_22413,N_21544);
xor U23926 (N_23926,N_22497,N_21901);
nor U23927 (N_23927,N_22416,N_21218);
or U23928 (N_23928,N_22464,N_21796);
xnor U23929 (N_23929,N_21495,N_22124);
xor U23930 (N_23930,N_21192,N_22020);
xnor U23931 (N_23931,N_21451,N_21892);
xnor U23932 (N_23932,N_21917,N_22117);
xnor U23933 (N_23933,N_21543,N_22288);
nand U23934 (N_23934,N_21201,N_22421);
and U23935 (N_23935,N_22231,N_21886);
nand U23936 (N_23936,N_21376,N_21713);
or U23937 (N_23937,N_21965,N_22476);
nor U23938 (N_23938,N_22348,N_21146);
nand U23939 (N_23939,N_21622,N_21560);
or U23940 (N_23940,N_22283,N_21899);
nand U23941 (N_23941,N_21478,N_21290);
nand U23942 (N_23942,N_21059,N_21268);
nor U23943 (N_23943,N_21669,N_21881);
nand U23944 (N_23944,N_21030,N_21950);
nand U23945 (N_23945,N_21643,N_21505);
and U23946 (N_23946,N_21322,N_22299);
or U23947 (N_23947,N_21621,N_22025);
nor U23948 (N_23948,N_22202,N_21198);
nand U23949 (N_23949,N_22209,N_22221);
or U23950 (N_23950,N_21927,N_21594);
or U23951 (N_23951,N_22142,N_21478);
or U23952 (N_23952,N_21847,N_21879);
and U23953 (N_23953,N_22246,N_22400);
nor U23954 (N_23954,N_21433,N_21202);
or U23955 (N_23955,N_21127,N_21365);
or U23956 (N_23956,N_22348,N_21957);
or U23957 (N_23957,N_21161,N_21856);
nor U23958 (N_23958,N_22045,N_22328);
nand U23959 (N_23959,N_21625,N_22107);
nand U23960 (N_23960,N_22231,N_21752);
xor U23961 (N_23961,N_22007,N_21275);
nand U23962 (N_23962,N_21234,N_21282);
or U23963 (N_23963,N_22304,N_22487);
xor U23964 (N_23964,N_21591,N_21571);
or U23965 (N_23965,N_22263,N_21781);
or U23966 (N_23966,N_21114,N_21579);
nor U23967 (N_23967,N_21540,N_21492);
or U23968 (N_23968,N_21479,N_21369);
nor U23969 (N_23969,N_21256,N_21401);
and U23970 (N_23970,N_21698,N_21210);
nor U23971 (N_23971,N_21146,N_22054);
and U23972 (N_23972,N_21004,N_22237);
nand U23973 (N_23973,N_21972,N_21347);
nor U23974 (N_23974,N_22129,N_21209);
and U23975 (N_23975,N_21060,N_21800);
xnor U23976 (N_23976,N_21055,N_21302);
nor U23977 (N_23977,N_21479,N_21376);
or U23978 (N_23978,N_21187,N_22246);
or U23979 (N_23979,N_22412,N_22370);
nor U23980 (N_23980,N_21765,N_21797);
or U23981 (N_23981,N_21490,N_22111);
nor U23982 (N_23982,N_21997,N_21255);
or U23983 (N_23983,N_22406,N_21579);
nor U23984 (N_23984,N_21365,N_21592);
or U23985 (N_23985,N_21425,N_21748);
and U23986 (N_23986,N_21111,N_22448);
or U23987 (N_23987,N_22303,N_22073);
or U23988 (N_23988,N_21920,N_21612);
nor U23989 (N_23989,N_21631,N_22012);
nor U23990 (N_23990,N_21308,N_21184);
or U23991 (N_23991,N_21062,N_21208);
and U23992 (N_23992,N_21873,N_21993);
or U23993 (N_23993,N_22151,N_21450);
nor U23994 (N_23994,N_21781,N_21663);
nand U23995 (N_23995,N_21723,N_21470);
nor U23996 (N_23996,N_22416,N_22279);
nand U23997 (N_23997,N_21398,N_21004);
xnor U23998 (N_23998,N_21401,N_22298);
and U23999 (N_23999,N_21796,N_21229);
nor U24000 (N_24000,N_22513,N_23044);
nor U24001 (N_24001,N_23782,N_23006);
xor U24002 (N_24002,N_23894,N_23027);
nor U24003 (N_24003,N_23973,N_23207);
nand U24004 (N_24004,N_23518,N_22609);
and U24005 (N_24005,N_23665,N_23466);
nor U24006 (N_24006,N_23406,N_23067);
or U24007 (N_24007,N_23639,N_23301);
or U24008 (N_24008,N_22624,N_23328);
nand U24009 (N_24009,N_23033,N_22934);
nand U24010 (N_24010,N_23870,N_22853);
or U24011 (N_24011,N_22715,N_23038);
and U24012 (N_24012,N_22680,N_23151);
or U24013 (N_24013,N_22518,N_22802);
or U24014 (N_24014,N_23650,N_23877);
or U24015 (N_24015,N_22866,N_23380);
xnor U24016 (N_24016,N_22943,N_23949);
nand U24017 (N_24017,N_22597,N_23911);
xnor U24018 (N_24018,N_23991,N_23239);
nor U24019 (N_24019,N_23288,N_23105);
nand U24020 (N_24020,N_23221,N_23429);
xnor U24021 (N_24021,N_23554,N_22595);
xor U24022 (N_24022,N_23420,N_23404);
and U24023 (N_24023,N_22588,N_23193);
nand U24024 (N_24024,N_23267,N_22623);
or U24025 (N_24025,N_22504,N_22817);
xnor U24026 (N_24026,N_23800,N_23352);
nand U24027 (N_24027,N_22948,N_23582);
nor U24028 (N_24028,N_22509,N_22613);
nor U24029 (N_24029,N_23369,N_22511);
nand U24030 (N_24030,N_22995,N_22753);
nor U24031 (N_24031,N_23141,N_23596);
nand U24032 (N_24032,N_22941,N_23290);
xor U24033 (N_24033,N_23892,N_22999);
and U24034 (N_24034,N_23299,N_22861);
nand U24035 (N_24035,N_23179,N_22606);
or U24036 (N_24036,N_23574,N_22694);
xnor U24037 (N_24037,N_23979,N_22614);
nand U24038 (N_24038,N_23543,N_23889);
nor U24039 (N_24039,N_22707,N_23424);
nor U24040 (N_24040,N_23696,N_22702);
or U24041 (N_24041,N_22611,N_23551);
and U24042 (N_24042,N_22988,N_22867);
and U24043 (N_24043,N_23592,N_22528);
or U24044 (N_24044,N_23920,N_22928);
nand U24045 (N_24045,N_23864,N_23212);
nor U24046 (N_24046,N_23855,N_22891);
or U24047 (N_24047,N_23148,N_22785);
or U24048 (N_24048,N_23536,N_22534);
xnor U24049 (N_24049,N_23116,N_23656);
and U24050 (N_24050,N_22514,N_23873);
nor U24051 (N_24051,N_23306,N_23760);
xnor U24052 (N_24052,N_23008,N_23707);
nor U24053 (N_24053,N_23679,N_23575);
xnor U24054 (N_24054,N_23617,N_22655);
nor U24055 (N_24055,N_23059,N_23515);
nand U24056 (N_24056,N_23524,N_23519);
nor U24057 (N_24057,N_23542,N_22505);
xnor U24058 (N_24058,N_22506,N_23478);
nand U24059 (N_24059,N_23337,N_23627);
and U24060 (N_24060,N_23032,N_22769);
nor U24061 (N_24061,N_22798,N_23324);
xnor U24062 (N_24062,N_23609,N_22708);
nor U24063 (N_24063,N_23937,N_22933);
and U24064 (N_24064,N_23928,N_23711);
and U24065 (N_24065,N_23427,N_23130);
nand U24066 (N_24066,N_22578,N_22716);
nor U24067 (N_24067,N_23079,N_23649);
or U24068 (N_24068,N_22766,N_23944);
and U24069 (N_24069,N_23190,N_23001);
or U24070 (N_24070,N_23454,N_22834);
and U24071 (N_24071,N_23635,N_23753);
xor U24072 (N_24072,N_23745,N_23110);
or U24073 (N_24073,N_23368,N_22627);
and U24074 (N_24074,N_23051,N_23218);
and U24075 (N_24075,N_22658,N_22846);
or U24076 (N_24076,N_22590,N_23568);
or U24077 (N_24077,N_22543,N_22758);
xor U24078 (N_24078,N_22521,N_23065);
nand U24079 (N_24079,N_22562,N_23255);
nor U24080 (N_24080,N_22664,N_23828);
nand U24081 (N_24081,N_23233,N_23164);
nor U24082 (N_24082,N_22951,N_23411);
or U24083 (N_24083,N_22987,N_23118);
and U24084 (N_24084,N_22932,N_22912);
xnor U24085 (N_24085,N_23201,N_23675);
nor U24086 (N_24086,N_23765,N_23375);
and U24087 (N_24087,N_23358,N_23175);
and U24088 (N_24088,N_23131,N_23136);
nand U24089 (N_24089,N_23532,N_22923);
nand U24090 (N_24090,N_23271,N_22617);
or U24091 (N_24091,N_23463,N_22974);
or U24092 (N_24092,N_23399,N_23492);
xnor U24093 (N_24093,N_23371,N_23234);
xor U24094 (N_24094,N_23822,N_22653);
and U24095 (N_24095,N_23719,N_23805);
and U24096 (N_24096,N_23419,N_22845);
nand U24097 (N_24097,N_23715,N_22537);
and U24098 (N_24098,N_22529,N_23260);
or U24099 (N_24099,N_23157,N_23872);
nand U24100 (N_24100,N_22795,N_23876);
xnor U24101 (N_24101,N_23701,N_23529);
or U24102 (N_24102,N_23899,N_22952);
nor U24103 (N_24103,N_23184,N_23390);
xor U24104 (N_24104,N_22905,N_23614);
nand U24105 (N_24105,N_23977,N_23552);
and U24106 (N_24106,N_23332,N_23245);
nor U24107 (N_24107,N_23476,N_23112);
and U24108 (N_24108,N_23169,N_23113);
xor U24109 (N_24109,N_23790,N_23231);
xnor U24110 (N_24110,N_23158,N_23653);
nor U24111 (N_24111,N_22575,N_23327);
nand U24112 (N_24112,N_22790,N_23600);
and U24113 (N_24113,N_23392,N_23633);
nor U24114 (N_24114,N_23481,N_22636);
nor U24115 (N_24115,N_23243,N_22897);
xnor U24116 (N_24116,N_22742,N_23764);
nor U24117 (N_24117,N_22593,N_23615);
and U24118 (N_24118,N_23263,N_23229);
nor U24119 (N_24119,N_23439,N_23559);
nand U24120 (N_24120,N_23452,N_23202);
and U24121 (N_24121,N_22589,N_23710);
xor U24122 (N_24122,N_23663,N_23171);
xnor U24123 (N_24123,N_23475,N_23856);
or U24124 (N_24124,N_22657,N_23250);
or U24125 (N_24125,N_22647,N_23569);
xor U24126 (N_24126,N_23848,N_23739);
or U24127 (N_24127,N_23793,N_22997);
nand U24128 (N_24128,N_22993,N_23882);
nor U24129 (N_24129,N_22972,N_23030);
or U24130 (N_24130,N_23692,N_23416);
nand U24131 (N_24131,N_23785,N_23311);
nor U24132 (N_24132,N_23125,N_23833);
or U24133 (N_24133,N_23520,N_23900);
xnor U24134 (N_24134,N_22918,N_23858);
nand U24135 (N_24135,N_23637,N_23455);
nor U24136 (N_24136,N_23350,N_22726);
nor U24137 (N_24137,N_23266,N_23984);
and U24138 (N_24138,N_23940,N_23581);
or U24139 (N_24139,N_23598,N_23382);
nor U24140 (N_24140,N_23082,N_23990);
nand U24141 (N_24141,N_22962,N_23307);
and U24142 (N_24142,N_23486,N_22629);
and U24143 (N_24143,N_22644,N_22828);
nand U24144 (N_24144,N_23694,N_23850);
xnor U24145 (N_24145,N_22904,N_23909);
nor U24146 (N_24146,N_23196,N_23448);
and U24147 (N_24147,N_23143,N_23908);
and U24148 (N_24148,N_22773,N_22699);
or U24149 (N_24149,N_23160,N_22931);
or U24150 (N_24150,N_22677,N_22901);
and U24151 (N_24151,N_23109,N_23622);
nand U24152 (N_24152,N_23686,N_23537);
nand U24153 (N_24153,N_22556,N_23487);
xor U24154 (N_24154,N_23535,N_22568);
xnor U24155 (N_24155,N_23323,N_23604);
xnor U24156 (N_24156,N_23253,N_23946);
or U24157 (N_24157,N_23036,N_23840);
nand U24158 (N_24158,N_22823,N_23821);
or U24159 (N_24159,N_23497,N_22605);
nand U24160 (N_24160,N_22973,N_23014);
nand U24161 (N_24161,N_23544,N_22608);
or U24162 (N_24162,N_23192,N_23580);
or U24163 (N_24163,N_23797,N_23688);
xnor U24164 (N_24164,N_23421,N_23781);
and U24165 (N_24165,N_23145,N_23733);
nand U24166 (N_24166,N_23824,N_23993);
or U24167 (N_24167,N_23312,N_22814);
or U24168 (N_24168,N_22693,N_23447);
or U24169 (N_24169,N_22807,N_22775);
or U24170 (N_24170,N_22570,N_23618);
and U24171 (N_24171,N_23256,N_23669);
and U24172 (N_24172,N_23778,N_22711);
nor U24173 (N_24173,N_22776,N_22573);
nor U24174 (N_24174,N_22820,N_23227);
and U24175 (N_24175,N_23788,N_22607);
and U24176 (N_24176,N_22908,N_23727);
or U24177 (N_24177,N_23837,N_23071);
or U24178 (N_24178,N_22851,N_23697);
and U24179 (N_24179,N_22937,N_22531);
and U24180 (N_24180,N_23225,N_23285);
or U24181 (N_24181,N_22586,N_22651);
and U24182 (N_24182,N_23440,N_23005);
xor U24183 (N_24183,N_23534,N_23444);
xnor U24184 (N_24184,N_23589,N_22947);
xor U24185 (N_24185,N_23955,N_22888);
xor U24186 (N_24186,N_23560,N_23351);
and U24187 (N_24187,N_23539,N_22770);
nor U24188 (N_24188,N_22811,N_23664);
xnor U24189 (N_24189,N_23122,N_23367);
nand U24190 (N_24190,N_22688,N_23956);
and U24191 (N_24191,N_22880,N_22641);
xor U24192 (N_24192,N_23803,N_23259);
nand U24193 (N_24193,N_23015,N_23579);
nand U24194 (N_24194,N_22519,N_22686);
and U24195 (N_24195,N_23340,N_23279);
xnor U24196 (N_24196,N_23771,N_23417);
xnor U24197 (N_24197,N_23126,N_23593);
or U24198 (N_24198,N_23249,N_22836);
nand U24199 (N_24199,N_23372,N_23210);
nor U24200 (N_24200,N_23456,N_23641);
xor U24201 (N_24201,N_22864,N_22990);
nor U24202 (N_24202,N_23680,N_23528);
nor U24203 (N_24203,N_23905,N_23446);
nor U24204 (N_24204,N_23523,N_23791);
and U24205 (N_24205,N_22965,N_23182);
xor U24206 (N_24206,N_22782,N_22916);
or U24207 (N_24207,N_23985,N_23017);
or U24208 (N_24208,N_22610,N_23055);
nor U24209 (N_24209,N_23572,N_22767);
nor U24210 (N_24210,N_22876,N_23296);
nand U24211 (N_24211,N_23999,N_23019);
nor U24212 (N_24212,N_23326,N_22849);
nand U24213 (N_24213,N_22789,N_23146);
or U24214 (N_24214,N_23414,N_23120);
nand U24215 (N_24215,N_23741,N_22522);
and U24216 (N_24216,N_23975,N_22827);
xor U24217 (N_24217,N_23860,N_22929);
and U24218 (N_24218,N_23499,N_23976);
xor U24219 (N_24219,N_23718,N_23958);
and U24220 (N_24220,N_22963,N_22899);
and U24221 (N_24221,N_23320,N_22700);
xor U24222 (N_24222,N_23964,N_23401);
and U24223 (N_24223,N_23366,N_22879);
and U24224 (N_24224,N_23965,N_23935);
or U24225 (N_24225,N_22895,N_23672);
xnor U24226 (N_24226,N_22865,N_23457);
and U24227 (N_24227,N_23379,N_23823);
nor U24228 (N_24228,N_22554,N_22631);
or U24229 (N_24229,N_23759,N_23098);
xor U24230 (N_24230,N_23652,N_23398);
nand U24231 (N_24231,N_23226,N_23303);
nor U24232 (N_24232,N_22885,N_22724);
nor U24233 (N_24233,N_22920,N_23467);
xor U24234 (N_24234,N_22924,N_23244);
nor U24235 (N_24235,N_23462,N_22898);
nand U24236 (N_24236,N_23220,N_23517);
and U24237 (N_24237,N_23359,N_23809);
and U24238 (N_24238,N_23717,N_22546);
and U24239 (N_24239,N_23738,N_23121);
nor U24240 (N_24240,N_22630,N_23063);
xnor U24241 (N_24241,N_22757,N_23504);
nand U24242 (N_24242,N_22825,N_23338);
and U24243 (N_24243,N_22859,N_23590);
xnor U24244 (N_24244,N_23029,N_23509);
nor U24245 (N_24245,N_22591,N_23871);
xor U24246 (N_24246,N_23325,N_22921);
nor U24247 (N_24247,N_22640,N_22894);
or U24248 (N_24248,N_22740,N_23838);
nor U24249 (N_24249,N_22500,N_22696);
nor U24250 (N_24250,N_23177,N_23625);
xnor U24251 (N_24251,N_22954,N_23655);
nor U24252 (N_24252,N_23150,N_23400);
xnor U24253 (N_24253,N_23674,N_23117);
and U24254 (N_24254,N_23932,N_22750);
and U24255 (N_24255,N_23153,N_23774);
or U24256 (N_24256,N_23996,N_23732);
xnor U24257 (N_24257,N_23770,N_22541);
and U24258 (N_24258,N_23197,N_23992);
nand U24259 (N_24259,N_23995,N_23951);
and U24260 (N_24260,N_22552,N_23237);
nand U24261 (N_24261,N_23070,N_22930);
xor U24262 (N_24262,N_23489,N_23431);
or U24263 (N_24263,N_23853,N_23751);
or U24264 (N_24264,N_23407,N_22792);
and U24265 (N_24265,N_23041,N_23094);
and U24266 (N_24266,N_22991,N_23302);
nor U24267 (N_24267,N_23780,N_22854);
nand U24268 (N_24268,N_23654,N_23018);
or U24269 (N_24269,N_23450,N_22871);
xor U24270 (N_24270,N_23361,N_23072);
nand U24271 (N_24271,N_22893,N_23045);
or U24272 (N_24272,N_23410,N_23247);
nor U24273 (N_24273,N_23586,N_23658);
xor U24274 (N_24274,N_23470,N_23695);
nand U24275 (N_24275,N_22622,N_22890);
nand U24276 (N_24276,N_23962,N_22542);
nor U24277 (N_24277,N_23046,N_23315);
and U24278 (N_24278,N_23709,N_23159);
and U24279 (N_24279,N_23630,N_23346);
xnor U24280 (N_24280,N_23083,N_22682);
xnor U24281 (N_24281,N_23383,N_23743);
nand U24282 (N_24282,N_23628,N_23161);
or U24283 (N_24283,N_22752,N_23128);
xor U24284 (N_24284,N_23566,N_22667);
and U24285 (N_24285,N_23522,N_23754);
nand U24286 (N_24286,N_22720,N_23847);
nor U24287 (N_24287,N_22967,N_23510);
nor U24288 (N_24288,N_23773,N_23806);
nor U24289 (N_24289,N_23123,N_23127);
nand U24290 (N_24290,N_23902,N_23835);
xor U24291 (N_24291,N_23960,N_22668);
or U24292 (N_24292,N_23648,N_23074);
and U24293 (N_24293,N_23099,N_22709);
and U24294 (N_24294,N_22692,N_22584);
nand U24295 (N_24295,N_23031,N_22783);
xor U24296 (N_24296,N_22632,N_23211);
nand U24297 (N_24297,N_22927,N_22648);
or U24298 (N_24298,N_23729,N_23353);
nand U24299 (N_24299,N_23103,N_22502);
or U24300 (N_24300,N_23493,N_22978);
or U24301 (N_24301,N_22594,N_23096);
and U24302 (N_24302,N_23297,N_23135);
nor U24303 (N_24303,N_23168,N_22882);
or U24304 (N_24304,N_23613,N_23119);
nor U24305 (N_24305,N_23483,N_22875);
nand U24306 (N_24306,N_23139,N_23418);
xnor U24307 (N_24307,N_23198,N_23922);
xnor U24308 (N_24308,N_23629,N_23336);
nand U24309 (N_24309,N_22723,N_22793);
nor U24310 (N_24310,N_23181,N_23740);
nor U24311 (N_24311,N_23278,N_23827);
nand U24312 (N_24312,N_23563,N_23144);
nor U24313 (N_24313,N_22571,N_23154);
nor U24314 (N_24314,N_22903,N_23721);
or U24315 (N_24315,N_23624,N_22714);
nand U24316 (N_24316,N_22966,N_23849);
or U24317 (N_24317,N_23281,N_23115);
or U24318 (N_24318,N_23028,N_22877);
nand U24319 (N_24319,N_23485,N_23636);
or U24320 (N_24320,N_23265,N_23866);
nor U24321 (N_24321,N_23091,N_23742);
and U24322 (N_24322,N_23792,N_23762);
and U24323 (N_24323,N_22910,N_23339);
nor U24324 (N_24324,N_22683,N_23508);
and U24325 (N_24325,N_22695,N_23562);
or U24326 (N_24326,N_22549,N_22544);
xor U24327 (N_24327,N_23310,N_22992);
or U24328 (N_24328,N_22772,N_23107);
nor U24329 (N_24329,N_23907,N_22887);
and U24330 (N_24330,N_22957,N_22625);
and U24331 (N_24331,N_23651,N_23254);
xnor U24332 (N_24332,N_23062,N_23132);
or U24333 (N_24333,N_23034,N_23086);
xnor U24334 (N_24334,N_22520,N_22751);
nor U24335 (N_24335,N_23183,N_22955);
nand U24336 (N_24336,N_22970,N_22730);
nand U24337 (N_24337,N_22652,N_23076);
nor U24338 (N_24338,N_23820,N_22975);
nor U24339 (N_24339,N_22710,N_23747);
or U24340 (N_24340,N_23058,N_22998);
nor U24341 (N_24341,N_22733,N_23378);
and U24342 (N_24342,N_23989,N_23166);
xnor U24343 (N_24343,N_22717,N_23966);
xor U24344 (N_24344,N_22796,N_22778);
nand U24345 (N_24345,N_23623,N_23722);
or U24346 (N_24346,N_22583,N_23863);
nand U24347 (N_24347,N_22684,N_22691);
xnor U24348 (N_24348,N_23769,N_23341);
nand U24349 (N_24349,N_23830,N_22536);
and U24350 (N_24350,N_23961,N_23587);
and U24351 (N_24351,N_23318,N_23564);
nand U24352 (N_24352,N_23904,N_22949);
xnor U24353 (N_24353,N_23251,N_23538);
nor U24354 (N_24354,N_23356,N_23605);
nor U24355 (N_24355,N_23084,N_23607);
nor U24356 (N_24356,N_23268,N_23316);
xor U24357 (N_24357,N_23917,N_22813);
nand U24358 (N_24358,N_22925,N_22615);
nand U24359 (N_24359,N_23437,N_22585);
nor U24360 (N_24360,N_22603,N_22808);
nand U24361 (N_24361,N_23736,N_23802);
or U24362 (N_24362,N_23496,N_23474);
nor U24363 (N_24363,N_22681,N_22824);
nor U24364 (N_24364,N_23248,N_22739);
and U24365 (N_24365,N_23801,N_23477);
and U24366 (N_24366,N_22831,N_22777);
nand U24367 (N_24367,N_22548,N_22780);
nand U24368 (N_24368,N_23918,N_22671);
and U24369 (N_24369,N_23408,N_23329);
and U24370 (N_24370,N_22958,N_23322);
xor U24371 (N_24371,N_22806,N_23494);
or U24372 (N_24372,N_23173,N_23436);
nor U24373 (N_24373,N_23502,N_23608);
or U24374 (N_24374,N_22977,N_23362);
xnor U24375 (N_24375,N_23576,N_23728);
nor U24376 (N_24376,N_23472,N_22530);
or U24377 (N_24377,N_23354,N_22968);
nor U24378 (N_24378,N_22857,N_22563);
or U24379 (N_24379,N_23595,N_22960);
or U24380 (N_24380,N_23947,N_23545);
xnor U24381 (N_24381,N_23730,N_23195);
nand U24382 (N_24382,N_23807,N_22832);
nand U24383 (N_24383,N_23152,N_23591);
nand U24384 (N_24384,N_23787,N_23088);
xnor U24385 (N_24385,N_23203,N_23355);
and U24386 (N_24386,N_23673,N_23693);
or U24387 (N_24387,N_23578,N_23540);
or U24388 (N_24388,N_22939,N_23364);
nor U24389 (N_24389,N_22889,N_22633);
and U24390 (N_24390,N_23558,N_22983);
xnor U24391 (N_24391,N_23441,N_23689);
and U24392 (N_24392,N_22580,N_22819);
nand U24393 (N_24393,N_23512,N_23621);
xnor U24394 (N_24394,N_23426,N_22533);
nand U24395 (N_24395,N_23343,N_23388);
and U24396 (N_24396,N_22674,N_23262);
nor U24397 (N_24397,N_23897,N_23443);
or U24398 (N_24398,N_23766,N_23808);
or U24399 (N_24399,N_23926,N_23189);
or U24400 (N_24400,N_23744,N_23549);
nand U24401 (N_24401,N_23165,N_22940);
nor U24402 (N_24402,N_23987,N_22713);
nor U24403 (N_24403,N_23373,N_22618);
nand U24404 (N_24404,N_22566,N_23895);
nand U24405 (N_24405,N_23829,N_23703);
xnor U24406 (N_24406,N_23402,N_23013);
nand U24407 (N_24407,N_23068,N_22612);
and U24408 (N_24408,N_23075,N_23464);
xnor U24409 (N_24409,N_22848,N_23000);
xnor U24410 (N_24410,N_23217,N_23513);
xnor U24411 (N_24411,N_23969,N_22516);
nor U24412 (N_24412,N_22768,N_23397);
nor U24413 (N_24413,N_23757,N_23186);
and U24414 (N_24414,N_23616,N_23490);
xnor U24415 (N_24415,N_22736,N_22656);
nor U24416 (N_24416,N_22560,N_23415);
xor U24417 (N_24417,N_23138,N_22804);
or U24418 (N_24418,N_22994,N_23097);
and U24419 (N_24419,N_23938,N_22685);
and U24420 (N_24420,N_22917,N_23275);
or U24421 (N_24421,N_23887,N_23445);
and U24422 (N_24422,N_23980,N_22964);
and U24423 (N_24423,N_23395,N_23533);
xnor U24424 (N_24424,N_22732,N_23915);
nand U24425 (N_24425,N_23242,N_23276);
and U24426 (N_24426,N_23804,N_22659);
xnor U24427 (N_24427,N_23691,N_22666);
or U24428 (N_24428,N_22749,N_23662);
and U24429 (N_24429,N_22689,N_23610);
nor U24430 (N_24430,N_23929,N_23022);
or U24431 (N_24431,N_23698,N_22805);
nand U24432 (N_24432,N_22762,N_23298);
nor U24433 (N_24433,N_22950,N_22788);
nor U24434 (N_24434,N_23933,N_23885);
or U24435 (N_24435,N_23571,N_23706);
or U24436 (N_24436,N_22971,N_22621);
xor U24437 (N_24437,N_23293,N_23156);
nand U24438 (N_24438,N_22855,N_23054);
or U24439 (N_24439,N_22914,N_22555);
nor U24440 (N_24440,N_23026,N_23205);
nor U24441 (N_24441,N_23289,N_23002);
nand U24442 (N_24442,N_23111,N_23037);
and U24443 (N_24443,N_23035,N_23606);
and U24444 (N_24444,N_23137,N_23506);
and U24445 (N_24445,N_22579,N_23064);
or U24446 (N_24446,N_23516,N_23039);
or U24447 (N_24447,N_22592,N_23347);
nor U24448 (N_24448,N_23982,N_23069);
nand U24449 (N_24449,N_23550,N_23547);
and U24450 (N_24450,N_22996,N_23716);
and U24451 (N_24451,N_23684,N_23188);
nor U24452 (N_24452,N_22842,N_23216);
and U24453 (N_24453,N_23313,N_23178);
nor U24454 (N_24454,N_22645,N_22512);
nor U24455 (N_24455,N_22705,N_23632);
nand U24456 (N_24456,N_23602,N_23875);
nand U24457 (N_24457,N_23282,N_23482);
nor U24458 (N_24458,N_23425,N_23505);
nor U24459 (N_24459,N_23387,N_22639);
and U24460 (N_24460,N_22665,N_23816);
nand U24461 (N_24461,N_23775,N_23913);
or U24462 (N_24462,N_22547,N_23546);
xor U24463 (N_24463,N_23057,N_23232);
or U24464 (N_24464,N_22794,N_23700);
nor U24465 (N_24465,N_22673,N_23106);
nor U24466 (N_24466,N_23852,N_22669);
or U24467 (N_24467,N_22856,N_22746);
and U24468 (N_24468,N_23836,N_23163);
and U24469 (N_24469,N_23270,N_23396);
or U24470 (N_24470,N_23024,N_23501);
nor U24471 (N_24471,N_23588,N_23720);
nand U24472 (N_24472,N_23080,N_22507);
xnor U24473 (N_24473,N_23174,N_23647);
and U24474 (N_24474,N_23772,N_23952);
and U24475 (N_24475,N_22900,N_23428);
nor U24476 (N_24476,N_22718,N_23180);
and U24477 (N_24477,N_22569,N_23142);
or U24478 (N_24478,N_22862,N_23573);
xnor U24479 (N_24479,N_23294,N_23868);
nand U24480 (N_24480,N_23813,N_22582);
or U24481 (N_24481,N_22508,N_23553);
xor U24482 (N_24482,N_23594,N_23500);
nor U24483 (N_24483,N_23898,N_22654);
xor U24484 (N_24484,N_23213,N_22872);
or U24485 (N_24485,N_23468,N_23129);
nand U24486 (N_24486,N_23789,N_23235);
and U24487 (N_24487,N_23831,N_23677);
nor U24488 (N_24488,N_23794,N_22599);
and U24489 (N_24489,N_23040,N_23678);
and U24490 (N_24490,N_23660,N_22841);
and U24491 (N_24491,N_23862,N_23705);
nor U24492 (N_24492,N_23643,N_22837);
or U24493 (N_24493,N_23810,N_23950);
nor U24494 (N_24494,N_23768,N_23095);
nor U24495 (N_24495,N_23971,N_23839);
xnor U24496 (N_24496,N_22719,N_23053);
xnor U24497 (N_24497,N_22911,N_23758);
nor U24498 (N_24498,N_23983,N_23304);
or U24499 (N_24499,N_23555,N_22833);
nand U24500 (N_24500,N_22881,N_23611);
or U24501 (N_24501,N_23584,N_23884);
nand U24502 (N_24502,N_23712,N_23878);
and U24503 (N_24503,N_22809,N_23011);
or U24504 (N_24504,N_23393,N_22517);
xor U24505 (N_24505,N_23597,N_22576);
and U24506 (N_24506,N_22902,N_22858);
and U24507 (N_24507,N_22884,N_23305);
and U24508 (N_24508,N_23089,N_23846);
xnor U24509 (N_24509,N_23147,N_23974);
or U24510 (N_24510,N_23585,N_22906);
and U24511 (N_24511,N_23252,N_23893);
xor U24512 (N_24512,N_23469,N_23646);
and U24513 (N_24513,N_23345,N_23682);
or U24514 (N_24514,N_23066,N_23104);
nand U24515 (N_24515,N_22701,N_22706);
and U24516 (N_24516,N_23430,N_23735);
nand U24517 (N_24517,N_23314,N_23713);
nand U24518 (N_24518,N_23459,N_23458);
xnor U24519 (N_24519,N_22524,N_23090);
and U24520 (N_24520,N_23357,N_23896);
nand U24521 (N_24521,N_23943,N_22821);
or U24522 (N_24522,N_23185,N_22734);
and U24523 (N_24523,N_22634,N_23619);
xnor U24524 (N_24524,N_23814,N_22527);
nor U24525 (N_24525,N_22852,N_22878);
nand U24526 (N_24526,N_22553,N_22635);
nor U24527 (N_24527,N_22926,N_22735);
xnor U24528 (N_24528,N_22535,N_23377);
or U24529 (N_24529,N_22907,N_23704);
nor U24530 (N_24530,N_23725,N_23799);
xor U24531 (N_24531,N_23230,N_22729);
or U24532 (N_24532,N_22815,N_22596);
or U24533 (N_24533,N_22860,N_23060);
and U24534 (N_24534,N_23925,N_23642);
xor U24535 (N_24535,N_23708,N_23087);
nand U24536 (N_24536,N_23498,N_23527);
or U24537 (N_24537,N_22979,N_22747);
and U24538 (N_24538,N_22980,N_23321);
nor U24539 (N_24539,N_23981,N_22938);
nand U24540 (N_24540,N_22587,N_23737);
nand U24541 (N_24541,N_22675,N_23200);
and U24542 (N_24542,N_23300,N_23016);
nor U24543 (N_24543,N_22679,N_22743);
xor U24544 (N_24544,N_23859,N_23204);
nor U24545 (N_24545,N_22915,N_22863);
or U24546 (N_24546,N_23910,N_23565);
nand U24547 (N_24547,N_23162,N_23687);
nor U24548 (N_24548,N_22501,N_23330);
nor U24549 (N_24549,N_23124,N_23874);
nand U24550 (N_24550,N_23280,N_22619);
nand U24551 (N_24551,N_23879,N_23284);
nand U24552 (N_24552,N_23025,N_23503);
nand U24553 (N_24553,N_23049,N_22830);
nor U24554 (N_24554,N_23750,N_22942);
or U24555 (N_24555,N_23890,N_23507);
and U24556 (N_24556,N_23967,N_23746);
nand U24557 (N_24557,N_22661,N_22558);
or U24558 (N_24558,N_22799,N_23667);
nand U24559 (N_24559,N_23714,N_23435);
and U24560 (N_24560,N_23644,N_23851);
or U24561 (N_24561,N_23078,N_23783);
xnor U24562 (N_24562,N_22985,N_23577);
xor U24563 (N_24563,N_22909,N_23798);
xnor U24564 (N_24564,N_22800,N_22976);
or U24565 (N_24565,N_23567,N_22981);
nor U24566 (N_24566,N_22919,N_22526);
xnor U24567 (N_24567,N_23349,N_22839);
nand U24568 (N_24568,N_23634,N_23434);
xor U24569 (N_24569,N_22755,N_22989);
nand U24570 (N_24570,N_22779,N_23761);
nand U24571 (N_24571,N_23945,N_22601);
or U24572 (N_24572,N_23342,N_23077);
nor U24573 (N_24573,N_23906,N_23149);
nand U24574 (N_24574,N_23335,N_22670);
and U24575 (N_24575,N_23948,N_23228);
or U24576 (N_24576,N_22628,N_23842);
nor U24577 (N_24577,N_22810,N_22759);
nor U24578 (N_24578,N_22602,N_23003);
nand U24579 (N_24579,N_23010,N_23274);
xnor U24580 (N_24580,N_23924,N_23108);
nand U24581 (N_24581,N_22774,N_23370);
nand U24582 (N_24582,N_23914,N_23214);
and U24583 (N_24583,N_23867,N_23394);
and U24584 (N_24584,N_23755,N_23385);
nand U24585 (N_24585,N_23681,N_22761);
or U24586 (N_24586,N_23916,N_23360);
and U24587 (N_24587,N_23854,N_23432);
nor U24588 (N_24588,N_22731,N_22797);
xnor U24589 (N_24589,N_22760,N_22984);
and U24590 (N_24590,N_23391,N_22784);
xor U24591 (N_24591,N_23936,N_23986);
nor U24592 (N_24592,N_23191,N_23841);
nor U24593 (N_24593,N_22886,N_23348);
and U24594 (N_24594,N_23570,N_23363);
nor U24595 (N_24595,N_22868,N_23812);
nand U24596 (N_24596,N_23796,N_23959);
nand U24597 (N_24597,N_23881,N_22559);
and U24598 (N_24598,N_23333,N_22835);
xor U24599 (N_24599,N_23903,N_23480);
or U24600 (N_24600,N_22944,N_22703);
nand U24601 (N_24601,N_22650,N_23521);
and U24602 (N_24602,N_23007,N_23413);
or U24603 (N_24603,N_23042,N_23626);
nand U24604 (N_24604,N_22748,N_23645);
nand U24605 (N_24605,N_22626,N_23465);
or U24606 (N_24606,N_23433,N_23931);
and U24607 (N_24607,N_22922,N_22786);
nor U24608 (N_24608,N_23557,N_23224);
xnor U24609 (N_24609,N_22791,N_23638);
nor U24610 (N_24610,N_22873,N_22616);
xnor U24611 (N_24611,N_23081,N_23389);
nand U24612 (N_24612,N_23934,N_22812);
nand U24613 (N_24613,N_23548,N_23919);
nor U24614 (N_24614,N_23939,N_23319);
nor U24615 (N_24615,N_22620,N_22803);
or U24616 (N_24616,N_23292,N_23530);
and U24617 (N_24617,N_23670,N_23777);
or U24618 (N_24618,N_23923,N_23222);
xnor U24619 (N_24619,N_23927,N_22764);
or U24620 (N_24620,N_23100,N_23998);
nor U24621 (N_24621,N_23690,N_22540);
nor U24622 (N_24622,N_23258,N_23246);
xnor U24623 (N_24623,N_23886,N_23666);
or U24624 (N_24624,N_22662,N_23269);
xor U24625 (N_24625,N_22869,N_22801);
nor U24626 (N_24626,N_22572,N_23009);
nand U24627 (N_24627,N_22577,N_23880);
xnor U24628 (N_24628,N_23047,N_22539);
and U24629 (N_24629,N_23734,N_22765);
nor U24630 (N_24630,N_22642,N_22676);
and U24631 (N_24631,N_22956,N_22523);
and U24632 (N_24632,N_22687,N_23187);
nor U24633 (N_24633,N_23381,N_23779);
nand U24634 (N_24634,N_22874,N_23376);
xnor U24635 (N_24635,N_23056,N_23818);
nor U24636 (N_24636,N_23451,N_22704);
nand U24637 (N_24637,N_23826,N_23215);
or U24638 (N_24638,N_23723,N_23620);
nor U24639 (N_24639,N_23921,N_23172);
nand U24640 (N_24640,N_22896,N_23219);
and U24641 (N_24641,N_22525,N_23073);
and U24642 (N_24642,N_22870,N_23048);
nand U24643 (N_24643,N_22561,N_23331);
nand U24644 (N_24644,N_23724,N_22600);
nor U24645 (N_24645,N_22532,N_23277);
nor U24646 (N_24646,N_22646,N_22557);
nor U24647 (N_24647,N_23978,N_22959);
nor U24648 (N_24648,N_23957,N_23726);
nand U24649 (N_24649,N_22781,N_23685);
nor U24650 (N_24650,N_22678,N_23473);
xnor U24651 (N_24651,N_23795,N_23287);
nor U24652 (N_24652,N_23832,N_23261);
xnor U24653 (N_24653,N_22844,N_22754);
nor U24654 (N_24654,N_23861,N_23968);
or U24655 (N_24655,N_22551,N_23170);
and U24656 (N_24656,N_23374,N_23988);
nor U24657 (N_24657,N_22745,N_23264);
nor U24658 (N_24658,N_22721,N_23479);
and U24659 (N_24659,N_22840,N_23869);
and U24660 (N_24660,N_23786,N_23941);
and U24661 (N_24661,N_23291,N_23963);
or U24662 (N_24662,N_23453,N_23155);
and U24663 (N_24663,N_23334,N_23901);
nor U24664 (N_24664,N_23811,N_23023);
or U24665 (N_24665,N_23206,N_22567);
and U24666 (N_24666,N_22604,N_22672);
xnor U24667 (N_24667,N_23384,N_22986);
and U24668 (N_24668,N_23683,N_23114);
xnor U24669 (N_24669,N_23972,N_23857);
xor U24670 (N_24670,N_23460,N_22936);
and U24671 (N_24671,N_23238,N_23541);
nand U24672 (N_24672,N_23661,N_23912);
or U24673 (N_24673,N_23133,N_22538);
nor U24674 (N_24674,N_23043,N_23756);
or U24675 (N_24675,N_23843,N_23930);
nor U24676 (N_24676,N_23449,N_22953);
or U24677 (N_24677,N_23484,N_23514);
and U24678 (N_24678,N_22961,N_23488);
nor U24679 (N_24679,N_22838,N_22763);
xnor U24680 (N_24680,N_22637,N_23491);
or U24681 (N_24681,N_23599,N_22565);
xnor U24682 (N_24682,N_23140,N_23819);
nor U24683 (N_24683,N_23405,N_23776);
and U24684 (N_24684,N_22850,N_23612);
or U24685 (N_24685,N_22737,N_23659);
nor U24686 (N_24686,N_22756,N_23583);
nor U24687 (N_24687,N_22787,N_23767);
nor U24688 (N_24688,N_23561,N_23702);
and U24689 (N_24689,N_23601,N_23194);
or U24690 (N_24690,N_23241,N_22550);
nand U24691 (N_24691,N_23236,N_22829);
and U24692 (N_24692,N_22728,N_23495);
or U24693 (N_24693,N_23442,N_23208);
xnor U24694 (N_24694,N_23556,N_23749);
nand U24695 (N_24695,N_23511,N_23942);
or U24696 (N_24696,N_22741,N_23748);
or U24697 (N_24697,N_22722,N_23526);
nor U24698 (N_24698,N_23344,N_22945);
and U24699 (N_24699,N_23020,N_23994);
xnor U24700 (N_24700,N_23422,N_22818);
nor U24701 (N_24701,N_23752,N_23052);
nand U24702 (N_24702,N_23295,N_22510);
or U24703 (N_24703,N_23438,N_23815);
nand U24704 (N_24704,N_22698,N_23531);
xor U24705 (N_24705,N_23092,N_22946);
nor U24706 (N_24706,N_23403,N_23257);
nand U24707 (N_24707,N_23223,N_22913);
and U24708 (N_24708,N_22515,N_23883);
nor U24709 (N_24709,N_23845,N_22744);
xnor U24710 (N_24710,N_23525,N_22545);
and U24711 (N_24711,N_23101,N_23834);
xnor U24712 (N_24712,N_23308,N_23102);
and U24713 (N_24713,N_23412,N_22690);
xnor U24714 (N_24714,N_22503,N_22816);
xnor U24715 (N_24715,N_22660,N_23409);
nor U24716 (N_24716,N_23004,N_23970);
xor U24717 (N_24717,N_23386,N_23423);
nor U24718 (N_24718,N_23365,N_23784);
and U24719 (N_24719,N_23657,N_23668);
and U24720 (N_24720,N_23093,N_23640);
nand U24721 (N_24721,N_22892,N_23061);
nor U24722 (N_24722,N_23461,N_23676);
and U24723 (N_24723,N_23309,N_22847);
nand U24724 (N_24724,N_23085,N_23603);
nor U24725 (N_24725,N_23731,N_23272);
xnor U24726 (N_24726,N_23167,N_22574);
xnor U24727 (N_24727,N_23209,N_23273);
and U24728 (N_24728,N_22727,N_22663);
or U24729 (N_24729,N_23888,N_23176);
xnor U24730 (N_24730,N_23997,N_23021);
nand U24731 (N_24731,N_22883,N_23240);
nand U24732 (N_24732,N_23471,N_23286);
nor U24733 (N_24733,N_22826,N_23953);
and U24734 (N_24734,N_22697,N_22643);
nor U24735 (N_24735,N_22771,N_23817);
nand U24736 (N_24736,N_22935,N_23865);
nor U24737 (N_24737,N_22822,N_22598);
xor U24738 (N_24738,N_23699,N_22969);
nand U24739 (N_24739,N_23012,N_22712);
or U24740 (N_24740,N_22843,N_22982);
nor U24741 (N_24741,N_23199,N_23763);
nor U24742 (N_24742,N_23671,N_23631);
or U24743 (N_24743,N_23825,N_23050);
nand U24744 (N_24744,N_22649,N_23283);
nand U24745 (N_24745,N_23134,N_22738);
nor U24746 (N_24746,N_23844,N_23317);
nand U24747 (N_24747,N_22638,N_23891);
nor U24748 (N_24748,N_22581,N_22725);
and U24749 (N_24749,N_22564,N_23954);
nand U24750 (N_24750,N_23541,N_23065);
xnor U24751 (N_24751,N_23202,N_23034);
xnor U24752 (N_24752,N_23415,N_22535);
nand U24753 (N_24753,N_23082,N_23795);
and U24754 (N_24754,N_23896,N_23973);
nand U24755 (N_24755,N_22706,N_22577);
nand U24756 (N_24756,N_23802,N_23168);
xnor U24757 (N_24757,N_22694,N_22582);
and U24758 (N_24758,N_23274,N_23115);
nand U24759 (N_24759,N_23868,N_23030);
xor U24760 (N_24760,N_22873,N_23775);
and U24761 (N_24761,N_23393,N_23595);
nor U24762 (N_24762,N_23198,N_22809);
or U24763 (N_24763,N_23116,N_23734);
xnor U24764 (N_24764,N_23513,N_23318);
nor U24765 (N_24765,N_23267,N_23349);
xor U24766 (N_24766,N_23601,N_23831);
or U24767 (N_24767,N_23342,N_23088);
or U24768 (N_24768,N_22509,N_23086);
xnor U24769 (N_24769,N_22558,N_23715);
or U24770 (N_24770,N_22709,N_23592);
xor U24771 (N_24771,N_22936,N_23556);
xor U24772 (N_24772,N_23889,N_23863);
and U24773 (N_24773,N_22548,N_23252);
nand U24774 (N_24774,N_23304,N_23280);
xnor U24775 (N_24775,N_22730,N_23580);
nor U24776 (N_24776,N_22768,N_23837);
or U24777 (N_24777,N_22747,N_23091);
xnor U24778 (N_24778,N_23520,N_23909);
nand U24779 (N_24779,N_22551,N_23096);
nor U24780 (N_24780,N_23238,N_22659);
and U24781 (N_24781,N_23533,N_23444);
nor U24782 (N_24782,N_22749,N_23003);
or U24783 (N_24783,N_23377,N_23548);
nor U24784 (N_24784,N_23164,N_23417);
xor U24785 (N_24785,N_22759,N_22580);
nor U24786 (N_24786,N_22563,N_22842);
or U24787 (N_24787,N_23366,N_23510);
or U24788 (N_24788,N_23322,N_22544);
nor U24789 (N_24789,N_23426,N_23314);
nor U24790 (N_24790,N_22574,N_23077);
and U24791 (N_24791,N_23682,N_23033);
nand U24792 (N_24792,N_23014,N_23235);
or U24793 (N_24793,N_23187,N_23914);
and U24794 (N_24794,N_23306,N_22618);
and U24795 (N_24795,N_22657,N_23411);
xor U24796 (N_24796,N_23556,N_23175);
or U24797 (N_24797,N_23138,N_23159);
nor U24798 (N_24798,N_23267,N_22606);
or U24799 (N_24799,N_23482,N_22668);
nand U24800 (N_24800,N_23960,N_23398);
or U24801 (N_24801,N_22516,N_23606);
nor U24802 (N_24802,N_23793,N_23112);
and U24803 (N_24803,N_23041,N_22834);
and U24804 (N_24804,N_23940,N_23528);
xnor U24805 (N_24805,N_23196,N_23296);
or U24806 (N_24806,N_22547,N_23751);
or U24807 (N_24807,N_23865,N_23201);
xor U24808 (N_24808,N_23997,N_23080);
nor U24809 (N_24809,N_22955,N_23539);
or U24810 (N_24810,N_22721,N_23079);
nand U24811 (N_24811,N_22927,N_22696);
and U24812 (N_24812,N_23804,N_22950);
nand U24813 (N_24813,N_23424,N_22858);
nor U24814 (N_24814,N_23300,N_23330);
and U24815 (N_24815,N_22720,N_23563);
or U24816 (N_24816,N_22878,N_23917);
or U24817 (N_24817,N_22668,N_23244);
or U24818 (N_24818,N_23896,N_22900);
or U24819 (N_24819,N_23403,N_22551);
and U24820 (N_24820,N_23238,N_23149);
nor U24821 (N_24821,N_22974,N_22978);
and U24822 (N_24822,N_23860,N_23025);
xor U24823 (N_24823,N_22832,N_23182);
or U24824 (N_24824,N_23875,N_23435);
and U24825 (N_24825,N_23419,N_23646);
and U24826 (N_24826,N_22841,N_23497);
nand U24827 (N_24827,N_23321,N_23210);
and U24828 (N_24828,N_23861,N_23571);
xnor U24829 (N_24829,N_23635,N_23990);
nor U24830 (N_24830,N_23140,N_23126);
and U24831 (N_24831,N_23956,N_23269);
nor U24832 (N_24832,N_22646,N_22664);
nand U24833 (N_24833,N_22857,N_22551);
nand U24834 (N_24834,N_22951,N_22736);
and U24835 (N_24835,N_23815,N_22520);
nor U24836 (N_24836,N_23084,N_22905);
nand U24837 (N_24837,N_23101,N_23343);
nand U24838 (N_24838,N_22760,N_23197);
or U24839 (N_24839,N_23206,N_23424);
nand U24840 (N_24840,N_23167,N_22799);
xor U24841 (N_24841,N_23951,N_23912);
or U24842 (N_24842,N_23274,N_22615);
and U24843 (N_24843,N_23082,N_23835);
nor U24844 (N_24844,N_22913,N_23965);
or U24845 (N_24845,N_22803,N_23438);
and U24846 (N_24846,N_23543,N_23520);
nand U24847 (N_24847,N_23515,N_23372);
or U24848 (N_24848,N_23738,N_23650);
or U24849 (N_24849,N_23014,N_23813);
nand U24850 (N_24850,N_23414,N_23010);
nor U24851 (N_24851,N_23514,N_22690);
or U24852 (N_24852,N_22637,N_23631);
or U24853 (N_24853,N_23674,N_23684);
xor U24854 (N_24854,N_22629,N_23285);
and U24855 (N_24855,N_23681,N_22774);
nor U24856 (N_24856,N_23041,N_23228);
xnor U24857 (N_24857,N_23355,N_23460);
nor U24858 (N_24858,N_23498,N_23048);
xor U24859 (N_24859,N_22954,N_23713);
or U24860 (N_24860,N_23270,N_23422);
nor U24861 (N_24861,N_23640,N_22624);
nor U24862 (N_24862,N_23616,N_22854);
nor U24863 (N_24863,N_22811,N_23283);
nor U24864 (N_24864,N_23100,N_23936);
nand U24865 (N_24865,N_23596,N_23844);
nor U24866 (N_24866,N_23405,N_22680);
nand U24867 (N_24867,N_22620,N_22813);
or U24868 (N_24868,N_23650,N_23923);
xor U24869 (N_24869,N_23091,N_22643);
xnor U24870 (N_24870,N_23958,N_22528);
xor U24871 (N_24871,N_23135,N_23310);
or U24872 (N_24872,N_23915,N_23213);
nor U24873 (N_24873,N_23125,N_22957);
nor U24874 (N_24874,N_23263,N_23308);
or U24875 (N_24875,N_23962,N_22565);
nand U24876 (N_24876,N_23433,N_23038);
and U24877 (N_24877,N_23668,N_23914);
xor U24878 (N_24878,N_23212,N_22508);
nand U24879 (N_24879,N_23477,N_23698);
nor U24880 (N_24880,N_23767,N_23800);
or U24881 (N_24881,N_23601,N_23739);
or U24882 (N_24882,N_22704,N_22683);
nor U24883 (N_24883,N_23016,N_23455);
nand U24884 (N_24884,N_23031,N_23812);
xor U24885 (N_24885,N_22770,N_23367);
xnor U24886 (N_24886,N_23733,N_22895);
and U24887 (N_24887,N_23645,N_23147);
nand U24888 (N_24888,N_23788,N_22582);
xnor U24889 (N_24889,N_22666,N_22727);
nand U24890 (N_24890,N_22764,N_23881);
xor U24891 (N_24891,N_23191,N_22944);
nand U24892 (N_24892,N_23956,N_22681);
and U24893 (N_24893,N_23954,N_22858);
xor U24894 (N_24894,N_22749,N_23066);
nor U24895 (N_24895,N_23352,N_22881);
or U24896 (N_24896,N_23883,N_22802);
xnor U24897 (N_24897,N_23914,N_23722);
or U24898 (N_24898,N_22582,N_22832);
xor U24899 (N_24899,N_22602,N_23145);
xor U24900 (N_24900,N_22669,N_23201);
nor U24901 (N_24901,N_23024,N_23922);
or U24902 (N_24902,N_22660,N_23497);
nor U24903 (N_24903,N_22832,N_22741);
or U24904 (N_24904,N_23817,N_23603);
nor U24905 (N_24905,N_23010,N_23520);
nand U24906 (N_24906,N_23706,N_22810);
xnor U24907 (N_24907,N_22569,N_23694);
or U24908 (N_24908,N_23582,N_23426);
nor U24909 (N_24909,N_23209,N_22703);
nand U24910 (N_24910,N_23582,N_23863);
and U24911 (N_24911,N_23144,N_23033);
nand U24912 (N_24912,N_23303,N_23569);
and U24913 (N_24913,N_22643,N_23709);
or U24914 (N_24914,N_23657,N_22718);
and U24915 (N_24915,N_22758,N_23255);
nand U24916 (N_24916,N_22811,N_22554);
xor U24917 (N_24917,N_23894,N_22673);
nand U24918 (N_24918,N_23881,N_22740);
nand U24919 (N_24919,N_23135,N_23545);
nand U24920 (N_24920,N_23064,N_23712);
nand U24921 (N_24921,N_23674,N_22664);
and U24922 (N_24922,N_23016,N_22930);
or U24923 (N_24923,N_23931,N_23026);
nor U24924 (N_24924,N_23688,N_22914);
and U24925 (N_24925,N_23257,N_23123);
or U24926 (N_24926,N_23426,N_22930);
or U24927 (N_24927,N_23074,N_22785);
nand U24928 (N_24928,N_23427,N_23577);
xor U24929 (N_24929,N_23051,N_22549);
xor U24930 (N_24930,N_23826,N_23271);
xor U24931 (N_24931,N_22772,N_23518);
or U24932 (N_24932,N_22796,N_23155);
xor U24933 (N_24933,N_23234,N_22719);
and U24934 (N_24934,N_23333,N_23206);
xnor U24935 (N_24935,N_23428,N_23691);
xor U24936 (N_24936,N_23428,N_22714);
nand U24937 (N_24937,N_23494,N_23551);
nor U24938 (N_24938,N_23105,N_22617);
or U24939 (N_24939,N_23805,N_23941);
nand U24940 (N_24940,N_23490,N_22753);
xor U24941 (N_24941,N_22649,N_23034);
and U24942 (N_24942,N_23598,N_23292);
and U24943 (N_24943,N_22670,N_23995);
xor U24944 (N_24944,N_22862,N_23565);
and U24945 (N_24945,N_22585,N_23397);
xnor U24946 (N_24946,N_22678,N_22946);
and U24947 (N_24947,N_23294,N_22514);
nor U24948 (N_24948,N_22631,N_23301);
and U24949 (N_24949,N_23287,N_23741);
nor U24950 (N_24950,N_23985,N_23386);
xor U24951 (N_24951,N_22708,N_23820);
xor U24952 (N_24952,N_23375,N_23130);
xnor U24953 (N_24953,N_23258,N_23406);
xnor U24954 (N_24954,N_23375,N_23588);
nor U24955 (N_24955,N_23494,N_23092);
and U24956 (N_24956,N_23730,N_23313);
or U24957 (N_24957,N_23919,N_23758);
xnor U24958 (N_24958,N_22613,N_23218);
nand U24959 (N_24959,N_23335,N_22632);
and U24960 (N_24960,N_23932,N_23361);
or U24961 (N_24961,N_23634,N_23911);
xnor U24962 (N_24962,N_23977,N_23008);
or U24963 (N_24963,N_23299,N_23609);
nand U24964 (N_24964,N_22971,N_23582);
nand U24965 (N_24965,N_23360,N_23888);
or U24966 (N_24966,N_23902,N_23969);
nor U24967 (N_24967,N_23046,N_23438);
xnor U24968 (N_24968,N_22775,N_23583);
or U24969 (N_24969,N_23390,N_23078);
nor U24970 (N_24970,N_23725,N_22895);
and U24971 (N_24971,N_23756,N_23410);
nor U24972 (N_24972,N_23200,N_23927);
xnor U24973 (N_24973,N_23245,N_23907);
and U24974 (N_24974,N_23866,N_23205);
xnor U24975 (N_24975,N_23815,N_23773);
nand U24976 (N_24976,N_23545,N_22909);
nor U24977 (N_24977,N_22857,N_22824);
nand U24978 (N_24978,N_23590,N_23860);
xnor U24979 (N_24979,N_22942,N_23809);
xor U24980 (N_24980,N_23269,N_23077);
xor U24981 (N_24981,N_22925,N_22834);
or U24982 (N_24982,N_22621,N_23018);
nand U24983 (N_24983,N_23285,N_23230);
nor U24984 (N_24984,N_23660,N_23924);
xor U24985 (N_24985,N_23427,N_23736);
xor U24986 (N_24986,N_23786,N_22834);
and U24987 (N_24987,N_23319,N_22789);
or U24988 (N_24988,N_23527,N_23946);
xnor U24989 (N_24989,N_23451,N_23982);
nor U24990 (N_24990,N_23723,N_22575);
and U24991 (N_24991,N_23795,N_23919);
nor U24992 (N_24992,N_23004,N_23331);
and U24993 (N_24993,N_23799,N_23997);
nand U24994 (N_24994,N_22692,N_22940);
nor U24995 (N_24995,N_23658,N_23212);
or U24996 (N_24996,N_22876,N_22947);
or U24997 (N_24997,N_22841,N_23043);
xnor U24998 (N_24998,N_23035,N_22610);
nor U24999 (N_24999,N_23587,N_23151);
nor U25000 (N_25000,N_22551,N_22678);
and U25001 (N_25001,N_23477,N_23404);
and U25002 (N_25002,N_22614,N_22701);
or U25003 (N_25003,N_23814,N_23472);
xnor U25004 (N_25004,N_23885,N_23690);
nor U25005 (N_25005,N_22878,N_22583);
nor U25006 (N_25006,N_22970,N_23645);
xnor U25007 (N_25007,N_22934,N_22659);
nand U25008 (N_25008,N_22778,N_23343);
nor U25009 (N_25009,N_23722,N_22574);
nand U25010 (N_25010,N_23247,N_23089);
and U25011 (N_25011,N_22580,N_23149);
nand U25012 (N_25012,N_23594,N_22864);
and U25013 (N_25013,N_23161,N_23022);
xor U25014 (N_25014,N_23422,N_22523);
and U25015 (N_25015,N_23368,N_22990);
nor U25016 (N_25016,N_22916,N_23320);
or U25017 (N_25017,N_23188,N_23128);
xor U25018 (N_25018,N_22878,N_22510);
and U25019 (N_25019,N_22506,N_22747);
nand U25020 (N_25020,N_23778,N_22787);
or U25021 (N_25021,N_22870,N_23523);
xnor U25022 (N_25022,N_23930,N_23871);
or U25023 (N_25023,N_22794,N_23043);
nor U25024 (N_25024,N_22963,N_23370);
nor U25025 (N_25025,N_23744,N_22599);
and U25026 (N_25026,N_23090,N_23449);
and U25027 (N_25027,N_22686,N_23018);
xor U25028 (N_25028,N_22742,N_22570);
and U25029 (N_25029,N_23309,N_23052);
or U25030 (N_25030,N_23076,N_23159);
or U25031 (N_25031,N_22501,N_22841);
nor U25032 (N_25032,N_22729,N_23404);
xor U25033 (N_25033,N_23157,N_23732);
and U25034 (N_25034,N_23501,N_23386);
or U25035 (N_25035,N_23566,N_23816);
xnor U25036 (N_25036,N_23938,N_23869);
and U25037 (N_25037,N_23213,N_23615);
xnor U25038 (N_25038,N_23645,N_23952);
xor U25039 (N_25039,N_23705,N_22951);
nand U25040 (N_25040,N_22853,N_23462);
nand U25041 (N_25041,N_22808,N_23828);
xnor U25042 (N_25042,N_22816,N_22502);
xnor U25043 (N_25043,N_23277,N_23418);
nand U25044 (N_25044,N_22561,N_23778);
nand U25045 (N_25045,N_22869,N_22854);
nor U25046 (N_25046,N_23490,N_23680);
nor U25047 (N_25047,N_23008,N_23100);
xnor U25048 (N_25048,N_23026,N_23071);
nor U25049 (N_25049,N_23085,N_23436);
and U25050 (N_25050,N_22628,N_23060);
xnor U25051 (N_25051,N_22571,N_23420);
nand U25052 (N_25052,N_23531,N_22552);
nand U25053 (N_25053,N_22583,N_23635);
nor U25054 (N_25054,N_22507,N_23890);
xnor U25055 (N_25055,N_23292,N_23063);
nor U25056 (N_25056,N_23570,N_22916);
or U25057 (N_25057,N_23849,N_23999);
nor U25058 (N_25058,N_23028,N_22919);
nor U25059 (N_25059,N_22554,N_23296);
and U25060 (N_25060,N_23276,N_22806);
or U25061 (N_25061,N_23644,N_23195);
nand U25062 (N_25062,N_22755,N_23435);
or U25063 (N_25063,N_23821,N_23165);
xor U25064 (N_25064,N_23640,N_23787);
nand U25065 (N_25065,N_23046,N_22567);
nand U25066 (N_25066,N_22619,N_23745);
nand U25067 (N_25067,N_23312,N_22824);
and U25068 (N_25068,N_23702,N_22566);
xor U25069 (N_25069,N_23862,N_23658);
xor U25070 (N_25070,N_23159,N_23010);
xor U25071 (N_25071,N_22846,N_23602);
xor U25072 (N_25072,N_23451,N_23840);
or U25073 (N_25073,N_23611,N_22734);
xnor U25074 (N_25074,N_23988,N_23928);
xor U25075 (N_25075,N_23497,N_22924);
xor U25076 (N_25076,N_23822,N_22899);
nand U25077 (N_25077,N_22869,N_22953);
or U25078 (N_25078,N_23402,N_23917);
nor U25079 (N_25079,N_23748,N_23266);
or U25080 (N_25080,N_23229,N_23775);
xor U25081 (N_25081,N_23924,N_23689);
or U25082 (N_25082,N_23539,N_23059);
and U25083 (N_25083,N_23616,N_23243);
nand U25084 (N_25084,N_23407,N_22561);
or U25085 (N_25085,N_23594,N_23532);
or U25086 (N_25086,N_22592,N_23466);
xor U25087 (N_25087,N_23374,N_23054);
nor U25088 (N_25088,N_23656,N_23583);
nand U25089 (N_25089,N_23444,N_22608);
or U25090 (N_25090,N_22750,N_22875);
nand U25091 (N_25091,N_23007,N_22902);
and U25092 (N_25092,N_23770,N_23929);
nor U25093 (N_25093,N_22875,N_23812);
or U25094 (N_25094,N_23540,N_23773);
nand U25095 (N_25095,N_23606,N_23412);
nand U25096 (N_25096,N_23673,N_22732);
or U25097 (N_25097,N_23634,N_22505);
nor U25098 (N_25098,N_22971,N_22781);
or U25099 (N_25099,N_23105,N_23277);
nor U25100 (N_25100,N_23702,N_23698);
xnor U25101 (N_25101,N_23917,N_22513);
xnor U25102 (N_25102,N_23471,N_22708);
or U25103 (N_25103,N_23690,N_23948);
nand U25104 (N_25104,N_23223,N_23444);
nor U25105 (N_25105,N_23589,N_22836);
or U25106 (N_25106,N_23538,N_23298);
or U25107 (N_25107,N_23275,N_23408);
xnor U25108 (N_25108,N_23789,N_23446);
xor U25109 (N_25109,N_23102,N_23725);
nand U25110 (N_25110,N_23372,N_23646);
xnor U25111 (N_25111,N_23557,N_23764);
nor U25112 (N_25112,N_23244,N_23061);
xnor U25113 (N_25113,N_23923,N_23106);
nor U25114 (N_25114,N_23474,N_23352);
or U25115 (N_25115,N_23703,N_22808);
and U25116 (N_25116,N_22665,N_23963);
or U25117 (N_25117,N_22800,N_23404);
xor U25118 (N_25118,N_23000,N_22943);
xnor U25119 (N_25119,N_23419,N_23881);
nand U25120 (N_25120,N_23348,N_22757);
nand U25121 (N_25121,N_23339,N_22869);
xnor U25122 (N_25122,N_22898,N_22826);
and U25123 (N_25123,N_22634,N_23709);
xnor U25124 (N_25124,N_22988,N_23131);
or U25125 (N_25125,N_23630,N_23132);
nand U25126 (N_25126,N_23325,N_22524);
xor U25127 (N_25127,N_23303,N_22936);
or U25128 (N_25128,N_23709,N_23639);
nand U25129 (N_25129,N_22806,N_23946);
nor U25130 (N_25130,N_22869,N_23197);
xor U25131 (N_25131,N_22989,N_23156);
nand U25132 (N_25132,N_23060,N_23538);
xnor U25133 (N_25133,N_22946,N_23466);
or U25134 (N_25134,N_22956,N_23522);
nand U25135 (N_25135,N_23366,N_23165);
nor U25136 (N_25136,N_22952,N_23803);
nor U25137 (N_25137,N_22843,N_23470);
and U25138 (N_25138,N_23836,N_22945);
and U25139 (N_25139,N_22694,N_23239);
nand U25140 (N_25140,N_23868,N_23307);
or U25141 (N_25141,N_23119,N_23267);
nor U25142 (N_25142,N_22775,N_23232);
or U25143 (N_25143,N_23331,N_23187);
or U25144 (N_25144,N_23721,N_22645);
nor U25145 (N_25145,N_23831,N_23504);
nor U25146 (N_25146,N_22722,N_23264);
xor U25147 (N_25147,N_22638,N_23866);
or U25148 (N_25148,N_23835,N_22996);
nor U25149 (N_25149,N_23665,N_22819);
nor U25150 (N_25150,N_22648,N_23173);
and U25151 (N_25151,N_22938,N_22996);
or U25152 (N_25152,N_23788,N_23885);
nor U25153 (N_25153,N_23252,N_22957);
xnor U25154 (N_25154,N_23445,N_22822);
and U25155 (N_25155,N_22661,N_22562);
nor U25156 (N_25156,N_22913,N_23805);
nand U25157 (N_25157,N_23153,N_23377);
xor U25158 (N_25158,N_22642,N_22952);
nand U25159 (N_25159,N_23532,N_23749);
xor U25160 (N_25160,N_23722,N_23519);
and U25161 (N_25161,N_22643,N_23190);
and U25162 (N_25162,N_23017,N_22663);
and U25163 (N_25163,N_23683,N_23557);
or U25164 (N_25164,N_23287,N_23909);
or U25165 (N_25165,N_23833,N_23715);
and U25166 (N_25166,N_22825,N_23736);
or U25167 (N_25167,N_23689,N_22537);
nor U25168 (N_25168,N_23207,N_22723);
or U25169 (N_25169,N_23587,N_23101);
or U25170 (N_25170,N_22886,N_22628);
and U25171 (N_25171,N_22634,N_22563);
xor U25172 (N_25172,N_23059,N_23895);
xor U25173 (N_25173,N_23806,N_23259);
xor U25174 (N_25174,N_23441,N_23921);
nand U25175 (N_25175,N_23063,N_23529);
nand U25176 (N_25176,N_22581,N_23598);
and U25177 (N_25177,N_22799,N_23673);
nand U25178 (N_25178,N_23929,N_23987);
and U25179 (N_25179,N_23989,N_22904);
nor U25180 (N_25180,N_23745,N_22556);
nor U25181 (N_25181,N_22597,N_22530);
nand U25182 (N_25182,N_22699,N_22635);
or U25183 (N_25183,N_22574,N_22693);
and U25184 (N_25184,N_22940,N_23087);
or U25185 (N_25185,N_23336,N_23900);
nor U25186 (N_25186,N_23822,N_22784);
nor U25187 (N_25187,N_23360,N_23643);
xnor U25188 (N_25188,N_23938,N_23086);
or U25189 (N_25189,N_23373,N_23914);
nor U25190 (N_25190,N_23652,N_22878);
nor U25191 (N_25191,N_23539,N_23906);
nand U25192 (N_25192,N_23987,N_23863);
and U25193 (N_25193,N_23582,N_23724);
xor U25194 (N_25194,N_23206,N_22658);
and U25195 (N_25195,N_23536,N_23921);
nor U25196 (N_25196,N_23749,N_23621);
and U25197 (N_25197,N_23619,N_23720);
or U25198 (N_25198,N_23670,N_22695);
nor U25199 (N_25199,N_23731,N_23063);
nand U25200 (N_25200,N_23558,N_22543);
nor U25201 (N_25201,N_22759,N_23440);
xnor U25202 (N_25202,N_23712,N_22944);
xor U25203 (N_25203,N_22540,N_22772);
nand U25204 (N_25204,N_23749,N_23302);
nor U25205 (N_25205,N_23628,N_23457);
xnor U25206 (N_25206,N_22593,N_22997);
nand U25207 (N_25207,N_23312,N_23754);
xnor U25208 (N_25208,N_23177,N_22800);
or U25209 (N_25209,N_23794,N_23233);
and U25210 (N_25210,N_23899,N_23472);
nor U25211 (N_25211,N_23429,N_23200);
xnor U25212 (N_25212,N_22513,N_23371);
xnor U25213 (N_25213,N_23903,N_23111);
nor U25214 (N_25214,N_23186,N_22728);
nand U25215 (N_25215,N_22711,N_22878);
and U25216 (N_25216,N_22867,N_22576);
or U25217 (N_25217,N_23730,N_23727);
or U25218 (N_25218,N_23116,N_22629);
and U25219 (N_25219,N_22787,N_23003);
nand U25220 (N_25220,N_23165,N_22829);
nand U25221 (N_25221,N_22900,N_23445);
nand U25222 (N_25222,N_22990,N_22554);
xnor U25223 (N_25223,N_22890,N_22727);
and U25224 (N_25224,N_23216,N_23501);
or U25225 (N_25225,N_23251,N_23635);
nand U25226 (N_25226,N_23844,N_23227);
xnor U25227 (N_25227,N_23789,N_23161);
nor U25228 (N_25228,N_23718,N_22759);
or U25229 (N_25229,N_23241,N_22732);
nand U25230 (N_25230,N_23989,N_22517);
and U25231 (N_25231,N_23152,N_23930);
or U25232 (N_25232,N_23612,N_23134);
nor U25233 (N_25233,N_23858,N_23806);
nand U25234 (N_25234,N_23515,N_23139);
or U25235 (N_25235,N_23481,N_23708);
nor U25236 (N_25236,N_22878,N_23266);
xor U25237 (N_25237,N_22952,N_22969);
nand U25238 (N_25238,N_22632,N_23053);
nor U25239 (N_25239,N_22839,N_23987);
nor U25240 (N_25240,N_23926,N_23521);
or U25241 (N_25241,N_22708,N_23623);
and U25242 (N_25242,N_23996,N_22790);
and U25243 (N_25243,N_23904,N_23515);
nand U25244 (N_25244,N_22506,N_23691);
nor U25245 (N_25245,N_23411,N_22921);
nand U25246 (N_25246,N_23036,N_23337);
and U25247 (N_25247,N_23427,N_23863);
xnor U25248 (N_25248,N_22513,N_23240);
xnor U25249 (N_25249,N_23027,N_22778);
xnor U25250 (N_25250,N_23678,N_23624);
nand U25251 (N_25251,N_23553,N_23979);
and U25252 (N_25252,N_23105,N_23503);
nor U25253 (N_25253,N_23825,N_23473);
or U25254 (N_25254,N_23901,N_22908);
and U25255 (N_25255,N_23536,N_23776);
and U25256 (N_25256,N_23650,N_23724);
or U25257 (N_25257,N_22703,N_23618);
nor U25258 (N_25258,N_22804,N_23259);
and U25259 (N_25259,N_23795,N_23371);
xnor U25260 (N_25260,N_22509,N_22535);
nand U25261 (N_25261,N_23728,N_23240);
and U25262 (N_25262,N_23932,N_23509);
nor U25263 (N_25263,N_23997,N_23342);
nand U25264 (N_25264,N_23788,N_23725);
xor U25265 (N_25265,N_23597,N_23466);
xor U25266 (N_25266,N_23414,N_23660);
nor U25267 (N_25267,N_23418,N_23934);
nand U25268 (N_25268,N_23634,N_23007);
xor U25269 (N_25269,N_23545,N_22598);
nor U25270 (N_25270,N_23396,N_23456);
or U25271 (N_25271,N_23012,N_22910);
and U25272 (N_25272,N_23521,N_23520);
and U25273 (N_25273,N_23737,N_23954);
xor U25274 (N_25274,N_22797,N_22831);
xor U25275 (N_25275,N_22588,N_23015);
and U25276 (N_25276,N_23110,N_23965);
or U25277 (N_25277,N_22739,N_23086);
xor U25278 (N_25278,N_23871,N_22736);
nor U25279 (N_25279,N_23659,N_23122);
or U25280 (N_25280,N_23751,N_23323);
nand U25281 (N_25281,N_23089,N_22983);
nor U25282 (N_25282,N_22626,N_22526);
or U25283 (N_25283,N_23682,N_22509);
or U25284 (N_25284,N_23541,N_23412);
or U25285 (N_25285,N_23079,N_22531);
nand U25286 (N_25286,N_22826,N_23926);
and U25287 (N_25287,N_22996,N_22742);
and U25288 (N_25288,N_23452,N_22974);
xor U25289 (N_25289,N_22981,N_22620);
and U25290 (N_25290,N_23428,N_22710);
xnor U25291 (N_25291,N_22977,N_22829);
or U25292 (N_25292,N_23160,N_22872);
and U25293 (N_25293,N_22531,N_23668);
or U25294 (N_25294,N_23793,N_23575);
or U25295 (N_25295,N_22575,N_23913);
xnor U25296 (N_25296,N_23273,N_23106);
xnor U25297 (N_25297,N_22827,N_22960);
and U25298 (N_25298,N_23917,N_22554);
and U25299 (N_25299,N_22883,N_22998);
xor U25300 (N_25300,N_22823,N_22975);
nand U25301 (N_25301,N_23973,N_23214);
xnor U25302 (N_25302,N_23006,N_23376);
nand U25303 (N_25303,N_22735,N_23619);
nor U25304 (N_25304,N_22666,N_23312);
nor U25305 (N_25305,N_23141,N_23842);
nor U25306 (N_25306,N_23814,N_23742);
and U25307 (N_25307,N_22971,N_22515);
and U25308 (N_25308,N_22558,N_23915);
xor U25309 (N_25309,N_23859,N_23583);
xnor U25310 (N_25310,N_23698,N_23998);
or U25311 (N_25311,N_23314,N_23575);
nor U25312 (N_25312,N_22541,N_23174);
nand U25313 (N_25313,N_23014,N_23684);
nand U25314 (N_25314,N_23413,N_22581);
nand U25315 (N_25315,N_23834,N_23637);
and U25316 (N_25316,N_23707,N_23007);
xor U25317 (N_25317,N_22663,N_22709);
or U25318 (N_25318,N_22953,N_22539);
xor U25319 (N_25319,N_23105,N_22654);
nand U25320 (N_25320,N_23204,N_22550);
and U25321 (N_25321,N_23846,N_22960);
and U25322 (N_25322,N_22957,N_23193);
nor U25323 (N_25323,N_22809,N_23367);
and U25324 (N_25324,N_23968,N_22555);
and U25325 (N_25325,N_23198,N_23390);
or U25326 (N_25326,N_22587,N_22820);
nand U25327 (N_25327,N_22963,N_23044);
and U25328 (N_25328,N_23272,N_23827);
nor U25329 (N_25329,N_23543,N_23249);
and U25330 (N_25330,N_23887,N_23986);
xor U25331 (N_25331,N_23595,N_23782);
xnor U25332 (N_25332,N_23508,N_23322);
or U25333 (N_25333,N_22948,N_23050);
or U25334 (N_25334,N_22894,N_23107);
nand U25335 (N_25335,N_22807,N_23214);
nand U25336 (N_25336,N_22593,N_23989);
and U25337 (N_25337,N_23875,N_22615);
nor U25338 (N_25338,N_23283,N_23691);
or U25339 (N_25339,N_23886,N_22804);
nor U25340 (N_25340,N_23852,N_23666);
nor U25341 (N_25341,N_23562,N_23266);
and U25342 (N_25342,N_23797,N_22979);
nand U25343 (N_25343,N_23444,N_23623);
nor U25344 (N_25344,N_23891,N_23587);
nand U25345 (N_25345,N_23269,N_23878);
or U25346 (N_25346,N_23967,N_22873);
nand U25347 (N_25347,N_23527,N_23592);
nand U25348 (N_25348,N_22728,N_23107);
xnor U25349 (N_25349,N_23848,N_22806);
and U25350 (N_25350,N_22724,N_22850);
nand U25351 (N_25351,N_23164,N_22910);
or U25352 (N_25352,N_23244,N_23821);
and U25353 (N_25353,N_23597,N_23601);
nor U25354 (N_25354,N_22613,N_23802);
or U25355 (N_25355,N_23880,N_23367);
nand U25356 (N_25356,N_23147,N_22776);
and U25357 (N_25357,N_22739,N_23894);
or U25358 (N_25358,N_23928,N_23775);
xnor U25359 (N_25359,N_22787,N_23383);
nor U25360 (N_25360,N_22680,N_23677);
or U25361 (N_25361,N_23402,N_22979);
nor U25362 (N_25362,N_22707,N_23231);
or U25363 (N_25363,N_23261,N_23783);
nand U25364 (N_25364,N_23429,N_23603);
nor U25365 (N_25365,N_23516,N_22581);
xor U25366 (N_25366,N_23722,N_22719);
xnor U25367 (N_25367,N_22933,N_23517);
or U25368 (N_25368,N_22593,N_23731);
or U25369 (N_25369,N_22500,N_23618);
and U25370 (N_25370,N_23453,N_23168);
nor U25371 (N_25371,N_23832,N_23052);
xnor U25372 (N_25372,N_23112,N_22702);
xnor U25373 (N_25373,N_23607,N_22877);
nand U25374 (N_25374,N_23674,N_23265);
xnor U25375 (N_25375,N_22872,N_23793);
or U25376 (N_25376,N_23118,N_23928);
and U25377 (N_25377,N_23685,N_22829);
nor U25378 (N_25378,N_23189,N_23009);
nand U25379 (N_25379,N_23557,N_22937);
nand U25380 (N_25380,N_22906,N_23954);
or U25381 (N_25381,N_23645,N_22852);
nor U25382 (N_25382,N_23463,N_23803);
and U25383 (N_25383,N_23525,N_22948);
nor U25384 (N_25384,N_23852,N_22730);
nor U25385 (N_25385,N_22924,N_23114);
nand U25386 (N_25386,N_23402,N_23956);
nand U25387 (N_25387,N_22530,N_23466);
nor U25388 (N_25388,N_22672,N_23235);
nand U25389 (N_25389,N_23682,N_23006);
xnor U25390 (N_25390,N_22837,N_22821);
and U25391 (N_25391,N_23124,N_22886);
or U25392 (N_25392,N_23353,N_23975);
or U25393 (N_25393,N_23131,N_23862);
or U25394 (N_25394,N_23839,N_22814);
and U25395 (N_25395,N_23790,N_22779);
nor U25396 (N_25396,N_22608,N_23106);
nand U25397 (N_25397,N_23156,N_22889);
nand U25398 (N_25398,N_23979,N_23253);
or U25399 (N_25399,N_23900,N_22782);
or U25400 (N_25400,N_23079,N_22972);
nor U25401 (N_25401,N_23730,N_23705);
xor U25402 (N_25402,N_23293,N_23429);
nor U25403 (N_25403,N_23181,N_23550);
nand U25404 (N_25404,N_23051,N_23084);
nand U25405 (N_25405,N_22839,N_23701);
nand U25406 (N_25406,N_22613,N_23493);
nand U25407 (N_25407,N_22610,N_23576);
and U25408 (N_25408,N_22761,N_23012);
or U25409 (N_25409,N_22915,N_23320);
nor U25410 (N_25410,N_22553,N_22928);
nand U25411 (N_25411,N_22945,N_23422);
xnor U25412 (N_25412,N_22794,N_23693);
nor U25413 (N_25413,N_23671,N_22889);
nand U25414 (N_25414,N_22887,N_23821);
nor U25415 (N_25415,N_23622,N_23254);
xnor U25416 (N_25416,N_23433,N_23456);
and U25417 (N_25417,N_23828,N_22846);
nand U25418 (N_25418,N_22730,N_22799);
or U25419 (N_25419,N_22913,N_22631);
nor U25420 (N_25420,N_23616,N_23408);
xor U25421 (N_25421,N_22623,N_23620);
nor U25422 (N_25422,N_22652,N_22625);
nor U25423 (N_25423,N_23125,N_22809);
nor U25424 (N_25424,N_23383,N_22833);
nor U25425 (N_25425,N_23871,N_22838);
or U25426 (N_25426,N_23577,N_23640);
nand U25427 (N_25427,N_23597,N_23836);
or U25428 (N_25428,N_23847,N_23739);
nand U25429 (N_25429,N_23694,N_23806);
and U25430 (N_25430,N_23547,N_22628);
or U25431 (N_25431,N_22876,N_23379);
and U25432 (N_25432,N_23769,N_22830);
nand U25433 (N_25433,N_22685,N_23822);
nand U25434 (N_25434,N_22773,N_23345);
nand U25435 (N_25435,N_22762,N_23392);
nand U25436 (N_25436,N_23321,N_22763);
and U25437 (N_25437,N_23076,N_22867);
nand U25438 (N_25438,N_23132,N_23798);
nor U25439 (N_25439,N_23627,N_23374);
xnor U25440 (N_25440,N_23691,N_23261);
nand U25441 (N_25441,N_23450,N_23627);
or U25442 (N_25442,N_22637,N_23505);
and U25443 (N_25443,N_23895,N_23003);
nand U25444 (N_25444,N_23436,N_23052);
or U25445 (N_25445,N_23767,N_23291);
nor U25446 (N_25446,N_23242,N_22663);
xnor U25447 (N_25447,N_22845,N_23623);
or U25448 (N_25448,N_23794,N_23651);
nand U25449 (N_25449,N_23262,N_22887);
xor U25450 (N_25450,N_23778,N_22740);
nand U25451 (N_25451,N_22840,N_22516);
or U25452 (N_25452,N_23422,N_23625);
or U25453 (N_25453,N_23304,N_23802);
nand U25454 (N_25454,N_22655,N_22919);
and U25455 (N_25455,N_22978,N_23195);
and U25456 (N_25456,N_23533,N_22884);
or U25457 (N_25457,N_23898,N_22923);
nor U25458 (N_25458,N_22819,N_22957);
and U25459 (N_25459,N_22848,N_23266);
nand U25460 (N_25460,N_23344,N_22865);
nand U25461 (N_25461,N_23351,N_23091);
xnor U25462 (N_25462,N_23306,N_23302);
nand U25463 (N_25463,N_23800,N_23419);
xor U25464 (N_25464,N_23953,N_22508);
xor U25465 (N_25465,N_22514,N_22685);
xor U25466 (N_25466,N_23233,N_22867);
xor U25467 (N_25467,N_22506,N_22889);
xnor U25468 (N_25468,N_23213,N_22611);
xor U25469 (N_25469,N_23353,N_23994);
nand U25470 (N_25470,N_22659,N_23739);
or U25471 (N_25471,N_23136,N_23249);
and U25472 (N_25472,N_23696,N_23277);
or U25473 (N_25473,N_23069,N_23551);
or U25474 (N_25474,N_23726,N_23221);
xor U25475 (N_25475,N_22793,N_22597);
and U25476 (N_25476,N_23444,N_22945);
nor U25477 (N_25477,N_23403,N_22769);
or U25478 (N_25478,N_22560,N_22736);
and U25479 (N_25479,N_23588,N_23489);
nor U25480 (N_25480,N_22950,N_22722);
and U25481 (N_25481,N_23790,N_22703);
and U25482 (N_25482,N_23837,N_23850);
xnor U25483 (N_25483,N_22969,N_23556);
xor U25484 (N_25484,N_23092,N_22644);
nor U25485 (N_25485,N_23235,N_23795);
nand U25486 (N_25486,N_23247,N_22894);
nor U25487 (N_25487,N_23240,N_22795);
or U25488 (N_25488,N_23486,N_23753);
and U25489 (N_25489,N_23954,N_22810);
nand U25490 (N_25490,N_23540,N_23198);
or U25491 (N_25491,N_22814,N_23512);
nor U25492 (N_25492,N_23524,N_22999);
and U25493 (N_25493,N_22846,N_22954);
nand U25494 (N_25494,N_23233,N_23785);
or U25495 (N_25495,N_22903,N_23261);
xor U25496 (N_25496,N_22656,N_23146);
nor U25497 (N_25497,N_23127,N_23563);
or U25498 (N_25498,N_22737,N_23365);
or U25499 (N_25499,N_22861,N_22988);
nand U25500 (N_25500,N_24393,N_24056);
and U25501 (N_25501,N_24374,N_25454);
nor U25502 (N_25502,N_24089,N_25010);
and U25503 (N_25503,N_24126,N_25402);
or U25504 (N_25504,N_24453,N_25433);
or U25505 (N_25505,N_24578,N_24308);
and U25506 (N_25506,N_24607,N_24432);
xnor U25507 (N_25507,N_24548,N_24492);
nand U25508 (N_25508,N_24654,N_24507);
xnor U25509 (N_25509,N_24159,N_25453);
and U25510 (N_25510,N_25340,N_25290);
and U25511 (N_25511,N_24029,N_24181);
nor U25512 (N_25512,N_24553,N_25445);
nand U25513 (N_25513,N_24883,N_24493);
and U25514 (N_25514,N_25456,N_24384);
xor U25515 (N_25515,N_24566,N_25094);
nor U25516 (N_25516,N_24331,N_24332);
xnor U25517 (N_25517,N_25351,N_24833);
nand U25518 (N_25518,N_24358,N_25328);
nor U25519 (N_25519,N_25493,N_24740);
nand U25520 (N_25520,N_24660,N_25278);
nand U25521 (N_25521,N_24219,N_24469);
nand U25522 (N_25522,N_25486,N_24301);
or U25523 (N_25523,N_24997,N_24665);
and U25524 (N_25524,N_25435,N_24719);
nor U25525 (N_25525,N_25246,N_25288);
and U25526 (N_25526,N_25177,N_24282);
or U25527 (N_25527,N_24437,N_25047);
and U25528 (N_25528,N_24972,N_25269);
nor U25529 (N_25529,N_24990,N_24976);
or U25530 (N_25530,N_25245,N_24125);
or U25531 (N_25531,N_24232,N_24956);
xor U25532 (N_25532,N_24193,N_24810);
or U25533 (N_25533,N_25065,N_24373);
nor U25534 (N_25534,N_24228,N_24173);
nor U25535 (N_25535,N_24354,N_24807);
xor U25536 (N_25536,N_24652,N_24072);
nor U25537 (N_25537,N_24310,N_25030);
nor U25538 (N_25538,N_24409,N_25172);
xnor U25539 (N_25539,N_25227,N_25239);
xnor U25540 (N_25540,N_24099,N_25299);
nand U25541 (N_25541,N_25281,N_24106);
or U25542 (N_25542,N_25021,N_24230);
nor U25543 (N_25543,N_25015,N_24682);
xor U25544 (N_25544,N_24641,N_25358);
nor U25545 (N_25545,N_24816,N_24555);
xor U25546 (N_25546,N_24890,N_24887);
or U25547 (N_25547,N_24508,N_24097);
and U25548 (N_25548,N_24010,N_25175);
nand U25549 (N_25549,N_24552,N_24852);
nor U25550 (N_25550,N_25184,N_24361);
nor U25551 (N_25551,N_25338,N_24382);
and U25552 (N_25552,N_24122,N_25482);
xor U25553 (N_25553,N_24520,N_25009);
nand U25554 (N_25554,N_24915,N_25032);
xor U25555 (N_25555,N_24454,N_25404);
xor U25556 (N_25556,N_24925,N_24467);
and U25557 (N_25557,N_24530,N_24789);
nor U25558 (N_25558,N_24580,N_24692);
nand U25559 (N_25559,N_25397,N_24535);
xor U25560 (N_25560,N_24819,N_24501);
nor U25561 (N_25561,N_25289,N_24055);
xnor U25562 (N_25562,N_25179,N_24762);
and U25563 (N_25563,N_24318,N_24919);
or U25564 (N_25564,N_25153,N_24563);
xor U25565 (N_25565,N_24522,N_24542);
nor U25566 (N_25566,N_24702,N_25162);
xnor U25567 (N_25567,N_25041,N_24662);
nand U25568 (N_25568,N_25183,N_25315);
nand U25569 (N_25569,N_25196,N_24827);
nor U25570 (N_25570,N_24325,N_24705);
and U25571 (N_25571,N_24567,N_24746);
xor U25572 (N_25572,N_24246,N_24250);
nor U25573 (N_25573,N_24775,N_24342);
xor U25574 (N_25574,N_24713,N_24823);
xnor U25575 (N_25575,N_25228,N_25220);
xor U25576 (N_25576,N_24212,N_24975);
nand U25577 (N_25577,N_24036,N_25400);
nand U25578 (N_25578,N_24054,N_25461);
nor U25579 (N_25579,N_25119,N_24770);
xnor U25580 (N_25580,N_24594,N_25398);
or U25581 (N_25581,N_24577,N_25255);
xnor U25582 (N_25582,N_25308,N_24281);
or U25583 (N_25583,N_24647,N_25320);
nand U25584 (N_25584,N_24289,N_24971);
or U25585 (N_25585,N_24004,N_24240);
and U25586 (N_25586,N_24486,N_24656);
and U25587 (N_25587,N_24120,N_24021);
nand U25588 (N_25588,N_25113,N_24529);
and U25589 (N_25589,N_25485,N_25084);
nor U25590 (N_25590,N_24397,N_25213);
nand U25591 (N_25591,N_24703,N_25440);
and U25592 (N_25592,N_24503,N_25182);
nor U25593 (N_25593,N_25495,N_24978);
nand U25594 (N_25594,N_24000,N_24020);
nor U25595 (N_25595,N_24188,N_25014);
xnor U25596 (N_25596,N_25173,N_24487);
nand U25597 (N_25597,N_25076,N_24715);
or U25598 (N_25598,N_24908,N_24119);
nor U25599 (N_25599,N_24375,N_24042);
and U25600 (N_25600,N_24627,N_24182);
and U25601 (N_25601,N_24366,N_24179);
and U25602 (N_25602,N_24778,N_25134);
nor U25603 (N_25603,N_24464,N_24693);
nor U25604 (N_25604,N_24950,N_24302);
and U25605 (N_25605,N_25035,N_24450);
and U25606 (N_25606,N_24988,N_24521);
nand U25607 (N_25607,N_25089,N_24076);
or U25608 (N_25608,N_25091,N_24628);
nor U25609 (N_25609,N_25250,N_25079);
and U25610 (N_25610,N_25294,N_24526);
and U25611 (N_25611,N_24668,N_25090);
and U25612 (N_25612,N_24401,N_24365);
xnor U25613 (N_25613,N_24792,N_24498);
nand U25614 (N_25614,N_24112,N_24345);
nand U25615 (N_25615,N_25307,N_24796);
xor U25616 (N_25616,N_24316,N_25092);
and U25617 (N_25617,N_24602,N_24635);
nand U25618 (N_25618,N_25459,N_24884);
and U25619 (N_25619,N_24273,N_24697);
nand U25620 (N_25620,N_24515,N_24002);
nand U25621 (N_25621,N_24839,N_24945);
nand U25622 (N_25622,N_24642,N_25152);
nor U25623 (N_25623,N_25163,N_25449);
nor U25624 (N_25624,N_24710,N_25253);
and U25625 (N_25625,N_25197,N_24428);
nand U25626 (N_25626,N_25023,N_24154);
or U25627 (N_25627,N_24413,N_25382);
or U25628 (N_25628,N_25463,N_24039);
and U25629 (N_25629,N_25011,N_25257);
nand U25630 (N_25630,N_25081,N_24234);
nand U25631 (N_25631,N_24914,N_25462);
xnor U25632 (N_25632,N_24894,N_24134);
or U25633 (N_25633,N_24573,N_24143);
and U25634 (N_25634,N_24528,N_25323);
nand U25635 (N_25635,N_24290,N_25161);
nand U25636 (N_25636,N_25284,N_25313);
or U25637 (N_25637,N_25359,N_24920);
and U25638 (N_25638,N_24330,N_24933);
nor U25639 (N_25639,N_24137,N_24438);
and U25640 (N_25640,N_24932,N_24136);
or U25641 (N_25641,N_25019,N_24747);
nand U25642 (N_25642,N_24032,N_24753);
or U25643 (N_25643,N_24203,N_24062);
nand U25644 (N_25644,N_24479,N_25037);
and U25645 (N_25645,N_24718,N_24673);
nand U25646 (N_25646,N_25038,N_25083);
or U25647 (N_25647,N_25329,N_25368);
or U25648 (N_25648,N_24221,N_25198);
nor U25649 (N_25649,N_24800,N_24699);
and U25650 (N_25650,N_24100,N_24574);
nor U25651 (N_25651,N_24296,N_24288);
nor U25652 (N_25652,N_24632,N_24116);
nand U25653 (N_25653,N_25258,N_24387);
nor U25654 (N_25654,N_24579,N_24617);
or U25655 (N_25655,N_24145,N_24306);
or U25656 (N_25656,N_24127,N_24340);
xnor U25657 (N_25657,N_25138,N_25276);
and U25658 (N_25658,N_24621,N_24830);
or U25659 (N_25659,N_24982,N_24672);
and U25660 (N_25660,N_24349,N_25249);
nor U25661 (N_25661,N_25355,N_24856);
nand U25662 (N_25662,N_24774,N_24451);
and U25663 (N_25663,N_25110,N_24944);
xor U25664 (N_25664,N_25251,N_25219);
xor U25665 (N_25665,N_25139,N_24645);
nand U25666 (N_25666,N_24601,N_24818);
nand U25667 (N_25667,N_24581,N_24410);
xnor U25668 (N_25668,N_24913,N_24108);
nand U25669 (N_25669,N_24995,N_24701);
nor U25670 (N_25670,N_24764,N_24168);
or U25671 (N_25671,N_25352,N_24786);
xnor U25672 (N_25672,N_25123,N_24284);
xor U25673 (N_25673,N_24423,N_24942);
xnor U25674 (N_25674,N_24675,N_24748);
xor U25675 (N_25675,N_24655,N_25200);
or U25676 (N_25676,N_24204,N_24691);
nand U25677 (N_25677,N_24155,N_25005);
or U25678 (N_25678,N_24756,N_25068);
or U25679 (N_25679,N_24322,N_24489);
nor U25680 (N_25680,N_25475,N_24892);
xor U25681 (N_25681,N_24977,N_24802);
nor U25682 (N_25682,N_24091,N_24257);
nand U25683 (N_25683,N_24805,N_24610);
and U25684 (N_25684,N_25260,N_25492);
or U25685 (N_25685,N_24554,N_25344);
nor U25686 (N_25686,N_25439,N_24556);
or U25687 (N_25687,N_24053,N_25121);
nand U25688 (N_25688,N_24663,N_24138);
nand U25689 (N_25689,N_25046,N_25059);
or U25690 (N_25690,N_24882,N_25303);
xnor U25691 (N_25691,N_24989,N_25469);
nor U25692 (N_25692,N_24721,N_24079);
or U25693 (N_25693,N_24880,N_25317);
nand U25694 (N_25694,N_24381,N_24772);
and U25695 (N_25695,N_24003,N_24419);
nand U25696 (N_25696,N_24456,N_25384);
nand U25697 (N_25697,N_24560,N_24139);
and U25698 (N_25698,N_24018,N_24092);
and U25699 (N_25699,N_25176,N_24376);
nand U25700 (N_25700,N_24031,N_24338);
or U25701 (N_25701,N_25088,N_25165);
or U25702 (N_25702,N_24429,N_24711);
nand U25703 (N_25703,N_24001,N_25054);
or U25704 (N_25704,N_25466,N_24534);
or U25705 (N_25705,N_25040,N_25056);
nand U25706 (N_25706,N_24620,N_25383);
xor U25707 (N_25707,N_24407,N_24446);
xor U25708 (N_25708,N_25008,N_24457);
and U25709 (N_25709,N_25471,N_24167);
xnor U25710 (N_25710,N_25286,N_25327);
or U25711 (N_25711,N_24133,N_24706);
and U25712 (N_25712,N_24047,N_24471);
nor U25713 (N_25713,N_25149,N_24545);
nor U25714 (N_25714,N_25018,N_24170);
nor U25715 (N_25715,N_25266,N_24861);
and U25716 (N_25716,N_24889,N_24795);
nor U25717 (N_25717,N_24941,N_24763);
xnor U25718 (N_25718,N_25264,N_24174);
and U25719 (N_25719,N_24938,N_24156);
nand U25720 (N_25720,N_24006,N_24847);
or U25721 (N_25721,N_24609,N_24356);
nand U25722 (N_25722,N_25222,N_24644);
nor U25723 (N_25723,N_25332,N_25272);
and U25724 (N_25724,N_24217,N_25248);
and U25725 (N_25725,N_24904,N_24911);
nor U25726 (N_25726,N_25016,N_24461);
xnor U25727 (N_25727,N_25434,N_24801);
nor U25728 (N_25728,N_24779,N_25424);
or U25729 (N_25729,N_24328,N_24983);
xnor U25730 (N_25730,N_24196,N_24160);
nor U25731 (N_25731,N_24252,N_24124);
nand U25732 (N_25732,N_24731,N_25298);
and U25733 (N_25733,N_24441,N_24996);
nor U25734 (N_25734,N_24439,N_24286);
and U25735 (N_25735,N_25007,N_25086);
or U25736 (N_25736,N_24618,N_24389);
nand U25737 (N_25737,N_24728,N_24040);
nand U25738 (N_25738,N_24192,N_24955);
nand U25739 (N_25739,N_24761,N_24336);
or U25740 (N_25740,N_24504,N_24038);
or U25741 (N_25741,N_24841,N_25418);
nor U25742 (N_25742,N_24750,N_25100);
or U25743 (N_25743,N_24992,N_24901);
and U25744 (N_25744,N_25311,N_25193);
and U25745 (N_25745,N_25326,N_24378);
or U25746 (N_25746,N_24448,N_24075);
nand U25747 (N_25747,N_25431,N_25033);
nand U25748 (N_25748,N_24631,N_24557);
nor U25749 (N_25749,N_25497,N_24478);
xor U25750 (N_25750,N_24392,N_24315);
xor U25751 (N_25751,N_25390,N_24667);
and U25752 (N_25752,N_24903,N_24958);
and U25753 (N_25753,N_24685,N_24900);
and U25754 (N_25754,N_25282,N_25131);
nand U25755 (N_25755,N_24591,N_24906);
nor U25756 (N_25756,N_25150,N_24200);
xor U25757 (N_25757,N_24050,N_25285);
nand U25758 (N_25758,N_25195,N_24538);
and U25759 (N_25759,N_24215,N_24590);
xnor U25760 (N_25760,N_25209,N_24482);
or U25761 (N_25761,N_24658,N_24071);
nand U25762 (N_25762,N_24837,N_25044);
nor U25763 (N_25763,N_25160,N_25136);
and U25764 (N_25764,N_24311,N_24164);
and U25765 (N_25765,N_24440,N_24060);
and U25766 (N_25766,N_24905,N_25167);
nor U25767 (N_25767,N_24371,N_25256);
or U25768 (N_25768,N_24473,N_24352);
nor U25769 (N_25769,N_25421,N_24277);
nor U25770 (N_25770,N_24386,N_24237);
xor U25771 (N_25771,N_24812,N_24576);
nand U25772 (N_25772,N_25247,N_24019);
or U25773 (N_25773,N_24659,N_24637);
nand U25774 (N_25774,N_24592,N_25448);
nor U25775 (N_25775,N_24611,N_24351);
or U25776 (N_25776,N_25204,N_24781);
nor U25777 (N_25777,N_24058,N_24926);
xnor U25778 (N_25778,N_25478,N_24022);
or U25779 (N_25779,N_24785,N_24085);
nor U25780 (N_25780,N_24109,N_24681);
nor U25781 (N_25781,N_24037,N_24649);
nor U25782 (N_25782,N_24803,N_24897);
or U25783 (N_25783,N_24811,N_24171);
nor U25784 (N_25784,N_25291,N_25498);
or U25785 (N_25785,N_24622,N_24863);
or U25786 (N_25786,N_24207,N_25034);
xnor U25787 (N_25787,N_24736,N_25292);
and U25788 (N_25788,N_25361,N_25186);
nor U25789 (N_25789,N_25096,N_24254);
nand U25790 (N_25790,N_24028,N_25302);
or U25791 (N_25791,N_24465,N_24688);
or U25792 (N_25792,N_24758,N_24524);
nor U25793 (N_25793,N_24981,N_24080);
nand U25794 (N_25794,N_24191,N_24095);
or U25795 (N_25795,N_24858,N_24166);
and U25796 (N_25796,N_25168,N_24025);
xnor U25797 (N_25797,N_25314,N_25104);
nor U25798 (N_25798,N_24488,N_24206);
xnor U25799 (N_25799,N_24829,N_24307);
xor U25800 (N_25800,N_25413,N_24474);
and U25801 (N_25801,N_25111,N_24293);
or U25802 (N_25802,N_24902,N_25262);
nor U25803 (N_25803,N_24113,N_24165);
nor U25804 (N_25804,N_24571,N_25004);
nor U25805 (N_25805,N_24225,N_24623);
nor U25806 (N_25806,N_24102,N_24074);
nor U25807 (N_25807,N_24712,N_24947);
or U25808 (N_25808,N_25267,N_24026);
nand U25809 (N_25809,N_24743,N_25191);
xnor U25810 (N_25810,N_24848,N_25367);
nor U25811 (N_25811,N_24210,N_25380);
or U25812 (N_25812,N_24633,N_25158);
nand U25813 (N_25813,N_24404,N_24238);
nor U25814 (N_25814,N_25305,N_24674);
nand U25815 (N_25815,N_24417,N_24783);
or U25816 (N_25816,N_25385,N_24999);
nor U25817 (N_25817,N_24013,N_24494);
nand U25818 (N_25818,N_24639,N_25487);
or U25819 (N_25819,N_24477,N_24549);
xor U25820 (N_25820,N_24023,N_24771);
nor U25821 (N_25821,N_24595,N_24634);
nand U25822 (N_25822,N_24510,N_25207);
nand U25823 (N_25823,N_24270,N_25364);
nand U25824 (N_25824,N_25379,N_24065);
xor U25825 (N_25825,N_24251,N_24888);
or U25826 (N_25826,N_25374,N_25316);
xnor U25827 (N_25827,N_24943,N_24421);
and U25828 (N_25828,N_24872,N_24436);
or U25829 (N_25829,N_24568,N_25097);
and U25830 (N_25830,N_25399,N_24247);
nor U25831 (N_25831,N_25318,N_24390);
nor U25832 (N_25832,N_25339,N_25000);
or U25833 (N_25833,N_24625,N_24248);
xnor U25834 (N_25834,N_24869,N_25169);
and U25835 (N_25835,N_25496,N_25429);
nor U25836 (N_25836,N_24271,N_24886);
nor U25837 (N_25837,N_25265,N_25401);
and U25838 (N_25838,N_24117,N_24757);
xor U25839 (N_25839,N_24317,N_24157);
nand U25840 (N_25840,N_25001,N_24445);
nand U25841 (N_25841,N_25140,N_24132);
or U25842 (N_25842,N_25042,N_25022);
nor U25843 (N_25843,N_24729,N_24853);
xnor U25844 (N_25844,N_24572,N_24149);
or U25845 (N_25845,N_25393,N_25052);
nand U25846 (N_25846,N_24733,N_24984);
or U25847 (N_25847,N_24460,N_24849);
nand U25848 (N_25848,N_24707,N_25093);
nand U25849 (N_25849,N_25066,N_24547);
and U25850 (N_25850,N_24312,N_24629);
nand U25851 (N_25851,N_25217,N_24496);
nor U25852 (N_25852,N_24426,N_24129);
and U25853 (N_25853,N_25129,N_24586);
and U25854 (N_25854,N_25109,N_25357);
xor U25855 (N_25855,N_25270,N_25408);
and U25856 (N_25856,N_24536,N_24924);
xor U25857 (N_25857,N_25263,N_24745);
nor U25858 (N_25858,N_24828,N_24323);
nor U25859 (N_25859,N_24544,N_25141);
or U25860 (N_25860,N_24049,N_25214);
nor U25861 (N_25861,N_24144,N_25166);
or U25862 (N_25862,N_25322,N_24222);
nand U25863 (N_25863,N_24388,N_25369);
nand U25864 (N_25864,N_24268,N_24497);
and U25865 (N_25865,N_25297,N_24940);
and U25866 (N_25866,N_24383,N_24636);
xnor U25867 (N_25867,N_24223,N_24135);
and U25868 (N_25868,N_24370,N_24430);
or U25869 (N_25869,N_24339,N_24295);
nor U25870 (N_25870,N_24612,N_24606);
nor U25871 (N_25871,N_25223,N_24261);
nand U25872 (N_25872,N_24015,N_24502);
and U25873 (N_25873,N_24648,N_25480);
and U25874 (N_25874,N_25230,N_24518);
nor U25875 (N_25875,N_24878,N_25127);
xor U25876 (N_25876,N_24831,N_24087);
or U25877 (N_25877,N_24584,N_25360);
or U25878 (N_25878,N_24422,N_24408);
and U25879 (N_25879,N_25238,N_24814);
and U25880 (N_25880,N_25447,N_24304);
xor U25881 (N_25881,N_25387,N_24798);
nor U25882 (N_25882,N_24103,N_24353);
nand U25883 (N_25883,N_25003,N_24073);
or U25884 (N_25884,N_24836,N_25375);
nor U25885 (N_25885,N_24511,N_25427);
xor U25886 (N_25886,N_25231,N_25101);
nand U25887 (N_25887,N_24414,N_24285);
nor U25888 (N_25888,N_25103,N_24259);
or U25889 (N_25889,N_24005,N_24499);
nand U25890 (N_25890,N_25268,N_24169);
nor U25891 (N_25891,N_25194,N_24817);
nand U25892 (N_25892,N_25406,N_24363);
xor U25893 (N_25893,N_25425,N_24041);
nand U25894 (N_25894,N_25178,N_24730);
nand U25895 (N_25895,N_25426,N_25414);
nand U25896 (N_25896,N_24776,N_25460);
or U25897 (N_25897,N_24813,N_24734);
nor U25898 (N_25898,N_24274,N_24367);
nor U25899 (N_25899,N_24162,N_24275);
nor U25900 (N_25900,N_25488,N_24550);
nor U25901 (N_25901,N_24677,N_25465);
nand U25902 (N_25902,N_25077,N_25403);
and U25903 (N_25903,N_25221,N_25412);
nor U25904 (N_25904,N_24090,N_24077);
nor U25905 (N_25905,N_24857,N_25189);
nand U25906 (N_25906,N_24186,N_24115);
and U25907 (N_25907,N_24030,N_24922);
xnor U25908 (N_25908,N_25132,N_25024);
nor U25909 (N_25909,N_25115,N_24939);
xnor U25910 (N_25910,N_25151,N_24141);
xor U25911 (N_25911,N_24359,N_24679);
xnor U25912 (N_25912,N_24724,N_24184);
nand U25913 (N_25913,N_24313,N_24434);
nor U25914 (N_25914,N_24185,N_24280);
or U25915 (N_25915,N_24993,N_24216);
xor U25916 (N_25916,N_24070,N_25451);
nor U25917 (N_25917,N_24333,N_24364);
nand U25918 (N_25918,N_24643,N_25107);
nand U25919 (N_25919,N_24509,N_24420);
nor U25920 (N_25920,N_24916,N_24597);
nand U25921 (N_25921,N_25287,N_24208);
nand U25922 (N_25922,N_24921,N_24431);
nor U25923 (N_25923,N_24418,N_24123);
and U25924 (N_25924,N_24344,N_24966);
xor U25925 (N_25925,N_25350,N_25055);
or U25926 (N_25926,N_24355,N_25409);
xor U25927 (N_25927,N_24394,N_24158);
or U25928 (N_25928,N_25283,N_24197);
xnor U25929 (N_25929,N_24279,N_24402);
xnor U25930 (N_25930,N_24088,N_24985);
nor U25931 (N_25931,N_24379,N_25330);
and U25932 (N_25932,N_24575,N_24176);
xnor U25933 (N_25933,N_24416,N_25117);
nor U25934 (N_25934,N_25063,N_25376);
and U25935 (N_25935,N_24303,N_25120);
nor U25936 (N_25936,N_24235,N_24415);
xnor U25937 (N_25937,N_25098,N_24403);
nand U25938 (N_25938,N_24128,N_25002);
nor U25939 (N_25939,N_24791,N_24787);
or U25940 (N_25940,N_25275,N_25325);
xor U25941 (N_25941,N_25244,N_24700);
nand U25942 (N_25942,N_24615,N_25061);
xnor U25943 (N_25943,N_24804,N_25225);
nand U25944 (N_25944,N_25036,N_24269);
or U25945 (N_25945,N_24797,N_24299);
xnor U25946 (N_25946,N_24016,N_24671);
nor U25947 (N_25947,N_24395,N_24287);
xor U25948 (N_25948,N_24458,N_24744);
nor U25949 (N_25949,N_24998,N_24199);
xor U25950 (N_25950,N_25411,N_24024);
or U25951 (N_25951,N_25174,N_24570);
and U25952 (N_25952,N_25026,N_25078);
nand U25953 (N_25953,N_24725,N_24427);
nor U25954 (N_25954,N_24959,N_24773);
nand U25955 (N_25955,N_25499,N_25490);
and U25956 (N_25956,N_24506,N_24650);
or U25957 (N_25957,N_24963,N_25025);
nand U25958 (N_25958,N_24098,N_25464);
nor U25959 (N_25959,N_24483,N_24893);
nand U25960 (N_25960,N_24033,N_24808);
and U25961 (N_25961,N_25452,N_25388);
or U25962 (N_25962,N_24832,N_24468);
or U25963 (N_25963,N_25199,N_25444);
nor U25964 (N_25964,N_24241,N_24582);
or U25965 (N_25965,N_25242,N_24569);
xor U25966 (N_25966,N_25277,N_25321);
nor U25967 (N_25967,N_24912,N_25389);
xnor U25968 (N_25968,N_24855,N_24399);
xor U25969 (N_25969,N_24840,N_25027);
and U25970 (N_25970,N_24824,N_24046);
nor U25971 (N_25971,N_24175,N_24011);
and U25972 (N_25972,N_24877,N_24505);
or U25973 (N_25973,N_24245,N_24873);
nand U25974 (N_25974,N_24537,N_24104);
xnor U25975 (N_25975,N_24107,N_25274);
and U25976 (N_25976,N_24096,N_24551);
nor U25977 (N_25977,N_24412,N_24968);
xor U25978 (N_25978,N_25210,N_24935);
nor U25979 (N_25979,N_24844,N_24953);
and U25980 (N_25980,N_24300,N_24640);
and U25981 (N_25981,N_24348,N_25342);
xnor U25982 (N_25982,N_24151,N_24346);
or U25983 (N_25983,N_25236,N_24646);
nor U25984 (N_25984,N_25337,N_24396);
nor U25985 (N_25985,N_24918,N_24183);
nor U25986 (N_25986,N_25353,N_24616);
nor U25987 (N_25987,N_25349,N_24201);
xor U25988 (N_25988,N_24979,N_24603);
or U25989 (N_25989,N_24604,N_24017);
or U25990 (N_25990,N_24531,N_25371);
xor U25991 (N_25991,N_24034,N_24084);
nand U25992 (N_25992,N_25407,N_25333);
or U25993 (N_25993,N_24444,N_24834);
nor U25994 (N_25994,N_25395,N_24140);
xor U25995 (N_25995,N_25112,N_25324);
xnor U25996 (N_25996,N_25192,N_24110);
nor U25997 (N_25997,N_24752,N_24907);
nand U25998 (N_25998,N_24854,N_24226);
and U25999 (N_25999,N_24875,N_24177);
or U26000 (N_26000,N_24626,N_24696);
nand U26001 (N_26001,N_25012,N_24256);
nor U26002 (N_26002,N_24562,N_24838);
or U26003 (N_26003,N_25484,N_25300);
nand U26004 (N_26004,N_25180,N_25457);
nor U26005 (N_26005,N_25483,N_24661);
and U26006 (N_26006,N_24741,N_24424);
xor U26007 (N_26007,N_25341,N_25187);
or U26008 (N_26008,N_24198,N_25336);
xnor U26009 (N_26009,N_24305,N_25377);
and U26010 (N_26010,N_25293,N_24891);
nand U26011 (N_26011,N_24951,N_25422);
xnor U26012 (N_26012,N_24881,N_25354);
nand U26013 (N_26013,N_25080,N_24224);
xor U26014 (N_26014,N_24964,N_25155);
xnor U26015 (N_26015,N_25334,N_24491);
or U26016 (N_26016,N_25416,N_25133);
nor U26017 (N_26017,N_24759,N_25212);
nand U26018 (N_26018,N_25105,N_24101);
xor U26019 (N_26019,N_25215,N_24083);
nand U26020 (N_26020,N_24868,N_24329);
xor U26021 (N_26021,N_24012,N_25203);
nor U26022 (N_26022,N_24064,N_25373);
xnor U26023 (N_26023,N_24263,N_24541);
xor U26024 (N_26024,N_24599,N_24686);
nand U26025 (N_26025,N_25396,N_24684);
nand U26026 (N_26026,N_24319,N_25280);
and U26027 (N_26027,N_25095,N_25345);
xor U26028 (N_26028,N_25450,N_24769);
nand U26029 (N_26029,N_24272,N_24455);
and U26030 (N_26030,N_24220,N_24716);
xnor U26031 (N_26031,N_24760,N_24987);
nor U26032 (N_26032,N_24533,N_25058);
xor U26033 (N_26033,N_24754,N_25020);
or U26034 (N_26034,N_24749,N_24879);
xor U26035 (N_26035,N_24600,N_24525);
and U26036 (N_26036,N_24044,N_24928);
xnor U26037 (N_26037,N_24267,N_25362);
nor U26038 (N_26038,N_25430,N_24057);
nand U26039 (N_26039,N_25128,N_24587);
nand U26040 (N_26040,N_24211,N_24561);
or U26041 (N_26041,N_24720,N_24068);
nand U26042 (N_26042,N_24243,N_24052);
nand U26043 (N_26043,N_24937,N_25108);
or U26044 (N_26044,N_25122,N_24742);
nor U26045 (N_26045,N_24689,N_24443);
and U26046 (N_26046,N_24266,N_24297);
or U26047 (N_26047,N_24147,N_25295);
xor U26048 (N_26048,N_25070,N_24860);
and U26049 (N_26049,N_25436,N_25147);
xor U26050 (N_26050,N_24683,N_24952);
or U26051 (N_26051,N_24727,N_24172);
nand U26052 (N_26052,N_24589,N_24276);
and U26053 (N_26053,N_24732,N_25356);
nor U26054 (N_26054,N_24481,N_25142);
nor U26055 (N_26055,N_25229,N_24695);
and U26056 (N_26056,N_25470,N_24253);
and U26057 (N_26057,N_25428,N_24957);
or U26058 (N_26058,N_24368,N_25130);
nor U26059 (N_26059,N_24898,N_25391);
nand U26060 (N_26060,N_24320,N_25423);
or U26061 (N_26061,N_24063,N_24846);
nand U26062 (N_26062,N_24564,N_25053);
xor U26063 (N_26063,N_25479,N_24826);
nand U26064 (N_26064,N_24954,N_24859);
nor U26065 (N_26065,N_25252,N_25312);
or U26066 (N_26066,N_24676,N_25082);
xor U26067 (N_26067,N_24842,N_24043);
nand U26068 (N_26068,N_24876,N_25386);
and U26069 (N_26069,N_25159,N_24835);
xor U26070 (N_26070,N_25415,N_25347);
nor U26071 (N_26071,N_24739,N_25442);
and U26072 (N_26072,N_25074,N_25346);
nor U26073 (N_26073,N_24755,N_25145);
nand U26074 (N_26074,N_24614,N_25211);
xor U26075 (N_26075,N_24082,N_24657);
or U26076 (N_26076,N_24283,N_24588);
or U26077 (N_26077,N_25392,N_25343);
nor U26078 (N_26078,N_25137,N_25243);
or U26079 (N_26079,N_24326,N_24400);
and U26080 (N_26080,N_24678,N_25156);
and U26081 (N_26081,N_24593,N_25048);
or U26082 (N_26082,N_24153,N_24398);
and U26083 (N_26083,N_24078,N_25208);
and U26084 (N_26084,N_24527,N_24517);
and U26085 (N_26085,N_24514,N_24209);
xor U26086 (N_26086,N_24061,N_24190);
and U26087 (N_26087,N_24086,N_24664);
or U26088 (N_26088,N_24146,N_25073);
nor U26089 (N_26089,N_24484,N_25241);
nand U26090 (N_26090,N_24093,N_24896);
xnor U26091 (N_26091,N_24008,N_24121);
nand U26092 (N_26092,N_24242,N_24485);
xor U26093 (N_26093,N_24341,N_24767);
nor U26094 (N_26094,N_25309,N_25443);
or U26095 (N_26095,N_25135,N_24213);
nand U26096 (N_26096,N_24864,N_25446);
nor U26097 (N_26097,N_24540,N_25372);
nor U26098 (N_26098,N_24680,N_25017);
xnor U26099 (N_26099,N_25467,N_24845);
nand U26100 (N_26100,N_24821,N_25261);
nor U26101 (N_26101,N_24726,N_24405);
and U26102 (N_26102,N_24111,N_25071);
xnor U26103 (N_26103,N_25335,N_24435);
or U26104 (N_26104,N_24899,N_24946);
nand U26105 (N_26105,N_24874,N_24452);
xnor U26106 (N_26106,N_24806,N_25474);
nor U26107 (N_26107,N_25218,N_25468);
or U26108 (N_26108,N_24969,N_24608);
and U26109 (N_26109,N_24466,N_24523);
or U26110 (N_26110,N_24009,N_24462);
nor U26111 (N_26111,N_25031,N_24513);
xnor U26112 (N_26112,N_24871,N_24327);
or U26113 (N_26113,N_24694,N_25075);
and U26114 (N_26114,N_25310,N_24708);
nand U26115 (N_26115,N_24927,N_25043);
xor U26116 (N_26116,N_24687,N_25226);
nor U26117 (N_26117,N_24051,N_24470);
nand U26118 (N_26118,N_24343,N_24027);
and U26119 (N_26119,N_24735,N_24965);
nor U26120 (N_26120,N_25154,N_25363);
and U26121 (N_26121,N_24784,N_24229);
and U26122 (N_26122,N_24495,N_24865);
nor U26123 (N_26123,N_24980,N_24931);
nand U26124 (N_26124,N_24380,N_24130);
or U26125 (N_26125,N_24596,N_25271);
nand U26126 (N_26126,N_25164,N_25437);
nand U26127 (N_26127,N_25381,N_25064);
and U26128 (N_26128,N_25124,N_24459);
nand U26129 (N_26129,N_24233,N_24391);
nand U26130 (N_26130,N_24360,N_24653);
and U26131 (N_26131,N_24048,N_24202);
nor U26132 (N_26132,N_24425,N_24619);
xor U26133 (N_26133,N_25206,N_24347);
xor U26134 (N_26134,N_25259,N_24059);
nand U26135 (N_26135,N_25472,N_24895);
nand U26136 (N_26136,N_24669,N_25494);
or U26137 (N_26137,N_25378,N_25365);
nand U26138 (N_26138,N_25273,N_24934);
and U26139 (N_26139,N_25458,N_25237);
nand U26140 (N_26140,N_24227,N_24558);
nor U26141 (N_26141,N_24780,N_25481);
xnor U26142 (N_26142,N_25477,N_24362);
and U26143 (N_26143,N_24377,N_24973);
nor U26144 (N_26144,N_24372,N_25157);
or U26145 (N_26145,N_25476,N_24150);
nand U26146 (N_26146,N_24264,N_25432);
nor U26147 (N_26147,N_24709,N_25050);
nand U26148 (N_26148,N_25170,N_24866);
nor U26149 (N_26149,N_24788,N_25144);
nand U26150 (N_26150,N_25232,N_25099);
or U26151 (N_26151,N_24258,N_24962);
or U26152 (N_26152,N_24782,N_25148);
nand U26153 (N_26153,N_25441,N_24178);
nor U26154 (N_26154,N_24163,N_25069);
xor U26155 (N_26155,N_24490,N_24532);
xnor U26156 (N_26156,N_24094,N_24986);
nor U26157 (N_26157,N_24974,N_24698);
and U26158 (N_26158,N_24476,N_24131);
and U26159 (N_26159,N_24670,N_24613);
xor U26160 (N_26160,N_24298,N_25279);
nand U26161 (N_26161,N_25114,N_24007);
or U26162 (N_26162,N_25006,N_24723);
nor U26163 (N_26163,N_24239,N_24794);
nor U26164 (N_26164,N_25301,N_24929);
and U26165 (N_26165,N_24624,N_25171);
and U26166 (N_26166,N_24867,N_24519);
nor U26167 (N_26167,N_24114,N_24214);
and U26168 (N_26168,N_24605,N_25106);
and U26169 (N_26169,N_24337,N_25405);
nor U26170 (N_26170,N_24142,N_25029);
and U26171 (N_26171,N_24930,N_24967);
and U26172 (N_26172,N_25051,N_24870);
or U26173 (N_26173,N_25240,N_24598);
xor U26174 (N_26174,N_25181,N_25116);
or U26175 (N_26175,N_25201,N_24194);
and U26176 (N_26176,N_24350,N_25489);
nand U26177 (N_26177,N_24815,N_24512);
xnor U26178 (N_26178,N_24357,N_24292);
xnor U26179 (N_26179,N_24949,N_24809);
or U26180 (N_26180,N_25394,N_24651);
or U26181 (N_26181,N_24189,N_25013);
and U26182 (N_26182,N_25205,N_24717);
or U26183 (N_26183,N_25126,N_24152);
nor U26184 (N_26184,N_24066,N_24751);
or U26185 (N_26185,N_24278,N_24406);
nor U26186 (N_26186,N_25072,N_24994);
nor U26187 (N_26187,N_24447,N_24069);
xnor U26188 (N_26188,N_24851,N_24936);
nand U26189 (N_26189,N_25028,N_25410);
or U26190 (N_26190,N_24294,N_24583);
xnor U26191 (N_26191,N_24411,N_24565);
and U26192 (N_26192,N_24433,N_24369);
nor U26193 (N_26193,N_25234,N_24585);
and U26194 (N_26194,N_24218,N_24910);
or U26195 (N_26195,N_24970,N_25045);
and U26196 (N_26196,N_24385,N_24249);
or U26197 (N_26197,N_25420,N_24738);
nor U26198 (N_26198,N_24768,N_24265);
and U26199 (N_26199,N_24081,N_24799);
or U26200 (N_26200,N_24255,N_24180);
or U26201 (N_26201,N_24793,N_24737);
and U26202 (N_26202,N_24885,N_25087);
nor U26203 (N_26203,N_24850,N_25438);
and U26204 (N_26204,N_24917,N_24335);
nand U26205 (N_26205,N_25419,N_25306);
nand U26206 (N_26206,N_25185,N_24067);
nand U26207 (N_26207,N_25216,N_25370);
and U26208 (N_26208,N_24500,N_24766);
nand U26209 (N_26209,N_25190,N_24324);
and U26210 (N_26210,N_25473,N_25188);
nor U26211 (N_26211,N_25331,N_25085);
and U26212 (N_26212,N_24472,N_25235);
nor U26213 (N_26213,N_24244,N_24463);
xor U26214 (N_26214,N_24923,N_24231);
xor U26215 (N_26215,N_24035,N_24045);
or U26216 (N_26216,N_24187,N_25417);
nand U26217 (N_26217,N_25366,N_24704);
or U26218 (N_26218,N_24991,N_24480);
nand U26219 (N_26219,N_25254,N_25348);
xnor U26220 (N_26220,N_25304,N_24714);
xor U26221 (N_26221,N_25067,N_25049);
nor U26222 (N_26222,N_24546,N_24777);
nand U26223 (N_26223,N_25060,N_25455);
nor U26224 (N_26224,N_24205,N_24666);
xnor U26225 (N_26225,N_24948,N_24260);
nand U26226 (N_26226,N_24195,N_24475);
nand U26227 (N_26227,N_25319,N_24961);
nor U26228 (N_26228,N_24820,N_24960);
nor U26229 (N_26229,N_25118,N_24334);
nor U26230 (N_26230,N_25102,N_25146);
nor U26231 (N_26231,N_25125,N_24822);
xnor U26232 (N_26232,N_24148,N_25039);
xnor U26233 (N_26233,N_24291,N_25491);
nand U26234 (N_26234,N_24449,N_24825);
or U26235 (N_26235,N_24516,N_24309);
nand U26236 (N_26236,N_24862,N_24321);
nand U26237 (N_26237,N_25143,N_24161);
xor U26238 (N_26238,N_25202,N_24690);
and U26239 (N_26239,N_24638,N_25057);
or U26240 (N_26240,N_25233,N_24105);
nor U26241 (N_26241,N_24262,N_25062);
or U26242 (N_26242,N_24630,N_24722);
nor U26243 (N_26243,N_25296,N_24118);
nor U26244 (N_26244,N_24843,N_24543);
xnor U26245 (N_26245,N_25224,N_24559);
nand U26246 (N_26246,N_24314,N_24909);
nor U26247 (N_26247,N_24442,N_24236);
or U26248 (N_26248,N_24790,N_24539);
xor U26249 (N_26249,N_24014,N_24765);
nor U26250 (N_26250,N_24941,N_25218);
or U26251 (N_26251,N_24704,N_24395);
xnor U26252 (N_26252,N_24557,N_24967);
nor U26253 (N_26253,N_24223,N_25237);
or U26254 (N_26254,N_24404,N_24999);
nand U26255 (N_26255,N_24544,N_24783);
and U26256 (N_26256,N_24728,N_24668);
and U26257 (N_26257,N_25462,N_25218);
xor U26258 (N_26258,N_25400,N_24936);
nor U26259 (N_26259,N_24029,N_25099);
nand U26260 (N_26260,N_25270,N_24469);
or U26261 (N_26261,N_24122,N_24402);
nand U26262 (N_26262,N_25454,N_24873);
or U26263 (N_26263,N_24273,N_24145);
and U26264 (N_26264,N_25122,N_25177);
nand U26265 (N_26265,N_24856,N_24199);
xor U26266 (N_26266,N_24834,N_25457);
and U26267 (N_26267,N_24590,N_24341);
nor U26268 (N_26268,N_24371,N_24109);
or U26269 (N_26269,N_24858,N_25325);
nor U26270 (N_26270,N_25351,N_25048);
or U26271 (N_26271,N_24551,N_24020);
nor U26272 (N_26272,N_24433,N_24372);
xnor U26273 (N_26273,N_24625,N_24643);
nor U26274 (N_26274,N_24663,N_24148);
nand U26275 (N_26275,N_25027,N_24025);
nand U26276 (N_26276,N_24164,N_25385);
or U26277 (N_26277,N_24480,N_24460);
and U26278 (N_26278,N_24003,N_25080);
nor U26279 (N_26279,N_24909,N_24823);
nor U26280 (N_26280,N_24161,N_25076);
nand U26281 (N_26281,N_24948,N_24938);
nand U26282 (N_26282,N_25065,N_24462);
or U26283 (N_26283,N_24369,N_25277);
nor U26284 (N_26284,N_24820,N_25317);
or U26285 (N_26285,N_24582,N_24508);
xor U26286 (N_26286,N_25153,N_25292);
nor U26287 (N_26287,N_25109,N_24308);
xor U26288 (N_26288,N_24398,N_25173);
and U26289 (N_26289,N_25194,N_24156);
or U26290 (N_26290,N_24920,N_25255);
nand U26291 (N_26291,N_24465,N_24540);
xnor U26292 (N_26292,N_25223,N_25008);
and U26293 (N_26293,N_25100,N_24428);
and U26294 (N_26294,N_25264,N_24352);
xor U26295 (N_26295,N_25483,N_24832);
xor U26296 (N_26296,N_24795,N_24572);
and U26297 (N_26297,N_24494,N_25317);
or U26298 (N_26298,N_24450,N_25244);
nor U26299 (N_26299,N_24803,N_24384);
nor U26300 (N_26300,N_24380,N_24987);
nand U26301 (N_26301,N_24165,N_25244);
or U26302 (N_26302,N_24629,N_25070);
and U26303 (N_26303,N_24166,N_24247);
or U26304 (N_26304,N_24809,N_25136);
nand U26305 (N_26305,N_24373,N_24100);
nand U26306 (N_26306,N_25289,N_25481);
nor U26307 (N_26307,N_24387,N_24467);
nand U26308 (N_26308,N_24321,N_24439);
or U26309 (N_26309,N_24776,N_24398);
nor U26310 (N_26310,N_24224,N_24046);
nand U26311 (N_26311,N_24157,N_25420);
nand U26312 (N_26312,N_25386,N_24416);
and U26313 (N_26313,N_24626,N_25179);
nand U26314 (N_26314,N_24727,N_24690);
xor U26315 (N_26315,N_24375,N_24415);
or U26316 (N_26316,N_24244,N_25173);
nor U26317 (N_26317,N_24157,N_24031);
nand U26318 (N_26318,N_25232,N_25167);
xnor U26319 (N_26319,N_24587,N_24060);
and U26320 (N_26320,N_24495,N_24395);
nand U26321 (N_26321,N_24128,N_24689);
nor U26322 (N_26322,N_25151,N_25227);
nand U26323 (N_26323,N_24963,N_25329);
xor U26324 (N_26324,N_24905,N_25340);
or U26325 (N_26325,N_24338,N_24501);
or U26326 (N_26326,N_25499,N_25242);
nor U26327 (N_26327,N_24726,N_24681);
nor U26328 (N_26328,N_24891,N_24552);
xnor U26329 (N_26329,N_24746,N_24975);
and U26330 (N_26330,N_25476,N_25022);
and U26331 (N_26331,N_24062,N_25388);
and U26332 (N_26332,N_25495,N_24135);
nor U26333 (N_26333,N_25063,N_24611);
or U26334 (N_26334,N_25033,N_24785);
nand U26335 (N_26335,N_24375,N_24773);
and U26336 (N_26336,N_25212,N_24963);
and U26337 (N_26337,N_24224,N_24764);
and U26338 (N_26338,N_25478,N_25105);
or U26339 (N_26339,N_24838,N_25209);
xnor U26340 (N_26340,N_24918,N_25085);
nor U26341 (N_26341,N_24464,N_24790);
or U26342 (N_26342,N_24679,N_24324);
or U26343 (N_26343,N_25053,N_24860);
nand U26344 (N_26344,N_25481,N_24838);
and U26345 (N_26345,N_24650,N_24573);
nor U26346 (N_26346,N_24267,N_24337);
nor U26347 (N_26347,N_25009,N_25031);
or U26348 (N_26348,N_24966,N_25115);
nor U26349 (N_26349,N_25477,N_24790);
nand U26350 (N_26350,N_24136,N_24636);
nand U26351 (N_26351,N_25318,N_24254);
and U26352 (N_26352,N_24929,N_24693);
or U26353 (N_26353,N_24363,N_25052);
or U26354 (N_26354,N_25015,N_25364);
nor U26355 (N_26355,N_25206,N_24550);
xnor U26356 (N_26356,N_24166,N_24121);
xor U26357 (N_26357,N_24420,N_25080);
nor U26358 (N_26358,N_25032,N_24870);
nand U26359 (N_26359,N_24997,N_25006);
or U26360 (N_26360,N_24666,N_25222);
and U26361 (N_26361,N_24542,N_24011);
xor U26362 (N_26362,N_25133,N_25484);
or U26363 (N_26363,N_24608,N_25251);
nand U26364 (N_26364,N_24042,N_24639);
nor U26365 (N_26365,N_24916,N_24245);
nand U26366 (N_26366,N_24566,N_24549);
nand U26367 (N_26367,N_24556,N_25299);
xor U26368 (N_26368,N_25320,N_25191);
nor U26369 (N_26369,N_24554,N_25122);
nor U26370 (N_26370,N_24560,N_25004);
nor U26371 (N_26371,N_25402,N_25103);
or U26372 (N_26372,N_24783,N_25001);
nor U26373 (N_26373,N_24658,N_24385);
nor U26374 (N_26374,N_24209,N_24999);
nor U26375 (N_26375,N_24068,N_24716);
nand U26376 (N_26376,N_24824,N_24362);
nor U26377 (N_26377,N_25337,N_24961);
nand U26378 (N_26378,N_24038,N_25322);
or U26379 (N_26379,N_24303,N_24164);
nor U26380 (N_26380,N_24353,N_24970);
nand U26381 (N_26381,N_25388,N_24302);
xor U26382 (N_26382,N_24617,N_24997);
nor U26383 (N_26383,N_24475,N_24298);
and U26384 (N_26384,N_24659,N_24145);
nand U26385 (N_26385,N_24377,N_24460);
nand U26386 (N_26386,N_25146,N_25301);
or U26387 (N_26387,N_25037,N_25226);
and U26388 (N_26388,N_25240,N_24543);
and U26389 (N_26389,N_24231,N_24177);
xnor U26390 (N_26390,N_25093,N_24112);
nand U26391 (N_26391,N_24370,N_24135);
or U26392 (N_26392,N_24130,N_25021);
nor U26393 (N_26393,N_24552,N_24464);
nand U26394 (N_26394,N_25222,N_24111);
xnor U26395 (N_26395,N_24944,N_24081);
xor U26396 (N_26396,N_25226,N_24681);
and U26397 (N_26397,N_24755,N_24330);
nor U26398 (N_26398,N_25083,N_24003);
xnor U26399 (N_26399,N_24350,N_25155);
and U26400 (N_26400,N_24750,N_25476);
xnor U26401 (N_26401,N_25292,N_24079);
xor U26402 (N_26402,N_24602,N_25094);
or U26403 (N_26403,N_25459,N_24132);
xnor U26404 (N_26404,N_25269,N_24967);
nand U26405 (N_26405,N_24418,N_24391);
and U26406 (N_26406,N_25362,N_25172);
nand U26407 (N_26407,N_25427,N_24721);
nand U26408 (N_26408,N_24740,N_24140);
nor U26409 (N_26409,N_24247,N_24941);
or U26410 (N_26410,N_25113,N_24368);
nand U26411 (N_26411,N_24920,N_24091);
or U26412 (N_26412,N_25213,N_24252);
or U26413 (N_26413,N_24853,N_25398);
nand U26414 (N_26414,N_25226,N_24432);
or U26415 (N_26415,N_24200,N_25138);
nand U26416 (N_26416,N_24523,N_24834);
or U26417 (N_26417,N_24808,N_24512);
and U26418 (N_26418,N_24034,N_25102);
nor U26419 (N_26419,N_24900,N_24936);
nand U26420 (N_26420,N_24459,N_25438);
nand U26421 (N_26421,N_24356,N_24876);
xor U26422 (N_26422,N_24207,N_24826);
or U26423 (N_26423,N_24959,N_24725);
nand U26424 (N_26424,N_24237,N_24210);
or U26425 (N_26425,N_25427,N_25256);
xnor U26426 (N_26426,N_24566,N_24844);
nand U26427 (N_26427,N_24990,N_24416);
and U26428 (N_26428,N_25485,N_24034);
nor U26429 (N_26429,N_24441,N_24092);
nor U26430 (N_26430,N_24726,N_25439);
nor U26431 (N_26431,N_24862,N_25308);
or U26432 (N_26432,N_25409,N_25429);
and U26433 (N_26433,N_24170,N_25477);
nand U26434 (N_26434,N_25025,N_24623);
and U26435 (N_26435,N_25145,N_25305);
xnor U26436 (N_26436,N_25381,N_24239);
or U26437 (N_26437,N_24498,N_24713);
and U26438 (N_26438,N_24405,N_25358);
nand U26439 (N_26439,N_24722,N_24645);
or U26440 (N_26440,N_24946,N_25021);
and U26441 (N_26441,N_24836,N_25234);
and U26442 (N_26442,N_24743,N_24887);
nand U26443 (N_26443,N_25090,N_25429);
nand U26444 (N_26444,N_24274,N_25036);
nand U26445 (N_26445,N_24706,N_25367);
and U26446 (N_26446,N_25118,N_24402);
nor U26447 (N_26447,N_24605,N_24609);
or U26448 (N_26448,N_24915,N_24475);
nand U26449 (N_26449,N_24095,N_24711);
and U26450 (N_26450,N_24182,N_24683);
and U26451 (N_26451,N_25393,N_24399);
and U26452 (N_26452,N_25044,N_25158);
xor U26453 (N_26453,N_25082,N_24608);
nor U26454 (N_26454,N_24766,N_24615);
or U26455 (N_26455,N_25059,N_25455);
xnor U26456 (N_26456,N_24397,N_24621);
nand U26457 (N_26457,N_24545,N_24252);
or U26458 (N_26458,N_25234,N_25409);
nor U26459 (N_26459,N_25036,N_25454);
nand U26460 (N_26460,N_24951,N_24884);
and U26461 (N_26461,N_25289,N_24893);
and U26462 (N_26462,N_25353,N_25034);
xor U26463 (N_26463,N_25265,N_25182);
and U26464 (N_26464,N_24905,N_24562);
nor U26465 (N_26465,N_25406,N_24709);
nand U26466 (N_26466,N_24418,N_25321);
nand U26467 (N_26467,N_25469,N_24829);
nand U26468 (N_26468,N_24287,N_24789);
nand U26469 (N_26469,N_25368,N_25097);
nor U26470 (N_26470,N_25039,N_25203);
and U26471 (N_26471,N_24121,N_24291);
and U26472 (N_26472,N_25052,N_24217);
nand U26473 (N_26473,N_24527,N_24998);
nand U26474 (N_26474,N_24222,N_24671);
nor U26475 (N_26475,N_24933,N_25153);
or U26476 (N_26476,N_24899,N_24301);
nor U26477 (N_26477,N_25216,N_24059);
xnor U26478 (N_26478,N_24574,N_24068);
nand U26479 (N_26479,N_24556,N_25458);
nand U26480 (N_26480,N_25261,N_25351);
nor U26481 (N_26481,N_24438,N_24123);
or U26482 (N_26482,N_25281,N_24050);
xnor U26483 (N_26483,N_24225,N_24233);
or U26484 (N_26484,N_25154,N_24615);
nor U26485 (N_26485,N_24055,N_24822);
and U26486 (N_26486,N_24872,N_24519);
nor U26487 (N_26487,N_24211,N_25198);
nand U26488 (N_26488,N_24272,N_24448);
and U26489 (N_26489,N_24231,N_25099);
nand U26490 (N_26490,N_24688,N_24988);
nor U26491 (N_26491,N_24605,N_24557);
or U26492 (N_26492,N_25323,N_24658);
or U26493 (N_26493,N_24337,N_25391);
xnor U26494 (N_26494,N_24850,N_24082);
nor U26495 (N_26495,N_25267,N_24116);
nand U26496 (N_26496,N_24404,N_24377);
xnor U26497 (N_26497,N_24672,N_25005);
xor U26498 (N_26498,N_24236,N_25348);
xor U26499 (N_26499,N_24652,N_24188);
xnor U26500 (N_26500,N_24359,N_24318);
xnor U26501 (N_26501,N_24461,N_24217);
or U26502 (N_26502,N_24880,N_25164);
or U26503 (N_26503,N_24651,N_25000);
or U26504 (N_26504,N_24559,N_25108);
xnor U26505 (N_26505,N_25336,N_24250);
nand U26506 (N_26506,N_24601,N_24600);
or U26507 (N_26507,N_24865,N_24490);
xnor U26508 (N_26508,N_24499,N_25363);
nand U26509 (N_26509,N_24171,N_24923);
xor U26510 (N_26510,N_25290,N_24980);
and U26511 (N_26511,N_24134,N_24760);
xor U26512 (N_26512,N_24649,N_25250);
nand U26513 (N_26513,N_25287,N_25449);
xor U26514 (N_26514,N_24145,N_24322);
xnor U26515 (N_26515,N_24078,N_24919);
nor U26516 (N_26516,N_25301,N_25466);
nand U26517 (N_26517,N_24445,N_24834);
nor U26518 (N_26518,N_25416,N_24885);
and U26519 (N_26519,N_24331,N_24892);
or U26520 (N_26520,N_25429,N_24896);
nand U26521 (N_26521,N_24360,N_24082);
or U26522 (N_26522,N_24549,N_24471);
and U26523 (N_26523,N_24992,N_24927);
nand U26524 (N_26524,N_24651,N_24586);
or U26525 (N_26525,N_25469,N_24550);
nor U26526 (N_26526,N_24782,N_24094);
xor U26527 (N_26527,N_24566,N_24407);
xnor U26528 (N_26528,N_25108,N_25313);
nand U26529 (N_26529,N_25469,N_24654);
xnor U26530 (N_26530,N_24501,N_24870);
xor U26531 (N_26531,N_24751,N_25276);
nor U26532 (N_26532,N_24010,N_25415);
xnor U26533 (N_26533,N_24299,N_24325);
nand U26534 (N_26534,N_25487,N_25481);
nand U26535 (N_26535,N_25165,N_24177);
and U26536 (N_26536,N_24742,N_24227);
or U26537 (N_26537,N_25065,N_24123);
and U26538 (N_26538,N_24421,N_24119);
nor U26539 (N_26539,N_24004,N_25178);
nor U26540 (N_26540,N_24339,N_24045);
nor U26541 (N_26541,N_24493,N_24917);
and U26542 (N_26542,N_24741,N_24410);
nand U26543 (N_26543,N_25252,N_25174);
or U26544 (N_26544,N_24465,N_24696);
xor U26545 (N_26545,N_24560,N_24402);
and U26546 (N_26546,N_24454,N_24772);
nand U26547 (N_26547,N_25428,N_24388);
xnor U26548 (N_26548,N_25229,N_25309);
and U26549 (N_26549,N_25240,N_25328);
nand U26550 (N_26550,N_25298,N_25362);
nor U26551 (N_26551,N_25112,N_25349);
nor U26552 (N_26552,N_24616,N_24167);
nand U26553 (N_26553,N_24173,N_24844);
nand U26554 (N_26554,N_24532,N_25491);
or U26555 (N_26555,N_25245,N_24165);
xnor U26556 (N_26556,N_24079,N_25299);
nor U26557 (N_26557,N_24425,N_25276);
nand U26558 (N_26558,N_24873,N_24105);
nand U26559 (N_26559,N_24304,N_24040);
and U26560 (N_26560,N_24668,N_25143);
and U26561 (N_26561,N_25483,N_24862);
nor U26562 (N_26562,N_24821,N_24692);
and U26563 (N_26563,N_24477,N_24940);
xor U26564 (N_26564,N_24680,N_24290);
nor U26565 (N_26565,N_24517,N_25399);
nand U26566 (N_26566,N_24271,N_24626);
or U26567 (N_26567,N_24866,N_24274);
or U26568 (N_26568,N_25268,N_24306);
nor U26569 (N_26569,N_24682,N_24721);
nand U26570 (N_26570,N_24710,N_25040);
and U26571 (N_26571,N_25136,N_24851);
nand U26572 (N_26572,N_24299,N_25435);
nor U26573 (N_26573,N_25139,N_24188);
nand U26574 (N_26574,N_24719,N_24180);
nand U26575 (N_26575,N_24874,N_24793);
nor U26576 (N_26576,N_24993,N_24785);
and U26577 (N_26577,N_25265,N_24699);
xnor U26578 (N_26578,N_24228,N_25135);
nand U26579 (N_26579,N_24887,N_24127);
and U26580 (N_26580,N_25103,N_25288);
xnor U26581 (N_26581,N_25169,N_24904);
or U26582 (N_26582,N_24649,N_24774);
and U26583 (N_26583,N_25025,N_24440);
nand U26584 (N_26584,N_24128,N_25418);
xor U26585 (N_26585,N_24930,N_24943);
xor U26586 (N_26586,N_24461,N_24013);
xor U26587 (N_26587,N_24317,N_24918);
nor U26588 (N_26588,N_24250,N_24641);
or U26589 (N_26589,N_25272,N_25271);
nor U26590 (N_26590,N_25070,N_24238);
or U26591 (N_26591,N_25494,N_25172);
nand U26592 (N_26592,N_24491,N_24055);
and U26593 (N_26593,N_24189,N_25205);
nand U26594 (N_26594,N_24771,N_24847);
or U26595 (N_26595,N_24390,N_24858);
nand U26596 (N_26596,N_24067,N_25180);
nand U26597 (N_26597,N_24015,N_24126);
and U26598 (N_26598,N_25352,N_25008);
or U26599 (N_26599,N_25110,N_25092);
or U26600 (N_26600,N_24451,N_24458);
nor U26601 (N_26601,N_24370,N_24961);
and U26602 (N_26602,N_24390,N_24833);
nand U26603 (N_26603,N_25302,N_25090);
xnor U26604 (N_26604,N_24041,N_24946);
nand U26605 (N_26605,N_24162,N_25478);
xor U26606 (N_26606,N_24749,N_24397);
nor U26607 (N_26607,N_25478,N_25176);
xnor U26608 (N_26608,N_25359,N_24402);
xnor U26609 (N_26609,N_25449,N_24948);
and U26610 (N_26610,N_24030,N_25203);
nand U26611 (N_26611,N_24104,N_24495);
and U26612 (N_26612,N_24069,N_24491);
nor U26613 (N_26613,N_24242,N_24415);
or U26614 (N_26614,N_24051,N_24642);
or U26615 (N_26615,N_24885,N_24362);
nand U26616 (N_26616,N_24567,N_24177);
or U26617 (N_26617,N_24621,N_24776);
or U26618 (N_26618,N_24004,N_24338);
or U26619 (N_26619,N_24135,N_24456);
nand U26620 (N_26620,N_25401,N_24287);
xnor U26621 (N_26621,N_24653,N_24198);
and U26622 (N_26622,N_24628,N_24898);
nand U26623 (N_26623,N_24936,N_24421);
or U26624 (N_26624,N_24725,N_25380);
nand U26625 (N_26625,N_24198,N_25256);
or U26626 (N_26626,N_25340,N_24733);
nor U26627 (N_26627,N_24496,N_24232);
and U26628 (N_26628,N_25005,N_25006);
or U26629 (N_26629,N_25456,N_25206);
nand U26630 (N_26630,N_24703,N_24726);
nand U26631 (N_26631,N_25149,N_24833);
nor U26632 (N_26632,N_24645,N_24888);
and U26633 (N_26633,N_25015,N_25244);
and U26634 (N_26634,N_24907,N_24353);
nand U26635 (N_26635,N_24324,N_24140);
xor U26636 (N_26636,N_24878,N_25418);
or U26637 (N_26637,N_24461,N_24660);
nor U26638 (N_26638,N_24566,N_24299);
nor U26639 (N_26639,N_24942,N_24028);
nand U26640 (N_26640,N_24985,N_24360);
xnor U26641 (N_26641,N_24658,N_24261);
nand U26642 (N_26642,N_25372,N_24596);
xnor U26643 (N_26643,N_24229,N_25036);
and U26644 (N_26644,N_25238,N_24946);
xor U26645 (N_26645,N_25316,N_24408);
and U26646 (N_26646,N_24840,N_25428);
xor U26647 (N_26647,N_25279,N_24162);
nor U26648 (N_26648,N_24022,N_25194);
xor U26649 (N_26649,N_24635,N_24118);
and U26650 (N_26650,N_25256,N_24413);
and U26651 (N_26651,N_25378,N_24324);
and U26652 (N_26652,N_25077,N_25489);
nor U26653 (N_26653,N_24479,N_24900);
and U26654 (N_26654,N_24648,N_24305);
nand U26655 (N_26655,N_25405,N_25240);
xor U26656 (N_26656,N_24776,N_24519);
xnor U26657 (N_26657,N_24391,N_24238);
nor U26658 (N_26658,N_25020,N_24693);
nand U26659 (N_26659,N_24760,N_25297);
nand U26660 (N_26660,N_24085,N_24772);
or U26661 (N_26661,N_24855,N_24909);
xnor U26662 (N_26662,N_24873,N_25032);
and U26663 (N_26663,N_24479,N_24308);
xnor U26664 (N_26664,N_25377,N_24593);
xnor U26665 (N_26665,N_24930,N_25086);
xnor U26666 (N_26666,N_24103,N_24294);
nor U26667 (N_26667,N_25263,N_24183);
or U26668 (N_26668,N_24235,N_25181);
and U26669 (N_26669,N_24162,N_24364);
and U26670 (N_26670,N_25029,N_24992);
or U26671 (N_26671,N_24627,N_24215);
nor U26672 (N_26672,N_24471,N_24334);
or U26673 (N_26673,N_24657,N_24443);
and U26674 (N_26674,N_24013,N_24119);
and U26675 (N_26675,N_24186,N_24269);
or U26676 (N_26676,N_24534,N_24336);
nand U26677 (N_26677,N_24876,N_25101);
nor U26678 (N_26678,N_25438,N_24764);
nand U26679 (N_26679,N_25324,N_24775);
or U26680 (N_26680,N_24418,N_24153);
and U26681 (N_26681,N_24828,N_24516);
nor U26682 (N_26682,N_24386,N_24279);
xnor U26683 (N_26683,N_25322,N_25314);
nor U26684 (N_26684,N_25235,N_25129);
nor U26685 (N_26685,N_24322,N_24767);
and U26686 (N_26686,N_25338,N_25456);
nand U26687 (N_26687,N_24881,N_24550);
nand U26688 (N_26688,N_24418,N_25319);
or U26689 (N_26689,N_25231,N_24288);
nor U26690 (N_26690,N_24629,N_25031);
nor U26691 (N_26691,N_24924,N_24853);
nand U26692 (N_26692,N_25272,N_24488);
nand U26693 (N_26693,N_25045,N_25163);
nor U26694 (N_26694,N_24566,N_25104);
or U26695 (N_26695,N_25389,N_24160);
nand U26696 (N_26696,N_25369,N_24382);
and U26697 (N_26697,N_24138,N_25337);
xnor U26698 (N_26698,N_24716,N_25360);
nor U26699 (N_26699,N_24357,N_24051);
nor U26700 (N_26700,N_25133,N_24644);
xnor U26701 (N_26701,N_25301,N_25199);
xnor U26702 (N_26702,N_24822,N_24133);
and U26703 (N_26703,N_24704,N_25255);
xor U26704 (N_26704,N_24624,N_25055);
xnor U26705 (N_26705,N_24105,N_24913);
and U26706 (N_26706,N_25470,N_24672);
xnor U26707 (N_26707,N_25197,N_24569);
nand U26708 (N_26708,N_24194,N_25089);
and U26709 (N_26709,N_25414,N_25158);
nor U26710 (N_26710,N_25315,N_24715);
nand U26711 (N_26711,N_25138,N_24233);
or U26712 (N_26712,N_25391,N_25481);
nand U26713 (N_26713,N_24928,N_24860);
and U26714 (N_26714,N_24247,N_24715);
and U26715 (N_26715,N_25240,N_24703);
xnor U26716 (N_26716,N_24620,N_24376);
nor U26717 (N_26717,N_25000,N_25287);
xor U26718 (N_26718,N_24486,N_24736);
xnor U26719 (N_26719,N_24465,N_24946);
or U26720 (N_26720,N_25297,N_24275);
and U26721 (N_26721,N_24852,N_24041);
xnor U26722 (N_26722,N_25277,N_25031);
or U26723 (N_26723,N_25366,N_25234);
and U26724 (N_26724,N_24391,N_24433);
nand U26725 (N_26725,N_25027,N_25322);
or U26726 (N_26726,N_25133,N_24101);
nor U26727 (N_26727,N_25291,N_24731);
nand U26728 (N_26728,N_24149,N_25448);
xnor U26729 (N_26729,N_24202,N_25003);
or U26730 (N_26730,N_25172,N_24956);
nor U26731 (N_26731,N_24761,N_24467);
xnor U26732 (N_26732,N_24783,N_24392);
nand U26733 (N_26733,N_24770,N_24101);
nand U26734 (N_26734,N_24500,N_24880);
nand U26735 (N_26735,N_24503,N_25087);
xnor U26736 (N_26736,N_24002,N_25466);
nand U26737 (N_26737,N_25265,N_24831);
nand U26738 (N_26738,N_24693,N_24308);
nand U26739 (N_26739,N_24678,N_24620);
and U26740 (N_26740,N_24687,N_24904);
nor U26741 (N_26741,N_25030,N_24978);
xnor U26742 (N_26742,N_25434,N_24532);
xnor U26743 (N_26743,N_24966,N_24676);
xor U26744 (N_26744,N_24956,N_25000);
nor U26745 (N_26745,N_24225,N_24515);
xor U26746 (N_26746,N_24974,N_24429);
xnor U26747 (N_26747,N_25362,N_25460);
and U26748 (N_26748,N_25264,N_25305);
and U26749 (N_26749,N_25485,N_24962);
nand U26750 (N_26750,N_24169,N_24726);
xnor U26751 (N_26751,N_24967,N_25149);
xor U26752 (N_26752,N_24199,N_25379);
or U26753 (N_26753,N_25140,N_24699);
and U26754 (N_26754,N_24435,N_24341);
nor U26755 (N_26755,N_24056,N_24368);
nor U26756 (N_26756,N_24476,N_24141);
nand U26757 (N_26757,N_25145,N_24031);
nor U26758 (N_26758,N_24587,N_24944);
or U26759 (N_26759,N_24223,N_25140);
nand U26760 (N_26760,N_24759,N_24851);
or U26761 (N_26761,N_24111,N_24069);
or U26762 (N_26762,N_24409,N_25495);
nor U26763 (N_26763,N_25332,N_25099);
nand U26764 (N_26764,N_24093,N_24177);
xnor U26765 (N_26765,N_24733,N_24136);
nor U26766 (N_26766,N_24819,N_24751);
nor U26767 (N_26767,N_24300,N_25415);
xnor U26768 (N_26768,N_25149,N_24097);
nor U26769 (N_26769,N_24795,N_25321);
and U26770 (N_26770,N_24956,N_25002);
nor U26771 (N_26771,N_24511,N_24113);
nand U26772 (N_26772,N_24969,N_24653);
nand U26773 (N_26773,N_24648,N_24566);
or U26774 (N_26774,N_24278,N_24641);
nand U26775 (N_26775,N_24117,N_24968);
or U26776 (N_26776,N_24114,N_24630);
nor U26777 (N_26777,N_25042,N_24034);
nand U26778 (N_26778,N_24338,N_24113);
nor U26779 (N_26779,N_24900,N_24117);
or U26780 (N_26780,N_24502,N_24610);
and U26781 (N_26781,N_25498,N_24825);
xnor U26782 (N_26782,N_24036,N_24144);
nand U26783 (N_26783,N_24587,N_24089);
and U26784 (N_26784,N_25088,N_24654);
nand U26785 (N_26785,N_25025,N_24966);
nand U26786 (N_26786,N_24111,N_24706);
and U26787 (N_26787,N_24709,N_24633);
nand U26788 (N_26788,N_25064,N_25382);
and U26789 (N_26789,N_24815,N_24103);
and U26790 (N_26790,N_24449,N_24457);
and U26791 (N_26791,N_24238,N_24150);
nor U26792 (N_26792,N_25328,N_25146);
nand U26793 (N_26793,N_25088,N_24848);
nor U26794 (N_26794,N_25389,N_25331);
nand U26795 (N_26795,N_25491,N_24722);
and U26796 (N_26796,N_25359,N_25175);
xnor U26797 (N_26797,N_25184,N_24409);
xnor U26798 (N_26798,N_25212,N_25000);
and U26799 (N_26799,N_24429,N_24936);
nor U26800 (N_26800,N_25295,N_25481);
xor U26801 (N_26801,N_25250,N_24544);
or U26802 (N_26802,N_24712,N_24418);
nand U26803 (N_26803,N_24653,N_24183);
nand U26804 (N_26804,N_24602,N_24654);
nand U26805 (N_26805,N_24881,N_24990);
xnor U26806 (N_26806,N_25277,N_25034);
xnor U26807 (N_26807,N_24885,N_24808);
nand U26808 (N_26808,N_25077,N_24523);
or U26809 (N_26809,N_24030,N_25257);
nand U26810 (N_26810,N_25375,N_24968);
nand U26811 (N_26811,N_24300,N_24816);
nor U26812 (N_26812,N_24580,N_25354);
xor U26813 (N_26813,N_24051,N_24527);
nor U26814 (N_26814,N_24539,N_24511);
xor U26815 (N_26815,N_24033,N_24410);
nand U26816 (N_26816,N_24517,N_25324);
nor U26817 (N_26817,N_24356,N_24090);
nor U26818 (N_26818,N_24119,N_25483);
and U26819 (N_26819,N_24011,N_24805);
xnor U26820 (N_26820,N_25004,N_25316);
and U26821 (N_26821,N_24663,N_24307);
xor U26822 (N_26822,N_24455,N_25492);
xnor U26823 (N_26823,N_24024,N_24323);
xor U26824 (N_26824,N_24306,N_24086);
xor U26825 (N_26825,N_25426,N_24224);
nand U26826 (N_26826,N_24399,N_24157);
nor U26827 (N_26827,N_24925,N_24962);
and U26828 (N_26828,N_24635,N_25451);
nor U26829 (N_26829,N_25355,N_24638);
xor U26830 (N_26830,N_24407,N_24592);
and U26831 (N_26831,N_25386,N_24724);
nand U26832 (N_26832,N_24172,N_25260);
xor U26833 (N_26833,N_24614,N_24592);
xor U26834 (N_26834,N_25384,N_25225);
and U26835 (N_26835,N_25090,N_25456);
nor U26836 (N_26836,N_24378,N_24248);
and U26837 (N_26837,N_24194,N_24058);
or U26838 (N_26838,N_24855,N_24763);
nor U26839 (N_26839,N_24195,N_25103);
nor U26840 (N_26840,N_25108,N_25269);
nor U26841 (N_26841,N_25397,N_24497);
nor U26842 (N_26842,N_24003,N_24796);
nand U26843 (N_26843,N_24325,N_25070);
or U26844 (N_26844,N_25389,N_24923);
nor U26845 (N_26845,N_24178,N_24246);
or U26846 (N_26846,N_24080,N_24633);
or U26847 (N_26847,N_24113,N_24868);
nor U26848 (N_26848,N_24835,N_24603);
and U26849 (N_26849,N_24928,N_24603);
nor U26850 (N_26850,N_24327,N_25226);
and U26851 (N_26851,N_24764,N_25376);
nand U26852 (N_26852,N_24508,N_25425);
xor U26853 (N_26853,N_24964,N_25308);
xor U26854 (N_26854,N_24539,N_24182);
nand U26855 (N_26855,N_24966,N_25244);
nand U26856 (N_26856,N_25351,N_25006);
or U26857 (N_26857,N_25422,N_24546);
xnor U26858 (N_26858,N_25465,N_25174);
nand U26859 (N_26859,N_24530,N_24152);
nand U26860 (N_26860,N_24722,N_25039);
nor U26861 (N_26861,N_24696,N_24944);
xnor U26862 (N_26862,N_24524,N_24307);
and U26863 (N_26863,N_25413,N_25278);
nor U26864 (N_26864,N_24140,N_24386);
nor U26865 (N_26865,N_24035,N_25434);
and U26866 (N_26866,N_25278,N_24090);
xnor U26867 (N_26867,N_24279,N_24145);
nor U26868 (N_26868,N_24699,N_24000);
and U26869 (N_26869,N_24342,N_24247);
or U26870 (N_26870,N_24757,N_24755);
nand U26871 (N_26871,N_24166,N_24084);
xnor U26872 (N_26872,N_25052,N_24589);
xnor U26873 (N_26873,N_24910,N_24445);
nand U26874 (N_26874,N_25395,N_25316);
or U26875 (N_26875,N_24286,N_24878);
or U26876 (N_26876,N_24816,N_25069);
nor U26877 (N_26877,N_24406,N_24775);
nand U26878 (N_26878,N_25348,N_24495);
xor U26879 (N_26879,N_25206,N_24046);
xnor U26880 (N_26880,N_25337,N_25026);
nand U26881 (N_26881,N_25097,N_25370);
or U26882 (N_26882,N_25269,N_25186);
nand U26883 (N_26883,N_25262,N_24530);
and U26884 (N_26884,N_25404,N_24038);
nand U26885 (N_26885,N_24291,N_25266);
nor U26886 (N_26886,N_24636,N_24242);
nor U26887 (N_26887,N_24298,N_24608);
nor U26888 (N_26888,N_24823,N_25037);
and U26889 (N_26889,N_24871,N_25311);
and U26890 (N_26890,N_24948,N_24249);
nor U26891 (N_26891,N_24871,N_24778);
nor U26892 (N_26892,N_25084,N_25317);
xor U26893 (N_26893,N_24599,N_25121);
nor U26894 (N_26894,N_25156,N_24529);
and U26895 (N_26895,N_25009,N_24964);
nand U26896 (N_26896,N_24843,N_25002);
nand U26897 (N_26897,N_24025,N_25457);
and U26898 (N_26898,N_24574,N_24900);
and U26899 (N_26899,N_25397,N_25462);
and U26900 (N_26900,N_24904,N_25043);
nor U26901 (N_26901,N_24777,N_24195);
nor U26902 (N_26902,N_24458,N_24614);
and U26903 (N_26903,N_24825,N_24987);
or U26904 (N_26904,N_25420,N_25448);
xnor U26905 (N_26905,N_24387,N_25447);
or U26906 (N_26906,N_24792,N_24775);
nor U26907 (N_26907,N_24689,N_24065);
nand U26908 (N_26908,N_24569,N_24212);
xnor U26909 (N_26909,N_24769,N_24914);
nor U26910 (N_26910,N_24303,N_25236);
nor U26911 (N_26911,N_24405,N_24803);
xnor U26912 (N_26912,N_25180,N_24211);
nand U26913 (N_26913,N_24097,N_25360);
and U26914 (N_26914,N_24196,N_24043);
or U26915 (N_26915,N_24420,N_24211);
xnor U26916 (N_26916,N_25282,N_24935);
and U26917 (N_26917,N_24617,N_24223);
or U26918 (N_26918,N_24397,N_24922);
and U26919 (N_26919,N_24055,N_24371);
nor U26920 (N_26920,N_24845,N_25121);
nand U26921 (N_26921,N_25404,N_24916);
xor U26922 (N_26922,N_25083,N_24496);
nand U26923 (N_26923,N_24031,N_24977);
xnor U26924 (N_26924,N_25314,N_24324);
nor U26925 (N_26925,N_25346,N_24430);
xnor U26926 (N_26926,N_25450,N_24521);
or U26927 (N_26927,N_24409,N_24444);
nor U26928 (N_26928,N_25478,N_24033);
and U26929 (N_26929,N_25278,N_24624);
and U26930 (N_26930,N_25345,N_24141);
nor U26931 (N_26931,N_25208,N_24079);
or U26932 (N_26932,N_24204,N_25015);
and U26933 (N_26933,N_24533,N_25269);
and U26934 (N_26934,N_24119,N_24494);
xnor U26935 (N_26935,N_24646,N_25453);
xnor U26936 (N_26936,N_24896,N_24973);
or U26937 (N_26937,N_24761,N_24107);
nor U26938 (N_26938,N_24648,N_24251);
xnor U26939 (N_26939,N_25041,N_25149);
xor U26940 (N_26940,N_24187,N_24002);
and U26941 (N_26941,N_24097,N_24811);
or U26942 (N_26942,N_24243,N_25183);
nand U26943 (N_26943,N_24981,N_24366);
nor U26944 (N_26944,N_24715,N_24320);
nor U26945 (N_26945,N_25236,N_24772);
nor U26946 (N_26946,N_24819,N_24149);
nor U26947 (N_26947,N_24276,N_25091);
xnor U26948 (N_26948,N_24670,N_24873);
nor U26949 (N_26949,N_24565,N_24266);
nand U26950 (N_26950,N_24774,N_25015);
and U26951 (N_26951,N_24163,N_24365);
xnor U26952 (N_26952,N_25074,N_24508);
nor U26953 (N_26953,N_24602,N_25232);
nor U26954 (N_26954,N_24659,N_25201);
or U26955 (N_26955,N_24863,N_24829);
nor U26956 (N_26956,N_25279,N_24767);
and U26957 (N_26957,N_24416,N_24240);
nand U26958 (N_26958,N_25290,N_24303);
or U26959 (N_26959,N_25028,N_24398);
nand U26960 (N_26960,N_24207,N_24147);
nand U26961 (N_26961,N_25173,N_24671);
and U26962 (N_26962,N_25284,N_24309);
nor U26963 (N_26963,N_25008,N_24984);
nand U26964 (N_26964,N_25015,N_24296);
nor U26965 (N_26965,N_25015,N_24002);
xnor U26966 (N_26966,N_24947,N_25402);
and U26967 (N_26967,N_24443,N_25204);
nor U26968 (N_26968,N_25471,N_24258);
xor U26969 (N_26969,N_25172,N_24078);
nor U26970 (N_26970,N_24749,N_24531);
or U26971 (N_26971,N_24714,N_25015);
nor U26972 (N_26972,N_25391,N_24114);
xnor U26973 (N_26973,N_25281,N_25096);
nand U26974 (N_26974,N_24621,N_24634);
and U26975 (N_26975,N_24560,N_24941);
or U26976 (N_26976,N_25412,N_25279);
nor U26977 (N_26977,N_24314,N_25190);
nor U26978 (N_26978,N_24384,N_24125);
xnor U26979 (N_26979,N_25410,N_24060);
nor U26980 (N_26980,N_24581,N_25496);
nor U26981 (N_26981,N_25231,N_24560);
xor U26982 (N_26982,N_24005,N_24519);
and U26983 (N_26983,N_25422,N_25402);
nor U26984 (N_26984,N_25446,N_25070);
nor U26985 (N_26985,N_24983,N_25397);
nor U26986 (N_26986,N_25203,N_24844);
nand U26987 (N_26987,N_24980,N_24575);
nand U26988 (N_26988,N_24980,N_24286);
nor U26989 (N_26989,N_25396,N_24144);
or U26990 (N_26990,N_24362,N_25220);
nor U26991 (N_26991,N_24220,N_25048);
nand U26992 (N_26992,N_24126,N_24028);
or U26993 (N_26993,N_24354,N_24245);
nor U26994 (N_26994,N_24126,N_24014);
or U26995 (N_26995,N_24497,N_24511);
xnor U26996 (N_26996,N_25085,N_25007);
nor U26997 (N_26997,N_24500,N_24545);
and U26998 (N_26998,N_24497,N_24372);
nand U26999 (N_26999,N_25249,N_25312);
and U27000 (N_27000,N_25649,N_26322);
nand U27001 (N_27001,N_26031,N_26096);
or U27002 (N_27002,N_25524,N_26425);
nand U27003 (N_27003,N_26368,N_26810);
nand U27004 (N_27004,N_25951,N_25804);
xor U27005 (N_27005,N_25675,N_26806);
nor U27006 (N_27006,N_26450,N_26674);
nor U27007 (N_27007,N_26835,N_26558);
or U27008 (N_27008,N_26588,N_26258);
nand U27009 (N_27009,N_26132,N_25686);
nand U27010 (N_27010,N_26242,N_25859);
xnor U27011 (N_27011,N_25693,N_26771);
or U27012 (N_27012,N_25714,N_25657);
or U27013 (N_27013,N_25729,N_26761);
xor U27014 (N_27014,N_26758,N_25909);
nor U27015 (N_27015,N_26897,N_26195);
xor U27016 (N_27016,N_26623,N_26513);
nor U27017 (N_27017,N_25728,N_25758);
xor U27018 (N_27018,N_25790,N_26615);
and U27019 (N_27019,N_26082,N_25533);
and U27020 (N_27020,N_26312,N_26553);
nand U27021 (N_27021,N_25960,N_26780);
and U27022 (N_27022,N_26916,N_25803);
and U27023 (N_27023,N_26966,N_25969);
or U27024 (N_27024,N_26795,N_26607);
xnor U27025 (N_27025,N_26975,N_25864);
nand U27026 (N_27026,N_26052,N_25702);
xnor U27027 (N_27027,N_26300,N_26363);
nand U27028 (N_27028,N_26816,N_26945);
nand U27029 (N_27029,N_26011,N_25906);
or U27030 (N_27030,N_26716,N_26562);
or U27031 (N_27031,N_26023,N_26579);
or U27032 (N_27032,N_25927,N_26569);
xor U27033 (N_27033,N_26419,N_26114);
nand U27034 (N_27034,N_26934,N_26888);
xor U27035 (N_27035,N_25796,N_25822);
nand U27036 (N_27036,N_26825,N_25881);
nand U27037 (N_27037,N_26552,N_26302);
xnor U27038 (N_27038,N_25833,N_26755);
nor U27039 (N_27039,N_25625,N_26701);
xor U27040 (N_27040,N_26563,N_26141);
xnor U27041 (N_27041,N_25886,N_25501);
xor U27042 (N_27042,N_26105,N_25628);
and U27043 (N_27043,N_26746,N_26478);
xnor U27044 (N_27044,N_26064,N_26852);
or U27045 (N_27045,N_26894,N_25579);
and U27046 (N_27046,N_26467,N_26914);
nor U27047 (N_27047,N_26753,N_26734);
and U27048 (N_27048,N_25954,N_25615);
or U27049 (N_27049,N_26048,N_26702);
and U27050 (N_27050,N_26620,N_25908);
nor U27051 (N_27051,N_25868,N_26338);
or U27052 (N_27052,N_26913,N_25654);
and U27053 (N_27053,N_26800,N_26733);
nor U27054 (N_27054,N_26074,N_26386);
xnor U27055 (N_27055,N_26005,N_26546);
and U27056 (N_27056,N_25737,N_26261);
and U27057 (N_27057,N_26818,N_26308);
nor U27058 (N_27058,N_26775,N_25583);
and U27059 (N_27059,N_26347,N_26687);
or U27060 (N_27060,N_26677,N_26531);
xor U27061 (N_27061,N_25571,N_25716);
or U27062 (N_27062,N_26429,N_25554);
xor U27063 (N_27063,N_25616,N_25867);
or U27064 (N_27064,N_26785,N_25592);
and U27065 (N_27065,N_26067,N_26808);
xnor U27066 (N_27066,N_26613,N_25650);
or U27067 (N_27067,N_26045,N_26221);
nand U27068 (N_27068,N_26153,N_26967);
xor U27069 (N_27069,N_26471,N_25919);
xnor U27070 (N_27070,N_25638,N_26621);
xor U27071 (N_27071,N_26051,N_26381);
nor U27072 (N_27072,N_26596,N_26653);
nand U27073 (N_27073,N_26255,N_25523);
nor U27074 (N_27074,N_25690,N_26732);
or U27075 (N_27075,N_25560,N_25842);
nor U27076 (N_27076,N_26744,N_26159);
xnor U27077 (N_27077,N_25752,N_26629);
nor U27078 (N_27078,N_26151,N_26044);
and U27079 (N_27079,N_26047,N_26887);
xnor U27080 (N_27080,N_26181,N_26752);
or U27081 (N_27081,N_26112,N_26778);
and U27082 (N_27082,N_26512,N_25931);
nor U27083 (N_27083,N_25572,N_26335);
and U27084 (N_27084,N_26978,N_26747);
nor U27085 (N_27085,N_26605,N_25713);
xor U27086 (N_27086,N_26526,N_25839);
xnor U27087 (N_27087,N_26352,N_26126);
nor U27088 (N_27088,N_26174,N_25725);
and U27089 (N_27089,N_26110,N_26911);
nor U27090 (N_27090,N_26492,N_25609);
xor U27091 (N_27091,N_25860,N_25639);
nand U27092 (N_27092,N_26533,N_25613);
or U27093 (N_27093,N_26509,N_26594);
xor U27094 (N_27094,N_25603,N_25514);
xor U27095 (N_27095,N_26718,N_25551);
and U27096 (N_27096,N_25937,N_26831);
nor U27097 (N_27097,N_26224,N_25669);
or U27098 (N_27098,N_26092,N_26198);
or U27099 (N_27099,N_25807,N_26611);
nor U27100 (N_27100,N_25917,N_26942);
nor U27101 (N_27101,N_25597,N_25971);
and U27102 (N_27102,N_25968,N_26903);
or U27103 (N_27103,N_26864,N_25838);
nor U27104 (N_27104,N_26637,N_26267);
nand U27105 (N_27105,N_26402,N_26560);
nor U27106 (N_27106,N_26028,N_26684);
xor U27107 (N_27107,N_26869,N_25990);
nand U27108 (N_27108,N_26061,N_26150);
xnor U27109 (N_27109,N_26206,N_26749);
nor U27110 (N_27110,N_26729,N_26708);
nor U27111 (N_27111,N_26403,N_26043);
xor U27112 (N_27112,N_26129,N_25707);
nor U27113 (N_27113,N_26644,N_25573);
nor U27114 (N_27114,N_26703,N_25832);
xnor U27115 (N_27115,N_25517,N_26514);
and U27116 (N_27116,N_26668,N_26090);
xor U27117 (N_27117,N_26858,N_26976);
nor U27118 (N_27118,N_26254,N_25903);
and U27119 (N_27119,N_26511,N_25784);
or U27120 (N_27120,N_25935,N_25594);
nand U27121 (N_27121,N_26275,N_26573);
or U27122 (N_27122,N_25856,N_25930);
nor U27123 (N_27123,N_25634,N_26669);
or U27124 (N_27124,N_25742,N_26710);
or U27125 (N_27125,N_25862,N_25845);
or U27126 (N_27126,N_25586,N_26582);
nor U27127 (N_27127,N_25595,N_26360);
nor U27128 (N_27128,N_26139,N_26018);
or U27129 (N_27129,N_26446,N_26457);
nor U27130 (N_27130,N_25801,N_25943);
or U27131 (N_27131,N_26544,N_26963);
and U27132 (N_27132,N_26086,N_26134);
and U27133 (N_27133,N_26177,N_26040);
xnor U27134 (N_27134,N_26205,N_26801);
nand U27135 (N_27135,N_25774,N_26304);
nand U27136 (N_27136,N_25827,N_26252);
and U27137 (N_27137,N_25666,N_25630);
and U27138 (N_27138,N_26237,N_26824);
nand U27139 (N_27139,N_26458,N_26279);
and U27140 (N_27140,N_26476,N_26313);
nand U27141 (N_27141,N_26422,N_26161);
nand U27142 (N_27142,N_26971,N_26367);
or U27143 (N_27143,N_26699,N_26389);
nor U27144 (N_27144,N_26010,N_26572);
xnor U27145 (N_27145,N_26507,N_26690);
and U27146 (N_27146,N_25948,N_25944);
or U27147 (N_27147,N_26245,N_25622);
and U27148 (N_27148,N_26137,N_25667);
or U27149 (N_27149,N_26902,N_26664);
or U27150 (N_27150,N_26575,N_26543);
and U27151 (N_27151,N_26817,N_26420);
nand U27152 (N_27152,N_26413,N_26626);
nand U27153 (N_27153,N_26953,N_26996);
xor U27154 (N_27154,N_26366,N_26763);
xor U27155 (N_27155,N_26908,N_26408);
or U27156 (N_27156,N_25763,N_26901);
nand U27157 (N_27157,N_26889,N_25826);
xnor U27158 (N_27158,N_25769,N_26979);
nand U27159 (N_27159,N_25522,N_26676);
nor U27160 (N_27160,N_26577,N_25687);
xor U27161 (N_27161,N_25646,N_26827);
and U27162 (N_27162,N_26004,N_26293);
xor U27163 (N_27163,N_26303,N_26548);
nand U27164 (N_27164,N_26725,N_26529);
or U27165 (N_27165,N_26097,N_26324);
and U27166 (N_27166,N_26371,N_26528);
nand U27167 (N_27167,N_26461,N_26712);
or U27168 (N_27168,N_26019,N_26649);
nand U27169 (N_27169,N_25670,N_26483);
or U27170 (N_27170,N_26223,N_25880);
nand U27171 (N_27171,N_25961,N_26183);
and U27172 (N_27172,N_26997,N_26355);
nor U27173 (N_27173,N_26142,N_26886);
or U27174 (N_27174,N_25818,N_25797);
xnor U27175 (N_27175,N_26792,N_26549);
nand U27176 (N_27176,N_26344,N_25815);
nand U27177 (N_27177,N_25734,N_26845);
nand U27178 (N_27178,N_26789,N_25976);
nor U27179 (N_27179,N_26186,N_25738);
or U27180 (N_27180,N_25962,N_25888);
nor U27181 (N_27181,N_25636,N_26091);
nand U27182 (N_27182,N_25889,N_26737);
or U27183 (N_27183,N_25882,N_26017);
or U27184 (N_27184,N_26561,N_26197);
xnor U27185 (N_27185,N_25967,N_26700);
and U27186 (N_27186,N_25910,N_25879);
nor U27187 (N_27187,N_26826,N_25559);
xor U27188 (N_27188,N_25662,N_26525);
and U27189 (N_27189,N_25537,N_25788);
nor U27190 (N_27190,N_26730,N_25525);
nand U27191 (N_27191,N_26000,N_26459);
nor U27192 (N_27192,N_26984,N_25538);
or U27193 (N_27193,N_26839,N_26414);
xor U27194 (N_27194,N_26184,N_26229);
nor U27195 (N_27195,N_25898,N_25979);
xnor U27196 (N_27196,N_26791,N_25664);
xor U27197 (N_27197,N_26247,N_26076);
nor U27198 (N_27198,N_26524,N_26833);
nand U27199 (N_27199,N_26609,N_26170);
nor U27200 (N_27200,N_26078,N_26297);
nand U27201 (N_27201,N_26962,N_26745);
and U27202 (N_27202,N_25706,N_25964);
xor U27203 (N_27203,N_26176,N_25743);
or U27204 (N_27204,N_26965,N_26721);
nand U27205 (N_27205,N_25590,N_26557);
or U27206 (N_27206,N_26204,N_25683);
xor U27207 (N_27207,N_26365,N_26764);
xnor U27208 (N_27208,N_26675,N_25697);
nor U27209 (N_27209,N_26390,N_26309);
nand U27210 (N_27210,N_25539,N_26412);
nor U27211 (N_27211,N_26372,N_25656);
or U27212 (N_27212,N_25722,N_26072);
or U27213 (N_27213,N_26906,N_26578);
nor U27214 (N_27214,N_26647,N_26416);
or U27215 (N_27215,N_26713,N_26232);
nor U27216 (N_27216,N_26188,N_25565);
or U27217 (N_27217,N_26027,N_26638);
or U27218 (N_27218,N_25527,N_25869);
xor U27219 (N_27219,N_25610,N_26940);
nor U27220 (N_27220,N_26504,N_26583);
nor U27221 (N_27221,N_26838,N_25512);
nor U27222 (N_27222,N_25721,N_25781);
nand U27223 (N_27223,N_25543,N_26014);
nand U27224 (N_27224,N_26180,N_25849);
and U27225 (N_27225,N_25791,N_25509);
nor U27226 (N_27226,N_26571,N_26256);
and U27227 (N_27227,N_25934,N_25552);
or U27228 (N_27228,N_26735,N_25651);
xnor U27229 (N_27229,N_26603,N_26325);
nor U27230 (N_27230,N_26738,N_26337);
xor U27231 (N_27231,N_26954,N_25566);
nor U27232 (N_27232,N_26301,N_26207);
and U27233 (N_27233,N_26270,N_26681);
and U27234 (N_27234,N_26427,N_26632);
nor U27235 (N_27235,N_25692,N_26794);
or U27236 (N_27236,N_26415,N_26821);
nor U27237 (N_27237,N_25553,N_26505);
nand U27238 (N_27238,N_26147,N_26099);
nor U27239 (N_27239,N_26958,N_25837);
xnor U27240 (N_27240,N_25872,N_25870);
or U27241 (N_27241,N_26506,N_26931);
nor U27242 (N_27242,N_26722,N_26202);
nor U27243 (N_27243,N_25907,N_25762);
and U27244 (N_27244,N_26863,N_25759);
or U27245 (N_27245,N_25998,N_26284);
nand U27246 (N_27246,N_26726,N_26435);
xnor U27247 (N_27247,N_25751,N_26243);
xor U27248 (N_27248,N_26597,N_26369);
xor U27249 (N_27249,N_26570,N_26989);
nand U27250 (N_27250,N_25732,N_26881);
nor U27251 (N_27251,N_26269,N_26055);
nand U27252 (N_27252,N_26073,N_26554);
xnor U27253 (N_27253,N_25808,N_26253);
and U27254 (N_27254,N_25782,N_26015);
xor U27255 (N_27255,N_26862,N_25585);
xnor U27256 (N_27256,N_25956,N_25526);
nor U27257 (N_27257,N_25545,N_25760);
xor U27258 (N_27258,N_26728,N_25618);
or U27259 (N_27259,N_26399,N_25581);
nor U27260 (N_27260,N_25564,N_26282);
xnor U27261 (N_27261,N_25661,N_25891);
nand U27262 (N_27262,N_26537,N_26037);
or U27263 (N_27263,N_26547,N_26851);
or U27264 (N_27264,N_26711,N_26782);
nand U27265 (N_27265,N_25865,N_25711);
nand U27266 (N_27266,N_26670,N_25733);
and U27267 (N_27267,N_25946,N_26316);
and U27268 (N_27268,N_26083,N_26550);
xor U27269 (N_27269,N_25556,N_25761);
or U27270 (N_27270,N_26856,N_26009);
xor U27271 (N_27271,N_26306,N_26356);
xnor U27272 (N_27272,N_26883,N_26036);
nand U27273 (N_27273,N_26465,N_26235);
nand U27274 (N_27274,N_25939,N_26790);
nor U27275 (N_27275,N_26636,N_26832);
nor U27276 (N_27276,N_25911,N_25720);
nor U27277 (N_27277,N_26030,N_26811);
or U27278 (N_27278,N_25570,N_26380);
xnor U27279 (N_27279,N_26006,N_26166);
and U27280 (N_27280,N_26796,N_26251);
nand U27281 (N_27281,N_26918,N_25994);
or U27282 (N_27282,N_26828,N_26264);
nor U27283 (N_27283,N_26317,N_25705);
and U27284 (N_27284,N_25844,N_25970);
xor U27285 (N_27285,N_25643,N_25633);
and U27286 (N_27286,N_26364,N_26591);
nand U27287 (N_27287,N_26879,N_26323);
or U27288 (N_27288,N_25812,N_26145);
nor U27289 (N_27289,N_25749,N_25996);
xor U27290 (N_27290,N_25647,N_26622);
xor U27291 (N_27291,N_26330,N_26157);
nor U27292 (N_27292,N_26873,N_26665);
or U27293 (N_27293,N_26936,N_25982);
nand U27294 (N_27294,N_25938,N_26717);
nand U27295 (N_27295,N_26119,N_25668);
and U27296 (N_27296,N_25770,N_26799);
nand U27297 (N_27297,N_25519,N_26238);
and U27298 (N_27298,N_26941,N_26651);
nor U27299 (N_27299,N_26866,N_26395);
nor U27300 (N_27300,N_26107,N_25850);
and U27301 (N_27301,N_26236,N_26510);
and U27302 (N_27302,N_26760,N_26213);
or U27303 (N_27303,N_25699,N_26877);
and U27304 (N_27304,N_26035,N_26248);
or U27305 (N_27305,N_26766,N_26436);
nor U27306 (N_27306,N_25975,N_25847);
nor U27307 (N_27307,N_25671,N_26156);
xnor U27308 (N_27308,N_26714,N_25767);
nand U27309 (N_27309,N_25963,N_26663);
or U27310 (N_27310,N_26567,N_25775);
nand U27311 (N_27311,N_26508,N_26468);
nand U27312 (N_27312,N_26972,N_25723);
and U27313 (N_27313,N_26391,N_26336);
or U27314 (N_27314,N_25730,N_25768);
and U27315 (N_27315,N_25875,N_26853);
nand U27316 (N_27316,N_26100,N_25981);
nor U27317 (N_27317,N_26441,N_26750);
nor U27318 (N_27318,N_26946,N_26173);
and U27319 (N_27319,N_26590,N_26884);
nand U27320 (N_27320,N_26757,N_26085);
nand U27321 (N_27321,N_26421,N_25606);
xnor U27322 (N_27322,N_26397,N_26354);
nand U27323 (N_27323,N_25952,N_26034);
nor U27324 (N_27324,N_26612,N_26444);
and U27325 (N_27325,N_25562,N_26103);
or U27326 (N_27326,N_26784,N_25915);
or U27327 (N_27327,N_26163,N_25648);
xnor U27328 (N_27328,N_25718,N_26185);
and U27329 (N_27329,N_26053,N_26350);
and U27330 (N_27330,N_25724,N_25793);
nand U27331 (N_27331,N_25691,N_25695);
nand U27332 (N_27332,N_26230,N_26199);
or U27333 (N_27333,N_26502,N_26109);
nand U27334 (N_27334,N_25698,N_26809);
nor U27335 (N_27335,N_25776,N_26069);
nor U27336 (N_27336,N_26219,N_26409);
and U27337 (N_27337,N_26374,N_26830);
xnor U27338 (N_27338,N_26585,N_25641);
xor U27339 (N_27339,N_25811,N_26541);
xnor U27340 (N_27340,N_26277,N_26222);
xor U27341 (N_27341,N_26305,N_26334);
nand U27342 (N_27342,N_26359,N_26228);
or U27343 (N_27343,N_25995,N_26262);
or U27344 (N_27344,N_26949,N_26379);
nor U27345 (N_27345,N_26731,N_25629);
nor U27346 (N_27346,N_26298,N_26475);
nor U27347 (N_27347,N_26280,N_26898);
or U27348 (N_27348,N_25905,N_26606);
nand U27349 (N_27349,N_26981,N_25973);
or U27350 (N_27350,N_25694,N_26445);
or U27351 (N_27351,N_26342,N_26314);
xor U27352 (N_27352,N_26628,N_26278);
and U27353 (N_27353,N_26307,N_25805);
and U27354 (N_27354,N_26233,N_26754);
and U27355 (N_27355,N_25861,N_25569);
nand U27356 (N_27356,N_25852,N_26633);
nor U27357 (N_27357,N_26417,N_26060);
and U27358 (N_27358,N_25999,N_26892);
or U27359 (N_27359,N_26056,N_25899);
or U27360 (N_27360,N_26662,N_25857);
nand U27361 (N_27361,N_25535,N_26480);
xnor U27362 (N_27362,N_25980,N_26135);
or U27363 (N_27363,N_26453,N_26857);
or U27364 (N_27364,N_25578,N_26042);
nand U27365 (N_27365,N_26319,N_26025);
xnor U27366 (N_27366,N_26026,N_25637);
and U27367 (N_27367,N_26815,N_26400);
xnor U27368 (N_27368,N_26178,N_25901);
nor U27369 (N_27369,N_25582,N_26385);
or U27370 (N_27370,N_25912,N_26196);
and U27371 (N_27371,N_25766,N_25949);
nor U27372 (N_27372,N_26617,N_26032);
nand U27373 (N_27373,N_25685,N_26635);
or U27374 (N_27374,N_25596,N_26604);
nor U27375 (N_27375,N_25736,N_25684);
xor U27376 (N_27376,N_26002,N_25500);
xor U27377 (N_27377,N_26783,N_26874);
xnor U27378 (N_27378,N_26382,N_26652);
nand U27379 (N_27379,N_25746,N_26172);
nor U27380 (N_27380,N_26589,N_26871);
nand U27381 (N_27381,N_26070,N_25810);
or U27382 (N_27382,N_26748,N_26117);
nor U27383 (N_27383,N_25914,N_26065);
and U27384 (N_27384,N_26239,N_25640);
nand U27385 (N_27385,N_26287,N_26281);
nand U27386 (N_27386,N_25704,N_26343);
and U27387 (N_27387,N_26285,N_26694);
xnor U27388 (N_27388,N_25557,N_26650);
nor U27389 (N_27389,N_26686,N_25588);
nor U27390 (N_27390,N_25604,N_25863);
or U27391 (N_27391,N_26639,N_26724);
or U27392 (N_27392,N_25885,N_26160);
and U27393 (N_27393,N_26926,N_26131);
or U27394 (N_27394,N_26767,N_26998);
xnor U27395 (N_27395,N_26938,N_26697);
and U27396 (N_27396,N_26426,N_26616);
and U27397 (N_27397,N_26268,N_25947);
nor U27398 (N_27398,N_26969,N_25877);
or U27399 (N_27399,N_26288,N_26265);
xor U27400 (N_27400,N_25819,N_26290);
and U27401 (N_27401,N_26574,N_26787);
and U27402 (N_27402,N_26234,N_26149);
or U27403 (N_27403,N_26580,N_26556);
and U27404 (N_27404,N_26688,N_26878);
xor U27405 (N_27405,N_25823,N_26904);
or U27406 (N_27406,N_26120,N_26671);
and U27407 (N_27407,N_26822,N_26793);
or U27408 (N_27408,N_25923,N_26434);
xnor U27409 (N_27409,N_26016,N_26250);
xnor U27410 (N_27410,N_26378,N_26602);
or U27411 (N_27411,N_25786,N_26487);
or U27412 (N_27412,N_25959,N_26672);
nand U27413 (N_27413,N_26486,N_25598);
nor U27414 (N_27414,N_26346,N_26765);
nor U27415 (N_27415,N_25544,N_25682);
and U27416 (N_27416,N_26407,N_26266);
or U27417 (N_27417,N_26460,N_26685);
nor U27418 (N_27418,N_26493,N_25587);
nand U27419 (N_27419,N_25918,N_26987);
or U27420 (N_27420,N_26679,N_26220);
or U27421 (N_27421,N_26715,N_26244);
or U27422 (N_27422,N_25676,N_26985);
and U27423 (N_27423,N_26263,N_26123);
xnor U27424 (N_27424,N_26349,N_26741);
and U27425 (N_27425,N_26376,N_26089);
or U27426 (N_27426,N_26861,N_26559);
and U27427 (N_27427,N_25813,N_26485);
nor U27428 (N_27428,N_26013,N_26843);
or U27429 (N_27429,N_26488,N_26829);
nand U27430 (N_27430,N_26723,N_26692);
xnor U27431 (N_27431,N_25828,N_25992);
nor U27432 (N_27432,N_26736,N_25620);
and U27433 (N_27433,N_26812,N_26693);
and U27434 (N_27434,N_26121,N_26656);
nand U27435 (N_27435,N_26551,N_25825);
and U27436 (N_27436,N_26294,N_26226);
nor U27437 (N_27437,N_26093,N_25611);
nor U27438 (N_27438,N_26891,N_25958);
and U27439 (N_27439,N_26977,N_26968);
nor U27440 (N_27440,N_25955,N_26068);
nand U27441 (N_27441,N_25505,N_25834);
or U27442 (N_27442,N_25726,N_26208);
xor U27443 (N_27443,N_26494,N_25653);
or U27444 (N_27444,N_26392,N_25926);
nand U27445 (N_27445,N_26454,N_26430);
or U27446 (N_27446,N_26803,N_26595);
and U27447 (N_27447,N_25717,N_26786);
or U27448 (N_27448,N_25904,N_25940);
and U27449 (N_27449,N_25515,N_26842);
or U27450 (N_27450,N_25617,N_25895);
nand U27451 (N_27451,N_25846,N_26432);
xnor U27452 (N_27452,N_25929,N_25753);
or U27453 (N_27453,N_26257,N_26707);
xnor U27454 (N_27454,N_25986,N_25502);
or U27455 (N_27455,N_25602,N_25672);
nand U27456 (N_27456,N_25983,N_26440);
nor U27457 (N_27457,N_25974,N_25941);
nand U27458 (N_27458,N_26071,N_26118);
and U27459 (N_27459,N_25658,N_26146);
or U27460 (N_27460,N_25874,N_26295);
xor U27461 (N_27461,N_26517,N_26720);
xnor U27462 (N_27462,N_26823,N_26933);
nor U27463 (N_27463,N_26565,N_26539);
and U27464 (N_27464,N_26875,N_26190);
nor U27465 (N_27465,N_25530,N_25550);
and U27466 (N_27466,N_26964,N_26116);
nand U27467 (N_27467,N_26848,N_26503);
and U27468 (N_27468,N_26489,N_25549);
nor U27469 (N_27469,N_25600,N_26080);
nor U27470 (N_27470,N_26740,N_25575);
and U27471 (N_27471,N_25506,N_25936);
nand U27472 (N_27472,N_26211,N_26154);
nand U27473 (N_27473,N_26384,N_26867);
nand U27474 (N_27474,N_25645,N_26104);
or U27475 (N_27475,N_26804,N_25851);
and U27476 (N_27476,N_26691,N_25679);
or U27477 (N_27477,N_26921,N_25508);
nor U27478 (N_27478,N_26568,N_26273);
nor U27479 (N_27479,N_26896,N_25984);
nand U27480 (N_27480,N_25599,N_25873);
and U27481 (N_27481,N_26944,N_26545);
or U27482 (N_27482,N_26431,N_26522);
nand U27483 (N_27483,N_26373,N_26581);
nand U27484 (N_27484,N_26847,N_26212);
and U27485 (N_27485,N_26532,N_26182);
nand U27486 (N_27486,N_25853,N_25740);
xnor U27487 (N_27487,N_26999,N_25681);
or U27488 (N_27488,N_26227,N_26937);
nand U27489 (N_27489,N_25892,N_26743);
nand U27490 (N_27490,N_26587,N_26296);
nand U27491 (N_27491,N_26138,N_26191);
nand U27492 (N_27492,N_25561,N_26555);
or U27493 (N_27493,N_25635,N_26327);
or U27494 (N_27494,N_26859,N_25624);
nor U27495 (N_27495,N_25950,N_26599);
nand U27496 (N_27496,N_26448,N_25841);
and U27497 (N_27497,N_25739,N_26576);
xnor U27498 (N_27498,N_25701,N_25985);
and U27499 (N_27499,N_26769,N_26405);
xor U27500 (N_27500,N_26915,N_25988);
nand U27501 (N_27501,N_26462,N_26592);
nor U27502 (N_27502,N_25589,N_25925);
nand U27503 (N_27503,N_26079,N_26630);
nor U27504 (N_27504,N_25848,N_26970);
nor U27505 (N_27505,N_26033,N_26739);
or U27506 (N_27506,N_26961,N_26643);
xnor U27507 (N_27507,N_26276,N_25757);
and U27508 (N_27508,N_26341,N_26704);
or U27509 (N_27509,N_25878,N_25591);
xnor U27510 (N_27510,N_26930,N_25689);
or U27511 (N_27511,N_26231,N_25655);
nand U27512 (N_27512,N_26923,N_26039);
and U27513 (N_27513,N_26660,N_26260);
nor U27514 (N_27514,N_26084,N_26340);
xor U27515 (N_27515,N_26952,N_26640);
nand U27516 (N_27516,N_25928,N_26927);
nor U27517 (N_27517,N_26187,N_25764);
nand U27518 (N_27518,N_25897,N_26192);
nor U27519 (N_27519,N_26564,N_26876);
nand U27520 (N_27520,N_25534,N_26496);
nor U27521 (N_27521,N_26950,N_26673);
or U27522 (N_27522,N_26566,N_26619);
nand U27523 (N_27523,N_26041,N_26846);
or U27524 (N_27524,N_26870,N_26860);
nand U27525 (N_27525,N_26169,N_25795);
or U27526 (N_27526,N_26274,N_26133);
nand U27527 (N_27527,N_25576,N_26956);
xnor U27528 (N_27528,N_26535,N_25748);
nand U27529 (N_27529,N_26943,N_26210);
or U27530 (N_27530,N_26534,N_26593);
or U27531 (N_27531,N_26900,N_26021);
or U27532 (N_27532,N_25829,N_26819);
nand U27533 (N_27533,N_26320,N_25887);
nor U27534 (N_27534,N_26209,N_26813);
nand U27535 (N_27535,N_25531,N_26907);
or U27536 (N_27536,N_25660,N_26536);
nor U27537 (N_27537,N_26136,N_26418);
nor U27538 (N_27538,N_25632,N_25712);
and U27539 (N_27539,N_25518,N_25765);
or U27540 (N_27540,N_25991,N_26929);
nand U27541 (N_27541,N_26655,N_26463);
xnor U27542 (N_27542,N_26709,N_26490);
nand U27543 (N_27543,N_26469,N_26411);
and U27544 (N_27544,N_26986,N_26917);
nor U27545 (N_27545,N_25972,N_26058);
and U27546 (N_27546,N_26925,N_25756);
nand U27547 (N_27547,N_26339,N_26951);
or U27548 (N_27548,N_26520,N_26844);
xnor U27549 (N_27549,N_26837,N_25902);
nand U27550 (N_27550,N_25778,N_25584);
nand U27551 (N_27551,N_26155,N_26905);
nand U27552 (N_27552,N_26868,N_25900);
nand U27553 (N_27553,N_26046,N_26601);
and U27554 (N_27554,N_25993,N_26608);
or U27555 (N_27555,N_25680,N_25816);
nor U27556 (N_27556,N_25866,N_26947);
or U27557 (N_27557,N_26271,N_26396);
and U27558 (N_27558,N_26909,N_25890);
or U27559 (N_27559,N_25820,N_25580);
nand U27560 (N_27560,N_26447,N_26893);
or U27561 (N_27561,N_26003,N_26115);
nand U27562 (N_27562,N_25800,N_26695);
nor U27563 (N_27563,N_25741,N_26497);
or U27564 (N_27564,N_26075,N_25965);
xor U27565 (N_27565,N_26854,N_25542);
xor U27566 (N_27566,N_26805,N_26610);
or U27567 (N_27567,N_26491,N_26329);
nand U27568 (N_27568,N_26624,N_26466);
or U27569 (N_27569,N_25727,N_26113);
nor U27570 (N_27570,N_26164,N_26162);
or U27571 (N_27571,N_26081,N_25787);
or U27572 (N_27572,N_26654,N_26988);
nor U27573 (N_27573,N_26175,N_25922);
xnor U27574 (N_27574,N_26326,N_25773);
nor U27575 (N_27575,N_25605,N_25916);
xor U27576 (N_27576,N_26143,N_25529);
nor U27577 (N_27577,N_25621,N_25708);
and U27578 (N_27578,N_26189,N_26477);
nand U27579 (N_27579,N_26530,N_26388);
nand U27580 (N_27580,N_26394,N_25798);
nand U27581 (N_27581,N_26456,N_25663);
and U27582 (N_27582,N_26836,N_25710);
nand U27583 (N_27583,N_26406,N_26659);
xnor U27584 (N_27584,N_26646,N_26500);
nand U27585 (N_27585,N_25989,N_26641);
or U27586 (N_27586,N_25612,N_25577);
nor U27587 (N_27587,N_25932,N_26678);
xor U27588 (N_27588,N_25623,N_25567);
nor U27589 (N_27589,N_26286,N_25709);
xnor U27590 (N_27590,N_26167,N_25843);
nor U27591 (N_27591,N_26957,N_26050);
nand U27592 (N_27592,N_25933,N_25978);
or U27593 (N_27593,N_25644,N_25607);
xnor U27594 (N_27594,N_26642,N_26059);
and U27595 (N_27595,N_25745,N_26474);
nand U27596 (N_27596,N_26614,N_26148);
nor U27597 (N_27597,N_26348,N_26470);
nor U27598 (N_27598,N_26658,N_26410);
nand U27599 (N_27599,N_26482,N_26727);
and U27600 (N_27600,N_25755,N_26377);
nand U27601 (N_27601,N_26982,N_25719);
or U27602 (N_27602,N_26479,N_26683);
or U27603 (N_27603,N_26020,N_26464);
or U27604 (N_27604,N_26001,N_26259);
nand U27605 (N_27605,N_26473,N_26240);
and U27606 (N_27606,N_26098,N_25855);
nor U27607 (N_27607,N_26974,N_26057);
or U27608 (N_27608,N_26960,N_26165);
xor U27609 (N_27609,N_26661,N_25896);
xor U27610 (N_27610,N_25854,N_26756);
and U27611 (N_27611,N_26855,N_25894);
nor U27612 (N_27612,N_25642,N_25824);
nand U27613 (N_27613,N_26179,N_25876);
and U27614 (N_27614,N_26124,N_26807);
or U27615 (N_27615,N_26973,N_25780);
xor U27616 (N_27616,N_26797,N_25700);
and U27617 (N_27617,N_26353,N_26841);
nor U27618 (N_27618,N_26087,N_25540);
nand U27619 (N_27619,N_25871,N_25987);
or U27620 (N_27620,N_26850,N_26993);
nor U27621 (N_27621,N_26994,N_26442);
nor U27622 (N_27622,N_26540,N_26899);
or U27623 (N_27623,N_25626,N_25814);
nand U27624 (N_27624,N_25809,N_25997);
xor U27625 (N_27625,N_26088,N_25789);
xor U27626 (N_27626,N_26443,N_26127);
and U27627 (N_27627,N_25677,N_26885);
nor U27628 (N_27628,N_25883,N_26193);
and U27629 (N_27629,N_25619,N_26292);
nor U27630 (N_27630,N_25715,N_26449);
nor U27631 (N_27631,N_25836,N_26600);
nor U27632 (N_27632,N_25546,N_25945);
or U27633 (N_27633,N_26542,N_26077);
and U27634 (N_27634,N_25659,N_26648);
or U27635 (N_27635,N_25821,N_26798);
xnor U27636 (N_27636,N_26959,N_26291);
nor U27637 (N_27637,N_26144,N_25513);
or U27638 (N_27638,N_25831,N_26404);
and U27639 (N_27639,N_26218,N_26895);
nand U27640 (N_27640,N_26433,N_25977);
or U27641 (N_27641,N_26880,N_26696);
xor U27642 (N_27642,N_25884,N_26249);
xnor U27643 (N_27643,N_26657,N_26049);
nand U27644 (N_27644,N_25674,N_25563);
or U27645 (N_27645,N_26521,N_26990);
xor U27646 (N_27646,N_26680,N_26401);
nand U27647 (N_27647,N_26438,N_25541);
and U27648 (N_27648,N_25688,N_26423);
xor U27649 (N_27649,N_26311,N_26772);
nand U27650 (N_27650,N_26631,N_26217);
nor U27651 (N_27651,N_26022,N_25921);
nor U27652 (N_27652,N_26495,N_25893);
or U27653 (N_27653,N_26007,N_26168);
nor U27654 (N_27654,N_26370,N_25510);
nand U27655 (N_27655,N_26667,N_25830);
and U27656 (N_27656,N_26038,N_26802);
nand U27657 (N_27657,N_26849,N_26499);
nor U27658 (N_27658,N_26770,N_25924);
nand U27659 (N_27659,N_26776,N_25532);
nor U27660 (N_27660,N_26634,N_26315);
or U27661 (N_27661,N_25665,N_25792);
nor U27662 (N_27662,N_26922,N_26216);
xor U27663 (N_27663,N_26106,N_26625);
and U27664 (N_27664,N_26125,N_26351);
or U27665 (N_27665,N_26948,N_25744);
nand U27666 (N_27666,N_26932,N_26452);
or U27667 (N_27667,N_25608,N_26774);
and U27668 (N_27668,N_25794,N_25799);
nand U27669 (N_27669,N_26762,N_26331);
and U27670 (N_27670,N_26920,N_26393);
nand U27671 (N_27671,N_26618,N_26584);
nand U27672 (N_27672,N_26928,N_25601);
nand U27673 (N_27673,N_26995,N_26814);
xor U27674 (N_27674,N_26283,N_25920);
nand U27675 (N_27675,N_26991,N_26054);
nor U27676 (N_27676,N_25835,N_26241);
xnor U27677 (N_27677,N_26383,N_26689);
or U27678 (N_27678,N_26742,N_26272);
or U27679 (N_27679,N_25511,N_26773);
nand U27680 (N_27680,N_25548,N_25747);
nor U27681 (N_27681,N_26598,N_26122);
nor U27682 (N_27682,N_25568,N_25516);
nor U27683 (N_27683,N_26439,N_26586);
and U27684 (N_27684,N_26924,N_25555);
xnor U27685 (N_27685,N_26910,N_26318);
nand U27686 (N_27686,N_26200,N_26481);
nand U27687 (N_27687,N_26140,N_26063);
nand U27688 (N_27688,N_26820,N_26246);
and U27689 (N_27689,N_26706,N_26424);
nand U27690 (N_27690,N_25503,N_26357);
or U27691 (N_27691,N_26102,N_26518);
and U27692 (N_27692,N_25558,N_26698);
nand U27693 (N_27693,N_25806,N_25521);
xnor U27694 (N_27694,N_26332,N_26779);
and U27695 (N_27695,N_26501,N_26865);
or U27696 (N_27696,N_26361,N_26203);
xor U27697 (N_27697,N_26939,N_25750);
nor U27698 (N_27698,N_26992,N_26130);
nand U27699 (N_27699,N_26328,N_26955);
nand U27700 (N_27700,N_25802,N_26362);
and U27701 (N_27701,N_25779,N_26214);
nor U27702 (N_27702,N_25547,N_26719);
xor U27703 (N_27703,N_26527,N_26062);
nand U27704 (N_27704,N_26768,N_25953);
nor U27705 (N_27705,N_26840,N_26111);
nand U27706 (N_27706,N_26108,N_26299);
or U27707 (N_27707,N_26627,N_26451);
and U27708 (N_27708,N_26158,N_26066);
xnor U27709 (N_27709,N_25754,N_25731);
xnor U27710 (N_27710,N_26705,N_26980);
nand U27711 (N_27711,N_26872,N_26321);
and U27712 (N_27712,N_26215,N_25777);
xor U27713 (N_27713,N_25536,N_26882);
and U27714 (N_27714,N_26834,N_26008);
nor U27715 (N_27715,N_25507,N_26194);
and U27716 (N_27716,N_25673,N_25966);
nand U27717 (N_27717,N_25783,N_26890);
nand U27718 (N_27718,N_26024,N_25840);
nor U27719 (N_27719,N_25652,N_26128);
xor U27720 (N_27720,N_25627,N_26375);
xnor U27721 (N_27721,N_26094,N_26788);
xnor U27722 (N_27722,N_26682,N_25703);
nand U27723 (N_27723,N_26428,N_26759);
xnor U27724 (N_27724,N_26751,N_26912);
nand U27725 (N_27725,N_26472,N_26484);
xor U27726 (N_27726,N_26538,N_26935);
or U27727 (N_27727,N_25735,N_26983);
or U27728 (N_27728,N_26498,N_25858);
nand U27729 (N_27729,N_25817,N_26201);
or U27730 (N_27730,N_26012,N_26225);
nor U27731 (N_27731,N_26523,N_26029);
and U27732 (N_27732,N_26387,N_26515);
nor U27733 (N_27733,N_26777,N_26519);
xor U27734 (N_27734,N_25696,N_26358);
nand U27735 (N_27735,N_25574,N_26645);
nand U27736 (N_27736,N_25913,N_26437);
or U27737 (N_27737,N_26101,N_25614);
nand U27738 (N_27738,N_25631,N_26289);
and U27739 (N_27739,N_26455,N_26333);
or U27740 (N_27740,N_25504,N_25593);
xnor U27741 (N_27741,N_25678,N_26516);
nand U27742 (N_27742,N_25520,N_26666);
and U27743 (N_27743,N_26919,N_25771);
nor U27744 (N_27744,N_25957,N_25528);
nand U27745 (N_27745,N_26398,N_25785);
xnor U27746 (N_27746,N_26781,N_26345);
or U27747 (N_27747,N_26171,N_25772);
nor U27748 (N_27748,N_26310,N_25942);
or U27749 (N_27749,N_26152,N_26095);
xor U27750 (N_27750,N_25667,N_25630);
and U27751 (N_27751,N_25609,N_26336);
or U27752 (N_27752,N_26451,N_26267);
nor U27753 (N_27753,N_26538,N_26302);
nor U27754 (N_27754,N_25878,N_26619);
or U27755 (N_27755,N_25827,N_25709);
or U27756 (N_27756,N_26797,N_26151);
xor U27757 (N_27757,N_26084,N_26549);
and U27758 (N_27758,N_25764,N_26993);
and U27759 (N_27759,N_26104,N_26432);
and U27760 (N_27760,N_26447,N_26988);
xor U27761 (N_27761,N_25995,N_26442);
nand U27762 (N_27762,N_26519,N_26124);
or U27763 (N_27763,N_26805,N_26067);
xor U27764 (N_27764,N_26280,N_26964);
and U27765 (N_27765,N_25654,N_25733);
nor U27766 (N_27766,N_26723,N_26629);
xnor U27767 (N_27767,N_26674,N_25618);
and U27768 (N_27768,N_26670,N_26710);
or U27769 (N_27769,N_25583,N_26190);
nor U27770 (N_27770,N_26054,N_25904);
nor U27771 (N_27771,N_26882,N_26722);
and U27772 (N_27772,N_25548,N_25799);
and U27773 (N_27773,N_26176,N_25635);
xor U27774 (N_27774,N_25620,N_26102);
xor U27775 (N_27775,N_25918,N_25864);
nor U27776 (N_27776,N_25734,N_26659);
or U27777 (N_27777,N_25598,N_26322);
xnor U27778 (N_27778,N_26435,N_25660);
nor U27779 (N_27779,N_26718,N_26106);
or U27780 (N_27780,N_26581,N_26525);
nand U27781 (N_27781,N_26565,N_26793);
nand U27782 (N_27782,N_26378,N_25812);
nand U27783 (N_27783,N_26533,N_25835);
xor U27784 (N_27784,N_25715,N_26605);
and U27785 (N_27785,N_25777,N_26319);
nor U27786 (N_27786,N_26830,N_26335);
xor U27787 (N_27787,N_26586,N_25771);
and U27788 (N_27788,N_26733,N_26481);
nand U27789 (N_27789,N_26819,N_26727);
nand U27790 (N_27790,N_26414,N_25861);
or U27791 (N_27791,N_26017,N_25618);
nand U27792 (N_27792,N_25860,N_25853);
xnor U27793 (N_27793,N_26958,N_26668);
nand U27794 (N_27794,N_25973,N_26871);
or U27795 (N_27795,N_26744,N_25635);
and U27796 (N_27796,N_25732,N_25776);
nor U27797 (N_27797,N_26703,N_25937);
xnor U27798 (N_27798,N_26154,N_26681);
xor U27799 (N_27799,N_26348,N_25527);
nor U27800 (N_27800,N_26492,N_25797);
nand U27801 (N_27801,N_26018,N_26261);
or U27802 (N_27802,N_26537,N_26572);
or U27803 (N_27803,N_26126,N_25630);
nand U27804 (N_27804,N_26264,N_26836);
or U27805 (N_27805,N_25827,N_25823);
nor U27806 (N_27806,N_26693,N_26091);
nand U27807 (N_27807,N_26186,N_26187);
xnor U27808 (N_27808,N_26834,N_25953);
or U27809 (N_27809,N_25721,N_26842);
xnor U27810 (N_27810,N_26748,N_25620);
nand U27811 (N_27811,N_26654,N_26359);
and U27812 (N_27812,N_26413,N_26792);
and U27813 (N_27813,N_26066,N_26343);
xnor U27814 (N_27814,N_25563,N_25546);
or U27815 (N_27815,N_26125,N_26059);
xnor U27816 (N_27816,N_26815,N_25799);
and U27817 (N_27817,N_26685,N_26378);
or U27818 (N_27818,N_26220,N_26062);
nand U27819 (N_27819,N_26585,N_26433);
nand U27820 (N_27820,N_26097,N_26024);
nor U27821 (N_27821,N_25817,N_25506);
or U27822 (N_27822,N_26359,N_26818);
or U27823 (N_27823,N_26505,N_25895);
xor U27824 (N_27824,N_26482,N_26532);
or U27825 (N_27825,N_26292,N_26186);
and U27826 (N_27826,N_26184,N_25751);
nand U27827 (N_27827,N_26153,N_26586);
nor U27828 (N_27828,N_26475,N_26121);
or U27829 (N_27829,N_26461,N_25547);
nand U27830 (N_27830,N_25578,N_26696);
nand U27831 (N_27831,N_25934,N_26545);
xor U27832 (N_27832,N_26808,N_25664);
and U27833 (N_27833,N_25716,N_26678);
or U27834 (N_27834,N_25610,N_26804);
and U27835 (N_27835,N_26130,N_26342);
and U27836 (N_27836,N_26586,N_26346);
nor U27837 (N_27837,N_26740,N_26688);
nor U27838 (N_27838,N_25996,N_25899);
xor U27839 (N_27839,N_25640,N_25536);
and U27840 (N_27840,N_25723,N_25610);
nor U27841 (N_27841,N_26409,N_26251);
and U27842 (N_27842,N_26109,N_26912);
nand U27843 (N_27843,N_26454,N_25964);
nand U27844 (N_27844,N_26849,N_25733);
xor U27845 (N_27845,N_26361,N_26175);
or U27846 (N_27846,N_26640,N_26242);
or U27847 (N_27847,N_26877,N_26157);
nor U27848 (N_27848,N_26076,N_25564);
xor U27849 (N_27849,N_25609,N_26412);
and U27850 (N_27850,N_26086,N_25557);
xnor U27851 (N_27851,N_26538,N_26032);
nand U27852 (N_27852,N_25751,N_26265);
nand U27853 (N_27853,N_25567,N_26708);
xnor U27854 (N_27854,N_26007,N_26108);
or U27855 (N_27855,N_25552,N_26660);
xnor U27856 (N_27856,N_26314,N_26173);
xor U27857 (N_27857,N_25539,N_26559);
and U27858 (N_27858,N_26994,N_25809);
xnor U27859 (N_27859,N_25556,N_26151);
xnor U27860 (N_27860,N_26714,N_26318);
or U27861 (N_27861,N_25912,N_25785);
and U27862 (N_27862,N_26151,N_26149);
nor U27863 (N_27863,N_26972,N_26483);
and U27864 (N_27864,N_26944,N_25997);
or U27865 (N_27865,N_26231,N_26468);
and U27866 (N_27866,N_26664,N_26050);
and U27867 (N_27867,N_26783,N_25736);
nand U27868 (N_27868,N_26273,N_26858);
xor U27869 (N_27869,N_26639,N_25869);
and U27870 (N_27870,N_26130,N_26244);
xor U27871 (N_27871,N_26803,N_26644);
nor U27872 (N_27872,N_26421,N_26520);
xnor U27873 (N_27873,N_25842,N_26074);
and U27874 (N_27874,N_26489,N_26902);
xor U27875 (N_27875,N_25616,N_26486);
and U27876 (N_27876,N_26460,N_26428);
or U27877 (N_27877,N_26632,N_25737);
xnor U27878 (N_27878,N_26086,N_26863);
nor U27879 (N_27879,N_25564,N_25745);
nor U27880 (N_27880,N_25787,N_26648);
nor U27881 (N_27881,N_26357,N_26446);
or U27882 (N_27882,N_25797,N_25960);
nor U27883 (N_27883,N_26487,N_26712);
or U27884 (N_27884,N_25850,N_26458);
nor U27885 (N_27885,N_26435,N_25727);
xnor U27886 (N_27886,N_26543,N_26138);
or U27887 (N_27887,N_26808,N_26802);
or U27888 (N_27888,N_25607,N_26634);
and U27889 (N_27889,N_26849,N_26255);
or U27890 (N_27890,N_25662,N_25992);
nor U27891 (N_27891,N_26987,N_26319);
or U27892 (N_27892,N_25736,N_26637);
and U27893 (N_27893,N_26340,N_26030);
nor U27894 (N_27894,N_26370,N_26323);
nand U27895 (N_27895,N_26875,N_26877);
and U27896 (N_27896,N_25628,N_25954);
and U27897 (N_27897,N_26176,N_26110);
or U27898 (N_27898,N_26269,N_25912);
or U27899 (N_27899,N_26777,N_26367);
nand U27900 (N_27900,N_26415,N_26544);
xor U27901 (N_27901,N_26099,N_25624);
nor U27902 (N_27902,N_25988,N_26721);
xnor U27903 (N_27903,N_26070,N_25948);
nand U27904 (N_27904,N_26010,N_25910);
nand U27905 (N_27905,N_26519,N_26622);
nand U27906 (N_27906,N_26418,N_26149);
and U27907 (N_27907,N_26854,N_26867);
or U27908 (N_27908,N_26238,N_26708);
xor U27909 (N_27909,N_25686,N_25627);
nor U27910 (N_27910,N_25977,N_26113);
or U27911 (N_27911,N_26303,N_25671);
nand U27912 (N_27912,N_25645,N_26718);
and U27913 (N_27913,N_26351,N_26302);
xor U27914 (N_27914,N_26640,N_25674);
or U27915 (N_27915,N_26118,N_26104);
nor U27916 (N_27916,N_25755,N_26304);
or U27917 (N_27917,N_26966,N_26183);
nand U27918 (N_27918,N_25708,N_26108);
or U27919 (N_27919,N_26424,N_26904);
nor U27920 (N_27920,N_26297,N_26030);
or U27921 (N_27921,N_26375,N_26603);
and U27922 (N_27922,N_26382,N_26717);
nor U27923 (N_27923,N_26620,N_25709);
nand U27924 (N_27924,N_25561,N_26330);
or U27925 (N_27925,N_25885,N_25950);
or U27926 (N_27926,N_26376,N_25937);
and U27927 (N_27927,N_26330,N_26328);
or U27928 (N_27928,N_25632,N_26203);
and U27929 (N_27929,N_25542,N_26355);
or U27930 (N_27930,N_26964,N_26787);
nor U27931 (N_27931,N_26818,N_26111);
and U27932 (N_27932,N_26940,N_26963);
or U27933 (N_27933,N_26507,N_26120);
and U27934 (N_27934,N_26209,N_26103);
and U27935 (N_27935,N_26066,N_26015);
nor U27936 (N_27936,N_26319,N_26814);
xnor U27937 (N_27937,N_25555,N_26368);
nand U27938 (N_27938,N_26290,N_26818);
and U27939 (N_27939,N_25582,N_26565);
or U27940 (N_27940,N_26655,N_25582);
nor U27941 (N_27941,N_26733,N_25961);
nor U27942 (N_27942,N_25581,N_26981);
nand U27943 (N_27943,N_26059,N_26131);
nand U27944 (N_27944,N_25630,N_25637);
xnor U27945 (N_27945,N_26399,N_26999);
nand U27946 (N_27946,N_26463,N_25727);
and U27947 (N_27947,N_25642,N_25854);
or U27948 (N_27948,N_26105,N_25999);
nand U27949 (N_27949,N_26130,N_26972);
nand U27950 (N_27950,N_26765,N_26784);
nand U27951 (N_27951,N_26512,N_26162);
nor U27952 (N_27952,N_26259,N_25537);
xnor U27953 (N_27953,N_25950,N_25831);
xor U27954 (N_27954,N_26862,N_26875);
xor U27955 (N_27955,N_26105,N_26312);
xnor U27956 (N_27956,N_26994,N_26949);
nor U27957 (N_27957,N_26570,N_26281);
or U27958 (N_27958,N_26910,N_26036);
or U27959 (N_27959,N_26504,N_25853);
xor U27960 (N_27960,N_26061,N_25551);
or U27961 (N_27961,N_26809,N_25608);
nand U27962 (N_27962,N_26234,N_25926);
nand U27963 (N_27963,N_25701,N_25572);
nor U27964 (N_27964,N_26827,N_26307);
xnor U27965 (N_27965,N_26622,N_25678);
nor U27966 (N_27966,N_25837,N_26629);
and U27967 (N_27967,N_25817,N_25819);
and U27968 (N_27968,N_26540,N_25730);
or U27969 (N_27969,N_26939,N_26223);
and U27970 (N_27970,N_25734,N_26647);
nor U27971 (N_27971,N_26641,N_26913);
nor U27972 (N_27972,N_26360,N_26151);
nor U27973 (N_27973,N_25559,N_26665);
nor U27974 (N_27974,N_26344,N_26100);
nand U27975 (N_27975,N_25668,N_25510);
and U27976 (N_27976,N_26408,N_26782);
nand U27977 (N_27977,N_26312,N_26774);
nor U27978 (N_27978,N_26711,N_26677);
xnor U27979 (N_27979,N_25735,N_26945);
nand U27980 (N_27980,N_26495,N_25898);
and U27981 (N_27981,N_26390,N_26691);
or U27982 (N_27982,N_26892,N_26225);
nand U27983 (N_27983,N_26813,N_25975);
xnor U27984 (N_27984,N_26492,N_26144);
nand U27985 (N_27985,N_25617,N_26590);
nor U27986 (N_27986,N_26157,N_26016);
nor U27987 (N_27987,N_26329,N_25802);
and U27988 (N_27988,N_26838,N_25973);
and U27989 (N_27989,N_25728,N_26255);
and U27990 (N_27990,N_25977,N_26791);
xor U27991 (N_27991,N_25612,N_26428);
nand U27992 (N_27992,N_26890,N_25620);
xor U27993 (N_27993,N_26599,N_26006);
nor U27994 (N_27994,N_26058,N_25625);
nand U27995 (N_27995,N_25544,N_26348);
nand U27996 (N_27996,N_26776,N_26904);
xor U27997 (N_27997,N_25796,N_26441);
xor U27998 (N_27998,N_26010,N_26816);
nand U27999 (N_27999,N_26635,N_26143);
and U28000 (N_28000,N_26080,N_25522);
nor U28001 (N_28001,N_26943,N_25524);
and U28002 (N_28002,N_26147,N_26684);
nand U28003 (N_28003,N_26499,N_26779);
xor U28004 (N_28004,N_26400,N_26257);
or U28005 (N_28005,N_26791,N_26829);
xor U28006 (N_28006,N_26266,N_26306);
or U28007 (N_28007,N_26327,N_26959);
and U28008 (N_28008,N_26310,N_26857);
xor U28009 (N_28009,N_26541,N_26738);
nand U28010 (N_28010,N_26071,N_25764);
nor U28011 (N_28011,N_26733,N_25867);
xor U28012 (N_28012,N_26096,N_26276);
and U28013 (N_28013,N_26227,N_25964);
xnor U28014 (N_28014,N_25884,N_26570);
and U28015 (N_28015,N_26772,N_26546);
and U28016 (N_28016,N_25932,N_26249);
or U28017 (N_28017,N_26220,N_26741);
xor U28018 (N_28018,N_26071,N_26690);
and U28019 (N_28019,N_25986,N_26729);
or U28020 (N_28020,N_26008,N_25972);
and U28021 (N_28021,N_25776,N_25930);
and U28022 (N_28022,N_26609,N_25903);
nand U28023 (N_28023,N_26372,N_25663);
and U28024 (N_28024,N_26331,N_25581);
or U28025 (N_28025,N_26486,N_25967);
and U28026 (N_28026,N_26073,N_25834);
nand U28027 (N_28027,N_26240,N_26504);
nand U28028 (N_28028,N_25716,N_25990);
nor U28029 (N_28029,N_26300,N_26187);
and U28030 (N_28030,N_25968,N_26261);
or U28031 (N_28031,N_25949,N_25546);
nor U28032 (N_28032,N_26634,N_25652);
nand U28033 (N_28033,N_25918,N_25750);
and U28034 (N_28034,N_26829,N_26345);
or U28035 (N_28035,N_26186,N_26836);
nand U28036 (N_28036,N_25874,N_25814);
xor U28037 (N_28037,N_26904,N_26046);
xnor U28038 (N_28038,N_26624,N_26610);
nand U28039 (N_28039,N_26918,N_25729);
xor U28040 (N_28040,N_26309,N_26886);
nor U28041 (N_28041,N_26754,N_26081);
xor U28042 (N_28042,N_26303,N_26649);
and U28043 (N_28043,N_25813,N_25881);
nand U28044 (N_28044,N_25615,N_26045);
and U28045 (N_28045,N_25727,N_26091);
xnor U28046 (N_28046,N_26605,N_26642);
and U28047 (N_28047,N_26326,N_26637);
and U28048 (N_28048,N_26354,N_25708);
and U28049 (N_28049,N_26048,N_25551);
and U28050 (N_28050,N_25790,N_26595);
nand U28051 (N_28051,N_26707,N_26411);
and U28052 (N_28052,N_25959,N_26390);
nand U28053 (N_28053,N_25582,N_26386);
or U28054 (N_28054,N_26545,N_25994);
or U28055 (N_28055,N_26890,N_26794);
nor U28056 (N_28056,N_25633,N_26133);
or U28057 (N_28057,N_25592,N_26040);
nand U28058 (N_28058,N_26303,N_26337);
nor U28059 (N_28059,N_26226,N_25647);
nand U28060 (N_28060,N_25688,N_25803);
and U28061 (N_28061,N_26200,N_26817);
nand U28062 (N_28062,N_26803,N_26670);
or U28063 (N_28063,N_26482,N_25761);
xor U28064 (N_28064,N_26912,N_25588);
xor U28065 (N_28065,N_26809,N_26690);
xor U28066 (N_28066,N_26333,N_26239);
xor U28067 (N_28067,N_26080,N_26968);
nand U28068 (N_28068,N_26049,N_26594);
nor U28069 (N_28069,N_26679,N_26379);
nand U28070 (N_28070,N_26534,N_26109);
nor U28071 (N_28071,N_26078,N_26907);
nand U28072 (N_28072,N_25804,N_26843);
and U28073 (N_28073,N_26365,N_26848);
xor U28074 (N_28074,N_26290,N_26554);
or U28075 (N_28075,N_26728,N_25752);
and U28076 (N_28076,N_25722,N_26486);
nand U28077 (N_28077,N_26591,N_26977);
and U28078 (N_28078,N_25658,N_26440);
or U28079 (N_28079,N_25721,N_26953);
nand U28080 (N_28080,N_26708,N_26337);
and U28081 (N_28081,N_25501,N_26883);
nand U28082 (N_28082,N_26762,N_26950);
and U28083 (N_28083,N_26554,N_26174);
and U28084 (N_28084,N_26886,N_26745);
and U28085 (N_28085,N_26048,N_26327);
xor U28086 (N_28086,N_25887,N_25942);
xor U28087 (N_28087,N_26632,N_26174);
or U28088 (N_28088,N_25624,N_26022);
xor U28089 (N_28089,N_25703,N_26665);
nand U28090 (N_28090,N_25637,N_26393);
or U28091 (N_28091,N_26213,N_26605);
or U28092 (N_28092,N_26030,N_26761);
nor U28093 (N_28093,N_25977,N_26411);
and U28094 (N_28094,N_26244,N_25830);
xnor U28095 (N_28095,N_26539,N_26984);
or U28096 (N_28096,N_26361,N_26652);
and U28097 (N_28097,N_26197,N_26495);
nand U28098 (N_28098,N_26462,N_25555);
nand U28099 (N_28099,N_26241,N_25744);
xor U28100 (N_28100,N_26419,N_26479);
nor U28101 (N_28101,N_26048,N_26018);
and U28102 (N_28102,N_26160,N_25934);
nor U28103 (N_28103,N_25973,N_25763);
nand U28104 (N_28104,N_26828,N_26625);
nor U28105 (N_28105,N_26730,N_26152);
nor U28106 (N_28106,N_25591,N_25934);
or U28107 (N_28107,N_25511,N_26190);
nor U28108 (N_28108,N_26151,N_26537);
or U28109 (N_28109,N_26712,N_25834);
and U28110 (N_28110,N_26755,N_26336);
nor U28111 (N_28111,N_26227,N_26576);
and U28112 (N_28112,N_26731,N_26549);
nand U28113 (N_28113,N_26607,N_26800);
xnor U28114 (N_28114,N_25577,N_26170);
xor U28115 (N_28115,N_26665,N_26699);
nor U28116 (N_28116,N_26269,N_25838);
nand U28117 (N_28117,N_26011,N_26335);
and U28118 (N_28118,N_26159,N_26213);
nor U28119 (N_28119,N_25913,N_26334);
nand U28120 (N_28120,N_25874,N_26634);
and U28121 (N_28121,N_26444,N_26360);
or U28122 (N_28122,N_25808,N_25506);
and U28123 (N_28123,N_25533,N_26372);
xor U28124 (N_28124,N_26997,N_26642);
and U28125 (N_28125,N_25616,N_25833);
and U28126 (N_28126,N_26929,N_25640);
nand U28127 (N_28127,N_26341,N_25535);
or U28128 (N_28128,N_26223,N_26698);
and U28129 (N_28129,N_25794,N_26320);
xnor U28130 (N_28130,N_25819,N_26282);
nand U28131 (N_28131,N_26724,N_26474);
or U28132 (N_28132,N_26539,N_25699);
xor U28133 (N_28133,N_25546,N_25737);
or U28134 (N_28134,N_26950,N_26515);
or U28135 (N_28135,N_26835,N_26517);
nor U28136 (N_28136,N_26783,N_26175);
and U28137 (N_28137,N_26676,N_26547);
nand U28138 (N_28138,N_26044,N_26957);
and U28139 (N_28139,N_26224,N_26358);
nand U28140 (N_28140,N_26671,N_25875);
and U28141 (N_28141,N_26878,N_26669);
and U28142 (N_28142,N_26725,N_26434);
nand U28143 (N_28143,N_26407,N_25521);
nand U28144 (N_28144,N_25910,N_26887);
and U28145 (N_28145,N_26605,N_25644);
and U28146 (N_28146,N_25639,N_26097);
nor U28147 (N_28147,N_26626,N_26910);
nand U28148 (N_28148,N_26561,N_26601);
nand U28149 (N_28149,N_25748,N_26216);
xor U28150 (N_28150,N_26317,N_26291);
and U28151 (N_28151,N_25582,N_25603);
nor U28152 (N_28152,N_25658,N_26659);
and U28153 (N_28153,N_25845,N_25824);
nand U28154 (N_28154,N_26190,N_26499);
and U28155 (N_28155,N_25676,N_26943);
or U28156 (N_28156,N_26973,N_25691);
nor U28157 (N_28157,N_26303,N_25892);
or U28158 (N_28158,N_25831,N_25990);
nor U28159 (N_28159,N_26202,N_26022);
or U28160 (N_28160,N_26364,N_26822);
nor U28161 (N_28161,N_26290,N_25776);
xor U28162 (N_28162,N_25679,N_25969);
and U28163 (N_28163,N_26499,N_26135);
and U28164 (N_28164,N_25836,N_26208);
or U28165 (N_28165,N_25970,N_25749);
nor U28166 (N_28166,N_25573,N_26773);
or U28167 (N_28167,N_25770,N_25854);
nor U28168 (N_28168,N_26770,N_26524);
nor U28169 (N_28169,N_25624,N_25625);
nand U28170 (N_28170,N_26149,N_25717);
nand U28171 (N_28171,N_26088,N_26348);
and U28172 (N_28172,N_26483,N_26702);
nor U28173 (N_28173,N_26935,N_26440);
and U28174 (N_28174,N_26183,N_26761);
and U28175 (N_28175,N_25513,N_26081);
nor U28176 (N_28176,N_25516,N_26208);
or U28177 (N_28177,N_26092,N_26993);
nor U28178 (N_28178,N_26389,N_26592);
and U28179 (N_28179,N_25970,N_26275);
xnor U28180 (N_28180,N_26295,N_26283);
xnor U28181 (N_28181,N_25646,N_25768);
and U28182 (N_28182,N_26022,N_25660);
nor U28183 (N_28183,N_26875,N_26336);
and U28184 (N_28184,N_26955,N_26216);
xor U28185 (N_28185,N_26334,N_25925);
nor U28186 (N_28186,N_25937,N_26467);
xor U28187 (N_28187,N_26901,N_26701);
nand U28188 (N_28188,N_26369,N_25611);
and U28189 (N_28189,N_26777,N_26479);
nand U28190 (N_28190,N_26680,N_26942);
and U28191 (N_28191,N_26251,N_25953);
or U28192 (N_28192,N_26483,N_26147);
nand U28193 (N_28193,N_26691,N_26864);
and U28194 (N_28194,N_26405,N_26995);
xnor U28195 (N_28195,N_26574,N_26446);
nand U28196 (N_28196,N_26028,N_25704);
xnor U28197 (N_28197,N_26849,N_26794);
xnor U28198 (N_28198,N_26605,N_25587);
or U28199 (N_28199,N_25698,N_26378);
nand U28200 (N_28200,N_26756,N_25617);
xor U28201 (N_28201,N_26772,N_26276);
and U28202 (N_28202,N_26140,N_25782);
nor U28203 (N_28203,N_25868,N_25974);
xor U28204 (N_28204,N_26426,N_25562);
or U28205 (N_28205,N_26553,N_25818);
and U28206 (N_28206,N_26558,N_26044);
nand U28207 (N_28207,N_26049,N_25834);
or U28208 (N_28208,N_26311,N_25884);
nor U28209 (N_28209,N_25787,N_25962);
nand U28210 (N_28210,N_26112,N_25801);
nand U28211 (N_28211,N_26921,N_26998);
xnor U28212 (N_28212,N_25705,N_26053);
xnor U28213 (N_28213,N_26028,N_25510);
and U28214 (N_28214,N_26939,N_26612);
or U28215 (N_28215,N_25956,N_26057);
nor U28216 (N_28216,N_25551,N_25997);
and U28217 (N_28217,N_26962,N_26463);
and U28218 (N_28218,N_26295,N_25564);
and U28219 (N_28219,N_25749,N_26497);
or U28220 (N_28220,N_25809,N_25799);
xnor U28221 (N_28221,N_25870,N_26508);
nand U28222 (N_28222,N_26085,N_26793);
and U28223 (N_28223,N_26927,N_25527);
and U28224 (N_28224,N_26017,N_25584);
or U28225 (N_28225,N_26762,N_26425);
nor U28226 (N_28226,N_26876,N_26412);
and U28227 (N_28227,N_26784,N_26858);
nor U28228 (N_28228,N_26803,N_26295);
nor U28229 (N_28229,N_26485,N_25677);
xor U28230 (N_28230,N_25534,N_26674);
nor U28231 (N_28231,N_25501,N_25836);
nand U28232 (N_28232,N_26469,N_25991);
or U28233 (N_28233,N_26595,N_26090);
or U28234 (N_28234,N_25503,N_26053);
and U28235 (N_28235,N_26576,N_26673);
or U28236 (N_28236,N_26250,N_26252);
or U28237 (N_28237,N_26073,N_26795);
and U28238 (N_28238,N_25573,N_25704);
and U28239 (N_28239,N_25706,N_26395);
or U28240 (N_28240,N_26691,N_26106);
and U28241 (N_28241,N_25653,N_26969);
nand U28242 (N_28242,N_26024,N_26908);
nor U28243 (N_28243,N_26591,N_26782);
nor U28244 (N_28244,N_26839,N_26821);
and U28245 (N_28245,N_25812,N_26338);
xor U28246 (N_28246,N_26631,N_26962);
or U28247 (N_28247,N_25862,N_26503);
nand U28248 (N_28248,N_25613,N_25706);
and U28249 (N_28249,N_26576,N_26120);
and U28250 (N_28250,N_25587,N_26792);
or U28251 (N_28251,N_25711,N_26868);
nor U28252 (N_28252,N_26427,N_26535);
or U28253 (N_28253,N_25624,N_25857);
nand U28254 (N_28254,N_26850,N_26776);
and U28255 (N_28255,N_26166,N_25601);
xor U28256 (N_28256,N_26476,N_25882);
and U28257 (N_28257,N_26705,N_25588);
nand U28258 (N_28258,N_26195,N_26191);
and U28259 (N_28259,N_25646,N_25819);
xor U28260 (N_28260,N_26849,N_26336);
nor U28261 (N_28261,N_26056,N_26832);
xor U28262 (N_28262,N_26462,N_26144);
nand U28263 (N_28263,N_25918,N_26050);
xnor U28264 (N_28264,N_26815,N_26291);
nor U28265 (N_28265,N_25637,N_25720);
xnor U28266 (N_28266,N_26444,N_26705);
or U28267 (N_28267,N_26435,N_26396);
nor U28268 (N_28268,N_26008,N_26259);
nor U28269 (N_28269,N_25516,N_25711);
or U28270 (N_28270,N_26921,N_26777);
and U28271 (N_28271,N_26002,N_26451);
nand U28272 (N_28272,N_26907,N_26412);
or U28273 (N_28273,N_26506,N_26127);
or U28274 (N_28274,N_26544,N_26668);
and U28275 (N_28275,N_26517,N_26230);
nor U28276 (N_28276,N_25633,N_26963);
nor U28277 (N_28277,N_26581,N_25788);
and U28278 (N_28278,N_25620,N_26901);
or U28279 (N_28279,N_26140,N_25951);
or U28280 (N_28280,N_26392,N_26878);
nor U28281 (N_28281,N_26252,N_26664);
xnor U28282 (N_28282,N_26533,N_26598);
or U28283 (N_28283,N_25831,N_26767);
nor U28284 (N_28284,N_25559,N_26040);
and U28285 (N_28285,N_25700,N_26823);
xnor U28286 (N_28286,N_26057,N_26110);
nand U28287 (N_28287,N_26031,N_25879);
nand U28288 (N_28288,N_26570,N_26756);
xnor U28289 (N_28289,N_26140,N_26620);
xor U28290 (N_28290,N_25660,N_26089);
xnor U28291 (N_28291,N_25713,N_25705);
xor U28292 (N_28292,N_26724,N_26027);
nor U28293 (N_28293,N_26213,N_25525);
nor U28294 (N_28294,N_26353,N_26057);
nor U28295 (N_28295,N_26801,N_25950);
or U28296 (N_28296,N_25670,N_25880);
and U28297 (N_28297,N_26146,N_26711);
or U28298 (N_28298,N_26598,N_26774);
nand U28299 (N_28299,N_26949,N_26632);
nand U28300 (N_28300,N_25950,N_26829);
or U28301 (N_28301,N_26311,N_26278);
or U28302 (N_28302,N_25800,N_25610);
nor U28303 (N_28303,N_25855,N_26985);
nand U28304 (N_28304,N_26205,N_25532);
and U28305 (N_28305,N_25566,N_25522);
nor U28306 (N_28306,N_25508,N_25554);
or U28307 (N_28307,N_26302,N_25897);
nor U28308 (N_28308,N_25804,N_26518);
nand U28309 (N_28309,N_25899,N_25869);
xor U28310 (N_28310,N_25637,N_26173);
and U28311 (N_28311,N_26201,N_26873);
or U28312 (N_28312,N_25673,N_26532);
or U28313 (N_28313,N_26281,N_26311);
nand U28314 (N_28314,N_26888,N_25873);
xor U28315 (N_28315,N_26916,N_26328);
nor U28316 (N_28316,N_26592,N_26092);
and U28317 (N_28317,N_26306,N_25875);
xnor U28318 (N_28318,N_26832,N_25994);
and U28319 (N_28319,N_26295,N_26185);
nand U28320 (N_28320,N_26155,N_25569);
or U28321 (N_28321,N_26438,N_26509);
and U28322 (N_28322,N_26552,N_26958);
nand U28323 (N_28323,N_25637,N_25851);
xnor U28324 (N_28324,N_26997,N_26779);
or U28325 (N_28325,N_25632,N_26800);
nand U28326 (N_28326,N_25906,N_26310);
xnor U28327 (N_28327,N_26577,N_26994);
nand U28328 (N_28328,N_25790,N_26760);
xnor U28329 (N_28329,N_26308,N_26730);
nand U28330 (N_28330,N_25687,N_26233);
xnor U28331 (N_28331,N_25952,N_25881);
nand U28332 (N_28332,N_26953,N_26604);
nand U28333 (N_28333,N_26767,N_26013);
nand U28334 (N_28334,N_25878,N_26152);
nand U28335 (N_28335,N_26528,N_25801);
xor U28336 (N_28336,N_26288,N_25872);
or U28337 (N_28337,N_25878,N_26087);
nand U28338 (N_28338,N_26490,N_25993);
nand U28339 (N_28339,N_25950,N_26056);
or U28340 (N_28340,N_25667,N_26458);
or U28341 (N_28341,N_26147,N_26003);
nand U28342 (N_28342,N_25837,N_25746);
xnor U28343 (N_28343,N_26970,N_26760);
nand U28344 (N_28344,N_25521,N_26843);
nor U28345 (N_28345,N_26783,N_26039);
and U28346 (N_28346,N_26901,N_26974);
or U28347 (N_28347,N_26737,N_26816);
or U28348 (N_28348,N_26148,N_26143);
or U28349 (N_28349,N_26841,N_26267);
nand U28350 (N_28350,N_25881,N_25910);
or U28351 (N_28351,N_26634,N_26072);
and U28352 (N_28352,N_26924,N_26184);
and U28353 (N_28353,N_26525,N_25772);
xor U28354 (N_28354,N_26634,N_25750);
nand U28355 (N_28355,N_26057,N_26402);
xnor U28356 (N_28356,N_25659,N_25790);
and U28357 (N_28357,N_26074,N_26318);
xnor U28358 (N_28358,N_26854,N_26811);
and U28359 (N_28359,N_26297,N_26893);
or U28360 (N_28360,N_26708,N_26549);
or U28361 (N_28361,N_25955,N_25883);
xor U28362 (N_28362,N_26152,N_25536);
nor U28363 (N_28363,N_25943,N_26733);
xnor U28364 (N_28364,N_25607,N_26008);
nand U28365 (N_28365,N_25846,N_26084);
and U28366 (N_28366,N_26670,N_26130);
and U28367 (N_28367,N_26926,N_26563);
and U28368 (N_28368,N_26364,N_26964);
nand U28369 (N_28369,N_26533,N_26719);
and U28370 (N_28370,N_26103,N_25703);
nand U28371 (N_28371,N_26214,N_25647);
nand U28372 (N_28372,N_25694,N_25739);
xnor U28373 (N_28373,N_26038,N_26464);
nand U28374 (N_28374,N_26486,N_26889);
or U28375 (N_28375,N_26119,N_26757);
nor U28376 (N_28376,N_25607,N_26505);
or U28377 (N_28377,N_26128,N_26467);
nand U28378 (N_28378,N_26519,N_26716);
nor U28379 (N_28379,N_26594,N_26381);
nor U28380 (N_28380,N_25969,N_26837);
nand U28381 (N_28381,N_25683,N_26941);
nor U28382 (N_28382,N_26133,N_25781);
nor U28383 (N_28383,N_26339,N_26783);
xnor U28384 (N_28384,N_26412,N_26180);
nand U28385 (N_28385,N_26107,N_25718);
and U28386 (N_28386,N_25859,N_26769);
nand U28387 (N_28387,N_26411,N_26598);
and U28388 (N_28388,N_26033,N_26670);
nand U28389 (N_28389,N_25958,N_26292);
or U28390 (N_28390,N_26646,N_25835);
or U28391 (N_28391,N_26025,N_26176);
and U28392 (N_28392,N_26808,N_25987);
nand U28393 (N_28393,N_26777,N_26418);
nor U28394 (N_28394,N_26200,N_25968);
nand U28395 (N_28395,N_26052,N_26162);
and U28396 (N_28396,N_26832,N_26909);
nand U28397 (N_28397,N_25780,N_26798);
and U28398 (N_28398,N_26077,N_26216);
xnor U28399 (N_28399,N_25903,N_26992);
nor U28400 (N_28400,N_26685,N_26790);
or U28401 (N_28401,N_26300,N_26621);
or U28402 (N_28402,N_26391,N_25963);
nor U28403 (N_28403,N_26356,N_25674);
nor U28404 (N_28404,N_26208,N_26657);
and U28405 (N_28405,N_25714,N_26765);
nand U28406 (N_28406,N_25959,N_25634);
nand U28407 (N_28407,N_25512,N_26639);
and U28408 (N_28408,N_26861,N_26069);
nor U28409 (N_28409,N_25848,N_26708);
nand U28410 (N_28410,N_25534,N_26776);
or U28411 (N_28411,N_26560,N_26916);
and U28412 (N_28412,N_26704,N_25835);
and U28413 (N_28413,N_26028,N_25981);
nor U28414 (N_28414,N_25781,N_26344);
nor U28415 (N_28415,N_26620,N_25660);
or U28416 (N_28416,N_25866,N_26110);
xor U28417 (N_28417,N_26759,N_25988);
nor U28418 (N_28418,N_26937,N_26172);
xor U28419 (N_28419,N_26152,N_26944);
nor U28420 (N_28420,N_25895,N_26098);
nor U28421 (N_28421,N_26574,N_25585);
nand U28422 (N_28422,N_25860,N_26232);
nand U28423 (N_28423,N_26552,N_26292);
and U28424 (N_28424,N_26451,N_25577);
and U28425 (N_28425,N_26783,N_26372);
or U28426 (N_28426,N_26250,N_25890);
and U28427 (N_28427,N_26795,N_26630);
nand U28428 (N_28428,N_26190,N_26774);
xnor U28429 (N_28429,N_26210,N_25836);
nor U28430 (N_28430,N_26258,N_26063);
or U28431 (N_28431,N_25566,N_26807);
nand U28432 (N_28432,N_26685,N_25856);
and U28433 (N_28433,N_25582,N_25806);
nand U28434 (N_28434,N_25798,N_26741);
nor U28435 (N_28435,N_25638,N_25661);
xnor U28436 (N_28436,N_25700,N_25960);
nand U28437 (N_28437,N_26476,N_25660);
nor U28438 (N_28438,N_26380,N_26180);
and U28439 (N_28439,N_26117,N_25669);
nor U28440 (N_28440,N_26548,N_25950);
and U28441 (N_28441,N_26797,N_26576);
or U28442 (N_28442,N_26765,N_26215);
or U28443 (N_28443,N_26938,N_26203);
or U28444 (N_28444,N_26061,N_26501);
and U28445 (N_28445,N_26120,N_26543);
nand U28446 (N_28446,N_25766,N_25792);
xor U28447 (N_28447,N_26016,N_25933);
nor U28448 (N_28448,N_25972,N_26492);
nor U28449 (N_28449,N_25686,N_26104);
nor U28450 (N_28450,N_26894,N_26380);
nor U28451 (N_28451,N_25898,N_26110);
nand U28452 (N_28452,N_26679,N_26974);
or U28453 (N_28453,N_25510,N_26739);
nor U28454 (N_28454,N_26806,N_26769);
or U28455 (N_28455,N_26698,N_26945);
or U28456 (N_28456,N_26321,N_25746);
nand U28457 (N_28457,N_26764,N_26572);
nand U28458 (N_28458,N_25900,N_25516);
nor U28459 (N_28459,N_25972,N_26095);
or U28460 (N_28460,N_26092,N_26454);
xnor U28461 (N_28461,N_25607,N_25591);
or U28462 (N_28462,N_26553,N_26070);
nand U28463 (N_28463,N_26668,N_26284);
nand U28464 (N_28464,N_25504,N_26652);
nor U28465 (N_28465,N_26369,N_26800);
nand U28466 (N_28466,N_26313,N_25807);
nor U28467 (N_28467,N_25855,N_26582);
and U28468 (N_28468,N_25714,N_26108);
or U28469 (N_28469,N_26241,N_25593);
nand U28470 (N_28470,N_26002,N_26120);
and U28471 (N_28471,N_26629,N_26421);
nor U28472 (N_28472,N_26644,N_26072);
xnor U28473 (N_28473,N_26112,N_25578);
nor U28474 (N_28474,N_25926,N_25687);
or U28475 (N_28475,N_26653,N_25651);
nand U28476 (N_28476,N_26609,N_26305);
nor U28477 (N_28477,N_26061,N_25825);
nand U28478 (N_28478,N_26977,N_26699);
nor U28479 (N_28479,N_26790,N_25566);
xnor U28480 (N_28480,N_26597,N_26673);
xor U28481 (N_28481,N_25650,N_26554);
or U28482 (N_28482,N_26368,N_25512);
or U28483 (N_28483,N_25912,N_26046);
and U28484 (N_28484,N_26363,N_25568);
or U28485 (N_28485,N_25624,N_26879);
nand U28486 (N_28486,N_25955,N_26849);
and U28487 (N_28487,N_25949,N_26034);
and U28488 (N_28488,N_25978,N_26195);
xnor U28489 (N_28489,N_26356,N_25602);
xnor U28490 (N_28490,N_26538,N_25528);
nand U28491 (N_28491,N_26381,N_26731);
nand U28492 (N_28492,N_26846,N_26348);
and U28493 (N_28493,N_26880,N_25838);
or U28494 (N_28494,N_25804,N_26812);
nand U28495 (N_28495,N_26715,N_26827);
nor U28496 (N_28496,N_26589,N_25628);
or U28497 (N_28497,N_26165,N_26020);
and U28498 (N_28498,N_26634,N_26807);
and U28499 (N_28499,N_26113,N_26362);
nand U28500 (N_28500,N_28312,N_27406);
nor U28501 (N_28501,N_28175,N_27989);
nor U28502 (N_28502,N_28195,N_27986);
and U28503 (N_28503,N_27946,N_27473);
or U28504 (N_28504,N_28329,N_28033);
nand U28505 (N_28505,N_27045,N_27896);
or U28506 (N_28506,N_28346,N_27366);
or U28507 (N_28507,N_27171,N_28478);
or U28508 (N_28508,N_28365,N_28088);
nand U28509 (N_28509,N_28288,N_27900);
nand U28510 (N_28510,N_27879,N_28093);
nor U28511 (N_28511,N_27584,N_28452);
nor U28512 (N_28512,N_28157,N_28462);
nand U28513 (N_28513,N_27567,N_27590);
or U28514 (N_28514,N_28366,N_27558);
or U28515 (N_28515,N_28274,N_27095);
and U28516 (N_28516,N_27904,N_27571);
xor U28517 (N_28517,N_27371,N_27310);
nor U28518 (N_28518,N_28063,N_28078);
xor U28519 (N_28519,N_27493,N_27538);
or U28520 (N_28520,N_27891,N_27942);
nor U28521 (N_28521,N_27856,N_28160);
or U28522 (N_28522,N_27870,N_27049);
nand U28523 (N_28523,N_27168,N_28412);
and U28524 (N_28524,N_28193,N_27104);
xnor U28525 (N_28525,N_28181,N_27597);
nor U28526 (N_28526,N_27144,N_27370);
nand U28527 (N_28527,N_28041,N_28013);
xnor U28528 (N_28528,N_27160,N_27350);
nor U28529 (N_28529,N_27710,N_27541);
and U28530 (N_28530,N_27809,N_27886);
or U28531 (N_28531,N_28451,N_27209);
and U28532 (N_28532,N_27062,N_27740);
or U28533 (N_28533,N_28330,N_27645);
or U28534 (N_28534,N_27549,N_28262);
nor U28535 (N_28535,N_27139,N_28189);
nand U28536 (N_28536,N_27253,N_28182);
xnor U28537 (N_28537,N_27353,N_28489);
or U28538 (N_28538,N_28018,N_27014);
xor U28539 (N_28539,N_27502,N_28048);
nor U28540 (N_28540,N_28449,N_28421);
and U28541 (N_28541,N_27529,N_27758);
nand U28542 (N_28542,N_27076,N_28126);
or U28543 (N_28543,N_28373,N_28153);
nand U28544 (N_28544,N_28315,N_27706);
nand U28545 (N_28545,N_28415,N_27823);
nand U28546 (N_28546,N_27179,N_27121);
nand U28547 (N_28547,N_28128,N_28375);
and U28548 (N_28548,N_27707,N_27781);
xnor U28549 (N_28549,N_28019,N_27734);
nand U28550 (N_28550,N_28463,N_28309);
xor U28551 (N_28551,N_27671,N_27569);
xnor U28552 (N_28552,N_27576,N_27991);
nor U28553 (N_28553,N_27196,N_28265);
nand U28554 (N_28554,N_28176,N_27820);
nand U28555 (N_28555,N_28453,N_28065);
and U28556 (N_28556,N_28227,N_27853);
nor U28557 (N_28557,N_27688,N_27336);
or U28558 (N_28558,N_27704,N_27197);
or U28559 (N_28559,N_27977,N_27928);
nand U28560 (N_28560,N_27507,N_28215);
xor U28561 (N_28561,N_27939,N_27323);
and U28562 (N_28562,N_28161,N_27804);
and U28563 (N_28563,N_27691,N_27627);
or U28564 (N_28564,N_27771,N_28199);
nand U28565 (N_28565,N_27748,N_27481);
nor U28566 (N_28566,N_27659,N_27960);
xnor U28567 (N_28567,N_27830,N_27134);
nor U28568 (N_28568,N_28214,N_27414);
xnor U28569 (N_28569,N_27916,N_27285);
and U28570 (N_28570,N_27772,N_27191);
nand U28571 (N_28571,N_27182,N_27093);
xor U28572 (N_28572,N_28276,N_27965);
and U28573 (N_28573,N_27317,N_28285);
or U28574 (N_28574,N_27511,N_27801);
and U28575 (N_28575,N_27954,N_27446);
or U28576 (N_28576,N_28247,N_28409);
and U28577 (N_28577,N_28235,N_28219);
xnor U28578 (N_28578,N_28370,N_27409);
nor U28579 (N_28579,N_27255,N_27447);
or U28580 (N_28580,N_27060,N_27193);
nand U28581 (N_28581,N_27633,N_27454);
xnor U28582 (N_28582,N_28258,N_27422);
or U28583 (N_28583,N_27556,N_28224);
xnor U28584 (N_28584,N_27925,N_28359);
nor U28585 (N_28585,N_28149,N_27485);
and U28586 (N_28586,N_27090,N_27848);
or U28587 (N_28587,N_27899,N_28143);
nand U28588 (N_28588,N_28098,N_27372);
and U28589 (N_28589,N_27073,N_27390);
and U28590 (N_28590,N_27222,N_27113);
nor U28591 (N_28591,N_28113,N_27137);
or U28592 (N_28592,N_28021,N_28269);
and U28593 (N_28593,N_27059,N_27037);
xor U28594 (N_28594,N_28356,N_27774);
nand U28595 (N_28595,N_27194,N_27387);
xor U28596 (N_28596,N_27973,N_27570);
xnor U28597 (N_28597,N_27015,N_27091);
nor U28598 (N_28598,N_28408,N_27933);
nor U28599 (N_28599,N_27065,N_27419);
xor U28600 (N_28600,N_27992,N_28164);
nor U28601 (N_28601,N_27302,N_27564);
xnor U28602 (N_28602,N_27079,N_27423);
nand U28603 (N_28603,N_27282,N_28147);
nor U28604 (N_28604,N_27509,N_28146);
or U28605 (N_28605,N_28395,N_27002);
and U28606 (N_28606,N_27996,N_28280);
xnor U28607 (N_28607,N_28135,N_27826);
or U28608 (N_28608,N_27180,N_27924);
or U28609 (N_28609,N_27273,N_27777);
nor U28610 (N_28610,N_27100,N_27554);
xnor U28611 (N_28611,N_27403,N_28349);
nor U28612 (N_28612,N_28045,N_27984);
xor U28613 (N_28613,N_28059,N_28180);
and U28614 (N_28614,N_27177,N_27382);
nand U28615 (N_28615,N_27877,N_27839);
and U28616 (N_28616,N_27822,N_28188);
xor U28617 (N_28617,N_27794,N_27543);
nand U28618 (N_28618,N_28350,N_27752);
xor U28619 (N_28619,N_27220,N_27525);
xor U28620 (N_28620,N_28481,N_27919);
nor U28621 (N_28621,N_27604,N_27985);
and U28622 (N_28622,N_28095,N_27724);
or U28623 (N_28623,N_27766,N_28191);
nor U28624 (N_28624,N_27844,N_27574);
xnor U28625 (N_28625,N_28005,N_28460);
xor U28626 (N_28626,N_27440,N_28347);
nand U28627 (N_28627,N_27813,N_27703);
nand U28628 (N_28628,N_27250,N_27239);
nand U28629 (N_28629,N_27467,N_28081);
or U28630 (N_28630,N_27845,N_27184);
nor U28631 (N_28631,N_28364,N_27269);
or U28632 (N_28632,N_27229,N_27640);
xor U28633 (N_28633,N_28355,N_27351);
or U28634 (N_28634,N_27270,N_27195);
and U28635 (N_28635,N_28301,N_27178);
nand U28636 (N_28636,N_28099,N_27625);
and U28637 (N_28637,N_28456,N_27666);
nand U28638 (N_28638,N_27782,N_28454);
xor U28639 (N_28639,N_27892,N_27364);
nor U28640 (N_28640,N_28084,N_27869);
xnor U28641 (N_28641,N_27593,N_27424);
and U28642 (N_28642,N_28000,N_27030);
nor U28643 (N_28643,N_27299,N_28020);
or U28644 (N_28644,N_27040,N_28290);
or U28645 (N_28645,N_27346,N_28251);
or U28646 (N_28646,N_28470,N_28034);
nor U28647 (N_28647,N_27316,N_27398);
xnor U28648 (N_28648,N_28233,N_27937);
and U28649 (N_28649,N_28402,N_28061);
or U28650 (N_28650,N_28232,N_27138);
nor U28651 (N_28651,N_28256,N_27715);
nand U28652 (N_28652,N_27594,N_27621);
or U28653 (N_28653,N_28221,N_28414);
nor U28654 (N_28654,N_27289,N_27784);
nand U28655 (N_28655,N_27235,N_28400);
nand U28656 (N_28656,N_27259,N_27321);
xor U28657 (N_28657,N_28142,N_27486);
nand U28658 (N_28658,N_27755,N_27940);
nand U28659 (N_28659,N_27871,N_27243);
nor U28660 (N_28660,N_28371,N_28319);
nor U28661 (N_28661,N_27808,N_27975);
and U28662 (N_28662,N_27341,N_28044);
or U28663 (N_28663,N_27883,N_27477);
nor U28664 (N_28664,N_27976,N_28039);
nand U28665 (N_28665,N_28066,N_27491);
nand U28666 (N_28666,N_27494,N_27663);
xnor U28667 (N_28667,N_27944,N_27320);
nor U28668 (N_28668,N_27544,N_28442);
xnor U28669 (N_28669,N_27585,N_27578);
nand U28670 (N_28670,N_28079,N_27212);
nand U28671 (N_28671,N_27034,N_27639);
or U28672 (N_28672,N_27022,N_28008);
nand U28673 (N_28673,N_28374,N_27327);
or U28674 (N_28674,N_27055,N_27797);
or U28675 (N_28675,N_28343,N_27990);
and U28676 (N_28676,N_27629,N_27394);
nand U28677 (N_28677,N_28060,N_28007);
and U28678 (N_28678,N_27747,N_28130);
and U28679 (N_28679,N_27611,N_27972);
nand U28680 (N_28680,N_27169,N_27967);
nor U28681 (N_28681,N_27118,N_27929);
nor U28682 (N_28682,N_27938,N_28255);
and U28683 (N_28683,N_27889,N_27651);
nor U28684 (N_28684,N_27729,N_27654);
nor U28685 (N_28685,N_28397,N_27648);
or U28686 (N_28686,N_27343,N_28268);
nor U28687 (N_28687,N_27738,N_27678);
nand U28688 (N_28688,N_28090,N_28448);
xor U28689 (N_28689,N_28390,N_28335);
nor U28690 (N_28690,N_27412,N_28138);
xnor U28691 (N_28691,N_27817,N_27769);
nor U28692 (N_28692,N_27070,N_27381);
xnor U28693 (N_28693,N_28393,N_27634);
xnor U28694 (N_28694,N_27218,N_28396);
nor U28695 (N_28695,N_27489,N_28302);
nor U28696 (N_28696,N_27643,N_28197);
nand U28697 (N_28697,N_27153,N_27162);
nand U28698 (N_28698,N_27997,N_27679);
xor U28699 (N_28699,N_27542,N_28417);
and U28700 (N_28700,N_28477,N_27515);
nand U28701 (N_28701,N_27921,N_27411);
or U28702 (N_28702,N_27290,N_27147);
xor U28703 (N_28703,N_27374,N_27264);
or U28704 (N_28704,N_27850,N_27297);
or U28705 (N_28705,N_28447,N_28002);
or U28706 (N_28706,N_27716,N_27665);
nand U28707 (N_28707,N_28490,N_27770);
nor U28708 (N_28708,N_28017,N_28497);
nor U28709 (N_28709,N_28245,N_27860);
or U28710 (N_28710,N_27741,N_27945);
and U28711 (N_28711,N_27257,N_27616);
nor U28712 (N_28712,N_27221,N_27893);
nor U28713 (N_28713,N_27814,N_27968);
nor U28714 (N_28714,N_27025,N_27623);
nor U28715 (N_28715,N_28201,N_27136);
nand U28716 (N_28716,N_28196,N_28441);
and U28717 (N_28717,N_27727,N_27119);
or U28718 (N_28718,N_28213,N_27154);
nand U28719 (N_28719,N_27789,N_28484);
xnor U28720 (N_28720,N_27956,N_27545);
nand U28721 (N_28721,N_28133,N_28054);
and U28722 (N_28722,N_28119,N_27152);
xor U28723 (N_28723,N_27677,N_28464);
or U28724 (N_28724,N_27547,N_27697);
xnor U28725 (N_28725,N_27488,N_27557);
nor U28726 (N_28726,N_27998,N_28023);
nand U28727 (N_28727,N_28275,N_28310);
nand U28728 (N_28728,N_28058,N_27818);
and U28729 (N_28729,N_27568,N_27686);
xnor U28730 (N_28730,N_28206,N_27628);
or U28731 (N_28731,N_27252,N_28291);
nor U28732 (N_28732,N_27463,N_28123);
or U28733 (N_28733,N_27490,N_27476);
nor U28734 (N_28734,N_27779,N_27081);
nand U28735 (N_28735,N_28073,N_27051);
nand U28736 (N_28736,N_27609,N_27334);
and U28737 (N_28737,N_27635,N_27834);
and U28738 (N_28738,N_28419,N_27452);
nand U28739 (N_28739,N_27895,N_27326);
and U28740 (N_28740,N_27456,N_28173);
nor U28741 (N_28741,N_28223,N_27167);
and U28742 (N_28742,N_27949,N_28218);
and U28743 (N_28743,N_28230,N_27805);
nor U28744 (N_28744,N_28372,N_28434);
nand U28745 (N_28745,N_27497,N_27393);
xnor U28746 (N_28746,N_27790,N_28340);
or U28747 (N_28747,N_27792,N_28498);
nand U28748 (N_28748,N_27248,N_27338);
xnor U28749 (N_28749,N_27237,N_28314);
xor U28750 (N_28750,N_27472,N_28328);
nand U28751 (N_28751,N_28381,N_27943);
and U28752 (N_28752,N_27052,N_28384);
and U28753 (N_28753,N_28169,N_28071);
and U28754 (N_28754,N_28234,N_28367);
xor U28755 (N_28755,N_28422,N_27001);
xnor U28756 (N_28756,N_27263,N_27355);
and U28757 (N_28757,N_27607,N_28237);
xor U28758 (N_28758,N_27254,N_28184);
nand U28759 (N_28759,N_27438,N_28363);
and U28760 (N_28760,N_27630,N_27032);
or U28761 (N_28761,N_28016,N_27717);
or U28762 (N_28762,N_28110,N_27133);
nand U28763 (N_28763,N_27934,N_27332);
nor U28764 (N_28764,N_27258,N_28420);
xnor U28765 (N_28765,N_28185,N_27961);
and U28766 (N_28766,N_27078,N_27386);
nor U28767 (N_28767,N_28103,N_28150);
nand U28768 (N_28768,N_28337,N_27425);
and U28769 (N_28769,N_27026,N_28287);
xnor U28770 (N_28770,N_28051,N_28226);
and U28771 (N_28771,N_27847,N_27760);
nor U28772 (N_28772,N_27508,N_27518);
nand U28773 (N_28773,N_27745,N_28010);
nor U28774 (N_28774,N_27329,N_27132);
and U28775 (N_28775,N_27385,N_27527);
or U28776 (N_28776,N_27214,N_27287);
or U28777 (N_28777,N_27474,N_28158);
or U28778 (N_28778,N_28148,N_27271);
xor U28779 (N_28779,N_27107,N_28012);
nor U28780 (N_28780,N_27711,N_27066);
nor U28781 (N_28781,N_27458,N_27009);
xnor U28782 (N_28782,N_27595,N_27783);
nand U28783 (N_28783,N_28487,N_27356);
or U28784 (N_28784,N_28488,N_27159);
nand U28785 (N_28785,N_28465,N_28125);
xor U28786 (N_28786,N_27999,N_27482);
or U28787 (N_28787,N_27101,N_27638);
xnor U28788 (N_28788,N_28202,N_28190);
or U28789 (N_28789,N_27471,N_28198);
or U28790 (N_28790,N_27097,N_28283);
nand U28791 (N_28791,N_28458,N_27964);
and U28792 (N_28792,N_27764,N_27314);
nand U28793 (N_28793,N_28252,N_27203);
and U28794 (N_28794,N_27459,N_28351);
nor U28795 (N_28795,N_28122,N_27156);
and U28796 (N_28796,N_27583,N_28222);
nor U28797 (N_28797,N_27714,N_27384);
xnor U28798 (N_28798,N_27658,N_27441);
nand U28799 (N_28799,N_27721,N_27106);
or U28800 (N_28800,N_28399,N_27242);
or U28801 (N_28801,N_28229,N_28433);
nand U28802 (N_28802,N_28004,N_27662);
nor U28803 (N_28803,N_27007,N_27068);
and U28804 (N_28804,N_28239,N_28286);
nand U28805 (N_28805,N_27085,N_27876);
and U28806 (N_28806,N_27033,N_27499);
or U28807 (N_28807,N_28425,N_27361);
nand U28808 (N_28808,N_27131,N_27448);
xnor U28809 (N_28809,N_27231,N_28140);
nand U28810 (N_28810,N_27575,N_27298);
and U28811 (N_28811,N_27580,N_28137);
nor U28812 (N_28812,N_28096,N_27039);
nand U28813 (N_28813,N_27276,N_27402);
nand U28814 (N_28814,N_27181,N_27827);
and U28815 (N_28815,N_27922,N_28313);
nor U28816 (N_28816,N_27735,N_27315);
and U28817 (N_28817,N_27852,N_28424);
nand U28818 (N_28818,N_27751,N_27465);
nor U28819 (N_28819,N_27552,N_27342);
xor U28820 (N_28820,N_27660,N_28210);
nor U28821 (N_28821,N_28134,N_28102);
xor U28822 (N_28822,N_27010,N_27731);
nor U28823 (N_28823,N_28294,N_27086);
xor U28824 (N_28824,N_27624,N_28032);
nand U28825 (N_28825,N_27176,N_27516);
nor U28826 (N_28826,N_27418,N_27140);
and U28827 (N_28827,N_27036,N_27466);
xor U28828 (N_28828,N_28411,N_28480);
nand U28829 (N_28829,N_28323,N_27931);
and U28830 (N_28830,N_27145,N_28334);
xnor U28831 (N_28831,N_27069,N_28388);
or U28832 (N_28832,N_28131,N_27498);
xnor U28833 (N_28833,N_27442,N_27056);
nand U28834 (N_28834,N_27304,N_27468);
nor U28835 (N_28835,N_27434,N_28357);
xor U28836 (N_28836,N_27786,N_27846);
and U28837 (N_28837,N_27027,N_28124);
and U28838 (N_28838,N_28220,N_27496);
or U28839 (N_28839,N_27071,N_28322);
and U28840 (N_28840,N_27701,N_27428);
or U28841 (N_28841,N_27200,N_27565);
nand U28842 (N_28842,N_27318,N_27331);
nand U28843 (N_28843,N_27513,N_28014);
xnor U28844 (N_28844,N_28321,N_27912);
and U28845 (N_28845,N_28423,N_27480);
xnor U28846 (N_28846,N_28459,N_27028);
xor U28847 (N_28847,N_28211,N_27275);
xnor U28848 (N_28848,N_27280,N_27308);
and U28849 (N_28849,N_28072,N_28391);
xor U28850 (N_28850,N_27105,N_27344);
or U28851 (N_28851,N_27533,N_27897);
xor U28852 (N_28852,N_27918,N_27395);
nand U28853 (N_28853,N_28281,N_28339);
xor U28854 (N_28854,N_27462,N_27043);
and U28855 (N_28855,N_27311,N_27828);
and U28856 (N_28856,N_27882,N_27894);
xnor U28857 (N_28857,N_27548,N_28295);
nor U28858 (N_28858,N_27358,N_27966);
nand U28859 (N_28859,N_27859,N_27146);
xor U28860 (N_28860,N_27802,N_27292);
nand U28861 (N_28861,N_28141,N_28368);
and U28862 (N_28862,N_27003,N_27560);
nand U28863 (N_28863,N_27608,N_28076);
nand U28864 (N_28864,N_27199,N_28426);
xor U28865 (N_28865,N_27941,N_27911);
and U28866 (N_28866,N_28022,N_27685);
xor U28867 (N_28867,N_27088,N_27713);
xnor U28868 (N_28868,N_27261,N_27019);
and U28869 (N_28869,N_27955,N_28062);
nor U28870 (N_28870,N_28431,N_28289);
nor U28871 (N_28871,N_27204,N_28109);
nor U28872 (N_28872,N_27504,N_27680);
xor U28873 (N_28873,N_27410,N_27413);
and U28874 (N_28874,N_27664,N_27301);
nand U28875 (N_28875,N_28293,N_27103);
and U28876 (N_28876,N_27234,N_27993);
or U28877 (N_28877,N_27572,N_27619);
xnor U28878 (N_28878,N_28476,N_27775);
and U28879 (N_28879,N_28491,N_28042);
and U28880 (N_28880,N_28468,N_28318);
nand U28881 (N_28881,N_27158,N_28435);
nor U28882 (N_28882,N_27464,N_27857);
or U28883 (N_28883,N_27247,N_27722);
nand U28884 (N_28884,N_27586,N_27682);
nor U28885 (N_28885,N_28485,N_28001);
nor U28886 (N_28886,N_27063,N_28474);
and U28887 (N_28887,N_27982,N_28067);
nor U28888 (N_28888,N_27155,N_27753);
or U28889 (N_28889,N_28087,N_27987);
xor U28890 (N_28890,N_27503,N_27469);
and U28891 (N_28891,N_28398,N_27267);
nor U28892 (N_28892,N_28111,N_27878);
xor U28893 (N_28893,N_27534,N_27436);
and U28894 (N_28894,N_28348,N_28244);
or U28895 (N_28895,N_28055,N_27661);
and U28896 (N_28896,N_27354,N_28186);
xor U28897 (N_28897,N_28483,N_27021);
nand U28898 (N_28898,N_27362,N_27487);
nand U28899 (N_28899,N_27072,N_27652);
or U28900 (N_28900,N_27401,N_27700);
nand U28901 (N_28901,N_27868,N_28282);
and U28902 (N_28902,N_27863,N_27453);
xor U28903 (N_28903,N_27577,N_27613);
and U28904 (N_28904,N_28404,N_27175);
and U28905 (N_28905,N_27127,N_28332);
nor U28906 (N_28906,N_27500,N_27189);
xor U28907 (N_28907,N_27192,N_27379);
nand U28908 (N_28908,N_27262,N_28106);
nand U28909 (N_28909,N_27008,N_27053);
and U28910 (N_28910,N_27683,N_28163);
xor U28911 (N_28911,N_27296,N_27979);
xor U28912 (N_28912,N_27884,N_28466);
xnor U28913 (N_28913,N_27368,N_27050);
or U28914 (N_28914,N_27305,N_27205);
xor U28915 (N_28915,N_27617,N_27404);
xnor U28916 (N_28916,N_27849,N_28246);
xor U28917 (N_28917,N_28089,N_27684);
or U28918 (N_28918,N_27018,N_28165);
and U28919 (N_28919,N_28212,N_28264);
and U28920 (N_28920,N_28139,N_27303);
or U28921 (N_28921,N_27631,N_27375);
or U28922 (N_28922,N_27274,N_27690);
nor U28923 (N_28923,N_27907,N_28405);
or U28924 (N_28924,N_27952,N_27978);
nand U28925 (N_28925,N_27125,N_27596);
nand U28926 (N_28926,N_27286,N_28338);
nor U28927 (N_28927,N_28410,N_27102);
or U28928 (N_28928,N_28192,N_27720);
nor U28929 (N_28929,N_28216,N_27759);
nand U28930 (N_28930,N_28317,N_28052);
nor U28931 (N_28931,N_27219,N_27444);
or U28932 (N_28932,N_28473,N_27730);
xor U28933 (N_28933,N_28241,N_27793);
or U28934 (N_28934,N_28151,N_28207);
nand U28935 (N_28935,N_28406,N_28177);
xor U28936 (N_28936,N_27475,N_27392);
or U28937 (N_28937,N_27673,N_27217);
and U28938 (N_28938,N_27913,N_27064);
and U28939 (N_28939,N_28438,N_27970);
nand U28940 (N_28940,N_27388,N_27359);
nor U28941 (N_28941,N_28116,N_27672);
xnor U28942 (N_28942,N_27562,N_28053);
nand U28943 (N_28943,N_27833,N_27732);
and U28944 (N_28944,N_27957,N_27898);
nand U28945 (N_28945,N_28171,N_28068);
nand U28946 (N_28946,N_27185,N_27719);
or U28947 (N_28947,N_27811,N_27902);
and U28948 (N_28948,N_27551,N_28430);
xnor U28949 (N_28949,N_27610,N_27561);
and U28950 (N_28950,N_28205,N_27130);
nand U28951 (N_28951,N_27825,N_28194);
and U28952 (N_28952,N_27872,N_28324);
and U28953 (N_28953,N_28209,N_27099);
nand U28954 (N_28954,N_27123,N_27373);
and U28955 (N_28955,N_27867,N_27116);
nand U28956 (N_28956,N_27540,N_27761);
and U28957 (N_28957,N_27950,N_27693);
nor U28958 (N_28958,N_27251,N_27689);
xor U28959 (N_28959,N_27492,N_28263);
nor U28960 (N_28960,N_28178,N_27294);
and U28961 (N_28961,N_27457,N_28077);
nor U28962 (N_28962,N_28311,N_28242);
nor U28963 (N_28963,N_27216,N_28037);
xor U28964 (N_28964,N_27512,N_28174);
or U28965 (N_28965,N_27166,N_27405);
nor U28966 (N_28966,N_28006,N_27582);
and U28967 (N_28967,N_27959,N_28046);
or U28968 (N_28968,N_28272,N_27708);
xnor U28969 (N_28969,N_27224,N_27926);
and U28970 (N_28970,N_28240,N_27519);
or U28971 (N_28971,N_27841,N_27378);
and U28972 (N_28972,N_27750,N_28080);
and U28973 (N_28973,N_28027,N_27958);
or U28974 (N_28974,N_27246,N_27389);
and U28975 (N_28975,N_27754,N_28117);
xnor U28976 (N_28976,N_27260,N_28166);
nand U28977 (N_28977,N_27363,N_27803);
and U28978 (N_28978,N_28091,N_27526);
nor U28979 (N_28979,N_27537,N_28386);
nor U28980 (N_28980,N_27749,N_27020);
nand U28981 (N_28981,N_27799,N_27330);
xor U28982 (N_28982,N_27426,N_28277);
nand U28983 (N_28983,N_27864,N_27328);
xor U28984 (N_28984,N_27161,N_28354);
nand U28985 (N_28985,N_27006,N_27550);
xnor U28986 (N_28986,N_27953,N_27031);
xnor U28987 (N_28987,N_28248,N_27909);
or U28988 (N_28988,N_27851,N_27888);
and U28989 (N_28989,N_28450,N_27762);
xnor U28990 (N_28990,N_27699,N_28273);
or U28991 (N_28991,N_28308,N_27279);
nand U28992 (N_28992,N_27129,N_27041);
nand U28993 (N_28993,N_28154,N_28494);
xor U28994 (N_28994,N_28187,N_27377);
or U28995 (N_28995,N_27521,N_28461);
or U28996 (N_28996,N_27058,N_28170);
xor U28997 (N_28997,N_27461,N_27213);
or U28998 (N_28998,N_28035,N_27670);
nand U28999 (N_28999,N_27000,N_27974);
or U29000 (N_29000,N_27520,N_27054);
and U29001 (N_29001,N_27245,N_27807);
xnor U29002 (N_29002,N_27187,N_28204);
and U29003 (N_29003,N_28394,N_27238);
nor U29004 (N_29004,N_27756,N_28432);
and U29005 (N_29005,N_28009,N_28376);
nand U29006 (N_29006,N_27215,N_27249);
or U29007 (N_29007,N_27449,N_27824);
xnor U29008 (N_29008,N_27380,N_27636);
or U29009 (N_29009,N_27591,N_28118);
nand U29010 (N_29010,N_27819,N_28443);
nand U29011 (N_29011,N_28025,N_28050);
xnor U29012 (N_29012,N_27046,N_28107);
and U29013 (N_29013,N_27995,N_28145);
or U29014 (N_29014,N_28026,N_28385);
xnor U29015 (N_29015,N_27906,N_27324);
or U29016 (N_29016,N_27650,N_27962);
xor U29017 (N_29017,N_27074,N_27620);
nand U29018 (N_29018,N_28307,N_28049);
nand U29019 (N_29019,N_27427,N_27173);
nand U29020 (N_29020,N_27932,N_28299);
xor U29021 (N_29021,N_27163,N_27695);
nor U29022 (N_29022,N_28352,N_27432);
and U29023 (N_29023,N_28467,N_27483);
nand U29024 (N_29024,N_27837,N_27044);
or U29025 (N_29025,N_27531,N_27865);
nor U29026 (N_29026,N_27908,N_27861);
xnor U29027 (N_29027,N_27687,N_27603);
nand U29028 (N_29028,N_27875,N_27005);
nor U29029 (N_29029,N_27035,N_27349);
nor U29030 (N_29030,N_27881,N_28416);
nor U29031 (N_29031,N_27587,N_28445);
nor U29032 (N_29032,N_27470,N_28361);
nor U29033 (N_29033,N_27528,N_28257);
nand U29034 (N_29034,N_27626,N_27559);
nor U29035 (N_29035,N_27098,N_27293);
nor U29036 (N_29036,N_27232,N_27082);
and U29037 (N_29037,N_28208,N_27935);
and U29038 (N_29038,N_28260,N_27675);
xnor U29039 (N_29039,N_27765,N_28378);
nand U29040 (N_29040,N_28493,N_27641);
xnor U29041 (N_29041,N_27357,N_27208);
nor U29042 (N_29042,N_28336,N_27903);
xnor U29043 (N_29043,N_28362,N_27347);
nand U29044 (N_29044,N_28389,N_28112);
or U29045 (N_29045,N_27694,N_27170);
nor U29046 (N_29046,N_27592,N_28475);
nor U29047 (N_29047,N_27223,N_28392);
and U29048 (N_29048,N_27495,N_27295);
nor U29049 (N_29049,N_27075,N_27435);
and U29050 (N_29050,N_28094,N_27810);
nor U29051 (N_29051,N_27244,N_27506);
xnor U29052 (N_29052,N_27573,N_27836);
nor U29053 (N_29053,N_27742,N_27451);
xor U29054 (N_29054,N_28344,N_28203);
or U29055 (N_29055,N_27816,N_27971);
nor U29056 (N_29056,N_27674,N_28057);
xnor U29057 (N_29057,N_27230,N_27739);
nand U29058 (N_29058,N_27268,N_27120);
nor U29059 (N_29059,N_28437,N_28407);
and U29060 (N_29060,N_27142,N_28379);
nor U29061 (N_29061,N_27815,N_28297);
nand U29062 (N_29062,N_27011,N_27080);
or U29063 (N_29063,N_27705,N_27637);
or U29064 (N_29064,N_27433,N_27352);
or U29065 (N_29065,N_28030,N_27606);
and U29066 (N_29066,N_27157,N_28086);
or U29067 (N_29067,N_27601,N_28105);
and U29068 (N_29068,N_28292,N_27084);
or U29069 (N_29069,N_27360,N_27581);
and U29070 (N_29070,N_27667,N_27602);
nor U29071 (N_29071,N_28486,N_27337);
xnor U29072 (N_29072,N_28092,N_28070);
or U29073 (N_29073,N_27599,N_27284);
xnor U29074 (N_29074,N_27057,N_27291);
and U29075 (N_29075,N_27450,N_28029);
xnor U29076 (N_29076,N_27460,N_27981);
xnor U29077 (N_29077,N_27164,N_27016);
or U29078 (N_29078,N_27763,N_27647);
nor U29079 (N_29079,N_27455,N_27951);
xor U29080 (N_29080,N_27148,N_28254);
nand U29081 (N_29081,N_27709,N_28296);
nor U29082 (N_29082,N_27345,N_27842);
xor U29083 (N_29083,N_28228,N_27281);
or U29084 (N_29084,N_27210,N_27702);
xor U29085 (N_29085,N_27743,N_28469);
or U29086 (N_29086,N_27905,N_28267);
xnor U29087 (N_29087,N_27421,N_27277);
or U29088 (N_29088,N_27910,N_27077);
xor U29089 (N_29089,N_28429,N_27383);
or U29090 (N_29090,N_28104,N_28120);
xnor U29091 (N_29091,N_27188,N_27150);
nor U29092 (N_29092,N_28427,N_28031);
xor U29093 (N_29093,N_27914,N_27319);
nor U29094 (N_29094,N_28200,N_27901);
nand U29095 (N_29095,N_27795,N_27798);
nor U29096 (N_29096,N_27087,N_27887);
nand U29097 (N_29097,N_27484,N_27927);
nand U29098 (N_29098,N_28168,N_28064);
nand U29099 (N_29099,N_27283,N_27873);
and U29100 (N_29100,N_27517,N_28325);
nand U29101 (N_29101,N_27067,N_27443);
xor U29102 (N_29102,N_27920,N_28278);
or U29103 (N_29103,N_27111,N_27838);
nor U29104 (N_29104,N_27539,N_27092);
or U29105 (N_29105,N_27831,N_28038);
or U29106 (N_29106,N_27198,N_27416);
xnor U29107 (N_29107,N_27445,N_28382);
nor U29108 (N_29108,N_28179,N_27397);
nand U29109 (N_29109,N_27535,N_27796);
or U29110 (N_29110,N_27530,N_27431);
and U29111 (N_29111,N_28284,N_27325);
xnor U29112 (N_29112,N_28496,N_27439);
xor U29113 (N_29113,N_27126,N_27012);
or U29114 (N_29114,N_27649,N_28320);
nand U29115 (N_29115,N_27874,N_28108);
and U29116 (N_29116,N_27038,N_27832);
nand U29117 (N_29117,N_27698,N_27644);
nor U29118 (N_29118,N_27190,N_27202);
and U29119 (N_29119,N_28156,N_28333);
and U29120 (N_29120,N_27785,N_28418);
nand U29121 (N_29121,N_27791,N_27256);
xnor U29122 (N_29122,N_27135,N_27312);
and U29123 (N_29123,N_27430,N_28115);
or U29124 (N_29124,N_27122,N_28015);
xor U29125 (N_29125,N_28069,N_27174);
nand U29126 (N_29126,N_27367,N_27128);
nand U29127 (N_29127,N_27108,N_27278);
or U29128 (N_29128,N_28377,N_27478);
and U29129 (N_29129,N_28326,N_27186);
or U29130 (N_29130,N_27042,N_28011);
nor U29131 (N_29131,N_28056,N_27307);
xnor U29132 (N_29132,N_27365,N_27980);
xnor U29133 (N_29133,N_27109,N_28028);
or U29134 (N_29134,N_28492,N_28479);
and U29135 (N_29135,N_27306,N_27736);
or U29136 (N_29136,N_27013,N_28217);
and U29137 (N_29137,N_28253,N_28144);
and U29138 (N_29138,N_28305,N_27930);
or U29139 (N_29139,N_27335,N_28121);
and U29140 (N_29140,N_27646,N_27115);
xor U29141 (N_29141,N_27555,N_28387);
xor U29142 (N_29142,N_27963,N_27532);
nor U29143 (N_29143,N_27692,N_27149);
and U29144 (N_29144,N_27348,N_27376);
or U29145 (N_29145,N_28413,N_27206);
and U29146 (N_29146,N_27725,N_27553);
and U29147 (N_29147,N_27642,N_27211);
and U29148 (N_29148,N_27096,N_27728);
xor U29149 (N_29149,N_28082,N_28369);
nor U29150 (N_29150,N_28353,N_28162);
nor U29151 (N_29151,N_28074,N_27023);
nand U29152 (N_29152,N_27437,N_27969);
or U29153 (N_29153,N_28043,N_28183);
nand U29154 (N_29154,N_27510,N_27110);
nor U29155 (N_29155,N_28114,N_27915);
or U29156 (N_29156,N_27201,N_27773);
and U29157 (N_29157,N_27563,N_27612);
nor U29158 (N_29158,N_28440,N_27618);
nand U29159 (N_29159,N_28303,N_27800);
nor U29160 (N_29160,N_27588,N_28085);
nand U29161 (N_29161,N_27890,N_27744);
xnor U29162 (N_29162,N_27225,N_27048);
xor U29163 (N_29163,N_28482,N_27429);
nand U29164 (N_29164,N_28401,N_27265);
nand U29165 (N_29165,N_27241,N_27313);
or U29166 (N_29166,N_28040,N_27757);
or U29167 (N_29167,N_27632,N_27536);
or U29168 (N_29168,N_27117,N_28455);
and U29169 (N_29169,N_28358,N_27718);
and U29170 (N_29170,N_27712,N_27821);
and U29171 (N_29171,N_27524,N_27083);
nand U29172 (N_29172,N_27207,N_27615);
or U29173 (N_29173,N_28261,N_27733);
nor U29174 (N_29174,N_28100,N_27523);
and U29175 (N_29175,N_27309,N_28316);
or U29176 (N_29176,N_27089,N_27668);
and U29177 (N_29177,N_28249,N_28075);
nor U29178 (N_29178,N_28083,N_28279);
and U29179 (N_29179,N_27917,N_28152);
xnor U29180 (N_29180,N_27369,N_27236);
or U29181 (N_29181,N_27340,N_27505);
nand U29182 (N_29182,N_27726,N_27479);
xor U29183 (N_29183,N_27840,N_27114);
xor U29184 (N_29184,N_28167,N_27233);
or U29185 (N_29185,N_27657,N_27272);
and U29186 (N_29186,N_28127,N_28457);
nor U29187 (N_29187,N_27047,N_28472);
and U29188 (N_29188,N_27420,N_28444);
xor U29189 (N_29189,N_27061,N_27681);
nand U29190 (N_29190,N_27885,N_28243);
xor U29191 (N_29191,N_28250,N_27566);
nor U29192 (N_29192,N_27947,N_28471);
xor U29193 (N_29193,N_27546,N_27780);
xnor U29194 (N_29194,N_27656,N_27948);
nand U29195 (N_29195,N_28446,N_27787);
nor U29196 (N_29196,N_27143,N_28495);
or U29197 (N_29197,N_27829,N_28341);
or U29198 (N_29198,N_28101,N_27165);
and U29199 (N_29199,N_28236,N_28428);
or U29200 (N_29200,N_27622,N_28436);
nor U29201 (N_29201,N_27768,N_27300);
nand U29202 (N_29202,N_28024,N_28383);
nand U29203 (N_29203,N_27141,N_28097);
and U29204 (N_29204,N_28259,N_27228);
xor U29205 (N_29205,N_28403,N_27339);
xor U29206 (N_29206,N_27400,N_27227);
xnor U29207 (N_29207,N_27767,N_28300);
and U29208 (N_29208,N_27778,N_28238);
nor U29209 (N_29209,N_27240,N_27094);
or U29210 (N_29210,N_27598,N_27746);
and U29211 (N_29211,N_28003,N_27866);
xnor U29212 (N_29212,N_27723,N_28327);
or U29213 (N_29213,N_27322,N_27589);
nand U29214 (N_29214,N_28360,N_27124);
xnor U29215 (N_29215,N_27605,N_28304);
xnor U29216 (N_29216,N_28129,N_27029);
or U29217 (N_29217,N_27862,N_27936);
nand U29218 (N_29218,N_28306,N_27501);
or U29219 (N_29219,N_27514,N_27669);
nor U29220 (N_29220,N_28036,N_28345);
and U29221 (N_29221,N_28136,N_27415);
xor U29222 (N_29222,N_27776,N_28298);
and U29223 (N_29223,N_28155,N_27288);
nand U29224 (N_29224,N_27994,N_27835);
nor U29225 (N_29225,N_27806,N_27151);
or U29226 (N_29226,N_28270,N_27988);
and U29227 (N_29227,N_27017,N_28331);
or U29228 (N_29228,N_27843,N_27266);
xor U29229 (N_29229,N_28159,N_28499);
nor U29230 (N_29230,N_27391,N_27172);
nand U29231 (N_29231,N_27112,N_27983);
xor U29232 (N_29232,N_28132,N_27880);
and U29233 (N_29233,N_27614,N_27676);
nor U29234 (N_29234,N_27408,N_27737);
nor U29235 (N_29235,N_27004,N_27333);
and U29236 (N_29236,N_27183,N_27696);
nand U29237 (N_29237,N_28225,N_27812);
xnor U29238 (N_29238,N_27579,N_28047);
and U29239 (N_29239,N_28231,N_27788);
xnor U29240 (N_29240,N_27923,N_27024);
nand U29241 (N_29241,N_28342,N_27653);
xor U29242 (N_29242,N_28439,N_27399);
nand U29243 (N_29243,N_27855,N_27858);
xnor U29244 (N_29244,N_27407,N_28172);
and U29245 (N_29245,N_27655,N_27854);
or U29246 (N_29246,N_28266,N_27522);
nor U29247 (N_29247,N_28271,N_27417);
xnor U29248 (N_29248,N_27396,N_28380);
nor U29249 (N_29249,N_27600,N_27226);
and U29250 (N_29250,N_28061,N_28334);
nand U29251 (N_29251,N_28288,N_27063);
and U29252 (N_29252,N_28273,N_27451);
nand U29253 (N_29253,N_27265,N_27063);
nand U29254 (N_29254,N_28407,N_27882);
nand U29255 (N_29255,N_27852,N_28297);
and U29256 (N_29256,N_28031,N_27485);
nand U29257 (N_29257,N_27689,N_27011);
nand U29258 (N_29258,N_27781,N_27030);
and U29259 (N_29259,N_28090,N_27907);
xor U29260 (N_29260,N_27030,N_27708);
nor U29261 (N_29261,N_27732,N_27469);
nand U29262 (N_29262,N_28492,N_28303);
xor U29263 (N_29263,N_27495,N_27603);
or U29264 (N_29264,N_27224,N_28118);
nand U29265 (N_29265,N_28107,N_27970);
or U29266 (N_29266,N_28361,N_27986);
and U29267 (N_29267,N_27917,N_28345);
and U29268 (N_29268,N_27720,N_27535);
nor U29269 (N_29269,N_27936,N_28334);
or U29270 (N_29270,N_27826,N_27950);
or U29271 (N_29271,N_28376,N_28409);
nor U29272 (N_29272,N_28215,N_27001);
nor U29273 (N_29273,N_27018,N_28281);
nor U29274 (N_29274,N_28330,N_28277);
or U29275 (N_29275,N_28454,N_28115);
xor U29276 (N_29276,N_27031,N_27035);
xor U29277 (N_29277,N_28077,N_27865);
or U29278 (N_29278,N_27520,N_27172);
or U29279 (N_29279,N_28098,N_27354);
xnor U29280 (N_29280,N_27015,N_27746);
and U29281 (N_29281,N_27910,N_27967);
nand U29282 (N_29282,N_27601,N_28101);
or U29283 (N_29283,N_27821,N_27661);
or U29284 (N_29284,N_28459,N_28456);
xor U29285 (N_29285,N_28001,N_27335);
nor U29286 (N_29286,N_27064,N_27307);
or U29287 (N_29287,N_27784,N_27756);
xnor U29288 (N_29288,N_28314,N_27311);
nor U29289 (N_29289,N_27817,N_27388);
or U29290 (N_29290,N_27494,N_27420);
xor U29291 (N_29291,N_28400,N_27445);
xnor U29292 (N_29292,N_27752,N_27619);
nor U29293 (N_29293,N_27097,N_27765);
and U29294 (N_29294,N_28406,N_27330);
or U29295 (N_29295,N_27982,N_27110);
nor U29296 (N_29296,N_28325,N_27338);
and U29297 (N_29297,N_27510,N_28215);
xnor U29298 (N_29298,N_27261,N_27599);
or U29299 (N_29299,N_27796,N_28120);
or U29300 (N_29300,N_27001,N_27557);
nand U29301 (N_29301,N_27614,N_27127);
xor U29302 (N_29302,N_27961,N_27000);
xor U29303 (N_29303,N_28343,N_28420);
nor U29304 (N_29304,N_27295,N_27695);
nand U29305 (N_29305,N_27755,N_27834);
and U29306 (N_29306,N_27085,N_28248);
nor U29307 (N_29307,N_27716,N_28428);
or U29308 (N_29308,N_27571,N_28444);
nand U29309 (N_29309,N_27980,N_28017);
xnor U29310 (N_29310,N_27704,N_27995);
xor U29311 (N_29311,N_28043,N_27973);
xor U29312 (N_29312,N_27823,N_27653);
or U29313 (N_29313,N_27024,N_28431);
nand U29314 (N_29314,N_28250,N_27875);
xnor U29315 (N_29315,N_27126,N_28410);
and U29316 (N_29316,N_28458,N_27189);
nand U29317 (N_29317,N_28462,N_28197);
and U29318 (N_29318,N_27270,N_28429);
xor U29319 (N_29319,N_28261,N_28277);
nand U29320 (N_29320,N_27071,N_28408);
xor U29321 (N_29321,N_28344,N_27262);
nand U29322 (N_29322,N_27713,N_27441);
nor U29323 (N_29323,N_27865,N_28266);
or U29324 (N_29324,N_27930,N_27717);
xor U29325 (N_29325,N_27085,N_27355);
xnor U29326 (N_29326,N_27884,N_28069);
nor U29327 (N_29327,N_28201,N_27679);
xnor U29328 (N_29328,N_28448,N_27979);
nand U29329 (N_29329,N_28426,N_27591);
nand U29330 (N_29330,N_28184,N_28054);
or U29331 (N_29331,N_28382,N_28390);
nor U29332 (N_29332,N_28477,N_27156);
or U29333 (N_29333,N_27070,N_27688);
nand U29334 (N_29334,N_27184,N_27033);
and U29335 (N_29335,N_28260,N_28244);
nor U29336 (N_29336,N_27724,N_28165);
or U29337 (N_29337,N_27889,N_27314);
xnor U29338 (N_29338,N_27922,N_28344);
or U29339 (N_29339,N_27064,N_27776);
nor U29340 (N_29340,N_27020,N_28214);
xor U29341 (N_29341,N_27224,N_27393);
or U29342 (N_29342,N_28176,N_27616);
nor U29343 (N_29343,N_27880,N_27760);
and U29344 (N_29344,N_27682,N_27075);
and U29345 (N_29345,N_28088,N_27281);
nor U29346 (N_29346,N_28269,N_28328);
nor U29347 (N_29347,N_27825,N_28168);
nand U29348 (N_29348,N_27211,N_27649);
nand U29349 (N_29349,N_27212,N_27391);
and U29350 (N_29350,N_27491,N_27796);
xnor U29351 (N_29351,N_28327,N_27058);
or U29352 (N_29352,N_27994,N_27580);
and U29353 (N_29353,N_27350,N_27988);
nand U29354 (N_29354,N_27781,N_27981);
nor U29355 (N_29355,N_28401,N_27342);
xnor U29356 (N_29356,N_27528,N_28444);
or U29357 (N_29357,N_27981,N_27218);
nor U29358 (N_29358,N_27097,N_27998);
nor U29359 (N_29359,N_28080,N_28273);
nand U29360 (N_29360,N_28366,N_27370);
and U29361 (N_29361,N_27399,N_28237);
or U29362 (N_29362,N_27770,N_27156);
nand U29363 (N_29363,N_28364,N_27873);
nor U29364 (N_29364,N_27930,N_27890);
and U29365 (N_29365,N_27185,N_27808);
nand U29366 (N_29366,N_28070,N_28416);
nor U29367 (N_29367,N_27214,N_27063);
nand U29368 (N_29368,N_27447,N_28301);
xnor U29369 (N_29369,N_27498,N_27054);
or U29370 (N_29370,N_27622,N_27480);
nand U29371 (N_29371,N_28185,N_28440);
and U29372 (N_29372,N_27367,N_27323);
xnor U29373 (N_29373,N_28279,N_27142);
xnor U29374 (N_29374,N_27367,N_28145);
xor U29375 (N_29375,N_27758,N_27807);
nand U29376 (N_29376,N_28490,N_28341);
or U29377 (N_29377,N_28064,N_28433);
nand U29378 (N_29378,N_28363,N_28349);
nor U29379 (N_29379,N_27007,N_27476);
or U29380 (N_29380,N_27382,N_27458);
or U29381 (N_29381,N_27416,N_28124);
xor U29382 (N_29382,N_27879,N_28446);
and U29383 (N_29383,N_28118,N_27631);
xnor U29384 (N_29384,N_27898,N_27706);
nand U29385 (N_29385,N_28268,N_27098);
or U29386 (N_29386,N_27213,N_27623);
nand U29387 (N_29387,N_28264,N_27116);
xor U29388 (N_29388,N_28184,N_27231);
nor U29389 (N_29389,N_27958,N_27995);
nand U29390 (N_29390,N_27646,N_27616);
xor U29391 (N_29391,N_27596,N_27058);
or U29392 (N_29392,N_27137,N_27174);
nand U29393 (N_29393,N_27825,N_27242);
nand U29394 (N_29394,N_27762,N_27097);
nor U29395 (N_29395,N_27371,N_27649);
and U29396 (N_29396,N_28452,N_27894);
nor U29397 (N_29397,N_27626,N_27963);
nand U29398 (N_29398,N_27480,N_27259);
xor U29399 (N_29399,N_27863,N_28104);
or U29400 (N_29400,N_27289,N_28132);
xnor U29401 (N_29401,N_27532,N_27245);
or U29402 (N_29402,N_28371,N_28184);
or U29403 (N_29403,N_27554,N_28256);
and U29404 (N_29404,N_27463,N_28117);
xnor U29405 (N_29405,N_27337,N_27847);
or U29406 (N_29406,N_27236,N_27536);
or U29407 (N_29407,N_28186,N_27766);
and U29408 (N_29408,N_27373,N_27177);
nor U29409 (N_29409,N_27365,N_27443);
and U29410 (N_29410,N_28170,N_27312);
xnor U29411 (N_29411,N_27256,N_27545);
xnor U29412 (N_29412,N_27395,N_28307);
xor U29413 (N_29413,N_27833,N_28070);
or U29414 (N_29414,N_27443,N_28118);
or U29415 (N_29415,N_27643,N_27042);
or U29416 (N_29416,N_27193,N_28117);
or U29417 (N_29417,N_27354,N_27746);
xnor U29418 (N_29418,N_28211,N_28410);
nand U29419 (N_29419,N_28209,N_28404);
or U29420 (N_29420,N_27522,N_28400);
xor U29421 (N_29421,N_27233,N_27452);
nand U29422 (N_29422,N_27855,N_27497);
xnor U29423 (N_29423,N_27418,N_28292);
xnor U29424 (N_29424,N_28108,N_28481);
or U29425 (N_29425,N_27884,N_28473);
and U29426 (N_29426,N_27477,N_27357);
nor U29427 (N_29427,N_27686,N_27962);
nor U29428 (N_29428,N_27427,N_27995);
nand U29429 (N_29429,N_28194,N_27576);
nand U29430 (N_29430,N_27953,N_28098);
and U29431 (N_29431,N_27337,N_27802);
nor U29432 (N_29432,N_28388,N_27541);
and U29433 (N_29433,N_27329,N_27125);
and U29434 (N_29434,N_28453,N_27140);
nand U29435 (N_29435,N_27624,N_28430);
nand U29436 (N_29436,N_27072,N_27279);
nor U29437 (N_29437,N_27185,N_28143);
or U29438 (N_29438,N_27417,N_27168);
nor U29439 (N_29439,N_27832,N_28375);
xor U29440 (N_29440,N_27334,N_27074);
or U29441 (N_29441,N_27385,N_27343);
xnor U29442 (N_29442,N_27823,N_27537);
nor U29443 (N_29443,N_27637,N_27853);
or U29444 (N_29444,N_27124,N_28039);
nand U29445 (N_29445,N_28063,N_28475);
nand U29446 (N_29446,N_28323,N_27813);
nand U29447 (N_29447,N_27266,N_27709);
nor U29448 (N_29448,N_27285,N_27473);
and U29449 (N_29449,N_27158,N_27773);
and U29450 (N_29450,N_27729,N_27097);
or U29451 (N_29451,N_28268,N_27045);
nor U29452 (N_29452,N_27697,N_28057);
and U29453 (N_29453,N_28352,N_28163);
nor U29454 (N_29454,N_27119,N_28292);
nand U29455 (N_29455,N_27080,N_27593);
or U29456 (N_29456,N_27334,N_28045);
nand U29457 (N_29457,N_27281,N_27269);
or U29458 (N_29458,N_28332,N_27755);
xnor U29459 (N_29459,N_27274,N_27955);
or U29460 (N_29460,N_27603,N_28143);
nor U29461 (N_29461,N_27240,N_28278);
xnor U29462 (N_29462,N_27192,N_28012);
or U29463 (N_29463,N_27624,N_27077);
nand U29464 (N_29464,N_27204,N_27928);
nor U29465 (N_29465,N_27343,N_27493);
and U29466 (N_29466,N_28108,N_27563);
nand U29467 (N_29467,N_28318,N_28368);
nor U29468 (N_29468,N_27283,N_27907);
xor U29469 (N_29469,N_27580,N_28451);
or U29470 (N_29470,N_27749,N_27488);
nor U29471 (N_29471,N_27395,N_28144);
nand U29472 (N_29472,N_27391,N_27575);
and U29473 (N_29473,N_28138,N_27862);
and U29474 (N_29474,N_27990,N_28191);
nand U29475 (N_29475,N_27076,N_28436);
or U29476 (N_29476,N_27445,N_27226);
or U29477 (N_29477,N_28453,N_27585);
nand U29478 (N_29478,N_27539,N_28069);
and U29479 (N_29479,N_28199,N_28315);
nand U29480 (N_29480,N_28009,N_28196);
or U29481 (N_29481,N_27272,N_27164);
and U29482 (N_29482,N_28034,N_27627);
and U29483 (N_29483,N_28450,N_28137);
or U29484 (N_29484,N_27067,N_28183);
and U29485 (N_29485,N_28477,N_27052);
nand U29486 (N_29486,N_27014,N_27985);
nand U29487 (N_29487,N_27191,N_27435);
nand U29488 (N_29488,N_27028,N_28257);
or U29489 (N_29489,N_27711,N_28048);
xor U29490 (N_29490,N_27717,N_27875);
nor U29491 (N_29491,N_27274,N_28412);
nand U29492 (N_29492,N_27049,N_27352);
or U29493 (N_29493,N_27165,N_28367);
xor U29494 (N_29494,N_27176,N_27799);
and U29495 (N_29495,N_27757,N_28392);
xnor U29496 (N_29496,N_28489,N_28416);
xnor U29497 (N_29497,N_27778,N_27067);
xnor U29498 (N_29498,N_27177,N_27735);
or U29499 (N_29499,N_28488,N_27779);
nand U29500 (N_29500,N_28499,N_27409);
and U29501 (N_29501,N_27296,N_28190);
or U29502 (N_29502,N_28360,N_27610);
nand U29503 (N_29503,N_28280,N_27116);
or U29504 (N_29504,N_27952,N_28004);
or U29505 (N_29505,N_27960,N_27900);
and U29506 (N_29506,N_27918,N_28459);
and U29507 (N_29507,N_28271,N_27201);
and U29508 (N_29508,N_27673,N_27529);
or U29509 (N_29509,N_27489,N_28165);
nor U29510 (N_29510,N_27198,N_28132);
xor U29511 (N_29511,N_28423,N_27531);
and U29512 (N_29512,N_28015,N_27267);
and U29513 (N_29513,N_27513,N_28290);
xnor U29514 (N_29514,N_27254,N_28099);
and U29515 (N_29515,N_27880,N_27081);
or U29516 (N_29516,N_27957,N_27725);
nor U29517 (N_29517,N_27227,N_27497);
nor U29518 (N_29518,N_27692,N_27393);
xor U29519 (N_29519,N_27179,N_27743);
xor U29520 (N_29520,N_27491,N_27436);
or U29521 (N_29521,N_27645,N_27108);
nor U29522 (N_29522,N_27762,N_27337);
and U29523 (N_29523,N_28048,N_27337);
and U29524 (N_29524,N_27460,N_27433);
nand U29525 (N_29525,N_27946,N_27577);
xnor U29526 (N_29526,N_28231,N_27322);
or U29527 (N_29527,N_28033,N_27512);
or U29528 (N_29528,N_27303,N_28124);
xnor U29529 (N_29529,N_28438,N_27000);
and U29530 (N_29530,N_28172,N_27418);
nor U29531 (N_29531,N_27671,N_27756);
or U29532 (N_29532,N_27801,N_27472);
nor U29533 (N_29533,N_27577,N_27045);
and U29534 (N_29534,N_27964,N_27991);
and U29535 (N_29535,N_27839,N_27292);
and U29536 (N_29536,N_28003,N_27232);
nor U29537 (N_29537,N_27791,N_27494);
nand U29538 (N_29538,N_27104,N_27858);
xnor U29539 (N_29539,N_27598,N_27675);
or U29540 (N_29540,N_27432,N_27626);
nand U29541 (N_29541,N_27666,N_28065);
or U29542 (N_29542,N_28006,N_27430);
nand U29543 (N_29543,N_27467,N_28269);
nor U29544 (N_29544,N_27577,N_27118);
nand U29545 (N_29545,N_27800,N_27556);
or U29546 (N_29546,N_27371,N_28222);
nor U29547 (N_29547,N_27962,N_27018);
xor U29548 (N_29548,N_28283,N_27811);
nor U29549 (N_29549,N_28190,N_27136);
nor U29550 (N_29550,N_27928,N_27569);
nand U29551 (N_29551,N_27157,N_27797);
xor U29552 (N_29552,N_27162,N_27806);
or U29553 (N_29553,N_28364,N_27856);
nand U29554 (N_29554,N_27694,N_27032);
or U29555 (N_29555,N_27841,N_28207);
nor U29556 (N_29556,N_27813,N_28076);
and U29557 (N_29557,N_27910,N_27345);
or U29558 (N_29558,N_28192,N_27006);
nand U29559 (N_29559,N_27063,N_27142);
nand U29560 (N_29560,N_28271,N_27600);
or U29561 (N_29561,N_28127,N_27430);
nand U29562 (N_29562,N_27481,N_27573);
nor U29563 (N_29563,N_27759,N_28059);
or U29564 (N_29564,N_27202,N_28446);
nor U29565 (N_29565,N_27253,N_28345);
nand U29566 (N_29566,N_28048,N_27178);
nor U29567 (N_29567,N_28011,N_27364);
nand U29568 (N_29568,N_27853,N_27968);
or U29569 (N_29569,N_27978,N_28321);
nand U29570 (N_29570,N_27686,N_27483);
nor U29571 (N_29571,N_27392,N_28236);
nor U29572 (N_29572,N_27908,N_27850);
nor U29573 (N_29573,N_27486,N_27758);
xor U29574 (N_29574,N_27739,N_27256);
nor U29575 (N_29575,N_27905,N_28118);
and U29576 (N_29576,N_27011,N_28315);
and U29577 (N_29577,N_27011,N_28082);
xnor U29578 (N_29578,N_27565,N_27128);
nor U29579 (N_29579,N_27878,N_27857);
xor U29580 (N_29580,N_27943,N_28407);
nand U29581 (N_29581,N_27568,N_28009);
nor U29582 (N_29582,N_27849,N_28103);
and U29583 (N_29583,N_28388,N_28411);
and U29584 (N_29584,N_28275,N_27038);
xor U29585 (N_29585,N_27024,N_27364);
nand U29586 (N_29586,N_28105,N_28015);
nor U29587 (N_29587,N_27998,N_27007);
or U29588 (N_29588,N_28423,N_27919);
or U29589 (N_29589,N_27621,N_27854);
nor U29590 (N_29590,N_27946,N_28359);
or U29591 (N_29591,N_27445,N_27095);
or U29592 (N_29592,N_28440,N_27126);
nor U29593 (N_29593,N_27124,N_27150);
or U29594 (N_29594,N_28195,N_27197);
nand U29595 (N_29595,N_27158,N_27426);
nand U29596 (N_29596,N_27179,N_27574);
nor U29597 (N_29597,N_27915,N_27026);
nor U29598 (N_29598,N_27886,N_27561);
and U29599 (N_29599,N_27864,N_27163);
and U29600 (N_29600,N_27619,N_27775);
nor U29601 (N_29601,N_27737,N_28252);
xor U29602 (N_29602,N_27529,N_27429);
or U29603 (N_29603,N_28116,N_28473);
xnor U29604 (N_29604,N_28210,N_28345);
nor U29605 (N_29605,N_27686,N_27582);
and U29606 (N_29606,N_27946,N_28029);
nor U29607 (N_29607,N_27739,N_28372);
nand U29608 (N_29608,N_27478,N_28290);
nand U29609 (N_29609,N_27274,N_27612);
and U29610 (N_29610,N_27150,N_27873);
and U29611 (N_29611,N_27068,N_27028);
or U29612 (N_29612,N_27715,N_27314);
nand U29613 (N_29613,N_28210,N_27312);
or U29614 (N_29614,N_28334,N_27360);
nor U29615 (N_29615,N_28315,N_27678);
nor U29616 (N_29616,N_27157,N_27997);
and U29617 (N_29617,N_27664,N_27118);
xor U29618 (N_29618,N_28039,N_28112);
nor U29619 (N_29619,N_27511,N_27862);
and U29620 (N_29620,N_27621,N_27850);
xnor U29621 (N_29621,N_27834,N_28336);
and U29622 (N_29622,N_27061,N_27181);
nor U29623 (N_29623,N_27918,N_28210);
xnor U29624 (N_29624,N_28355,N_27861);
nor U29625 (N_29625,N_28476,N_27781);
nand U29626 (N_29626,N_27231,N_27045);
xor U29627 (N_29627,N_28116,N_27331);
or U29628 (N_29628,N_27989,N_27382);
nor U29629 (N_29629,N_27884,N_27997);
nand U29630 (N_29630,N_27452,N_28001);
nand U29631 (N_29631,N_28104,N_28359);
nand U29632 (N_29632,N_28062,N_27327);
nand U29633 (N_29633,N_27936,N_28295);
or U29634 (N_29634,N_27785,N_27371);
xor U29635 (N_29635,N_27316,N_28398);
and U29636 (N_29636,N_27389,N_27553);
xnor U29637 (N_29637,N_27702,N_28194);
xnor U29638 (N_29638,N_27109,N_27404);
nand U29639 (N_29639,N_27578,N_27161);
or U29640 (N_29640,N_27937,N_28497);
nor U29641 (N_29641,N_28030,N_27018);
nand U29642 (N_29642,N_27332,N_27649);
or U29643 (N_29643,N_27275,N_27486);
nor U29644 (N_29644,N_27237,N_27836);
nor U29645 (N_29645,N_28332,N_28311);
and U29646 (N_29646,N_28095,N_27158);
or U29647 (N_29647,N_27456,N_27546);
or U29648 (N_29648,N_28483,N_27239);
xnor U29649 (N_29649,N_28223,N_28228);
nor U29650 (N_29650,N_27390,N_28048);
or U29651 (N_29651,N_27168,N_27933);
and U29652 (N_29652,N_27352,N_27463);
xnor U29653 (N_29653,N_28094,N_27302);
nor U29654 (N_29654,N_27433,N_27888);
or U29655 (N_29655,N_27426,N_27723);
nand U29656 (N_29656,N_28201,N_27952);
xor U29657 (N_29657,N_28350,N_28143);
or U29658 (N_29658,N_28078,N_27946);
xor U29659 (N_29659,N_27070,N_28300);
or U29660 (N_29660,N_28036,N_27420);
nand U29661 (N_29661,N_27926,N_28044);
nand U29662 (N_29662,N_28133,N_27396);
nand U29663 (N_29663,N_27964,N_27487);
and U29664 (N_29664,N_28288,N_28323);
nor U29665 (N_29665,N_27281,N_28269);
and U29666 (N_29666,N_27034,N_27428);
or U29667 (N_29667,N_27367,N_27465);
nand U29668 (N_29668,N_27902,N_27230);
nand U29669 (N_29669,N_27303,N_27801);
or U29670 (N_29670,N_27692,N_27610);
or U29671 (N_29671,N_27197,N_27415);
and U29672 (N_29672,N_28035,N_27597);
or U29673 (N_29673,N_27591,N_28444);
or U29674 (N_29674,N_27436,N_27986);
xor U29675 (N_29675,N_28059,N_27923);
and U29676 (N_29676,N_27728,N_27505);
nand U29677 (N_29677,N_27026,N_27179);
nand U29678 (N_29678,N_27175,N_27939);
nor U29679 (N_29679,N_28146,N_28341);
nor U29680 (N_29680,N_28144,N_27575);
nand U29681 (N_29681,N_27890,N_27728);
nand U29682 (N_29682,N_27637,N_27141);
nor U29683 (N_29683,N_28139,N_27853);
nor U29684 (N_29684,N_27255,N_28012);
and U29685 (N_29685,N_28067,N_28149);
or U29686 (N_29686,N_28140,N_28453);
or U29687 (N_29687,N_28483,N_28463);
nand U29688 (N_29688,N_28343,N_27892);
xor U29689 (N_29689,N_28438,N_28139);
nand U29690 (N_29690,N_27076,N_27778);
xor U29691 (N_29691,N_27784,N_27158);
or U29692 (N_29692,N_28229,N_28238);
and U29693 (N_29693,N_27498,N_27553);
and U29694 (N_29694,N_27857,N_28190);
and U29695 (N_29695,N_27341,N_27270);
and U29696 (N_29696,N_27674,N_27967);
nor U29697 (N_29697,N_27511,N_27092);
and U29698 (N_29698,N_27127,N_28306);
and U29699 (N_29699,N_28374,N_28359);
and U29700 (N_29700,N_28134,N_27062);
or U29701 (N_29701,N_28281,N_27453);
xnor U29702 (N_29702,N_27433,N_27894);
or U29703 (N_29703,N_27800,N_27660);
nor U29704 (N_29704,N_27304,N_27865);
and U29705 (N_29705,N_27410,N_27816);
nor U29706 (N_29706,N_27895,N_27005);
or U29707 (N_29707,N_27192,N_27932);
xnor U29708 (N_29708,N_27274,N_27835);
and U29709 (N_29709,N_27181,N_27542);
nand U29710 (N_29710,N_28086,N_28120);
or U29711 (N_29711,N_28473,N_27702);
nand U29712 (N_29712,N_27027,N_28210);
or U29713 (N_29713,N_27984,N_28292);
nand U29714 (N_29714,N_28057,N_28097);
nand U29715 (N_29715,N_27420,N_27715);
or U29716 (N_29716,N_27599,N_28302);
xnor U29717 (N_29717,N_27561,N_28322);
xnor U29718 (N_29718,N_28373,N_27319);
and U29719 (N_29719,N_28352,N_28202);
nand U29720 (N_29720,N_27744,N_28115);
nor U29721 (N_29721,N_27667,N_27586);
nor U29722 (N_29722,N_28314,N_27641);
nand U29723 (N_29723,N_27545,N_27715);
and U29724 (N_29724,N_28320,N_27355);
xor U29725 (N_29725,N_27151,N_28057);
xor U29726 (N_29726,N_27760,N_27448);
or U29727 (N_29727,N_28266,N_28478);
nand U29728 (N_29728,N_28393,N_27513);
nor U29729 (N_29729,N_28389,N_28081);
and U29730 (N_29730,N_27026,N_27266);
and U29731 (N_29731,N_27280,N_28158);
xnor U29732 (N_29732,N_27291,N_27253);
xor U29733 (N_29733,N_27269,N_28390);
and U29734 (N_29734,N_27714,N_27754);
or U29735 (N_29735,N_27168,N_27772);
nor U29736 (N_29736,N_27864,N_27952);
nor U29737 (N_29737,N_27573,N_27461);
and U29738 (N_29738,N_27843,N_27326);
xnor U29739 (N_29739,N_27932,N_27404);
or U29740 (N_29740,N_27459,N_27227);
or U29741 (N_29741,N_27290,N_27931);
or U29742 (N_29742,N_27967,N_27112);
xnor U29743 (N_29743,N_27864,N_27336);
and U29744 (N_29744,N_27428,N_27736);
and U29745 (N_29745,N_27016,N_27716);
xor U29746 (N_29746,N_27492,N_28267);
or U29747 (N_29747,N_27023,N_27601);
and U29748 (N_29748,N_28352,N_27278);
nor U29749 (N_29749,N_27214,N_27293);
or U29750 (N_29750,N_27533,N_27481);
xor U29751 (N_29751,N_27736,N_27782);
nor U29752 (N_29752,N_27950,N_28287);
xnor U29753 (N_29753,N_28413,N_27011);
nand U29754 (N_29754,N_27539,N_28451);
nand U29755 (N_29755,N_27936,N_27204);
nand U29756 (N_29756,N_28436,N_27424);
nand U29757 (N_29757,N_27092,N_27220);
xor U29758 (N_29758,N_28452,N_27658);
xnor U29759 (N_29759,N_27454,N_27309);
xnor U29760 (N_29760,N_27219,N_27342);
or U29761 (N_29761,N_27166,N_27731);
or U29762 (N_29762,N_27044,N_27349);
xor U29763 (N_29763,N_28160,N_28236);
and U29764 (N_29764,N_28354,N_28438);
or U29765 (N_29765,N_27382,N_28059);
nand U29766 (N_29766,N_28074,N_27989);
xor U29767 (N_29767,N_28385,N_27094);
xor U29768 (N_29768,N_28225,N_27145);
nand U29769 (N_29769,N_27297,N_27542);
or U29770 (N_29770,N_27297,N_27706);
nand U29771 (N_29771,N_28231,N_27542);
and U29772 (N_29772,N_27040,N_27246);
nand U29773 (N_29773,N_27041,N_27032);
nand U29774 (N_29774,N_27937,N_28380);
nor U29775 (N_29775,N_27413,N_27099);
nand U29776 (N_29776,N_27520,N_27903);
nor U29777 (N_29777,N_27545,N_27090);
nor U29778 (N_29778,N_27979,N_27428);
xor U29779 (N_29779,N_28337,N_27286);
xor U29780 (N_29780,N_27803,N_27449);
or U29781 (N_29781,N_27855,N_28008);
and U29782 (N_29782,N_27839,N_27345);
xor U29783 (N_29783,N_27304,N_27347);
xnor U29784 (N_29784,N_27192,N_27586);
or U29785 (N_29785,N_27089,N_27591);
or U29786 (N_29786,N_27050,N_28219);
nand U29787 (N_29787,N_27329,N_28258);
and U29788 (N_29788,N_27352,N_28147);
nand U29789 (N_29789,N_27382,N_27042);
nor U29790 (N_29790,N_28224,N_28211);
xor U29791 (N_29791,N_28139,N_27500);
xnor U29792 (N_29792,N_27186,N_27425);
and U29793 (N_29793,N_27350,N_27345);
nor U29794 (N_29794,N_27553,N_27155);
nand U29795 (N_29795,N_27352,N_27969);
nor U29796 (N_29796,N_28456,N_27095);
nor U29797 (N_29797,N_27080,N_27463);
nor U29798 (N_29798,N_27059,N_27347);
nand U29799 (N_29799,N_27307,N_27833);
and U29800 (N_29800,N_28420,N_28327);
xor U29801 (N_29801,N_27645,N_27750);
or U29802 (N_29802,N_27532,N_27266);
xor U29803 (N_29803,N_27139,N_27004);
and U29804 (N_29804,N_27199,N_27417);
xnor U29805 (N_29805,N_28138,N_27982);
nand U29806 (N_29806,N_27621,N_27702);
and U29807 (N_29807,N_27868,N_27828);
and U29808 (N_29808,N_27576,N_27739);
and U29809 (N_29809,N_27924,N_28084);
xnor U29810 (N_29810,N_27056,N_27297);
nand U29811 (N_29811,N_27777,N_28202);
and U29812 (N_29812,N_28441,N_27189);
nor U29813 (N_29813,N_28490,N_27779);
nor U29814 (N_29814,N_27508,N_28100);
or U29815 (N_29815,N_27063,N_27131);
or U29816 (N_29816,N_28215,N_27416);
and U29817 (N_29817,N_27263,N_27991);
xor U29818 (N_29818,N_27621,N_27469);
nor U29819 (N_29819,N_27822,N_27762);
xor U29820 (N_29820,N_28024,N_27739);
xnor U29821 (N_29821,N_27521,N_27320);
nor U29822 (N_29822,N_28072,N_27647);
nand U29823 (N_29823,N_27014,N_28005);
or U29824 (N_29824,N_27993,N_27522);
or U29825 (N_29825,N_27075,N_27691);
nand U29826 (N_29826,N_27948,N_27578);
nand U29827 (N_29827,N_28406,N_27134);
xnor U29828 (N_29828,N_27644,N_28066);
xor U29829 (N_29829,N_27927,N_27994);
nor U29830 (N_29830,N_27292,N_27459);
nor U29831 (N_29831,N_27025,N_27011);
or U29832 (N_29832,N_28283,N_28208);
or U29833 (N_29833,N_28136,N_28224);
nor U29834 (N_29834,N_27869,N_27922);
nor U29835 (N_29835,N_27449,N_27274);
nor U29836 (N_29836,N_27481,N_27360);
and U29837 (N_29837,N_27037,N_27862);
and U29838 (N_29838,N_27880,N_27277);
or U29839 (N_29839,N_28358,N_27581);
or U29840 (N_29840,N_28470,N_27493);
and U29841 (N_29841,N_27026,N_27292);
or U29842 (N_29842,N_27984,N_27837);
and U29843 (N_29843,N_27725,N_27422);
xor U29844 (N_29844,N_28037,N_27776);
and U29845 (N_29845,N_28405,N_28234);
and U29846 (N_29846,N_27836,N_28182);
nor U29847 (N_29847,N_27735,N_27844);
or U29848 (N_29848,N_27057,N_27626);
nand U29849 (N_29849,N_27470,N_27167);
xnor U29850 (N_29850,N_27481,N_27256);
nor U29851 (N_29851,N_28222,N_27140);
nor U29852 (N_29852,N_28177,N_27029);
and U29853 (N_29853,N_27330,N_28459);
and U29854 (N_29854,N_27295,N_27265);
xnor U29855 (N_29855,N_28031,N_27828);
nand U29856 (N_29856,N_27771,N_28027);
and U29857 (N_29857,N_27497,N_27604);
or U29858 (N_29858,N_27479,N_27940);
nand U29859 (N_29859,N_27780,N_27612);
nand U29860 (N_29860,N_27377,N_27797);
xnor U29861 (N_29861,N_27179,N_27116);
nor U29862 (N_29862,N_27545,N_28339);
and U29863 (N_29863,N_27924,N_28282);
and U29864 (N_29864,N_27750,N_27589);
xor U29865 (N_29865,N_27797,N_27633);
nand U29866 (N_29866,N_27922,N_27875);
xor U29867 (N_29867,N_27031,N_28125);
or U29868 (N_29868,N_28054,N_28151);
nand U29869 (N_29869,N_28287,N_28498);
xnor U29870 (N_29870,N_27309,N_28219);
or U29871 (N_29871,N_27222,N_28329);
xnor U29872 (N_29872,N_27442,N_28258);
and U29873 (N_29873,N_27977,N_28190);
nor U29874 (N_29874,N_27404,N_27118);
and U29875 (N_29875,N_28381,N_28314);
xnor U29876 (N_29876,N_27763,N_28163);
nand U29877 (N_29877,N_27933,N_27348);
nand U29878 (N_29878,N_27809,N_28177);
or U29879 (N_29879,N_27374,N_27296);
xor U29880 (N_29880,N_27495,N_27065);
xnor U29881 (N_29881,N_27882,N_27521);
nand U29882 (N_29882,N_27975,N_27428);
or U29883 (N_29883,N_27774,N_27088);
xor U29884 (N_29884,N_27738,N_27411);
xor U29885 (N_29885,N_28323,N_27633);
or U29886 (N_29886,N_27708,N_27753);
xnor U29887 (N_29887,N_27084,N_28168);
and U29888 (N_29888,N_28347,N_28416);
and U29889 (N_29889,N_27175,N_27023);
nor U29890 (N_29890,N_28070,N_27973);
nand U29891 (N_29891,N_27819,N_28483);
or U29892 (N_29892,N_27821,N_27381);
xnor U29893 (N_29893,N_28319,N_27279);
nor U29894 (N_29894,N_27655,N_27594);
nand U29895 (N_29895,N_27273,N_27878);
or U29896 (N_29896,N_28337,N_27926);
nor U29897 (N_29897,N_27106,N_27664);
nand U29898 (N_29898,N_27290,N_27802);
or U29899 (N_29899,N_27693,N_27478);
xor U29900 (N_29900,N_27631,N_27338);
and U29901 (N_29901,N_27646,N_27057);
nor U29902 (N_29902,N_27104,N_27057);
nand U29903 (N_29903,N_28225,N_27300);
nand U29904 (N_29904,N_27566,N_27363);
nor U29905 (N_29905,N_27362,N_27097);
nand U29906 (N_29906,N_27807,N_28460);
or U29907 (N_29907,N_27903,N_27154);
xor U29908 (N_29908,N_28011,N_27015);
or U29909 (N_29909,N_28256,N_27105);
xor U29910 (N_29910,N_27953,N_28411);
nand U29911 (N_29911,N_27838,N_28109);
and U29912 (N_29912,N_28122,N_28217);
and U29913 (N_29913,N_27217,N_27380);
or U29914 (N_29914,N_28212,N_28167);
nor U29915 (N_29915,N_28391,N_28487);
and U29916 (N_29916,N_27079,N_27740);
nand U29917 (N_29917,N_28046,N_27923);
nor U29918 (N_29918,N_27319,N_28367);
and U29919 (N_29919,N_27970,N_27052);
or U29920 (N_29920,N_27125,N_27609);
nand U29921 (N_29921,N_27813,N_27956);
nor U29922 (N_29922,N_27595,N_27687);
nand U29923 (N_29923,N_27601,N_27452);
nand U29924 (N_29924,N_27806,N_28344);
xnor U29925 (N_29925,N_27859,N_28045);
and U29926 (N_29926,N_27135,N_28108);
or U29927 (N_29927,N_28033,N_28111);
and U29928 (N_29928,N_27386,N_27303);
and U29929 (N_29929,N_27728,N_28066);
nor U29930 (N_29930,N_27333,N_27960);
and U29931 (N_29931,N_28278,N_28285);
or U29932 (N_29932,N_27051,N_28244);
or U29933 (N_29933,N_27013,N_28207);
xor U29934 (N_29934,N_27694,N_27253);
nor U29935 (N_29935,N_27045,N_27507);
nand U29936 (N_29936,N_28204,N_27679);
nor U29937 (N_29937,N_27349,N_28354);
or U29938 (N_29938,N_28462,N_28426);
nand U29939 (N_29939,N_27557,N_27062);
nand U29940 (N_29940,N_27815,N_27358);
xor U29941 (N_29941,N_27851,N_27352);
and U29942 (N_29942,N_27337,N_27694);
or U29943 (N_29943,N_27056,N_27337);
nand U29944 (N_29944,N_27555,N_27262);
nor U29945 (N_29945,N_27685,N_27506);
nand U29946 (N_29946,N_27143,N_28018);
nand U29947 (N_29947,N_27051,N_28400);
xor U29948 (N_29948,N_28213,N_27919);
and U29949 (N_29949,N_28177,N_27519);
nor U29950 (N_29950,N_27177,N_28172);
xnor U29951 (N_29951,N_28414,N_27994);
and U29952 (N_29952,N_28124,N_27319);
nor U29953 (N_29953,N_27701,N_27932);
xor U29954 (N_29954,N_27633,N_27985);
nor U29955 (N_29955,N_27021,N_27566);
nand U29956 (N_29956,N_27766,N_28220);
nand U29957 (N_29957,N_27809,N_27579);
and U29958 (N_29958,N_28307,N_27198);
and U29959 (N_29959,N_28019,N_27588);
nand U29960 (N_29960,N_27640,N_28285);
and U29961 (N_29961,N_27082,N_28365);
nand U29962 (N_29962,N_28319,N_27040);
xor U29963 (N_29963,N_27668,N_27814);
and U29964 (N_29964,N_27805,N_28439);
and U29965 (N_29965,N_28363,N_27497);
nor U29966 (N_29966,N_27876,N_28353);
and U29967 (N_29967,N_27185,N_27937);
and U29968 (N_29968,N_28345,N_27894);
and U29969 (N_29969,N_27211,N_28275);
xnor U29970 (N_29970,N_27198,N_27337);
nand U29971 (N_29971,N_28045,N_27263);
xor U29972 (N_29972,N_27109,N_27816);
nand U29973 (N_29973,N_28000,N_27753);
nand U29974 (N_29974,N_27824,N_27129);
nor U29975 (N_29975,N_28284,N_27327);
xor U29976 (N_29976,N_27204,N_27138);
nand U29977 (N_29977,N_28385,N_27335);
nor U29978 (N_29978,N_28188,N_28006);
or U29979 (N_29979,N_27406,N_27424);
and U29980 (N_29980,N_27763,N_27292);
xor U29981 (N_29981,N_27385,N_27708);
nand U29982 (N_29982,N_27822,N_27494);
and U29983 (N_29983,N_27763,N_28419);
and U29984 (N_29984,N_28425,N_27665);
or U29985 (N_29985,N_27322,N_27320);
nor U29986 (N_29986,N_27090,N_27982);
nor U29987 (N_29987,N_27445,N_27350);
xor U29988 (N_29988,N_27366,N_27468);
nor U29989 (N_29989,N_27513,N_27085);
and U29990 (N_29990,N_28142,N_28478);
or U29991 (N_29991,N_27920,N_28279);
nand U29992 (N_29992,N_27702,N_27027);
xor U29993 (N_29993,N_27698,N_27024);
nand U29994 (N_29994,N_27247,N_28242);
nand U29995 (N_29995,N_28276,N_27641);
and U29996 (N_29996,N_28417,N_27529);
and U29997 (N_29997,N_27832,N_27903);
and U29998 (N_29998,N_28263,N_28449);
and U29999 (N_29999,N_28492,N_27270);
nor UO_0 (O_0,N_29220,N_29433);
nor UO_1 (O_1,N_28591,N_29556);
xnor UO_2 (O_2,N_29628,N_29047);
or UO_3 (O_3,N_28540,N_29744);
or UO_4 (O_4,N_29666,N_28626);
nand UO_5 (O_5,N_29037,N_29261);
and UO_6 (O_6,N_29411,N_29956);
nor UO_7 (O_7,N_29819,N_28682);
xnor UO_8 (O_8,N_29729,N_28895);
nor UO_9 (O_9,N_29098,N_29310);
nand UO_10 (O_10,N_28872,N_29686);
nand UO_11 (O_11,N_28772,N_29318);
nor UO_12 (O_12,N_29592,N_29152);
nor UO_13 (O_13,N_29947,N_29428);
or UO_14 (O_14,N_28880,N_29174);
xnor UO_15 (O_15,N_29466,N_29732);
and UO_16 (O_16,N_28551,N_28806);
and UO_17 (O_17,N_29724,N_29972);
nor UO_18 (O_18,N_29312,N_29386);
and UO_19 (O_19,N_28810,N_28592);
nor UO_20 (O_20,N_29024,N_29429);
xnor UO_21 (O_21,N_29752,N_29055);
xor UO_22 (O_22,N_29532,N_29927);
nor UO_23 (O_23,N_28614,N_28501);
or UO_24 (O_24,N_28522,N_29427);
xnor UO_25 (O_25,N_29909,N_29269);
and UO_26 (O_26,N_29562,N_29499);
nor UO_27 (O_27,N_29706,N_29151);
nand UO_28 (O_28,N_29767,N_29528);
or UO_29 (O_29,N_29383,N_29449);
nand UO_30 (O_30,N_28555,N_28726);
or UO_31 (O_31,N_29825,N_29863);
and UO_32 (O_32,N_29406,N_28918);
nor UO_33 (O_33,N_28815,N_29604);
and UO_34 (O_34,N_29622,N_29665);
nand UO_35 (O_35,N_29064,N_29038);
and UO_36 (O_36,N_28889,N_28640);
nor UO_37 (O_37,N_28808,N_29831);
nor UO_38 (O_38,N_28990,N_28693);
and UO_39 (O_39,N_28803,N_29274);
nand UO_40 (O_40,N_28809,N_28517);
xor UO_41 (O_41,N_29679,N_29451);
xor UO_42 (O_42,N_29390,N_28790);
nand UO_43 (O_43,N_29086,N_29896);
or UO_44 (O_44,N_29516,N_29177);
and UO_45 (O_45,N_28960,N_29892);
and UO_46 (O_46,N_29273,N_29755);
xor UO_47 (O_47,N_29631,N_29072);
or UO_48 (O_48,N_29566,N_29176);
or UO_49 (O_49,N_28535,N_28929);
or UO_50 (O_50,N_29534,N_29304);
xnor UO_51 (O_51,N_29696,N_29568);
nand UO_52 (O_52,N_28845,N_29749);
nor UO_53 (O_53,N_29469,N_29789);
and UO_54 (O_54,N_29053,N_28792);
or UO_55 (O_55,N_29302,N_29475);
or UO_56 (O_56,N_29702,N_29114);
or UO_57 (O_57,N_29019,N_28746);
xor UO_58 (O_58,N_29860,N_28589);
and UO_59 (O_59,N_28745,N_29366);
and UO_60 (O_60,N_29093,N_28516);
and UO_61 (O_61,N_28839,N_28694);
or UO_62 (O_62,N_28903,N_28852);
or UO_63 (O_63,N_29125,N_29751);
nand UO_64 (O_64,N_28628,N_29911);
and UO_65 (O_65,N_28964,N_29605);
xor UO_66 (O_66,N_29746,N_29058);
nand UO_67 (O_67,N_29349,N_29658);
nand UO_68 (O_68,N_29317,N_28921);
and UO_69 (O_69,N_29106,N_29527);
or UO_70 (O_70,N_28877,N_29398);
or UO_71 (O_71,N_29472,N_29889);
and UO_72 (O_72,N_28734,N_28612);
or UO_73 (O_73,N_28527,N_29336);
xor UO_74 (O_74,N_28637,N_29803);
nor UO_75 (O_75,N_28621,N_29922);
nand UO_76 (O_76,N_29593,N_29197);
or UO_77 (O_77,N_29680,N_29089);
nand UO_78 (O_78,N_29669,N_29776);
nand UO_79 (O_79,N_29589,N_28630);
nor UO_80 (O_80,N_28727,N_29163);
or UO_81 (O_81,N_29657,N_29172);
xnor UO_82 (O_82,N_28579,N_29278);
and UO_83 (O_83,N_29063,N_29613);
and UO_84 (O_84,N_29888,N_29950);
and UO_85 (O_85,N_29136,N_29337);
xor UO_86 (O_86,N_29090,N_28563);
nand UO_87 (O_87,N_29999,N_28798);
and UO_88 (O_88,N_29581,N_29768);
nor UO_89 (O_89,N_28751,N_28641);
nand UO_90 (O_90,N_29540,N_29756);
xor UO_91 (O_91,N_29832,N_29387);
nand UO_92 (O_92,N_29004,N_29655);
xor UO_93 (O_93,N_28847,N_29365);
and UO_94 (O_94,N_28971,N_29200);
nor UO_95 (O_95,N_28666,N_29097);
nor UO_96 (O_96,N_29033,N_29710);
and UO_97 (O_97,N_29573,N_28862);
xor UO_98 (O_98,N_29786,N_29866);
and UO_99 (O_99,N_29775,N_29112);
and UO_100 (O_100,N_29798,N_29073);
nor UO_101 (O_101,N_28660,N_29692);
or UO_102 (O_102,N_28785,N_28654);
nor UO_103 (O_103,N_29695,N_29096);
nand UO_104 (O_104,N_29632,N_29627);
xor UO_105 (O_105,N_28677,N_29480);
and UO_106 (O_106,N_28504,N_29837);
nand UO_107 (O_107,N_29564,N_29194);
or UO_108 (O_108,N_29476,N_29862);
nor UO_109 (O_109,N_28565,N_29121);
or UO_110 (O_110,N_29027,N_28566);
nor UO_111 (O_111,N_29462,N_28663);
or UO_112 (O_112,N_29915,N_29659);
and UO_113 (O_113,N_28568,N_28793);
or UO_114 (O_114,N_28529,N_28577);
and UO_115 (O_115,N_29691,N_29223);
and UO_116 (O_116,N_29973,N_28635);
nand UO_117 (O_117,N_28986,N_29653);
or UO_118 (O_118,N_29687,N_29968);
and UO_119 (O_119,N_29967,N_28992);
xor UO_120 (O_120,N_29629,N_29512);
and UO_121 (O_121,N_28689,N_28943);
xnor UO_122 (O_122,N_29330,N_29638);
nand UO_123 (O_123,N_28908,N_28993);
nand UO_124 (O_124,N_29062,N_29298);
or UO_125 (O_125,N_29236,N_29539);
and UO_126 (O_126,N_29974,N_28781);
and UO_127 (O_127,N_29234,N_29519);
nor UO_128 (O_128,N_29893,N_29331);
xor UO_129 (O_129,N_29128,N_28538);
nand UO_130 (O_130,N_29554,N_29407);
nand UO_131 (O_131,N_29282,N_29319);
xor UO_132 (O_132,N_28818,N_29815);
nand UO_133 (O_133,N_28837,N_29906);
xor UO_134 (O_134,N_29017,N_28850);
xor UO_135 (O_135,N_29471,N_29118);
nand UO_136 (O_136,N_28776,N_28899);
or UO_137 (O_137,N_29596,N_28933);
or UO_138 (O_138,N_29671,N_29391);
nand UO_139 (O_139,N_28795,N_29087);
xnor UO_140 (O_140,N_28981,N_29182);
nor UO_141 (O_141,N_28824,N_29738);
nand UO_142 (O_142,N_29230,N_29148);
xor UO_143 (O_143,N_28710,N_28557);
or UO_144 (O_144,N_28548,N_28757);
and UO_145 (O_145,N_29711,N_28890);
nor UO_146 (O_146,N_28878,N_28584);
xor UO_147 (O_147,N_29035,N_28705);
nand UO_148 (O_148,N_29328,N_28636);
and UO_149 (O_149,N_28728,N_29771);
or UO_150 (O_150,N_29849,N_28658);
nor UO_151 (O_151,N_29885,N_28915);
xnor UO_152 (O_152,N_28999,N_28729);
nand UO_153 (O_153,N_29676,N_29457);
and UO_154 (O_154,N_29621,N_28860);
nor UO_155 (O_155,N_29697,N_29161);
nand UO_156 (O_156,N_29934,N_29699);
nand UO_157 (O_157,N_29708,N_29907);
nand UO_158 (O_158,N_29456,N_29714);
nor UO_159 (O_159,N_29464,N_29198);
or UO_160 (O_160,N_29742,N_28683);
and UO_161 (O_161,N_28593,N_28619);
or UO_162 (O_162,N_29508,N_29928);
xnor UO_163 (O_163,N_29061,N_29162);
and UO_164 (O_164,N_29681,N_29529);
and UO_165 (O_165,N_29716,N_29381);
and UO_166 (O_166,N_29216,N_28920);
nand UO_167 (O_167,N_29279,N_29802);
and UO_168 (O_168,N_29690,N_29984);
or UO_169 (O_169,N_29455,N_29662);
nand UO_170 (O_170,N_29419,N_28972);
and UO_171 (O_171,N_29651,N_29044);
xor UO_172 (O_172,N_29010,N_29203);
nor UO_173 (O_173,N_29232,N_29715);
or UO_174 (O_174,N_28714,N_29809);
nand UO_175 (O_175,N_29853,N_29856);
and UO_176 (O_176,N_29685,N_29770);
xnor UO_177 (O_177,N_28639,N_29287);
nor UO_178 (O_178,N_29436,N_29667);
nor UO_179 (O_179,N_28969,N_29886);
nor UO_180 (O_180,N_29268,N_29007);
and UO_181 (O_181,N_28595,N_28668);
or UO_182 (O_182,N_28703,N_29313);
nor UO_183 (O_183,N_29293,N_28622);
nand UO_184 (O_184,N_29835,N_28644);
nor UO_185 (O_185,N_29231,N_29897);
and UO_186 (O_186,N_29481,N_29498);
or UO_187 (O_187,N_29066,N_28788);
nor UO_188 (O_188,N_29649,N_29076);
nor UO_189 (O_189,N_28913,N_28934);
nand UO_190 (O_190,N_28773,N_28843);
and UO_191 (O_191,N_29022,N_28708);
nor UO_192 (O_192,N_29341,N_28676);
and UO_193 (O_193,N_29818,N_29080);
nand UO_194 (O_194,N_28725,N_28740);
nor UO_195 (O_195,N_29294,N_29343);
nor UO_196 (O_196,N_28875,N_29202);
nand UO_197 (O_197,N_28927,N_28859);
and UO_198 (O_198,N_29624,N_28506);
nor UO_199 (O_199,N_29535,N_28946);
or UO_200 (O_200,N_29421,N_29167);
and UO_201 (O_201,N_29397,N_29726);
or UO_202 (O_202,N_28713,N_29990);
or UO_203 (O_203,N_29473,N_28684);
and UO_204 (O_204,N_29969,N_29590);
xnor UO_205 (O_205,N_29355,N_29213);
and UO_206 (O_206,N_29130,N_29673);
or UO_207 (O_207,N_28616,N_28893);
xnor UO_208 (O_208,N_29447,N_28755);
nand UO_209 (O_209,N_29143,N_28980);
xnor UO_210 (O_210,N_29595,N_29487);
nand UO_211 (O_211,N_29424,N_29500);
or UO_212 (O_212,N_29981,N_29542);
nand UO_213 (O_213,N_29065,N_29762);
or UO_214 (O_214,N_29208,N_29851);
xnor UO_215 (O_215,N_28864,N_29159);
or UO_216 (O_216,N_29147,N_29448);
or UO_217 (O_217,N_28573,N_29942);
and UO_218 (O_218,N_29545,N_29980);
nor UO_219 (O_219,N_29102,N_29575);
or UO_220 (O_220,N_29727,N_28873);
or UO_221 (O_221,N_29871,N_29354);
or UO_222 (O_222,N_29737,N_29538);
nor UO_223 (O_223,N_29021,N_29260);
nand UO_224 (O_224,N_28581,N_29619);
nand UO_225 (O_225,N_29547,N_28602);
and UO_226 (O_226,N_29895,N_29070);
nor UO_227 (O_227,N_29083,N_28937);
xor UO_228 (O_228,N_29808,N_29369);
xnor UO_229 (O_229,N_29914,N_28756);
nor UO_230 (O_230,N_29393,N_29637);
nor UO_231 (O_231,N_29747,N_28603);
nand UO_232 (O_232,N_29926,N_28554);
xor UO_233 (O_233,N_29694,N_29205);
nand UO_234 (O_234,N_28503,N_29485);
nand UO_235 (O_235,N_28995,N_29943);
or UO_236 (O_236,N_28816,N_28704);
and UO_237 (O_237,N_28904,N_29241);
or UO_238 (O_238,N_29426,N_29016);
nand UO_239 (O_239,N_29578,N_29109);
or UO_240 (O_240,N_29401,N_29859);
xnor UO_241 (O_241,N_29413,N_28505);
nor UO_242 (O_242,N_29765,N_28580);
or UO_243 (O_243,N_29192,N_29122);
and UO_244 (O_244,N_29249,N_29002);
nor UO_245 (O_245,N_29992,N_28894);
xor UO_246 (O_246,N_29790,N_29396);
xor UO_247 (O_247,N_29602,N_29647);
or UO_248 (O_248,N_28970,N_29993);
and UO_249 (O_249,N_29222,N_29142);
nor UO_250 (O_250,N_29733,N_28987);
xnor UO_251 (O_251,N_28779,N_29403);
xnor UO_252 (O_252,N_29041,N_29156);
or UO_253 (O_253,N_28748,N_29700);
or UO_254 (O_254,N_29555,N_29215);
nand UO_255 (O_255,N_28968,N_29614);
or UO_256 (O_256,N_28783,N_29842);
or UO_257 (O_257,N_29067,N_29190);
or UO_258 (O_258,N_28978,N_28536);
or UO_259 (O_259,N_29625,N_29404);
nand UO_260 (O_260,N_29830,N_29826);
xnor UO_261 (O_261,N_28962,N_28907);
xnor UO_262 (O_262,N_29858,N_29281);
xor UO_263 (O_263,N_28617,N_28784);
or UO_264 (O_264,N_29930,N_29560);
or UO_265 (O_265,N_29865,N_29346);
or UO_266 (O_266,N_29546,N_28802);
nor UO_267 (O_267,N_29378,N_29445);
nand UO_268 (O_268,N_28928,N_29582);
xor UO_269 (O_269,N_28975,N_28782);
or UO_270 (O_270,N_29431,N_29339);
xnor UO_271 (O_271,N_29434,N_29759);
and UO_272 (O_272,N_28743,N_28631);
nand UO_273 (O_273,N_29848,N_28819);
and UO_274 (O_274,N_29878,N_29875);
and UO_275 (O_275,N_29777,N_29502);
and UO_276 (O_276,N_29259,N_29263);
nor UO_277 (O_277,N_28508,N_28511);
nand UO_278 (O_278,N_29201,N_28645);
or UO_279 (O_279,N_28530,N_29437);
nor UO_280 (O_280,N_29039,N_28896);
nand UO_281 (O_281,N_28923,N_28547);
xnor UO_282 (O_282,N_29359,N_28825);
nand UO_283 (O_283,N_28605,N_29739);
xor UO_284 (O_284,N_29633,N_29368);
xnor UO_285 (O_285,N_28855,N_29996);
or UO_286 (O_286,N_29841,N_29001);
or UO_287 (O_287,N_28897,N_29029);
xor UO_288 (O_288,N_29049,N_29876);
nand UO_289 (O_289,N_29266,N_28738);
nand UO_290 (O_290,N_29115,N_29218);
and UO_291 (O_291,N_29301,N_29412);
and UO_292 (O_292,N_29600,N_28752);
nor UO_293 (O_293,N_29827,N_29873);
xnor UO_294 (O_294,N_29408,N_29214);
nand UO_295 (O_295,N_28601,N_28853);
nor UO_296 (O_296,N_29243,N_29085);
nor UO_297 (O_297,N_29908,N_29988);
xnor UO_298 (O_298,N_28537,N_28868);
xnor UO_299 (O_299,N_29845,N_28510);
nand UO_300 (O_300,N_28789,N_28966);
xnor UO_301 (O_301,N_29843,N_28791);
or UO_302 (O_302,N_29548,N_28754);
and UO_303 (O_303,N_29536,N_29601);
or UO_304 (O_304,N_29482,N_28940);
nor UO_305 (O_305,N_29454,N_28932);
nor UO_306 (O_306,N_29913,N_29077);
xnor UO_307 (O_307,N_28892,N_28556);
xnor UO_308 (O_308,N_29418,N_29489);
nand UO_309 (O_309,N_29006,N_29394);
xor UO_310 (O_310,N_29013,N_29509);
nand UO_311 (O_311,N_28874,N_29682);
nand UO_312 (O_312,N_28515,N_29854);
or UO_313 (O_313,N_29634,N_29674);
xnor UO_314 (O_314,N_28925,N_28935);
xnor UO_315 (O_315,N_29183,N_29193);
nor UO_316 (O_316,N_29840,N_29290);
or UO_317 (O_317,N_28749,N_29636);
nor UO_318 (O_318,N_29763,N_29423);
xor UO_319 (O_319,N_29844,N_29584);
nor UO_320 (O_320,N_29654,N_29551);
or UO_321 (O_321,N_28849,N_29146);
or UO_322 (O_322,N_29116,N_28623);
xnor UO_323 (O_323,N_28587,N_28611);
nand UO_324 (O_324,N_28659,N_29361);
and UO_325 (O_325,N_29552,N_29285);
or UO_326 (O_326,N_29821,N_29299);
xor UO_327 (O_327,N_29617,N_29371);
and UO_328 (O_328,N_29779,N_28513);
or UO_329 (O_329,N_29558,N_29253);
nor UO_330 (O_330,N_28553,N_29363);
or UO_331 (O_331,N_29518,N_29945);
and UO_332 (O_332,N_29663,N_29233);
nand UO_333 (O_333,N_28866,N_29874);
nor UO_334 (O_334,N_29565,N_29367);
nor UO_335 (O_335,N_29170,N_29311);
xor UO_336 (O_336,N_29987,N_28811);
or UO_337 (O_337,N_28902,N_29166);
xor UO_338 (O_338,N_29661,N_29958);
xor UO_339 (O_339,N_29280,N_29126);
xnor UO_340 (O_340,N_28898,N_29957);
and UO_341 (O_341,N_28807,N_29414);
and UO_342 (O_342,N_29348,N_28730);
xor UO_343 (O_343,N_29828,N_29292);
xor UO_344 (O_344,N_29051,N_29375);
nor UO_345 (O_345,N_28680,N_29940);
and UO_346 (O_346,N_29497,N_29571);
xor UO_347 (O_347,N_29157,N_29150);
or UO_348 (O_348,N_28732,N_29164);
nand UO_349 (O_349,N_29944,N_28858);
nand UO_350 (O_350,N_28833,N_29916);
nor UO_351 (O_351,N_28741,N_29490);
nand UO_352 (O_352,N_29415,N_29890);
xor UO_353 (O_353,N_29158,N_29537);
and UO_354 (O_354,N_29515,N_29320);
xor UO_355 (O_355,N_29219,N_28952);
xor UO_356 (O_356,N_28838,N_28576);
nand UO_357 (O_357,N_29553,N_29432);
xor UO_358 (O_358,N_29797,N_29884);
xor UO_359 (O_359,N_28716,N_29678);
xor UO_360 (O_360,N_29606,N_28914);
xor UO_361 (O_361,N_29664,N_29787);
and UO_362 (O_362,N_28844,N_28761);
nor UO_363 (O_363,N_28590,N_28531);
nand UO_364 (O_364,N_29296,N_28922);
nand UO_365 (O_365,N_29899,N_28883);
and UO_366 (O_366,N_29054,N_28686);
xor UO_367 (O_367,N_28957,N_29081);
or UO_368 (O_368,N_29675,N_28608);
nand UO_369 (O_369,N_29823,N_29785);
nand UO_370 (O_370,N_29982,N_28888);
or UO_371 (O_371,N_29199,N_29530);
and UO_372 (O_372,N_28744,N_29640);
and UO_373 (O_373,N_29074,N_28820);
or UO_374 (O_374,N_29506,N_28528);
nand UO_375 (O_375,N_28953,N_29948);
or UO_376 (O_376,N_28560,N_29869);
and UO_377 (O_377,N_29250,N_29356);
and UO_378 (O_378,N_28674,N_29898);
nor UO_379 (O_379,N_29479,N_29373);
and UO_380 (O_380,N_29683,N_28620);
nand UO_381 (O_381,N_29392,N_29439);
or UO_382 (O_382,N_29486,N_29782);
or UO_383 (O_383,N_29740,N_28656);
nor UO_384 (O_384,N_29879,N_29872);
xnor UO_385 (O_385,N_29703,N_28780);
and UO_386 (O_386,N_28707,N_28836);
and UO_387 (O_387,N_28613,N_29141);
nand UO_388 (O_388,N_29474,N_29730);
nand UO_389 (O_389,N_29719,N_29283);
nand UO_390 (O_390,N_29069,N_29275);
nand UO_391 (O_391,N_28724,N_29184);
nand UO_392 (O_392,N_28588,N_28854);
nor UO_393 (O_393,N_29607,N_29023);
xnor UO_394 (O_394,N_29855,N_29224);
xnor UO_395 (O_395,N_29015,N_29824);
and UO_396 (O_396,N_29652,N_29329);
xnor UO_397 (O_397,N_28692,N_29570);
nand UO_398 (O_398,N_29920,N_28669);
xnor UO_399 (O_399,N_28766,N_29501);
or UO_400 (O_400,N_29389,N_29399);
nand UO_401 (O_401,N_29068,N_29376);
and UO_402 (O_402,N_29806,N_29258);
nor UO_403 (O_403,N_29995,N_28646);
and UO_404 (O_404,N_28760,N_29971);
or UO_405 (O_405,N_29861,N_28687);
xor UO_406 (O_406,N_29923,N_29611);
nand UO_407 (O_407,N_29882,N_29377);
and UO_408 (O_408,N_29020,N_29894);
nand UO_409 (O_409,N_29094,N_29970);
or UO_410 (O_410,N_29810,N_29082);
nor UO_411 (O_411,N_29154,N_29327);
nand UO_412 (O_412,N_29405,N_29416);
and UO_413 (O_413,N_28984,N_29623);
nor UO_414 (O_414,N_29977,N_28985);
nand UO_415 (O_415,N_28998,N_28884);
and UO_416 (O_416,N_29478,N_29936);
or UO_417 (O_417,N_29598,N_29251);
nand UO_418 (O_418,N_28721,N_28550);
nand UO_419 (O_419,N_28685,N_29340);
nor UO_420 (O_420,N_28930,N_29100);
nand UO_421 (O_421,N_29795,N_28558);
xor UO_422 (O_422,N_29380,N_28632);
nor UO_423 (O_423,N_29769,N_28649);
nand UO_424 (O_424,N_28712,N_29395);
xnor UO_425 (O_425,N_29731,N_28828);
nand UO_426 (O_426,N_28545,N_29129);
nand UO_427 (O_427,N_29324,N_29422);
xor UO_428 (O_428,N_29758,N_29326);
nand UO_429 (O_429,N_29748,N_28831);
or UO_430 (O_430,N_29991,N_29983);
xor UO_431 (O_431,N_28701,N_28696);
nor UO_432 (O_432,N_29180,N_29493);
or UO_433 (O_433,N_29496,N_29839);
nor UO_434 (O_434,N_29075,N_29347);
and UO_435 (O_435,N_29712,N_28690);
and UO_436 (O_436,N_29783,N_29402);
nor UO_437 (O_437,N_29921,N_28643);
nor UO_438 (O_438,N_29985,N_29736);
and UO_439 (O_439,N_28861,N_29117);
and UO_440 (O_440,N_29484,N_29059);
or UO_441 (O_441,N_29847,N_29955);
nand UO_442 (O_442,N_28762,N_29240);
xnor UO_443 (O_443,N_28570,N_29919);
and UO_444 (O_444,N_29071,N_29288);
nand UO_445 (O_445,N_28846,N_29800);
and UO_446 (O_446,N_29206,N_29468);
nand UO_447 (O_447,N_29227,N_29134);
nand UO_448 (O_448,N_29435,N_28801);
and UO_449 (O_449,N_28519,N_28821);
or UO_450 (O_450,N_29244,N_29887);
nand UO_451 (O_451,N_29549,N_29211);
nor UO_452 (O_452,N_29931,N_28768);
and UO_453 (O_453,N_29505,N_29780);
or UO_454 (O_454,N_28769,N_28830);
xnor UO_455 (O_455,N_29668,N_29757);
and UO_456 (O_456,N_29734,N_29791);
and UO_457 (O_457,N_29814,N_29559);
nor UO_458 (O_458,N_28735,N_29781);
nand UO_459 (O_459,N_29175,N_29979);
xnor UO_460 (O_460,N_29352,N_28642);
xor UO_461 (O_461,N_28650,N_28597);
xor UO_462 (O_462,N_29084,N_29760);
xor UO_463 (O_463,N_28917,N_29264);
and UO_464 (O_464,N_29901,N_29588);
xnor UO_465 (O_465,N_28722,N_28552);
xnor UO_466 (O_466,N_29026,N_29254);
nand UO_467 (O_467,N_29149,N_28610);
xor UO_468 (O_468,N_29812,N_28634);
nand UO_469 (O_469,N_28879,N_29221);
xnor UO_470 (O_470,N_28931,N_29891);
and UO_471 (O_471,N_29764,N_29195);
or UO_472 (O_472,N_29574,N_28607);
or UO_473 (O_473,N_28829,N_28512);
nor UO_474 (O_474,N_29409,N_29181);
xor UO_475 (O_475,N_29333,N_29514);
nor UO_476 (O_476,N_29441,N_28651);
and UO_477 (O_477,N_29009,N_29018);
nor UO_478 (O_478,N_29228,N_28906);
nor UO_479 (O_479,N_29838,N_29725);
nand UO_480 (O_480,N_28544,N_29978);
xnor UO_481 (O_481,N_28594,N_28700);
xnor UO_482 (O_482,N_29091,N_28799);
or UO_483 (O_483,N_29079,N_29179);
nor UO_484 (O_484,N_28662,N_28835);
or UO_485 (O_485,N_28814,N_29171);
and UO_486 (O_486,N_28882,N_28842);
and UO_487 (O_487,N_29212,N_29030);
nand UO_488 (O_488,N_29829,N_28675);
nor UO_489 (O_489,N_28822,N_29962);
nand UO_490 (O_490,N_29822,N_28891);
xor UO_491 (O_491,N_28653,N_29513);
nand UO_492 (O_492,N_28955,N_28678);
and UO_493 (O_493,N_28956,N_29550);
and UO_494 (O_494,N_28977,N_28759);
and UO_495 (O_495,N_28509,N_28876);
and UO_496 (O_496,N_29295,N_29951);
nor UO_497 (O_497,N_28647,N_28994);
or UO_498 (O_498,N_28942,N_29857);
or UO_499 (O_499,N_28681,N_29511);
nand UO_500 (O_500,N_29591,N_28961);
and UO_501 (O_501,N_29976,N_29103);
xnor UO_502 (O_502,N_29133,N_29120);
nand UO_503 (O_503,N_29937,N_28912);
or UO_504 (O_504,N_29963,N_29772);
or UO_505 (O_505,N_29188,N_29495);
or UO_506 (O_506,N_29155,N_28950);
or UO_507 (O_507,N_29168,N_29693);
xnor UO_508 (O_508,N_29521,N_28758);
nand UO_509 (O_509,N_29095,N_29639);
or UO_510 (O_510,N_29544,N_29332);
xnor UO_511 (O_511,N_28887,N_28599);
xor UO_512 (O_512,N_29483,N_29774);
nor UO_513 (O_513,N_29576,N_28947);
nor UO_514 (O_514,N_28869,N_28870);
nand UO_515 (O_515,N_28667,N_29052);
or UO_516 (O_516,N_29989,N_28688);
xnor UO_517 (O_517,N_29569,N_29003);
xnor UO_518 (O_518,N_28598,N_29056);
nor UO_519 (O_519,N_28747,N_28936);
xnor UO_520 (O_520,N_29262,N_28702);
nand UO_521 (O_521,N_28723,N_29226);
nand UO_522 (O_522,N_29543,N_29105);
nand UO_523 (O_523,N_29272,N_29289);
xnor UO_524 (O_524,N_29941,N_29965);
nor UO_525 (O_525,N_28804,N_29910);
and UO_526 (O_526,N_28737,N_28582);
nor UO_527 (O_527,N_29510,N_29314);
xnor UO_528 (O_528,N_28518,N_29586);
and UO_529 (O_529,N_28965,N_29960);
nand UO_530 (O_530,N_28996,N_28857);
and UO_531 (O_531,N_29925,N_28963);
and UO_532 (O_532,N_28575,N_29717);
nor UO_533 (O_533,N_28796,N_29850);
and UO_534 (O_534,N_29111,N_29357);
nand UO_535 (O_535,N_29458,N_29784);
or UO_536 (O_536,N_29488,N_29964);
nand UO_537 (O_537,N_29609,N_28549);
nand UO_538 (O_538,N_28812,N_28697);
and UO_539 (O_539,N_29975,N_29046);
and UO_540 (O_540,N_29612,N_29688);
nand UO_541 (O_541,N_28542,N_29867);
xnor UO_542 (O_542,N_28983,N_28564);
and UO_543 (O_543,N_28736,N_28764);
nand UO_544 (O_544,N_29788,N_29594);
or UO_545 (O_545,N_28502,N_28534);
xor UO_546 (O_546,N_28572,N_29463);
and UO_547 (O_547,N_29043,N_29078);
nor UO_548 (O_548,N_29477,N_29316);
xnor UO_549 (O_549,N_28805,N_28767);
nand UO_550 (O_550,N_28585,N_29104);
nand UO_551 (O_551,N_29754,N_29881);
and UO_552 (O_552,N_28941,N_28774);
nand UO_553 (O_553,N_28665,N_29522);
or UO_554 (O_554,N_28944,N_29417);
xor UO_555 (O_555,N_29338,N_28797);
or UO_556 (O_556,N_29804,N_28661);
xor UO_557 (O_557,N_29265,N_29599);
nor UO_558 (O_558,N_29031,N_29246);
or UO_559 (O_559,N_29905,N_29323);
and UO_560 (O_560,N_28911,N_29836);
nor UO_561 (O_561,N_29709,N_28596);
xor UO_562 (O_562,N_29904,N_28771);
nor UO_563 (O_563,N_29608,N_29286);
and UO_564 (O_564,N_28840,N_28698);
xor UO_565 (O_565,N_29745,N_28856);
and UO_566 (O_566,N_29245,N_29229);
or UO_567 (O_567,N_29132,N_29092);
nand UO_568 (O_568,N_29721,N_29267);
and UO_569 (O_569,N_29953,N_28664);
nor UO_570 (O_570,N_28718,N_29603);
or UO_571 (O_571,N_29620,N_29342);
and UO_572 (O_572,N_29032,N_29572);
nand UO_573 (O_573,N_29291,N_29935);
or UO_574 (O_574,N_28532,N_28520);
xnor UO_575 (O_575,N_29846,N_29099);
or UO_576 (O_576,N_28525,N_28562);
xor UO_577 (O_577,N_29470,N_29811);
nand UO_578 (O_578,N_29185,N_28910);
xor UO_579 (O_579,N_28826,N_29938);
and UO_580 (O_580,N_29137,N_28989);
xor UO_581 (O_581,N_29110,N_29531);
nor UO_582 (O_582,N_28567,N_29191);
nand UO_583 (O_583,N_29656,N_28938);
or UO_584 (O_584,N_29303,N_28709);
and UO_585 (O_585,N_28739,N_28841);
and UO_586 (O_586,N_28720,N_28982);
nor UO_587 (O_587,N_29577,N_29225);
nand UO_588 (O_588,N_29646,N_28750);
or UO_589 (O_589,N_29954,N_29520);
xnor UO_590 (O_590,N_29325,N_28867);
nand UO_591 (O_591,N_29060,N_29277);
xor UO_592 (O_592,N_29817,N_28673);
and UO_593 (O_593,N_29048,N_29169);
nor UO_594 (O_594,N_28945,N_28753);
or UO_595 (O_595,N_29207,N_28546);
nand UO_596 (O_596,N_28919,N_29644);
nand UO_597 (O_597,N_29986,N_28578);
and UO_598 (O_598,N_28625,N_29807);
or UO_599 (O_599,N_29503,N_29670);
xor UO_600 (O_600,N_29643,N_29933);
or UO_601 (O_601,N_29883,N_29443);
nand UO_602 (O_602,N_29276,N_28823);
or UO_603 (O_603,N_29040,N_29308);
xor UO_604 (O_604,N_29459,N_28974);
xnor UO_605 (O_605,N_29902,N_29580);
nor UO_606 (O_606,N_28976,N_29966);
nor UO_607 (O_607,N_29360,N_28905);
nand UO_608 (O_608,N_29239,N_29541);
nand UO_609 (O_609,N_28900,N_29722);
and UO_610 (O_610,N_29880,N_28574);
and UO_611 (O_611,N_28997,N_28916);
or UO_612 (O_612,N_29561,N_28794);
xor UO_613 (O_613,N_28786,N_29334);
and UO_614 (O_614,N_29959,N_29796);
nor UO_615 (O_615,N_29350,N_28954);
and UO_616 (O_616,N_29833,N_28670);
nand UO_617 (O_617,N_29635,N_29138);
xor UO_618 (O_618,N_28813,N_28615);
and UO_619 (O_619,N_29045,N_29641);
nand UO_620 (O_620,N_28500,N_29189);
nor UO_621 (O_621,N_29583,N_29305);
and UO_622 (O_622,N_28731,N_29335);
xnor UO_623 (O_623,N_28652,N_29799);
nor UO_624 (O_624,N_28507,N_28848);
nor UO_625 (O_625,N_29813,N_28733);
xnor UO_626 (O_626,N_29452,N_29952);
nand UO_627 (O_627,N_29107,N_29140);
or UO_628 (O_628,N_28539,N_29723);
nor UO_629 (O_629,N_28924,N_28777);
nor UO_630 (O_630,N_29677,N_29707);
nand UO_631 (O_631,N_28926,N_28909);
nor UO_632 (O_632,N_29315,N_29309);
nand UO_633 (O_633,N_29400,N_28817);
or UO_634 (O_634,N_29135,N_29900);
and UO_635 (O_635,N_29820,N_28827);
nor UO_636 (O_636,N_29028,N_29322);
nor UO_637 (O_637,N_29247,N_29660);
and UO_638 (O_638,N_29460,N_29533);
nand UO_639 (O_639,N_28571,N_29187);
and UO_640 (O_640,N_28604,N_29877);
and UO_641 (O_641,N_28526,N_28719);
xnor UO_642 (O_642,N_29504,N_29864);
nor UO_643 (O_643,N_28901,N_29597);
xor UO_644 (O_644,N_29430,N_28959);
xor UO_645 (O_645,N_28514,N_29217);
nand UO_646 (O_646,N_29364,N_29008);
nand UO_647 (O_647,N_29494,N_29297);
and UO_648 (O_648,N_28967,N_29257);
nor UO_649 (O_649,N_28715,N_29718);
nor UO_650 (O_650,N_28832,N_29626);
nand UO_651 (O_651,N_29425,N_28979);
xnor UO_652 (O_652,N_28871,N_29123);
xor UO_653 (O_653,N_29912,N_28951);
xnor UO_654 (O_654,N_29237,N_28949);
nand UO_655 (O_655,N_29160,N_29794);
and UO_656 (O_656,N_29994,N_29353);
or UO_657 (O_657,N_28671,N_29204);
nand UO_658 (O_658,N_28533,N_29924);
or UO_659 (O_659,N_29036,N_29618);
nor UO_660 (O_660,N_29145,N_29351);
nand UO_661 (O_661,N_29949,N_28778);
xnor UO_662 (O_662,N_29642,N_28775);
nand UO_663 (O_663,N_29388,N_29672);
and UO_664 (O_664,N_28885,N_28973);
nand UO_665 (O_665,N_29173,N_28706);
or UO_666 (O_666,N_28865,N_28851);
nor UO_667 (O_667,N_29379,N_28765);
or UO_668 (O_668,N_29563,N_29057);
xnor UO_669 (O_669,N_28606,N_28699);
xor UO_670 (O_670,N_28541,N_29778);
nor UO_671 (O_671,N_29567,N_29753);
nand UO_672 (O_672,N_29307,N_29209);
and UO_673 (O_673,N_29384,N_28800);
nor UO_674 (O_674,N_29698,N_29793);
xor UO_675 (O_675,N_29235,N_28521);
and UO_676 (O_676,N_28624,N_29701);
xor UO_677 (O_677,N_28695,N_29801);
nor UO_678 (O_678,N_29196,N_29034);
nand UO_679 (O_679,N_29248,N_29374);
and UO_680 (O_680,N_28679,N_29645);
xor UO_681 (O_681,N_29650,N_29186);
nand UO_682 (O_682,N_29610,N_28742);
nor UO_683 (O_683,N_28711,N_29932);
nor UO_684 (O_684,N_29321,N_28834);
and UO_685 (O_685,N_29689,N_29442);
nor UO_686 (O_686,N_28988,N_29524);
nand UO_687 (O_687,N_29616,N_29465);
nor UO_688 (O_688,N_28583,N_28648);
xnor UO_689 (O_689,N_29773,N_29720);
nor UO_690 (O_690,N_29750,N_28939);
or UO_691 (O_691,N_28770,N_29903);
or UO_692 (O_692,N_28691,N_28717);
and UO_693 (O_693,N_29119,N_29050);
xnor UO_694 (O_694,N_28672,N_29101);
xnor UO_695 (O_695,N_29805,N_29523);
or UO_696 (O_696,N_29238,N_29728);
nor UO_697 (O_697,N_29615,N_28609);
xor UO_698 (O_698,N_29300,N_29526);
and UO_699 (O_699,N_29713,N_28958);
or UO_700 (O_700,N_28638,N_29255);
or UO_701 (O_701,N_29587,N_29382);
nor UO_702 (O_702,N_28881,N_28627);
nand UO_703 (O_703,N_28618,N_29420);
nor UO_704 (O_704,N_29270,N_28600);
nor UO_705 (O_705,N_29385,N_29440);
nand UO_706 (O_706,N_29648,N_29792);
nor UO_707 (O_707,N_29946,N_29852);
xnor UO_708 (O_708,N_28655,N_29917);
or UO_709 (O_709,N_29131,N_29557);
or UO_710 (O_710,N_28543,N_29362);
nand UO_711 (O_711,N_29410,N_29005);
nand UO_712 (O_712,N_28763,N_29868);
and UO_713 (O_713,N_29870,N_29306);
nor UO_714 (O_714,N_28569,N_29741);
and UO_715 (O_715,N_29467,N_29372);
nand UO_716 (O_716,N_29113,N_29834);
nor UO_717 (O_717,N_29242,N_29000);
nand UO_718 (O_718,N_28586,N_29743);
nand UO_719 (O_719,N_28948,N_29997);
and UO_720 (O_720,N_29144,N_29014);
nor UO_721 (O_721,N_29124,N_29684);
nand UO_722 (O_722,N_29284,N_29153);
and UO_723 (O_723,N_28633,N_29178);
nor UO_724 (O_724,N_29210,N_28991);
and UO_725 (O_725,N_29345,N_28629);
or UO_726 (O_726,N_29088,N_28523);
nor UO_727 (O_727,N_29929,N_29735);
xnor UO_728 (O_728,N_29012,N_28524);
xor UO_729 (O_729,N_29492,N_29579);
nor UO_730 (O_730,N_29491,N_29939);
nand UO_731 (O_731,N_29816,N_28886);
nand UO_732 (O_732,N_29108,N_29517);
and UO_733 (O_733,N_29704,N_29358);
xor UO_734 (O_734,N_29525,N_29450);
or UO_735 (O_735,N_29461,N_29252);
nor UO_736 (O_736,N_29271,N_29011);
or UO_737 (O_737,N_29761,N_28863);
and UO_738 (O_738,N_29127,N_29344);
nand UO_739 (O_739,N_28559,N_29998);
nand UO_740 (O_740,N_29370,N_29444);
and UO_741 (O_741,N_29961,N_29165);
and UO_742 (O_742,N_29438,N_29630);
nand UO_743 (O_743,N_29025,N_29507);
xnor UO_744 (O_744,N_28657,N_28787);
nor UO_745 (O_745,N_29918,N_29453);
nand UO_746 (O_746,N_29585,N_29042);
or UO_747 (O_747,N_29256,N_29766);
nand UO_748 (O_748,N_29446,N_29139);
or UO_749 (O_749,N_29705,N_28561);
xnor UO_750 (O_750,N_28628,N_28992);
xor UO_751 (O_751,N_28894,N_28542);
xnor UO_752 (O_752,N_29576,N_29298);
nand UO_753 (O_753,N_29742,N_29631);
and UO_754 (O_754,N_28977,N_29928);
or UO_755 (O_755,N_28578,N_29054);
xor UO_756 (O_756,N_29766,N_29668);
xor UO_757 (O_757,N_29961,N_29785);
nor UO_758 (O_758,N_29343,N_29418);
xor UO_759 (O_759,N_29263,N_29715);
nand UO_760 (O_760,N_29445,N_28651);
nor UO_761 (O_761,N_29117,N_29536);
nand UO_762 (O_762,N_29258,N_29228);
or UO_763 (O_763,N_29995,N_29342);
or UO_764 (O_764,N_29337,N_29140);
nor UO_765 (O_765,N_28690,N_29285);
nand UO_766 (O_766,N_29575,N_29763);
xor UO_767 (O_767,N_29603,N_29702);
and UO_768 (O_768,N_28947,N_29030);
nor UO_769 (O_769,N_29969,N_28674);
nor UO_770 (O_770,N_28849,N_29960);
nand UO_771 (O_771,N_28618,N_29773);
nor UO_772 (O_772,N_29341,N_29122);
or UO_773 (O_773,N_29498,N_29001);
or UO_774 (O_774,N_28909,N_29851);
nand UO_775 (O_775,N_29229,N_29887);
nor UO_776 (O_776,N_28870,N_28677);
nand UO_777 (O_777,N_29686,N_28768);
nand UO_778 (O_778,N_29517,N_28717);
xor UO_779 (O_779,N_28883,N_29634);
xnor UO_780 (O_780,N_29340,N_28871);
nand UO_781 (O_781,N_29846,N_29216);
xnor UO_782 (O_782,N_29783,N_29988);
nor UO_783 (O_783,N_28894,N_29521);
nand UO_784 (O_784,N_28824,N_29141);
or UO_785 (O_785,N_29648,N_29894);
nor UO_786 (O_786,N_29551,N_28605);
xnor UO_787 (O_787,N_29917,N_28649);
or UO_788 (O_788,N_28891,N_29057);
nor UO_789 (O_789,N_29645,N_28778);
nor UO_790 (O_790,N_29609,N_29041);
nand UO_791 (O_791,N_28534,N_29631);
and UO_792 (O_792,N_28703,N_29353);
or UO_793 (O_793,N_29141,N_29007);
nor UO_794 (O_794,N_28553,N_28638);
or UO_795 (O_795,N_29961,N_28538);
xnor UO_796 (O_796,N_29855,N_28779);
nor UO_797 (O_797,N_29261,N_28706);
and UO_798 (O_798,N_28698,N_28500);
nand UO_799 (O_799,N_29808,N_29704);
or UO_800 (O_800,N_29730,N_28717);
nor UO_801 (O_801,N_29154,N_29241);
nor UO_802 (O_802,N_29763,N_29592);
xor UO_803 (O_803,N_28764,N_28513);
or UO_804 (O_804,N_29516,N_29351);
and UO_805 (O_805,N_28778,N_28858);
and UO_806 (O_806,N_28860,N_29620);
xor UO_807 (O_807,N_28766,N_29789);
nand UO_808 (O_808,N_28564,N_29490);
xor UO_809 (O_809,N_29253,N_29627);
nor UO_810 (O_810,N_29809,N_29879);
nor UO_811 (O_811,N_29100,N_29682);
xor UO_812 (O_812,N_29650,N_28622);
nand UO_813 (O_813,N_29807,N_29833);
or UO_814 (O_814,N_29394,N_28922);
nand UO_815 (O_815,N_28839,N_28594);
or UO_816 (O_816,N_29577,N_29428);
or UO_817 (O_817,N_29969,N_28562);
nor UO_818 (O_818,N_29351,N_29450);
nand UO_819 (O_819,N_29931,N_28705);
nor UO_820 (O_820,N_29886,N_29220);
and UO_821 (O_821,N_29673,N_28909);
xor UO_822 (O_822,N_29489,N_29390);
xnor UO_823 (O_823,N_29221,N_29882);
xnor UO_824 (O_824,N_28958,N_29634);
or UO_825 (O_825,N_28813,N_29913);
xnor UO_826 (O_826,N_29426,N_29701);
nor UO_827 (O_827,N_29622,N_28696);
and UO_828 (O_828,N_29472,N_29389);
nor UO_829 (O_829,N_28892,N_29624);
or UO_830 (O_830,N_29420,N_29017);
xnor UO_831 (O_831,N_28769,N_28919);
nor UO_832 (O_832,N_29080,N_28916);
xnor UO_833 (O_833,N_29801,N_29558);
and UO_834 (O_834,N_28955,N_28505);
nor UO_835 (O_835,N_28589,N_29935);
and UO_836 (O_836,N_29255,N_29375);
nand UO_837 (O_837,N_29453,N_29149);
xor UO_838 (O_838,N_29178,N_28934);
xor UO_839 (O_839,N_28522,N_28923);
and UO_840 (O_840,N_28818,N_29051);
nand UO_841 (O_841,N_28928,N_29194);
nor UO_842 (O_842,N_29241,N_29326);
nor UO_843 (O_843,N_28980,N_28578);
nor UO_844 (O_844,N_29424,N_29306);
xor UO_845 (O_845,N_28595,N_28746);
nor UO_846 (O_846,N_29211,N_29755);
or UO_847 (O_847,N_29249,N_29037);
and UO_848 (O_848,N_28887,N_29663);
and UO_849 (O_849,N_29497,N_28805);
or UO_850 (O_850,N_29636,N_29687);
nand UO_851 (O_851,N_29879,N_29548);
or UO_852 (O_852,N_29253,N_28720);
nand UO_853 (O_853,N_29155,N_28927);
or UO_854 (O_854,N_29072,N_29299);
and UO_855 (O_855,N_28761,N_29127);
nand UO_856 (O_856,N_29415,N_29586);
and UO_857 (O_857,N_29152,N_28778);
nor UO_858 (O_858,N_29679,N_29699);
and UO_859 (O_859,N_28827,N_28606);
and UO_860 (O_860,N_28749,N_29851);
nor UO_861 (O_861,N_28537,N_29178);
nand UO_862 (O_862,N_29331,N_29461);
xnor UO_863 (O_863,N_28787,N_29111);
nor UO_864 (O_864,N_28992,N_29618);
and UO_865 (O_865,N_29500,N_28717);
nor UO_866 (O_866,N_28620,N_29614);
or UO_867 (O_867,N_28676,N_29114);
or UO_868 (O_868,N_29794,N_28591);
xnor UO_869 (O_869,N_28557,N_28776);
and UO_870 (O_870,N_29983,N_29821);
xor UO_871 (O_871,N_28678,N_29845);
or UO_872 (O_872,N_28580,N_28984);
nor UO_873 (O_873,N_29246,N_29793);
nor UO_874 (O_874,N_29422,N_29076);
or UO_875 (O_875,N_29181,N_28907);
xnor UO_876 (O_876,N_29842,N_28965);
and UO_877 (O_877,N_29643,N_29297);
xnor UO_878 (O_878,N_28863,N_28647);
xnor UO_879 (O_879,N_29525,N_29168);
xor UO_880 (O_880,N_29620,N_28934);
nand UO_881 (O_881,N_29754,N_29194);
nand UO_882 (O_882,N_28731,N_29711);
nand UO_883 (O_883,N_29191,N_29478);
or UO_884 (O_884,N_29973,N_28607);
xor UO_885 (O_885,N_28832,N_29185);
nand UO_886 (O_886,N_28677,N_29576);
and UO_887 (O_887,N_29779,N_29550);
xnor UO_888 (O_888,N_28959,N_29770);
nand UO_889 (O_889,N_28987,N_29099);
xnor UO_890 (O_890,N_29646,N_29529);
xor UO_891 (O_891,N_28921,N_29719);
or UO_892 (O_892,N_29387,N_29736);
and UO_893 (O_893,N_29889,N_29851);
nand UO_894 (O_894,N_28512,N_29054);
nand UO_895 (O_895,N_29192,N_29016);
nor UO_896 (O_896,N_28512,N_28984);
nand UO_897 (O_897,N_29878,N_28942);
and UO_898 (O_898,N_29037,N_29947);
nand UO_899 (O_899,N_29042,N_29320);
or UO_900 (O_900,N_29277,N_29440);
and UO_901 (O_901,N_29040,N_29013);
nor UO_902 (O_902,N_28694,N_29568);
and UO_903 (O_903,N_28915,N_29792);
or UO_904 (O_904,N_29444,N_29860);
and UO_905 (O_905,N_28946,N_28832);
xor UO_906 (O_906,N_28863,N_29854);
xnor UO_907 (O_907,N_29506,N_28623);
nor UO_908 (O_908,N_29564,N_29440);
xor UO_909 (O_909,N_29025,N_29631);
nand UO_910 (O_910,N_29540,N_29587);
and UO_911 (O_911,N_29652,N_28652);
or UO_912 (O_912,N_29481,N_29935);
xor UO_913 (O_913,N_29852,N_29685);
or UO_914 (O_914,N_29102,N_28990);
nand UO_915 (O_915,N_28800,N_28678);
and UO_916 (O_916,N_28651,N_29399);
xnor UO_917 (O_917,N_29537,N_29562);
and UO_918 (O_918,N_28612,N_29009);
xnor UO_919 (O_919,N_29065,N_29753);
or UO_920 (O_920,N_28962,N_29854);
and UO_921 (O_921,N_29624,N_29619);
or UO_922 (O_922,N_29981,N_29308);
xor UO_923 (O_923,N_29299,N_28712);
xnor UO_924 (O_924,N_29141,N_28726);
or UO_925 (O_925,N_29136,N_29304);
nand UO_926 (O_926,N_29512,N_29942);
and UO_927 (O_927,N_28932,N_28961);
xnor UO_928 (O_928,N_29037,N_29032);
nand UO_929 (O_929,N_29782,N_29468);
or UO_930 (O_930,N_28599,N_29482);
nand UO_931 (O_931,N_29473,N_29696);
xor UO_932 (O_932,N_29422,N_28866);
nor UO_933 (O_933,N_29667,N_28825);
nor UO_934 (O_934,N_28911,N_28549);
or UO_935 (O_935,N_29052,N_28570);
or UO_936 (O_936,N_29007,N_28509);
or UO_937 (O_937,N_28848,N_29180);
xor UO_938 (O_938,N_29462,N_29736);
and UO_939 (O_939,N_29523,N_29328);
or UO_940 (O_940,N_28713,N_29135);
and UO_941 (O_941,N_29992,N_29326);
nor UO_942 (O_942,N_29633,N_29192);
xor UO_943 (O_943,N_28829,N_29862);
nand UO_944 (O_944,N_28684,N_29666);
xnor UO_945 (O_945,N_29097,N_29544);
nor UO_946 (O_946,N_29970,N_29228);
and UO_947 (O_947,N_29982,N_29182);
xor UO_948 (O_948,N_29136,N_29310);
or UO_949 (O_949,N_29960,N_28985);
nand UO_950 (O_950,N_29763,N_29831);
or UO_951 (O_951,N_28597,N_29638);
nor UO_952 (O_952,N_28770,N_29221);
and UO_953 (O_953,N_28717,N_29944);
or UO_954 (O_954,N_29337,N_29889);
nor UO_955 (O_955,N_28667,N_29988);
or UO_956 (O_956,N_28540,N_28788);
or UO_957 (O_957,N_29058,N_29896);
nor UO_958 (O_958,N_29572,N_29468);
or UO_959 (O_959,N_29159,N_29602);
nor UO_960 (O_960,N_28746,N_29363);
nor UO_961 (O_961,N_29595,N_29773);
and UO_962 (O_962,N_29205,N_29726);
or UO_963 (O_963,N_28800,N_29805);
and UO_964 (O_964,N_28606,N_29863);
nor UO_965 (O_965,N_28782,N_29679);
nand UO_966 (O_966,N_29673,N_29067);
xnor UO_967 (O_967,N_28604,N_28837);
and UO_968 (O_968,N_29037,N_29235);
nand UO_969 (O_969,N_29057,N_28610);
xor UO_970 (O_970,N_28596,N_28831);
or UO_971 (O_971,N_29160,N_29802);
or UO_972 (O_972,N_29200,N_29385);
or UO_973 (O_973,N_29524,N_28694);
and UO_974 (O_974,N_29769,N_29488);
or UO_975 (O_975,N_29654,N_29124);
or UO_976 (O_976,N_29759,N_29528);
xor UO_977 (O_977,N_29193,N_29347);
and UO_978 (O_978,N_28580,N_29573);
and UO_979 (O_979,N_29161,N_28511);
nand UO_980 (O_980,N_28719,N_29738);
and UO_981 (O_981,N_28827,N_28807);
or UO_982 (O_982,N_28534,N_29696);
nor UO_983 (O_983,N_29332,N_29952);
nand UO_984 (O_984,N_29315,N_28904);
nor UO_985 (O_985,N_29881,N_29270);
or UO_986 (O_986,N_29228,N_29033);
nor UO_987 (O_987,N_28942,N_28720);
xnor UO_988 (O_988,N_29615,N_29979);
and UO_989 (O_989,N_29487,N_29718);
nand UO_990 (O_990,N_28523,N_29799);
nor UO_991 (O_991,N_28956,N_28580);
or UO_992 (O_992,N_29359,N_29972);
nand UO_993 (O_993,N_29487,N_29102);
nand UO_994 (O_994,N_29145,N_28530);
nand UO_995 (O_995,N_29028,N_29849);
nand UO_996 (O_996,N_29654,N_29247);
xnor UO_997 (O_997,N_28647,N_29924);
nand UO_998 (O_998,N_29915,N_28647);
xnor UO_999 (O_999,N_29669,N_28636);
and UO_1000 (O_1000,N_29383,N_29824);
and UO_1001 (O_1001,N_29771,N_28599);
nor UO_1002 (O_1002,N_29741,N_28537);
nand UO_1003 (O_1003,N_29480,N_29815);
xor UO_1004 (O_1004,N_28587,N_28583);
and UO_1005 (O_1005,N_28636,N_29234);
and UO_1006 (O_1006,N_29190,N_29768);
xnor UO_1007 (O_1007,N_29562,N_28729);
xor UO_1008 (O_1008,N_29380,N_29763);
or UO_1009 (O_1009,N_28819,N_29756);
and UO_1010 (O_1010,N_28534,N_29449);
xor UO_1011 (O_1011,N_28579,N_29632);
xnor UO_1012 (O_1012,N_29325,N_29081);
and UO_1013 (O_1013,N_29731,N_28898);
nor UO_1014 (O_1014,N_29773,N_29829);
and UO_1015 (O_1015,N_28543,N_29186);
or UO_1016 (O_1016,N_28701,N_29107);
or UO_1017 (O_1017,N_29061,N_29708);
or UO_1018 (O_1018,N_28577,N_28836);
nand UO_1019 (O_1019,N_28894,N_29999);
and UO_1020 (O_1020,N_29678,N_28638);
nand UO_1021 (O_1021,N_29988,N_29572);
xnor UO_1022 (O_1022,N_28751,N_28657);
or UO_1023 (O_1023,N_28752,N_29888);
and UO_1024 (O_1024,N_28888,N_29340);
nand UO_1025 (O_1025,N_29004,N_29772);
xor UO_1026 (O_1026,N_29747,N_28511);
and UO_1027 (O_1027,N_29467,N_28822);
xnor UO_1028 (O_1028,N_29025,N_29256);
xnor UO_1029 (O_1029,N_28634,N_28774);
nor UO_1030 (O_1030,N_29508,N_29807);
and UO_1031 (O_1031,N_29455,N_29751);
nand UO_1032 (O_1032,N_29756,N_29059);
and UO_1033 (O_1033,N_29200,N_29424);
or UO_1034 (O_1034,N_28718,N_28541);
and UO_1035 (O_1035,N_29217,N_29509);
nand UO_1036 (O_1036,N_29359,N_29683);
nand UO_1037 (O_1037,N_28643,N_29014);
xor UO_1038 (O_1038,N_28799,N_29607);
or UO_1039 (O_1039,N_29762,N_28680);
and UO_1040 (O_1040,N_28964,N_28630);
or UO_1041 (O_1041,N_29356,N_28757);
and UO_1042 (O_1042,N_28675,N_29232);
and UO_1043 (O_1043,N_28899,N_28871);
nor UO_1044 (O_1044,N_29906,N_29434);
xor UO_1045 (O_1045,N_29103,N_28867);
nor UO_1046 (O_1046,N_28806,N_29612);
nor UO_1047 (O_1047,N_28652,N_29800);
or UO_1048 (O_1048,N_29459,N_29207);
nand UO_1049 (O_1049,N_29043,N_29705);
nand UO_1050 (O_1050,N_28769,N_28936);
and UO_1051 (O_1051,N_29012,N_29363);
and UO_1052 (O_1052,N_28680,N_28876);
or UO_1053 (O_1053,N_29632,N_28571);
nor UO_1054 (O_1054,N_28793,N_28882);
or UO_1055 (O_1055,N_29082,N_29086);
nor UO_1056 (O_1056,N_28967,N_29263);
or UO_1057 (O_1057,N_28547,N_29928);
or UO_1058 (O_1058,N_28793,N_28706);
nand UO_1059 (O_1059,N_29082,N_29909);
xor UO_1060 (O_1060,N_29387,N_29914);
or UO_1061 (O_1061,N_28741,N_29827);
nor UO_1062 (O_1062,N_29439,N_29306);
and UO_1063 (O_1063,N_29264,N_28887);
nor UO_1064 (O_1064,N_29875,N_29121);
or UO_1065 (O_1065,N_28530,N_28723);
xor UO_1066 (O_1066,N_28798,N_29145);
and UO_1067 (O_1067,N_29550,N_29169);
or UO_1068 (O_1068,N_29399,N_28620);
nand UO_1069 (O_1069,N_29645,N_29900);
and UO_1070 (O_1070,N_28888,N_28848);
xnor UO_1071 (O_1071,N_29003,N_29264);
nand UO_1072 (O_1072,N_28926,N_29534);
nor UO_1073 (O_1073,N_29248,N_29195);
and UO_1074 (O_1074,N_28736,N_28700);
nand UO_1075 (O_1075,N_29374,N_28929);
nor UO_1076 (O_1076,N_28949,N_29238);
xnor UO_1077 (O_1077,N_28926,N_29908);
or UO_1078 (O_1078,N_29739,N_29146);
nand UO_1079 (O_1079,N_29060,N_28510);
and UO_1080 (O_1080,N_29632,N_28816);
and UO_1081 (O_1081,N_28821,N_29407);
or UO_1082 (O_1082,N_29942,N_29035);
nand UO_1083 (O_1083,N_29928,N_29794);
or UO_1084 (O_1084,N_29979,N_29400);
and UO_1085 (O_1085,N_29525,N_29070);
and UO_1086 (O_1086,N_29051,N_29116);
or UO_1087 (O_1087,N_29535,N_29570);
xor UO_1088 (O_1088,N_29316,N_28740);
and UO_1089 (O_1089,N_29983,N_29386);
or UO_1090 (O_1090,N_29549,N_29410);
or UO_1091 (O_1091,N_29061,N_28801);
and UO_1092 (O_1092,N_29289,N_28737);
nand UO_1093 (O_1093,N_28941,N_29911);
nand UO_1094 (O_1094,N_29265,N_28733);
or UO_1095 (O_1095,N_29129,N_29382);
nand UO_1096 (O_1096,N_29749,N_28760);
and UO_1097 (O_1097,N_29355,N_28744);
or UO_1098 (O_1098,N_29225,N_29622);
or UO_1099 (O_1099,N_29452,N_29937);
nor UO_1100 (O_1100,N_29468,N_28754);
or UO_1101 (O_1101,N_29193,N_28703);
nor UO_1102 (O_1102,N_28771,N_28593);
nand UO_1103 (O_1103,N_29074,N_28804);
nor UO_1104 (O_1104,N_29758,N_29468);
and UO_1105 (O_1105,N_28939,N_29085);
xnor UO_1106 (O_1106,N_29743,N_29097);
nor UO_1107 (O_1107,N_29192,N_29274);
nor UO_1108 (O_1108,N_29584,N_29278);
and UO_1109 (O_1109,N_29456,N_29904);
or UO_1110 (O_1110,N_29267,N_28659);
nand UO_1111 (O_1111,N_29212,N_29767);
nor UO_1112 (O_1112,N_29851,N_29663);
and UO_1113 (O_1113,N_28646,N_29807);
nand UO_1114 (O_1114,N_29787,N_29542);
and UO_1115 (O_1115,N_29268,N_29591);
or UO_1116 (O_1116,N_28806,N_29582);
or UO_1117 (O_1117,N_29840,N_29315);
xnor UO_1118 (O_1118,N_29452,N_29601);
xnor UO_1119 (O_1119,N_28633,N_29136);
nand UO_1120 (O_1120,N_29245,N_29748);
or UO_1121 (O_1121,N_28597,N_29674);
xor UO_1122 (O_1122,N_29961,N_28783);
nor UO_1123 (O_1123,N_29682,N_29400);
and UO_1124 (O_1124,N_29155,N_29190);
nor UO_1125 (O_1125,N_29861,N_28820);
and UO_1126 (O_1126,N_28868,N_29883);
or UO_1127 (O_1127,N_29129,N_29782);
xnor UO_1128 (O_1128,N_29665,N_28571);
nor UO_1129 (O_1129,N_28973,N_29140);
nand UO_1130 (O_1130,N_28639,N_28887);
xor UO_1131 (O_1131,N_28921,N_29221);
nand UO_1132 (O_1132,N_29006,N_29264);
or UO_1133 (O_1133,N_29897,N_29517);
xnor UO_1134 (O_1134,N_29260,N_29002);
xnor UO_1135 (O_1135,N_29908,N_28682);
or UO_1136 (O_1136,N_29634,N_28551);
and UO_1137 (O_1137,N_29913,N_29617);
nor UO_1138 (O_1138,N_28903,N_28546);
xor UO_1139 (O_1139,N_29873,N_28838);
nand UO_1140 (O_1140,N_28569,N_29554);
and UO_1141 (O_1141,N_28928,N_29265);
xor UO_1142 (O_1142,N_28967,N_29530);
nor UO_1143 (O_1143,N_28893,N_28693);
xnor UO_1144 (O_1144,N_28758,N_29043);
xnor UO_1145 (O_1145,N_28915,N_28938);
or UO_1146 (O_1146,N_29696,N_29285);
or UO_1147 (O_1147,N_29054,N_29483);
or UO_1148 (O_1148,N_29779,N_28572);
nor UO_1149 (O_1149,N_29558,N_29757);
and UO_1150 (O_1150,N_29212,N_29851);
and UO_1151 (O_1151,N_29692,N_29688);
nor UO_1152 (O_1152,N_29031,N_28867);
xnor UO_1153 (O_1153,N_28969,N_29602);
and UO_1154 (O_1154,N_29267,N_29230);
and UO_1155 (O_1155,N_29725,N_29392);
and UO_1156 (O_1156,N_28542,N_29666);
and UO_1157 (O_1157,N_28586,N_29389);
or UO_1158 (O_1158,N_29519,N_29609);
and UO_1159 (O_1159,N_29879,N_29756);
nand UO_1160 (O_1160,N_29725,N_29026);
and UO_1161 (O_1161,N_29649,N_28912);
xor UO_1162 (O_1162,N_29875,N_29773);
nor UO_1163 (O_1163,N_29878,N_28934);
and UO_1164 (O_1164,N_29465,N_28859);
xor UO_1165 (O_1165,N_28658,N_29062);
nand UO_1166 (O_1166,N_28945,N_29008);
nand UO_1167 (O_1167,N_29190,N_28920);
nand UO_1168 (O_1168,N_29477,N_29400);
nor UO_1169 (O_1169,N_29108,N_28819);
nand UO_1170 (O_1170,N_28693,N_29134);
nand UO_1171 (O_1171,N_29320,N_29481);
nand UO_1172 (O_1172,N_29305,N_29165);
nor UO_1173 (O_1173,N_29695,N_29610);
nor UO_1174 (O_1174,N_29175,N_29456);
nand UO_1175 (O_1175,N_29740,N_28767);
xor UO_1176 (O_1176,N_28790,N_28557);
or UO_1177 (O_1177,N_29362,N_29516);
nor UO_1178 (O_1178,N_28516,N_29929);
nor UO_1179 (O_1179,N_29990,N_28779);
or UO_1180 (O_1180,N_28708,N_29662);
and UO_1181 (O_1181,N_28512,N_28835);
nor UO_1182 (O_1182,N_29843,N_29535);
and UO_1183 (O_1183,N_29532,N_29260);
xnor UO_1184 (O_1184,N_29143,N_28616);
nor UO_1185 (O_1185,N_29388,N_29964);
or UO_1186 (O_1186,N_29418,N_28786);
nor UO_1187 (O_1187,N_29106,N_28644);
xor UO_1188 (O_1188,N_29688,N_29203);
nor UO_1189 (O_1189,N_28637,N_29655);
xnor UO_1190 (O_1190,N_29625,N_29830);
nor UO_1191 (O_1191,N_28601,N_28596);
nor UO_1192 (O_1192,N_29244,N_28509);
and UO_1193 (O_1193,N_28872,N_28669);
or UO_1194 (O_1194,N_29380,N_29754);
or UO_1195 (O_1195,N_28968,N_29763);
xnor UO_1196 (O_1196,N_29591,N_29449);
and UO_1197 (O_1197,N_29976,N_29925);
nand UO_1198 (O_1198,N_29370,N_28613);
nand UO_1199 (O_1199,N_28906,N_28587);
or UO_1200 (O_1200,N_29652,N_28818);
or UO_1201 (O_1201,N_29289,N_29566);
nand UO_1202 (O_1202,N_29240,N_29930);
nand UO_1203 (O_1203,N_28724,N_29744);
xor UO_1204 (O_1204,N_28522,N_29263);
nand UO_1205 (O_1205,N_28649,N_29787);
or UO_1206 (O_1206,N_28916,N_28999);
xnor UO_1207 (O_1207,N_29822,N_29782);
nor UO_1208 (O_1208,N_28592,N_29551);
or UO_1209 (O_1209,N_28545,N_29134);
or UO_1210 (O_1210,N_28722,N_28549);
nor UO_1211 (O_1211,N_29243,N_29689);
xnor UO_1212 (O_1212,N_28790,N_29353);
nor UO_1213 (O_1213,N_29048,N_28840);
or UO_1214 (O_1214,N_29294,N_28650);
and UO_1215 (O_1215,N_29431,N_28926);
and UO_1216 (O_1216,N_28784,N_28796);
nor UO_1217 (O_1217,N_29008,N_28881);
nand UO_1218 (O_1218,N_28715,N_29791);
and UO_1219 (O_1219,N_29398,N_29603);
or UO_1220 (O_1220,N_29356,N_28957);
xnor UO_1221 (O_1221,N_28903,N_29212);
or UO_1222 (O_1222,N_28698,N_28859);
nand UO_1223 (O_1223,N_29828,N_29326);
nand UO_1224 (O_1224,N_29435,N_28527);
and UO_1225 (O_1225,N_29805,N_28557);
and UO_1226 (O_1226,N_28941,N_28790);
nor UO_1227 (O_1227,N_29790,N_28745);
and UO_1228 (O_1228,N_28584,N_28708);
and UO_1229 (O_1229,N_28540,N_28713);
and UO_1230 (O_1230,N_28517,N_29312);
or UO_1231 (O_1231,N_29298,N_29330);
and UO_1232 (O_1232,N_28770,N_28682);
and UO_1233 (O_1233,N_29665,N_29606);
and UO_1234 (O_1234,N_29654,N_29743);
xnor UO_1235 (O_1235,N_28908,N_29158);
nand UO_1236 (O_1236,N_29195,N_29482);
and UO_1237 (O_1237,N_29036,N_29665);
nand UO_1238 (O_1238,N_29536,N_29359);
nand UO_1239 (O_1239,N_29554,N_29692);
nand UO_1240 (O_1240,N_29014,N_28626);
nand UO_1241 (O_1241,N_29931,N_28653);
nor UO_1242 (O_1242,N_29046,N_29316);
or UO_1243 (O_1243,N_28689,N_29671);
nor UO_1244 (O_1244,N_28980,N_29955);
or UO_1245 (O_1245,N_29961,N_29831);
xnor UO_1246 (O_1246,N_29652,N_28923);
or UO_1247 (O_1247,N_28717,N_28871);
nor UO_1248 (O_1248,N_29728,N_28556);
nand UO_1249 (O_1249,N_29440,N_29704);
nor UO_1250 (O_1250,N_28681,N_29430);
or UO_1251 (O_1251,N_29591,N_29083);
or UO_1252 (O_1252,N_29588,N_29788);
or UO_1253 (O_1253,N_29481,N_28772);
nand UO_1254 (O_1254,N_29722,N_29755);
and UO_1255 (O_1255,N_29280,N_28862);
nor UO_1256 (O_1256,N_28521,N_29959);
xnor UO_1257 (O_1257,N_28991,N_29846);
xnor UO_1258 (O_1258,N_28933,N_29567);
nand UO_1259 (O_1259,N_29012,N_29239);
and UO_1260 (O_1260,N_29192,N_29468);
and UO_1261 (O_1261,N_28562,N_29675);
and UO_1262 (O_1262,N_29460,N_29868);
and UO_1263 (O_1263,N_28582,N_28855);
nor UO_1264 (O_1264,N_28599,N_29535);
xnor UO_1265 (O_1265,N_28702,N_29698);
and UO_1266 (O_1266,N_29854,N_29567);
and UO_1267 (O_1267,N_28868,N_29116);
or UO_1268 (O_1268,N_28658,N_29225);
and UO_1269 (O_1269,N_28949,N_28670);
nor UO_1270 (O_1270,N_28894,N_29426);
or UO_1271 (O_1271,N_29928,N_29856);
xnor UO_1272 (O_1272,N_29267,N_28549);
or UO_1273 (O_1273,N_28962,N_29535);
nor UO_1274 (O_1274,N_28513,N_29836);
nor UO_1275 (O_1275,N_29362,N_29232);
nor UO_1276 (O_1276,N_29918,N_28504);
or UO_1277 (O_1277,N_29869,N_29186);
and UO_1278 (O_1278,N_29351,N_28564);
and UO_1279 (O_1279,N_29047,N_28999);
nand UO_1280 (O_1280,N_28567,N_29574);
and UO_1281 (O_1281,N_28760,N_29092);
and UO_1282 (O_1282,N_29419,N_29738);
nor UO_1283 (O_1283,N_29089,N_28881);
nand UO_1284 (O_1284,N_29982,N_29725);
and UO_1285 (O_1285,N_29927,N_29392);
nand UO_1286 (O_1286,N_28814,N_29750);
xor UO_1287 (O_1287,N_29941,N_28785);
nor UO_1288 (O_1288,N_29687,N_28611);
xor UO_1289 (O_1289,N_29339,N_29258);
xor UO_1290 (O_1290,N_29636,N_29539);
nor UO_1291 (O_1291,N_28740,N_29896);
nor UO_1292 (O_1292,N_29816,N_29328);
xnor UO_1293 (O_1293,N_29756,N_29235);
nand UO_1294 (O_1294,N_29353,N_29215);
nor UO_1295 (O_1295,N_29553,N_29491);
or UO_1296 (O_1296,N_29926,N_29997);
or UO_1297 (O_1297,N_28816,N_29585);
nor UO_1298 (O_1298,N_28660,N_29456);
nand UO_1299 (O_1299,N_29022,N_29782);
nand UO_1300 (O_1300,N_29562,N_29563);
xnor UO_1301 (O_1301,N_28957,N_28565);
nand UO_1302 (O_1302,N_29119,N_28764);
or UO_1303 (O_1303,N_29733,N_29523);
xor UO_1304 (O_1304,N_29005,N_28617);
xnor UO_1305 (O_1305,N_28572,N_29503);
xnor UO_1306 (O_1306,N_29178,N_29022);
and UO_1307 (O_1307,N_28992,N_29865);
xnor UO_1308 (O_1308,N_29001,N_29414);
or UO_1309 (O_1309,N_29498,N_28948);
and UO_1310 (O_1310,N_29417,N_28644);
and UO_1311 (O_1311,N_28950,N_28874);
nand UO_1312 (O_1312,N_29904,N_29506);
xor UO_1313 (O_1313,N_28853,N_29975);
and UO_1314 (O_1314,N_29210,N_28755);
nand UO_1315 (O_1315,N_29698,N_28751);
nand UO_1316 (O_1316,N_29521,N_28986);
nand UO_1317 (O_1317,N_29956,N_28868);
nor UO_1318 (O_1318,N_28580,N_29816);
nor UO_1319 (O_1319,N_28830,N_29346);
nor UO_1320 (O_1320,N_28801,N_29556);
or UO_1321 (O_1321,N_29123,N_29113);
or UO_1322 (O_1322,N_29542,N_29508);
nand UO_1323 (O_1323,N_28801,N_29775);
xor UO_1324 (O_1324,N_29390,N_29083);
nand UO_1325 (O_1325,N_29686,N_29777);
or UO_1326 (O_1326,N_28519,N_29955);
and UO_1327 (O_1327,N_29054,N_29096);
nor UO_1328 (O_1328,N_29951,N_29317);
and UO_1329 (O_1329,N_29457,N_29488);
or UO_1330 (O_1330,N_29813,N_29927);
xor UO_1331 (O_1331,N_28928,N_29823);
xor UO_1332 (O_1332,N_29351,N_29029);
or UO_1333 (O_1333,N_29900,N_28651);
or UO_1334 (O_1334,N_28974,N_29680);
and UO_1335 (O_1335,N_28803,N_29600);
xnor UO_1336 (O_1336,N_29282,N_28720);
nand UO_1337 (O_1337,N_29035,N_28514);
nand UO_1338 (O_1338,N_29816,N_28531);
nor UO_1339 (O_1339,N_28945,N_29356);
nand UO_1340 (O_1340,N_29776,N_29264);
nand UO_1341 (O_1341,N_29923,N_28788);
nand UO_1342 (O_1342,N_29700,N_28642);
nand UO_1343 (O_1343,N_29351,N_28619);
nand UO_1344 (O_1344,N_29323,N_29770);
xnor UO_1345 (O_1345,N_28596,N_28970);
or UO_1346 (O_1346,N_29145,N_29594);
or UO_1347 (O_1347,N_29503,N_29057);
nor UO_1348 (O_1348,N_29589,N_29920);
and UO_1349 (O_1349,N_29439,N_29427);
nand UO_1350 (O_1350,N_29393,N_29674);
and UO_1351 (O_1351,N_29506,N_28542);
xnor UO_1352 (O_1352,N_29839,N_29488);
nand UO_1353 (O_1353,N_29713,N_28589);
nand UO_1354 (O_1354,N_29453,N_28856);
or UO_1355 (O_1355,N_29786,N_28697);
xor UO_1356 (O_1356,N_29157,N_29701);
nand UO_1357 (O_1357,N_29167,N_29910);
xnor UO_1358 (O_1358,N_28936,N_29468);
nor UO_1359 (O_1359,N_29740,N_28605);
nor UO_1360 (O_1360,N_28673,N_28761);
xor UO_1361 (O_1361,N_29048,N_28682);
nor UO_1362 (O_1362,N_28575,N_29320);
xnor UO_1363 (O_1363,N_29311,N_28971);
xnor UO_1364 (O_1364,N_29677,N_29768);
xor UO_1365 (O_1365,N_28985,N_28731);
nand UO_1366 (O_1366,N_28714,N_29277);
xnor UO_1367 (O_1367,N_29550,N_29483);
and UO_1368 (O_1368,N_29863,N_29851);
nand UO_1369 (O_1369,N_29535,N_29086);
nand UO_1370 (O_1370,N_29426,N_29873);
and UO_1371 (O_1371,N_29192,N_28711);
and UO_1372 (O_1372,N_29404,N_28553);
and UO_1373 (O_1373,N_28819,N_29018);
nand UO_1374 (O_1374,N_29873,N_28672);
xor UO_1375 (O_1375,N_29201,N_28796);
xor UO_1376 (O_1376,N_29271,N_29038);
and UO_1377 (O_1377,N_29515,N_29856);
nand UO_1378 (O_1378,N_28783,N_28968);
and UO_1379 (O_1379,N_28603,N_29099);
xor UO_1380 (O_1380,N_28589,N_29801);
nor UO_1381 (O_1381,N_28977,N_28579);
nand UO_1382 (O_1382,N_28638,N_29689);
nand UO_1383 (O_1383,N_28593,N_29537);
xor UO_1384 (O_1384,N_29415,N_29289);
nor UO_1385 (O_1385,N_29737,N_28948);
or UO_1386 (O_1386,N_29399,N_28598);
nand UO_1387 (O_1387,N_29368,N_29619);
or UO_1388 (O_1388,N_28865,N_28504);
nand UO_1389 (O_1389,N_29311,N_29490);
or UO_1390 (O_1390,N_29985,N_28548);
nor UO_1391 (O_1391,N_29786,N_29208);
nand UO_1392 (O_1392,N_28713,N_29580);
xnor UO_1393 (O_1393,N_28805,N_28532);
nand UO_1394 (O_1394,N_29858,N_29233);
nor UO_1395 (O_1395,N_28974,N_29249);
nor UO_1396 (O_1396,N_29804,N_28899);
xnor UO_1397 (O_1397,N_29777,N_28749);
or UO_1398 (O_1398,N_29864,N_29771);
nor UO_1399 (O_1399,N_29709,N_29978);
nor UO_1400 (O_1400,N_29354,N_28695);
or UO_1401 (O_1401,N_29161,N_29680);
nand UO_1402 (O_1402,N_29235,N_29225);
or UO_1403 (O_1403,N_29461,N_29109);
nand UO_1404 (O_1404,N_28543,N_29169);
nand UO_1405 (O_1405,N_29001,N_29206);
or UO_1406 (O_1406,N_29811,N_28752);
or UO_1407 (O_1407,N_29549,N_29616);
or UO_1408 (O_1408,N_29863,N_29524);
and UO_1409 (O_1409,N_29986,N_28881);
or UO_1410 (O_1410,N_29771,N_28778);
and UO_1411 (O_1411,N_29501,N_29181);
xor UO_1412 (O_1412,N_29673,N_29135);
and UO_1413 (O_1413,N_28742,N_29840);
and UO_1414 (O_1414,N_29063,N_29889);
nor UO_1415 (O_1415,N_29836,N_29973);
and UO_1416 (O_1416,N_29793,N_29268);
nor UO_1417 (O_1417,N_28800,N_29498);
nor UO_1418 (O_1418,N_28515,N_29723);
xor UO_1419 (O_1419,N_29135,N_28839);
and UO_1420 (O_1420,N_29893,N_28630);
xor UO_1421 (O_1421,N_29390,N_29496);
nor UO_1422 (O_1422,N_29093,N_29774);
or UO_1423 (O_1423,N_28796,N_28834);
nor UO_1424 (O_1424,N_28926,N_29680);
or UO_1425 (O_1425,N_28666,N_29821);
xnor UO_1426 (O_1426,N_29583,N_29618);
or UO_1427 (O_1427,N_29637,N_28693);
xor UO_1428 (O_1428,N_28750,N_28804);
nand UO_1429 (O_1429,N_29126,N_28897);
xor UO_1430 (O_1430,N_29584,N_28604);
or UO_1431 (O_1431,N_28742,N_29263);
and UO_1432 (O_1432,N_28569,N_28978);
nand UO_1433 (O_1433,N_29104,N_28546);
nand UO_1434 (O_1434,N_29277,N_29425);
nand UO_1435 (O_1435,N_29254,N_29086);
or UO_1436 (O_1436,N_29227,N_29566);
and UO_1437 (O_1437,N_29925,N_28752);
xor UO_1438 (O_1438,N_29493,N_28579);
and UO_1439 (O_1439,N_29276,N_29241);
and UO_1440 (O_1440,N_28544,N_29446);
or UO_1441 (O_1441,N_28693,N_29607);
or UO_1442 (O_1442,N_29226,N_29258);
and UO_1443 (O_1443,N_29273,N_29328);
and UO_1444 (O_1444,N_29292,N_29859);
nor UO_1445 (O_1445,N_29914,N_29647);
nor UO_1446 (O_1446,N_29156,N_29605);
nor UO_1447 (O_1447,N_28882,N_29320);
nor UO_1448 (O_1448,N_29414,N_28547);
nand UO_1449 (O_1449,N_28621,N_29265);
and UO_1450 (O_1450,N_29168,N_29635);
nand UO_1451 (O_1451,N_28818,N_29584);
xnor UO_1452 (O_1452,N_29715,N_29156);
xor UO_1453 (O_1453,N_29945,N_28676);
and UO_1454 (O_1454,N_28886,N_29780);
nor UO_1455 (O_1455,N_29058,N_29304);
nor UO_1456 (O_1456,N_28691,N_29463);
xnor UO_1457 (O_1457,N_29146,N_28543);
and UO_1458 (O_1458,N_29637,N_29069);
and UO_1459 (O_1459,N_29338,N_29852);
xnor UO_1460 (O_1460,N_28875,N_29581);
or UO_1461 (O_1461,N_29444,N_28582);
and UO_1462 (O_1462,N_29910,N_29544);
or UO_1463 (O_1463,N_29576,N_28639);
nand UO_1464 (O_1464,N_28916,N_28507);
nor UO_1465 (O_1465,N_29143,N_29831);
xnor UO_1466 (O_1466,N_29367,N_29458);
nand UO_1467 (O_1467,N_29128,N_28665);
nand UO_1468 (O_1468,N_29135,N_29468);
and UO_1469 (O_1469,N_29880,N_29886);
or UO_1470 (O_1470,N_28791,N_28762);
nor UO_1471 (O_1471,N_28535,N_28899);
nor UO_1472 (O_1472,N_29504,N_29808);
and UO_1473 (O_1473,N_29957,N_29137);
nand UO_1474 (O_1474,N_29554,N_28921);
or UO_1475 (O_1475,N_29389,N_28526);
nand UO_1476 (O_1476,N_28541,N_28883);
nor UO_1477 (O_1477,N_29657,N_29069);
or UO_1478 (O_1478,N_29455,N_29201);
nor UO_1479 (O_1479,N_29736,N_29599);
nor UO_1480 (O_1480,N_28942,N_29415);
or UO_1481 (O_1481,N_29559,N_29134);
or UO_1482 (O_1482,N_29477,N_29806);
nand UO_1483 (O_1483,N_29602,N_29351);
nor UO_1484 (O_1484,N_29025,N_29024);
and UO_1485 (O_1485,N_28593,N_28562);
and UO_1486 (O_1486,N_28831,N_29756);
or UO_1487 (O_1487,N_29946,N_29224);
xor UO_1488 (O_1488,N_28584,N_29032);
or UO_1489 (O_1489,N_28800,N_29465);
or UO_1490 (O_1490,N_29857,N_28752);
and UO_1491 (O_1491,N_29615,N_29430);
xnor UO_1492 (O_1492,N_28780,N_29252);
xor UO_1493 (O_1493,N_29044,N_29104);
nor UO_1494 (O_1494,N_29244,N_29246);
xnor UO_1495 (O_1495,N_29778,N_28860);
or UO_1496 (O_1496,N_29818,N_29985);
nor UO_1497 (O_1497,N_28805,N_28958);
nor UO_1498 (O_1498,N_29394,N_28933);
xnor UO_1499 (O_1499,N_29026,N_29671);
and UO_1500 (O_1500,N_28636,N_28528);
and UO_1501 (O_1501,N_29540,N_28539);
and UO_1502 (O_1502,N_29188,N_29616);
and UO_1503 (O_1503,N_29100,N_28901);
and UO_1504 (O_1504,N_28526,N_29367);
nor UO_1505 (O_1505,N_29123,N_29308);
and UO_1506 (O_1506,N_29816,N_28692);
nand UO_1507 (O_1507,N_28696,N_28773);
nor UO_1508 (O_1508,N_28810,N_29244);
and UO_1509 (O_1509,N_28849,N_28571);
and UO_1510 (O_1510,N_29648,N_28758);
and UO_1511 (O_1511,N_29345,N_28568);
or UO_1512 (O_1512,N_28923,N_29571);
xnor UO_1513 (O_1513,N_29408,N_28737);
nor UO_1514 (O_1514,N_29953,N_29092);
nand UO_1515 (O_1515,N_28982,N_28718);
nand UO_1516 (O_1516,N_28590,N_28829);
and UO_1517 (O_1517,N_29477,N_28563);
nand UO_1518 (O_1518,N_29714,N_28567);
and UO_1519 (O_1519,N_29838,N_29935);
xor UO_1520 (O_1520,N_28909,N_29142);
nor UO_1521 (O_1521,N_29193,N_29783);
nand UO_1522 (O_1522,N_28990,N_29241);
nor UO_1523 (O_1523,N_29190,N_29875);
and UO_1524 (O_1524,N_28828,N_29412);
or UO_1525 (O_1525,N_28899,N_28724);
and UO_1526 (O_1526,N_28631,N_29201);
xnor UO_1527 (O_1527,N_29626,N_28819);
or UO_1528 (O_1528,N_29966,N_28940);
or UO_1529 (O_1529,N_29967,N_29040);
and UO_1530 (O_1530,N_29740,N_29530);
and UO_1531 (O_1531,N_29140,N_29625);
xnor UO_1532 (O_1532,N_29659,N_29151);
and UO_1533 (O_1533,N_28652,N_29233);
nand UO_1534 (O_1534,N_29829,N_28633);
or UO_1535 (O_1535,N_29273,N_29074);
nor UO_1536 (O_1536,N_28581,N_28899);
or UO_1537 (O_1537,N_29423,N_29318);
xor UO_1538 (O_1538,N_29678,N_29724);
xor UO_1539 (O_1539,N_28642,N_29639);
or UO_1540 (O_1540,N_28794,N_28551);
xor UO_1541 (O_1541,N_29286,N_29364);
and UO_1542 (O_1542,N_28974,N_29752);
or UO_1543 (O_1543,N_28565,N_29754);
nand UO_1544 (O_1544,N_28528,N_29906);
and UO_1545 (O_1545,N_29200,N_29434);
nand UO_1546 (O_1546,N_29791,N_29584);
nand UO_1547 (O_1547,N_28671,N_29252);
nor UO_1548 (O_1548,N_28677,N_28504);
xnor UO_1549 (O_1549,N_28516,N_29664);
and UO_1550 (O_1550,N_28621,N_28732);
nor UO_1551 (O_1551,N_28628,N_29260);
and UO_1552 (O_1552,N_29673,N_28613);
nand UO_1553 (O_1553,N_28580,N_29450);
nor UO_1554 (O_1554,N_29185,N_29831);
and UO_1555 (O_1555,N_28578,N_29066);
and UO_1556 (O_1556,N_28558,N_29946);
nand UO_1557 (O_1557,N_29769,N_29348);
or UO_1558 (O_1558,N_29137,N_29427);
nand UO_1559 (O_1559,N_28639,N_28539);
xor UO_1560 (O_1560,N_29081,N_28912);
or UO_1561 (O_1561,N_29152,N_29154);
nor UO_1562 (O_1562,N_29012,N_29260);
xor UO_1563 (O_1563,N_28698,N_29495);
nand UO_1564 (O_1564,N_29160,N_29862);
and UO_1565 (O_1565,N_28643,N_29951);
and UO_1566 (O_1566,N_29725,N_28673);
and UO_1567 (O_1567,N_29442,N_29559);
nand UO_1568 (O_1568,N_29552,N_28595);
xnor UO_1569 (O_1569,N_29586,N_29818);
nor UO_1570 (O_1570,N_28968,N_28924);
nor UO_1571 (O_1571,N_29699,N_29100);
xor UO_1572 (O_1572,N_29181,N_29803);
and UO_1573 (O_1573,N_29130,N_29147);
nor UO_1574 (O_1574,N_28983,N_28725);
nor UO_1575 (O_1575,N_29415,N_29845);
nor UO_1576 (O_1576,N_29611,N_29325);
and UO_1577 (O_1577,N_29527,N_29949);
nand UO_1578 (O_1578,N_29063,N_28557);
nor UO_1579 (O_1579,N_28678,N_28740);
and UO_1580 (O_1580,N_29533,N_28945);
or UO_1581 (O_1581,N_28501,N_29369);
and UO_1582 (O_1582,N_28661,N_29595);
or UO_1583 (O_1583,N_28998,N_28692);
nand UO_1584 (O_1584,N_28961,N_28942);
and UO_1585 (O_1585,N_28508,N_29408);
xnor UO_1586 (O_1586,N_29932,N_29027);
xor UO_1587 (O_1587,N_29594,N_29733);
nand UO_1588 (O_1588,N_29149,N_29918);
xnor UO_1589 (O_1589,N_29883,N_29540);
nor UO_1590 (O_1590,N_29982,N_28503);
xor UO_1591 (O_1591,N_29055,N_28909);
and UO_1592 (O_1592,N_28675,N_28573);
and UO_1593 (O_1593,N_28629,N_28789);
nor UO_1594 (O_1594,N_29352,N_28560);
xnor UO_1595 (O_1595,N_29716,N_29670);
and UO_1596 (O_1596,N_29844,N_29291);
xnor UO_1597 (O_1597,N_28616,N_29781);
or UO_1598 (O_1598,N_29929,N_29681);
nand UO_1599 (O_1599,N_29479,N_28818);
or UO_1600 (O_1600,N_29467,N_28717);
and UO_1601 (O_1601,N_29030,N_29593);
xor UO_1602 (O_1602,N_29433,N_28538);
nand UO_1603 (O_1603,N_29040,N_28889);
or UO_1604 (O_1604,N_29658,N_29242);
nor UO_1605 (O_1605,N_29930,N_29912);
nor UO_1606 (O_1606,N_28906,N_28931);
nand UO_1607 (O_1607,N_29339,N_29976);
nand UO_1608 (O_1608,N_29480,N_29856);
or UO_1609 (O_1609,N_29328,N_29391);
nand UO_1610 (O_1610,N_29725,N_29386);
xor UO_1611 (O_1611,N_29540,N_29304);
xnor UO_1612 (O_1612,N_28878,N_29060);
and UO_1613 (O_1613,N_28634,N_29648);
nand UO_1614 (O_1614,N_29530,N_29903);
xnor UO_1615 (O_1615,N_29023,N_28577);
or UO_1616 (O_1616,N_29935,N_29705);
or UO_1617 (O_1617,N_28563,N_28966);
nor UO_1618 (O_1618,N_29523,N_29894);
nor UO_1619 (O_1619,N_29150,N_28567);
or UO_1620 (O_1620,N_28692,N_28559);
nand UO_1621 (O_1621,N_28812,N_29988);
and UO_1622 (O_1622,N_28840,N_29375);
or UO_1623 (O_1623,N_29547,N_28742);
nand UO_1624 (O_1624,N_29637,N_28906);
nor UO_1625 (O_1625,N_28780,N_28983);
nand UO_1626 (O_1626,N_29374,N_29237);
and UO_1627 (O_1627,N_29728,N_29345);
nand UO_1628 (O_1628,N_29284,N_29478);
xnor UO_1629 (O_1629,N_28997,N_28570);
and UO_1630 (O_1630,N_29952,N_29764);
nand UO_1631 (O_1631,N_29992,N_29274);
nand UO_1632 (O_1632,N_28967,N_29527);
xnor UO_1633 (O_1633,N_28589,N_29188);
or UO_1634 (O_1634,N_29581,N_29614);
xor UO_1635 (O_1635,N_29862,N_29258);
and UO_1636 (O_1636,N_28802,N_29177);
and UO_1637 (O_1637,N_29777,N_28587);
nor UO_1638 (O_1638,N_28937,N_28902);
xnor UO_1639 (O_1639,N_28598,N_29024);
or UO_1640 (O_1640,N_29057,N_29557);
or UO_1641 (O_1641,N_29509,N_28985);
nand UO_1642 (O_1642,N_29807,N_29733);
or UO_1643 (O_1643,N_29207,N_29037);
and UO_1644 (O_1644,N_28685,N_28888);
nand UO_1645 (O_1645,N_29652,N_29822);
nor UO_1646 (O_1646,N_29640,N_29497);
xnor UO_1647 (O_1647,N_29399,N_29658);
nand UO_1648 (O_1648,N_29424,N_29058);
nand UO_1649 (O_1649,N_28548,N_29894);
and UO_1650 (O_1650,N_29946,N_29896);
or UO_1651 (O_1651,N_29464,N_29658);
and UO_1652 (O_1652,N_29562,N_29491);
nor UO_1653 (O_1653,N_29606,N_28865);
xnor UO_1654 (O_1654,N_29692,N_29538);
and UO_1655 (O_1655,N_28904,N_29089);
nor UO_1656 (O_1656,N_29365,N_28993);
xor UO_1657 (O_1657,N_29619,N_29266);
and UO_1658 (O_1658,N_29258,N_29208);
nand UO_1659 (O_1659,N_29481,N_29068);
or UO_1660 (O_1660,N_29066,N_29877);
nor UO_1661 (O_1661,N_29819,N_29334);
and UO_1662 (O_1662,N_29953,N_28699);
nor UO_1663 (O_1663,N_28535,N_29676);
nand UO_1664 (O_1664,N_29483,N_29604);
or UO_1665 (O_1665,N_29820,N_29518);
and UO_1666 (O_1666,N_28598,N_29706);
xor UO_1667 (O_1667,N_28777,N_29199);
and UO_1668 (O_1668,N_28767,N_29734);
xnor UO_1669 (O_1669,N_29524,N_29859);
xnor UO_1670 (O_1670,N_29966,N_28543);
nor UO_1671 (O_1671,N_29939,N_28854);
or UO_1672 (O_1672,N_29199,N_29520);
or UO_1673 (O_1673,N_28764,N_29968);
nand UO_1674 (O_1674,N_28553,N_28992);
xnor UO_1675 (O_1675,N_29838,N_29351);
and UO_1676 (O_1676,N_29746,N_29189);
nor UO_1677 (O_1677,N_29381,N_28542);
or UO_1678 (O_1678,N_29613,N_28711);
or UO_1679 (O_1679,N_29024,N_28937);
nand UO_1680 (O_1680,N_29737,N_28766);
or UO_1681 (O_1681,N_29697,N_28721);
and UO_1682 (O_1682,N_29499,N_29039);
nor UO_1683 (O_1683,N_29088,N_29863);
xor UO_1684 (O_1684,N_29933,N_28624);
and UO_1685 (O_1685,N_29210,N_28888);
or UO_1686 (O_1686,N_29146,N_29394);
nand UO_1687 (O_1687,N_29772,N_29650);
xnor UO_1688 (O_1688,N_29915,N_29156);
and UO_1689 (O_1689,N_29591,N_29852);
xor UO_1690 (O_1690,N_29844,N_29551);
nor UO_1691 (O_1691,N_29365,N_29679);
nor UO_1692 (O_1692,N_29526,N_29986);
xnor UO_1693 (O_1693,N_29738,N_28782);
or UO_1694 (O_1694,N_29804,N_29078);
or UO_1695 (O_1695,N_29067,N_29235);
nand UO_1696 (O_1696,N_29897,N_29571);
nor UO_1697 (O_1697,N_29639,N_28711);
xnor UO_1698 (O_1698,N_29218,N_28658);
nor UO_1699 (O_1699,N_29626,N_29916);
nor UO_1700 (O_1700,N_29558,N_28507);
and UO_1701 (O_1701,N_29461,N_28683);
nand UO_1702 (O_1702,N_29878,N_29856);
or UO_1703 (O_1703,N_28557,N_28903);
xnor UO_1704 (O_1704,N_28530,N_29410);
xnor UO_1705 (O_1705,N_28787,N_29207);
nand UO_1706 (O_1706,N_29409,N_29754);
or UO_1707 (O_1707,N_28764,N_29692);
or UO_1708 (O_1708,N_29234,N_29302);
nor UO_1709 (O_1709,N_29420,N_28970);
and UO_1710 (O_1710,N_29176,N_29107);
or UO_1711 (O_1711,N_28829,N_28791);
nor UO_1712 (O_1712,N_29962,N_28583);
xor UO_1713 (O_1713,N_29470,N_28610);
nor UO_1714 (O_1714,N_29466,N_29464);
or UO_1715 (O_1715,N_29269,N_28718);
xor UO_1716 (O_1716,N_29911,N_29625);
nand UO_1717 (O_1717,N_28568,N_29927);
nor UO_1718 (O_1718,N_29081,N_29356);
xnor UO_1719 (O_1719,N_28500,N_29772);
and UO_1720 (O_1720,N_28596,N_29269);
nand UO_1721 (O_1721,N_29818,N_29117);
nand UO_1722 (O_1722,N_29877,N_28732);
nand UO_1723 (O_1723,N_29217,N_29247);
xor UO_1724 (O_1724,N_29712,N_29871);
nor UO_1725 (O_1725,N_29543,N_28966);
or UO_1726 (O_1726,N_29397,N_28912);
nand UO_1727 (O_1727,N_29647,N_29877);
nor UO_1728 (O_1728,N_28677,N_28643);
nand UO_1729 (O_1729,N_29473,N_28744);
or UO_1730 (O_1730,N_29143,N_28682);
and UO_1731 (O_1731,N_28616,N_29459);
nand UO_1732 (O_1732,N_28816,N_29451);
and UO_1733 (O_1733,N_29751,N_29218);
nor UO_1734 (O_1734,N_29238,N_29626);
xnor UO_1735 (O_1735,N_28524,N_29513);
xnor UO_1736 (O_1736,N_28570,N_29574);
nor UO_1737 (O_1737,N_29435,N_29609);
or UO_1738 (O_1738,N_29235,N_29282);
or UO_1739 (O_1739,N_29973,N_28764);
xnor UO_1740 (O_1740,N_29995,N_28950);
or UO_1741 (O_1741,N_29021,N_29207);
xnor UO_1742 (O_1742,N_29936,N_28795);
nor UO_1743 (O_1743,N_29605,N_29135);
nor UO_1744 (O_1744,N_29843,N_28950);
or UO_1745 (O_1745,N_29397,N_28767);
nand UO_1746 (O_1746,N_29674,N_29663);
or UO_1747 (O_1747,N_29301,N_28605);
nand UO_1748 (O_1748,N_29968,N_29952);
or UO_1749 (O_1749,N_29089,N_29854);
nor UO_1750 (O_1750,N_29246,N_29518);
nand UO_1751 (O_1751,N_29800,N_29267);
nor UO_1752 (O_1752,N_28967,N_28774);
xnor UO_1753 (O_1753,N_29929,N_28539);
nand UO_1754 (O_1754,N_28665,N_28803);
or UO_1755 (O_1755,N_29716,N_28662);
nand UO_1756 (O_1756,N_28714,N_28993);
nor UO_1757 (O_1757,N_29080,N_28803);
nand UO_1758 (O_1758,N_29100,N_29786);
or UO_1759 (O_1759,N_29126,N_29421);
nor UO_1760 (O_1760,N_28851,N_29242);
xor UO_1761 (O_1761,N_29858,N_28605);
nor UO_1762 (O_1762,N_29710,N_29571);
nor UO_1763 (O_1763,N_29473,N_28867);
xnor UO_1764 (O_1764,N_28739,N_28652);
or UO_1765 (O_1765,N_29421,N_29525);
and UO_1766 (O_1766,N_28658,N_28976);
and UO_1767 (O_1767,N_29829,N_29450);
nand UO_1768 (O_1768,N_28585,N_29320);
nand UO_1769 (O_1769,N_29681,N_28559);
and UO_1770 (O_1770,N_29225,N_28815);
nand UO_1771 (O_1771,N_28693,N_29752);
and UO_1772 (O_1772,N_28735,N_28559);
or UO_1773 (O_1773,N_29592,N_28710);
and UO_1774 (O_1774,N_29455,N_28801);
or UO_1775 (O_1775,N_29583,N_28776);
and UO_1776 (O_1776,N_29328,N_29389);
or UO_1777 (O_1777,N_28615,N_29921);
and UO_1778 (O_1778,N_28637,N_29787);
or UO_1779 (O_1779,N_29213,N_29943);
xor UO_1780 (O_1780,N_28944,N_28911);
xnor UO_1781 (O_1781,N_29667,N_29620);
and UO_1782 (O_1782,N_29487,N_28598);
nor UO_1783 (O_1783,N_29803,N_28687);
nor UO_1784 (O_1784,N_28853,N_28505);
nor UO_1785 (O_1785,N_29706,N_28984);
or UO_1786 (O_1786,N_29100,N_29298);
and UO_1787 (O_1787,N_28600,N_29754);
nor UO_1788 (O_1788,N_29363,N_28720);
xnor UO_1789 (O_1789,N_28816,N_28864);
nand UO_1790 (O_1790,N_29533,N_29306);
xnor UO_1791 (O_1791,N_29291,N_29963);
or UO_1792 (O_1792,N_28576,N_29746);
nand UO_1793 (O_1793,N_29947,N_29799);
and UO_1794 (O_1794,N_29849,N_29062);
or UO_1795 (O_1795,N_29374,N_29950);
nor UO_1796 (O_1796,N_28750,N_29743);
nor UO_1797 (O_1797,N_29252,N_29839);
or UO_1798 (O_1798,N_29867,N_29359);
xor UO_1799 (O_1799,N_29372,N_29900);
or UO_1800 (O_1800,N_29768,N_29536);
xor UO_1801 (O_1801,N_29384,N_28734);
or UO_1802 (O_1802,N_29432,N_28945);
nor UO_1803 (O_1803,N_28907,N_29648);
nand UO_1804 (O_1804,N_28522,N_29180);
and UO_1805 (O_1805,N_29091,N_28625);
or UO_1806 (O_1806,N_29813,N_29090);
nor UO_1807 (O_1807,N_29718,N_28675);
and UO_1808 (O_1808,N_29284,N_29499);
nand UO_1809 (O_1809,N_29301,N_28762);
and UO_1810 (O_1810,N_29660,N_28963);
or UO_1811 (O_1811,N_29194,N_29579);
xnor UO_1812 (O_1812,N_29002,N_29584);
xor UO_1813 (O_1813,N_29845,N_28874);
or UO_1814 (O_1814,N_28551,N_29853);
xor UO_1815 (O_1815,N_29246,N_28699);
or UO_1816 (O_1816,N_29979,N_29362);
xor UO_1817 (O_1817,N_28855,N_28688);
and UO_1818 (O_1818,N_29891,N_28545);
or UO_1819 (O_1819,N_29590,N_28528);
nand UO_1820 (O_1820,N_29425,N_29866);
nand UO_1821 (O_1821,N_29141,N_29907);
or UO_1822 (O_1822,N_29768,N_28928);
nand UO_1823 (O_1823,N_28500,N_29735);
nand UO_1824 (O_1824,N_29074,N_29562);
nand UO_1825 (O_1825,N_29014,N_29774);
or UO_1826 (O_1826,N_28607,N_28510);
or UO_1827 (O_1827,N_28867,N_29416);
xor UO_1828 (O_1828,N_29647,N_29567);
or UO_1829 (O_1829,N_29701,N_29186);
or UO_1830 (O_1830,N_28541,N_28698);
nand UO_1831 (O_1831,N_28803,N_29221);
and UO_1832 (O_1832,N_29815,N_29449);
nand UO_1833 (O_1833,N_29123,N_29881);
nand UO_1834 (O_1834,N_28930,N_29173);
nand UO_1835 (O_1835,N_29608,N_28646);
or UO_1836 (O_1836,N_28973,N_29112);
xor UO_1837 (O_1837,N_29222,N_29402);
nand UO_1838 (O_1838,N_28895,N_28861);
nor UO_1839 (O_1839,N_28806,N_29648);
and UO_1840 (O_1840,N_29893,N_28779);
and UO_1841 (O_1841,N_28921,N_29019);
or UO_1842 (O_1842,N_29689,N_28502);
and UO_1843 (O_1843,N_29918,N_29223);
xnor UO_1844 (O_1844,N_28739,N_28672);
or UO_1845 (O_1845,N_28951,N_28892);
nand UO_1846 (O_1846,N_29747,N_28989);
nand UO_1847 (O_1847,N_29677,N_29644);
or UO_1848 (O_1848,N_29386,N_28613);
xor UO_1849 (O_1849,N_29888,N_29756);
nand UO_1850 (O_1850,N_29243,N_29861);
nand UO_1851 (O_1851,N_28704,N_29179);
nor UO_1852 (O_1852,N_29690,N_29853);
nand UO_1853 (O_1853,N_29159,N_29301);
or UO_1854 (O_1854,N_29753,N_29974);
or UO_1855 (O_1855,N_29777,N_29275);
nor UO_1856 (O_1856,N_28560,N_29569);
and UO_1857 (O_1857,N_29852,N_29022);
nor UO_1858 (O_1858,N_28580,N_28873);
and UO_1859 (O_1859,N_28609,N_29319);
nand UO_1860 (O_1860,N_29863,N_29666);
nand UO_1861 (O_1861,N_28530,N_28737);
nand UO_1862 (O_1862,N_29704,N_29748);
nand UO_1863 (O_1863,N_29638,N_28998);
and UO_1864 (O_1864,N_29104,N_29167);
or UO_1865 (O_1865,N_29448,N_28593);
nor UO_1866 (O_1866,N_29659,N_29981);
nor UO_1867 (O_1867,N_29966,N_29571);
xnor UO_1868 (O_1868,N_28806,N_29701);
and UO_1869 (O_1869,N_29449,N_29245);
nand UO_1870 (O_1870,N_29345,N_29933);
and UO_1871 (O_1871,N_28538,N_29157);
xnor UO_1872 (O_1872,N_28715,N_29377);
or UO_1873 (O_1873,N_29931,N_29654);
xnor UO_1874 (O_1874,N_29336,N_29487);
or UO_1875 (O_1875,N_29847,N_29708);
nor UO_1876 (O_1876,N_29692,N_29466);
nand UO_1877 (O_1877,N_29981,N_29157);
nand UO_1878 (O_1878,N_29858,N_29388);
xor UO_1879 (O_1879,N_29417,N_28863);
nor UO_1880 (O_1880,N_29418,N_28923);
nor UO_1881 (O_1881,N_29758,N_28875);
or UO_1882 (O_1882,N_28963,N_29943);
nor UO_1883 (O_1883,N_28861,N_29093);
xnor UO_1884 (O_1884,N_29651,N_28660);
nand UO_1885 (O_1885,N_29572,N_29440);
xor UO_1886 (O_1886,N_29825,N_29014);
nor UO_1887 (O_1887,N_29551,N_28999);
nor UO_1888 (O_1888,N_28761,N_29401);
and UO_1889 (O_1889,N_28544,N_28796);
nor UO_1890 (O_1890,N_28986,N_29528);
nor UO_1891 (O_1891,N_29747,N_29488);
and UO_1892 (O_1892,N_28794,N_29148);
and UO_1893 (O_1893,N_29748,N_28623);
nor UO_1894 (O_1894,N_29279,N_28988);
nor UO_1895 (O_1895,N_29675,N_29212);
and UO_1896 (O_1896,N_29188,N_29768);
nand UO_1897 (O_1897,N_29961,N_29522);
nor UO_1898 (O_1898,N_28757,N_29104);
and UO_1899 (O_1899,N_28854,N_28532);
nand UO_1900 (O_1900,N_28986,N_29683);
nor UO_1901 (O_1901,N_29447,N_28526);
or UO_1902 (O_1902,N_29833,N_29428);
or UO_1903 (O_1903,N_29980,N_29426);
nor UO_1904 (O_1904,N_28945,N_28957);
nand UO_1905 (O_1905,N_29935,N_29716);
or UO_1906 (O_1906,N_29110,N_28741);
nand UO_1907 (O_1907,N_29274,N_29887);
and UO_1908 (O_1908,N_29037,N_28951);
nor UO_1909 (O_1909,N_29907,N_28502);
xor UO_1910 (O_1910,N_29769,N_29775);
nor UO_1911 (O_1911,N_29009,N_29457);
xor UO_1912 (O_1912,N_28857,N_28626);
nand UO_1913 (O_1913,N_28985,N_29369);
or UO_1914 (O_1914,N_29274,N_28832);
xnor UO_1915 (O_1915,N_28600,N_29999);
nor UO_1916 (O_1916,N_28649,N_29422);
xnor UO_1917 (O_1917,N_29568,N_29758);
and UO_1918 (O_1918,N_28687,N_28603);
nand UO_1919 (O_1919,N_28781,N_29395);
xor UO_1920 (O_1920,N_29658,N_28532);
nand UO_1921 (O_1921,N_29652,N_29925);
and UO_1922 (O_1922,N_28680,N_29612);
or UO_1923 (O_1923,N_28998,N_28586);
nand UO_1924 (O_1924,N_28799,N_28599);
nand UO_1925 (O_1925,N_29802,N_28711);
xnor UO_1926 (O_1926,N_29265,N_29784);
xor UO_1927 (O_1927,N_29096,N_28636);
or UO_1928 (O_1928,N_29473,N_29979);
nand UO_1929 (O_1929,N_29411,N_29205);
xnor UO_1930 (O_1930,N_28528,N_29229);
or UO_1931 (O_1931,N_28523,N_29669);
nor UO_1932 (O_1932,N_29974,N_29118);
nor UO_1933 (O_1933,N_29619,N_28796);
nor UO_1934 (O_1934,N_29382,N_29710);
or UO_1935 (O_1935,N_29308,N_29085);
xnor UO_1936 (O_1936,N_29576,N_29072);
xor UO_1937 (O_1937,N_28739,N_29492);
or UO_1938 (O_1938,N_29338,N_29111);
and UO_1939 (O_1939,N_29382,N_28575);
nand UO_1940 (O_1940,N_29781,N_29201);
nor UO_1941 (O_1941,N_29218,N_29935);
nor UO_1942 (O_1942,N_28858,N_28905);
and UO_1943 (O_1943,N_29120,N_29206);
nand UO_1944 (O_1944,N_29077,N_28556);
nand UO_1945 (O_1945,N_28593,N_29009);
or UO_1946 (O_1946,N_29273,N_29765);
xor UO_1947 (O_1947,N_29204,N_29739);
nand UO_1948 (O_1948,N_29203,N_28895);
and UO_1949 (O_1949,N_28633,N_28822);
nor UO_1950 (O_1950,N_29227,N_29876);
and UO_1951 (O_1951,N_29430,N_29579);
nand UO_1952 (O_1952,N_29176,N_29123);
or UO_1953 (O_1953,N_28892,N_28971);
or UO_1954 (O_1954,N_29376,N_28674);
nand UO_1955 (O_1955,N_29901,N_29458);
nand UO_1956 (O_1956,N_29644,N_28923);
nand UO_1957 (O_1957,N_29861,N_29308);
and UO_1958 (O_1958,N_29496,N_28942);
nor UO_1959 (O_1959,N_28895,N_29193);
and UO_1960 (O_1960,N_29680,N_28574);
nand UO_1961 (O_1961,N_28902,N_29127);
or UO_1962 (O_1962,N_29658,N_29564);
xor UO_1963 (O_1963,N_29785,N_29067);
nor UO_1964 (O_1964,N_29664,N_29352);
and UO_1965 (O_1965,N_28653,N_29486);
nor UO_1966 (O_1966,N_28940,N_28531);
xor UO_1967 (O_1967,N_29984,N_28791);
or UO_1968 (O_1968,N_29242,N_29317);
and UO_1969 (O_1969,N_28565,N_29368);
or UO_1970 (O_1970,N_28946,N_28788);
nor UO_1971 (O_1971,N_29680,N_28962);
or UO_1972 (O_1972,N_29745,N_29141);
and UO_1973 (O_1973,N_29962,N_29482);
or UO_1974 (O_1974,N_28559,N_28912);
nor UO_1975 (O_1975,N_29314,N_28788);
xnor UO_1976 (O_1976,N_29207,N_29211);
xor UO_1977 (O_1977,N_29118,N_29619);
or UO_1978 (O_1978,N_28550,N_29745);
or UO_1979 (O_1979,N_28809,N_29449);
and UO_1980 (O_1980,N_29619,N_29089);
xor UO_1981 (O_1981,N_28612,N_28804);
nor UO_1982 (O_1982,N_29715,N_29972);
xnor UO_1983 (O_1983,N_29805,N_28601);
nand UO_1984 (O_1984,N_28608,N_29711);
nor UO_1985 (O_1985,N_29111,N_28752);
nand UO_1986 (O_1986,N_28600,N_29227);
nand UO_1987 (O_1987,N_29619,N_29847);
or UO_1988 (O_1988,N_29160,N_29062);
nor UO_1989 (O_1989,N_29992,N_29853);
and UO_1990 (O_1990,N_28719,N_28926);
or UO_1991 (O_1991,N_28521,N_29286);
nand UO_1992 (O_1992,N_28875,N_29612);
and UO_1993 (O_1993,N_29964,N_29844);
nor UO_1994 (O_1994,N_29028,N_28905);
nand UO_1995 (O_1995,N_28945,N_29028);
or UO_1996 (O_1996,N_28595,N_29309);
xnor UO_1997 (O_1997,N_28899,N_29529);
xnor UO_1998 (O_1998,N_28903,N_29909);
xor UO_1999 (O_1999,N_29849,N_28680);
nand UO_2000 (O_2000,N_29518,N_29232);
xnor UO_2001 (O_2001,N_29993,N_29695);
or UO_2002 (O_2002,N_28852,N_29334);
or UO_2003 (O_2003,N_29495,N_29590);
nor UO_2004 (O_2004,N_29245,N_28641);
xor UO_2005 (O_2005,N_28576,N_29110);
or UO_2006 (O_2006,N_28919,N_29827);
or UO_2007 (O_2007,N_28592,N_29044);
and UO_2008 (O_2008,N_28574,N_28547);
nor UO_2009 (O_2009,N_29174,N_29659);
nor UO_2010 (O_2010,N_28974,N_29352);
nand UO_2011 (O_2011,N_29264,N_28649);
or UO_2012 (O_2012,N_28607,N_29430);
and UO_2013 (O_2013,N_29670,N_29759);
xor UO_2014 (O_2014,N_28949,N_28895);
nand UO_2015 (O_2015,N_29152,N_29765);
nor UO_2016 (O_2016,N_29783,N_29813);
nand UO_2017 (O_2017,N_29383,N_29430);
nand UO_2018 (O_2018,N_29138,N_29135);
or UO_2019 (O_2019,N_29181,N_29180);
nand UO_2020 (O_2020,N_28570,N_29609);
xor UO_2021 (O_2021,N_28974,N_29537);
and UO_2022 (O_2022,N_29933,N_29378);
nand UO_2023 (O_2023,N_29113,N_28549);
nand UO_2024 (O_2024,N_28623,N_29740);
nand UO_2025 (O_2025,N_29925,N_28817);
and UO_2026 (O_2026,N_29120,N_28913);
xnor UO_2027 (O_2027,N_29689,N_29280);
and UO_2028 (O_2028,N_28819,N_29912);
or UO_2029 (O_2029,N_29617,N_28605);
and UO_2030 (O_2030,N_28983,N_29791);
nand UO_2031 (O_2031,N_29000,N_29575);
nand UO_2032 (O_2032,N_28764,N_28709);
nand UO_2033 (O_2033,N_28546,N_28827);
xnor UO_2034 (O_2034,N_29066,N_28785);
or UO_2035 (O_2035,N_28634,N_29386);
or UO_2036 (O_2036,N_28549,N_29819);
or UO_2037 (O_2037,N_29344,N_28758);
and UO_2038 (O_2038,N_28601,N_29029);
or UO_2039 (O_2039,N_29425,N_28611);
and UO_2040 (O_2040,N_28684,N_28737);
and UO_2041 (O_2041,N_29153,N_29684);
nand UO_2042 (O_2042,N_29682,N_29966);
xnor UO_2043 (O_2043,N_29719,N_28657);
xnor UO_2044 (O_2044,N_29810,N_28729);
xnor UO_2045 (O_2045,N_28743,N_29732);
nor UO_2046 (O_2046,N_29862,N_29315);
or UO_2047 (O_2047,N_29737,N_29749);
or UO_2048 (O_2048,N_28647,N_29864);
or UO_2049 (O_2049,N_28605,N_28532);
nor UO_2050 (O_2050,N_29893,N_28584);
xnor UO_2051 (O_2051,N_28965,N_29078);
or UO_2052 (O_2052,N_29778,N_29418);
nand UO_2053 (O_2053,N_29333,N_29371);
nand UO_2054 (O_2054,N_29271,N_29974);
xnor UO_2055 (O_2055,N_29415,N_29900);
xnor UO_2056 (O_2056,N_28823,N_28800);
xnor UO_2057 (O_2057,N_29715,N_29803);
nor UO_2058 (O_2058,N_29960,N_29301);
nor UO_2059 (O_2059,N_29642,N_29765);
nand UO_2060 (O_2060,N_29230,N_29837);
xor UO_2061 (O_2061,N_29484,N_29137);
or UO_2062 (O_2062,N_29258,N_28668);
and UO_2063 (O_2063,N_29560,N_28735);
xor UO_2064 (O_2064,N_28608,N_29318);
nor UO_2065 (O_2065,N_28786,N_29799);
nor UO_2066 (O_2066,N_28839,N_29126);
and UO_2067 (O_2067,N_29072,N_29747);
and UO_2068 (O_2068,N_29198,N_29760);
or UO_2069 (O_2069,N_29627,N_29695);
or UO_2070 (O_2070,N_29992,N_28952);
xnor UO_2071 (O_2071,N_28858,N_29213);
or UO_2072 (O_2072,N_29443,N_29729);
nor UO_2073 (O_2073,N_28797,N_29712);
or UO_2074 (O_2074,N_28732,N_28504);
nor UO_2075 (O_2075,N_29564,N_28723);
and UO_2076 (O_2076,N_29556,N_29331);
or UO_2077 (O_2077,N_28684,N_28946);
and UO_2078 (O_2078,N_28848,N_29984);
and UO_2079 (O_2079,N_29576,N_29810);
and UO_2080 (O_2080,N_29140,N_29269);
nor UO_2081 (O_2081,N_29902,N_28828);
and UO_2082 (O_2082,N_29376,N_29253);
and UO_2083 (O_2083,N_29215,N_29225);
and UO_2084 (O_2084,N_28565,N_28521);
nand UO_2085 (O_2085,N_29434,N_29140);
nor UO_2086 (O_2086,N_29403,N_29654);
xor UO_2087 (O_2087,N_28970,N_29786);
and UO_2088 (O_2088,N_29765,N_29231);
and UO_2089 (O_2089,N_29253,N_28666);
and UO_2090 (O_2090,N_28624,N_29532);
or UO_2091 (O_2091,N_29168,N_29000);
nor UO_2092 (O_2092,N_29904,N_29651);
or UO_2093 (O_2093,N_29832,N_29764);
and UO_2094 (O_2094,N_28883,N_29123);
nor UO_2095 (O_2095,N_29101,N_29817);
and UO_2096 (O_2096,N_28522,N_29659);
or UO_2097 (O_2097,N_29791,N_29647);
nand UO_2098 (O_2098,N_29844,N_28715);
nand UO_2099 (O_2099,N_28655,N_29199);
nand UO_2100 (O_2100,N_28751,N_29279);
nor UO_2101 (O_2101,N_28734,N_29343);
nor UO_2102 (O_2102,N_29458,N_29456);
nand UO_2103 (O_2103,N_29769,N_29217);
nor UO_2104 (O_2104,N_29373,N_29076);
and UO_2105 (O_2105,N_28569,N_29045);
and UO_2106 (O_2106,N_29371,N_28724);
nor UO_2107 (O_2107,N_29287,N_28520);
nor UO_2108 (O_2108,N_28958,N_29793);
nor UO_2109 (O_2109,N_29055,N_29600);
and UO_2110 (O_2110,N_29422,N_28597);
nor UO_2111 (O_2111,N_29852,N_28929);
nand UO_2112 (O_2112,N_29095,N_29119);
xor UO_2113 (O_2113,N_28909,N_29849);
nand UO_2114 (O_2114,N_29856,N_29941);
xnor UO_2115 (O_2115,N_29406,N_29428);
and UO_2116 (O_2116,N_29660,N_28929);
nand UO_2117 (O_2117,N_29619,N_28522);
xor UO_2118 (O_2118,N_28556,N_29381);
or UO_2119 (O_2119,N_28906,N_29674);
xor UO_2120 (O_2120,N_29732,N_28591);
xor UO_2121 (O_2121,N_29957,N_28508);
xnor UO_2122 (O_2122,N_28650,N_29623);
and UO_2123 (O_2123,N_29219,N_29660);
or UO_2124 (O_2124,N_29724,N_29531);
and UO_2125 (O_2125,N_29356,N_28529);
and UO_2126 (O_2126,N_29046,N_29563);
nor UO_2127 (O_2127,N_28786,N_29140);
or UO_2128 (O_2128,N_29392,N_28587);
nand UO_2129 (O_2129,N_28864,N_29878);
xnor UO_2130 (O_2130,N_29626,N_29851);
nor UO_2131 (O_2131,N_29488,N_29677);
and UO_2132 (O_2132,N_28595,N_29274);
xor UO_2133 (O_2133,N_28938,N_29548);
xor UO_2134 (O_2134,N_29929,N_29321);
nor UO_2135 (O_2135,N_28618,N_28595);
nor UO_2136 (O_2136,N_28513,N_29420);
nand UO_2137 (O_2137,N_29374,N_29512);
nand UO_2138 (O_2138,N_29074,N_29836);
or UO_2139 (O_2139,N_29851,N_29355);
xnor UO_2140 (O_2140,N_29190,N_29802);
nor UO_2141 (O_2141,N_29787,N_28634);
xor UO_2142 (O_2142,N_29558,N_28505);
and UO_2143 (O_2143,N_28927,N_28521);
and UO_2144 (O_2144,N_29824,N_28935);
xnor UO_2145 (O_2145,N_29363,N_28517);
nand UO_2146 (O_2146,N_29995,N_29198);
nand UO_2147 (O_2147,N_29649,N_29828);
or UO_2148 (O_2148,N_29931,N_29507);
nand UO_2149 (O_2149,N_29088,N_29726);
xor UO_2150 (O_2150,N_29582,N_29276);
nand UO_2151 (O_2151,N_29136,N_28936);
or UO_2152 (O_2152,N_28719,N_28870);
or UO_2153 (O_2153,N_29235,N_29289);
xor UO_2154 (O_2154,N_28555,N_28986);
nor UO_2155 (O_2155,N_29656,N_29954);
xnor UO_2156 (O_2156,N_29773,N_29601);
xor UO_2157 (O_2157,N_29079,N_28958);
or UO_2158 (O_2158,N_29144,N_29691);
or UO_2159 (O_2159,N_29119,N_28668);
and UO_2160 (O_2160,N_28502,N_28656);
xnor UO_2161 (O_2161,N_28870,N_29313);
xnor UO_2162 (O_2162,N_28717,N_29001);
or UO_2163 (O_2163,N_28839,N_29199);
nor UO_2164 (O_2164,N_29058,N_29573);
nor UO_2165 (O_2165,N_29052,N_29975);
xnor UO_2166 (O_2166,N_29095,N_28529);
and UO_2167 (O_2167,N_28518,N_29688);
nor UO_2168 (O_2168,N_29954,N_28644);
xnor UO_2169 (O_2169,N_29687,N_29571);
xnor UO_2170 (O_2170,N_29970,N_29609);
nand UO_2171 (O_2171,N_29009,N_28881);
nand UO_2172 (O_2172,N_29703,N_29699);
nor UO_2173 (O_2173,N_29225,N_29264);
and UO_2174 (O_2174,N_29304,N_28602);
or UO_2175 (O_2175,N_29579,N_29328);
and UO_2176 (O_2176,N_29602,N_29969);
or UO_2177 (O_2177,N_29730,N_29514);
nand UO_2178 (O_2178,N_28798,N_28628);
and UO_2179 (O_2179,N_29501,N_29710);
and UO_2180 (O_2180,N_29988,N_28814);
or UO_2181 (O_2181,N_29144,N_29556);
xnor UO_2182 (O_2182,N_28689,N_28922);
nand UO_2183 (O_2183,N_29216,N_29110);
nor UO_2184 (O_2184,N_29687,N_28586);
nand UO_2185 (O_2185,N_29337,N_29107);
or UO_2186 (O_2186,N_29957,N_29615);
nor UO_2187 (O_2187,N_29401,N_29515);
or UO_2188 (O_2188,N_29293,N_28651);
or UO_2189 (O_2189,N_29650,N_29456);
nor UO_2190 (O_2190,N_29464,N_28787);
or UO_2191 (O_2191,N_29315,N_28601);
and UO_2192 (O_2192,N_29664,N_29384);
nor UO_2193 (O_2193,N_29289,N_29088);
and UO_2194 (O_2194,N_29324,N_29726);
xnor UO_2195 (O_2195,N_29526,N_29608);
nand UO_2196 (O_2196,N_28756,N_29007);
and UO_2197 (O_2197,N_28767,N_29593);
or UO_2198 (O_2198,N_28782,N_29421);
nor UO_2199 (O_2199,N_29128,N_29312);
xor UO_2200 (O_2200,N_29906,N_28749);
nor UO_2201 (O_2201,N_29275,N_29669);
nor UO_2202 (O_2202,N_29769,N_29841);
nor UO_2203 (O_2203,N_29876,N_28860);
or UO_2204 (O_2204,N_29400,N_29178);
nor UO_2205 (O_2205,N_28530,N_29955);
or UO_2206 (O_2206,N_28786,N_29909);
nor UO_2207 (O_2207,N_29726,N_29139);
nand UO_2208 (O_2208,N_28642,N_29742);
and UO_2209 (O_2209,N_29877,N_29822);
and UO_2210 (O_2210,N_29334,N_28813);
xnor UO_2211 (O_2211,N_29052,N_29426);
or UO_2212 (O_2212,N_29379,N_28695);
and UO_2213 (O_2213,N_29617,N_28611);
nand UO_2214 (O_2214,N_29317,N_29149);
or UO_2215 (O_2215,N_28886,N_29871);
nand UO_2216 (O_2216,N_29588,N_29023);
xnor UO_2217 (O_2217,N_29143,N_29255);
or UO_2218 (O_2218,N_29337,N_29435);
or UO_2219 (O_2219,N_29917,N_29527);
or UO_2220 (O_2220,N_29612,N_29486);
or UO_2221 (O_2221,N_28615,N_29653);
xor UO_2222 (O_2222,N_29623,N_28983);
nand UO_2223 (O_2223,N_28996,N_29266);
or UO_2224 (O_2224,N_29340,N_29008);
or UO_2225 (O_2225,N_29602,N_29293);
or UO_2226 (O_2226,N_29633,N_29747);
and UO_2227 (O_2227,N_28945,N_29833);
nor UO_2228 (O_2228,N_29395,N_29291);
xor UO_2229 (O_2229,N_29864,N_29595);
xor UO_2230 (O_2230,N_28901,N_29569);
and UO_2231 (O_2231,N_28803,N_28540);
nor UO_2232 (O_2232,N_29537,N_29274);
xnor UO_2233 (O_2233,N_29620,N_28801);
nand UO_2234 (O_2234,N_29181,N_28503);
nand UO_2235 (O_2235,N_28589,N_28993);
xnor UO_2236 (O_2236,N_29067,N_28846);
and UO_2237 (O_2237,N_29214,N_28839);
and UO_2238 (O_2238,N_29779,N_28566);
and UO_2239 (O_2239,N_29309,N_29982);
nand UO_2240 (O_2240,N_28829,N_28712);
and UO_2241 (O_2241,N_28909,N_29624);
nand UO_2242 (O_2242,N_29180,N_29771);
nor UO_2243 (O_2243,N_29782,N_29333);
and UO_2244 (O_2244,N_29612,N_28975);
nor UO_2245 (O_2245,N_28927,N_28976);
or UO_2246 (O_2246,N_28881,N_29819);
and UO_2247 (O_2247,N_29682,N_29115);
and UO_2248 (O_2248,N_29834,N_29609);
nand UO_2249 (O_2249,N_28798,N_29892);
nand UO_2250 (O_2250,N_29299,N_29381);
nor UO_2251 (O_2251,N_29939,N_29728);
and UO_2252 (O_2252,N_28867,N_29912);
nand UO_2253 (O_2253,N_29963,N_29129);
xor UO_2254 (O_2254,N_29610,N_29466);
xor UO_2255 (O_2255,N_29475,N_29203);
nand UO_2256 (O_2256,N_29262,N_28613);
nand UO_2257 (O_2257,N_29521,N_29967);
or UO_2258 (O_2258,N_29524,N_28926);
xor UO_2259 (O_2259,N_29818,N_29042);
nor UO_2260 (O_2260,N_29290,N_29320);
or UO_2261 (O_2261,N_28519,N_28741);
nor UO_2262 (O_2262,N_29021,N_29834);
nor UO_2263 (O_2263,N_29214,N_29736);
nor UO_2264 (O_2264,N_29553,N_29948);
or UO_2265 (O_2265,N_29275,N_28966);
nand UO_2266 (O_2266,N_29744,N_29050);
and UO_2267 (O_2267,N_28543,N_28664);
nand UO_2268 (O_2268,N_28860,N_28628);
nor UO_2269 (O_2269,N_29907,N_29725);
nor UO_2270 (O_2270,N_29850,N_28735);
xnor UO_2271 (O_2271,N_29658,N_29144);
or UO_2272 (O_2272,N_29279,N_29617);
nand UO_2273 (O_2273,N_29371,N_28704);
and UO_2274 (O_2274,N_28972,N_28845);
xnor UO_2275 (O_2275,N_28774,N_29357);
and UO_2276 (O_2276,N_29925,N_29358);
xor UO_2277 (O_2277,N_28807,N_28804);
or UO_2278 (O_2278,N_29260,N_29222);
and UO_2279 (O_2279,N_28806,N_28804);
and UO_2280 (O_2280,N_29662,N_29496);
nor UO_2281 (O_2281,N_29786,N_29189);
nor UO_2282 (O_2282,N_29795,N_29588);
nand UO_2283 (O_2283,N_29264,N_28862);
nand UO_2284 (O_2284,N_29721,N_29180);
xor UO_2285 (O_2285,N_28794,N_28660);
xnor UO_2286 (O_2286,N_29914,N_28788);
xnor UO_2287 (O_2287,N_29014,N_28894);
and UO_2288 (O_2288,N_29671,N_29001);
nor UO_2289 (O_2289,N_29114,N_28640);
nand UO_2290 (O_2290,N_29980,N_28749);
nand UO_2291 (O_2291,N_28906,N_29553);
nor UO_2292 (O_2292,N_29687,N_29743);
or UO_2293 (O_2293,N_29845,N_28956);
or UO_2294 (O_2294,N_29445,N_29736);
nor UO_2295 (O_2295,N_29742,N_28551);
xnor UO_2296 (O_2296,N_29246,N_29094);
nor UO_2297 (O_2297,N_28762,N_28555);
nand UO_2298 (O_2298,N_28862,N_29697);
nor UO_2299 (O_2299,N_29893,N_29877);
and UO_2300 (O_2300,N_28822,N_29563);
nor UO_2301 (O_2301,N_29699,N_28801);
nand UO_2302 (O_2302,N_29094,N_29956);
nor UO_2303 (O_2303,N_29552,N_28778);
xnor UO_2304 (O_2304,N_28783,N_29944);
nor UO_2305 (O_2305,N_29380,N_28920);
xor UO_2306 (O_2306,N_28930,N_29670);
nor UO_2307 (O_2307,N_28505,N_29053);
xor UO_2308 (O_2308,N_29963,N_29981);
xnor UO_2309 (O_2309,N_29360,N_29930);
and UO_2310 (O_2310,N_29674,N_29771);
nor UO_2311 (O_2311,N_29375,N_29770);
and UO_2312 (O_2312,N_28791,N_29396);
nor UO_2313 (O_2313,N_29910,N_28508);
nor UO_2314 (O_2314,N_29174,N_29353);
or UO_2315 (O_2315,N_28910,N_29497);
xnor UO_2316 (O_2316,N_28771,N_29571);
xor UO_2317 (O_2317,N_29521,N_29935);
or UO_2318 (O_2318,N_29150,N_28538);
or UO_2319 (O_2319,N_29935,N_29415);
nor UO_2320 (O_2320,N_29505,N_28649);
xnor UO_2321 (O_2321,N_29330,N_28509);
xnor UO_2322 (O_2322,N_28858,N_29263);
nor UO_2323 (O_2323,N_29250,N_29901);
nand UO_2324 (O_2324,N_29319,N_29507);
and UO_2325 (O_2325,N_29560,N_29465);
or UO_2326 (O_2326,N_28587,N_28543);
nor UO_2327 (O_2327,N_29917,N_29737);
nand UO_2328 (O_2328,N_28774,N_29684);
or UO_2329 (O_2329,N_29764,N_29136);
or UO_2330 (O_2330,N_29796,N_28684);
and UO_2331 (O_2331,N_29586,N_29206);
and UO_2332 (O_2332,N_29209,N_28794);
or UO_2333 (O_2333,N_28550,N_28570);
or UO_2334 (O_2334,N_29825,N_29086);
or UO_2335 (O_2335,N_29953,N_29711);
xnor UO_2336 (O_2336,N_29466,N_29285);
nand UO_2337 (O_2337,N_29499,N_29161);
and UO_2338 (O_2338,N_29557,N_29678);
or UO_2339 (O_2339,N_29146,N_29323);
nand UO_2340 (O_2340,N_29736,N_29223);
or UO_2341 (O_2341,N_29635,N_29391);
xnor UO_2342 (O_2342,N_29659,N_29239);
and UO_2343 (O_2343,N_28707,N_28879);
or UO_2344 (O_2344,N_29878,N_29366);
and UO_2345 (O_2345,N_29577,N_28586);
and UO_2346 (O_2346,N_28994,N_29717);
or UO_2347 (O_2347,N_28739,N_28982);
xnor UO_2348 (O_2348,N_28858,N_29783);
nor UO_2349 (O_2349,N_29268,N_28578);
or UO_2350 (O_2350,N_29304,N_29372);
nor UO_2351 (O_2351,N_29842,N_28968);
xor UO_2352 (O_2352,N_29799,N_29009);
and UO_2353 (O_2353,N_29519,N_28818);
and UO_2354 (O_2354,N_28980,N_28732);
xor UO_2355 (O_2355,N_28818,N_28857);
or UO_2356 (O_2356,N_29551,N_28825);
and UO_2357 (O_2357,N_29322,N_28519);
xor UO_2358 (O_2358,N_29259,N_29639);
and UO_2359 (O_2359,N_29122,N_28598);
nand UO_2360 (O_2360,N_29507,N_28510);
xnor UO_2361 (O_2361,N_29932,N_28713);
or UO_2362 (O_2362,N_28602,N_29225);
nand UO_2363 (O_2363,N_29731,N_29541);
and UO_2364 (O_2364,N_29026,N_28684);
nor UO_2365 (O_2365,N_28645,N_28593);
and UO_2366 (O_2366,N_29677,N_28840);
nand UO_2367 (O_2367,N_29886,N_29630);
nor UO_2368 (O_2368,N_29349,N_29631);
or UO_2369 (O_2369,N_29106,N_29941);
and UO_2370 (O_2370,N_29860,N_29383);
or UO_2371 (O_2371,N_29090,N_29738);
and UO_2372 (O_2372,N_29318,N_28667);
or UO_2373 (O_2373,N_29189,N_28758);
xnor UO_2374 (O_2374,N_29733,N_29485);
or UO_2375 (O_2375,N_28794,N_28937);
nor UO_2376 (O_2376,N_28771,N_29287);
nand UO_2377 (O_2377,N_29681,N_29306);
nand UO_2378 (O_2378,N_29804,N_29930);
or UO_2379 (O_2379,N_29839,N_28929);
and UO_2380 (O_2380,N_29659,N_29643);
nand UO_2381 (O_2381,N_28582,N_28651);
nor UO_2382 (O_2382,N_28737,N_28800);
xor UO_2383 (O_2383,N_28548,N_28916);
nor UO_2384 (O_2384,N_29547,N_29185);
nand UO_2385 (O_2385,N_29821,N_28966);
or UO_2386 (O_2386,N_28569,N_29597);
and UO_2387 (O_2387,N_28664,N_28657);
xor UO_2388 (O_2388,N_29634,N_28584);
and UO_2389 (O_2389,N_28908,N_29360);
nor UO_2390 (O_2390,N_29555,N_29850);
nor UO_2391 (O_2391,N_29349,N_29110);
xor UO_2392 (O_2392,N_28590,N_29940);
and UO_2393 (O_2393,N_28543,N_29979);
nand UO_2394 (O_2394,N_28744,N_29137);
or UO_2395 (O_2395,N_29063,N_28840);
nor UO_2396 (O_2396,N_28722,N_29169);
nor UO_2397 (O_2397,N_29507,N_29996);
xor UO_2398 (O_2398,N_28969,N_29427);
or UO_2399 (O_2399,N_29603,N_28916);
and UO_2400 (O_2400,N_28821,N_28867);
and UO_2401 (O_2401,N_29259,N_29172);
nand UO_2402 (O_2402,N_29942,N_29049);
or UO_2403 (O_2403,N_29354,N_28883);
or UO_2404 (O_2404,N_29028,N_29627);
and UO_2405 (O_2405,N_28872,N_29142);
and UO_2406 (O_2406,N_29487,N_29212);
and UO_2407 (O_2407,N_29576,N_28664);
xor UO_2408 (O_2408,N_28889,N_28612);
or UO_2409 (O_2409,N_29937,N_29429);
and UO_2410 (O_2410,N_29900,N_29755);
nand UO_2411 (O_2411,N_29330,N_29689);
and UO_2412 (O_2412,N_29961,N_28556);
nor UO_2413 (O_2413,N_29930,N_28550);
nor UO_2414 (O_2414,N_29964,N_29793);
xor UO_2415 (O_2415,N_29153,N_29231);
nand UO_2416 (O_2416,N_28772,N_28655);
nor UO_2417 (O_2417,N_28914,N_29509);
nand UO_2418 (O_2418,N_29038,N_28814);
nor UO_2419 (O_2419,N_29133,N_29739);
nand UO_2420 (O_2420,N_29723,N_28805);
nor UO_2421 (O_2421,N_29719,N_28775);
and UO_2422 (O_2422,N_29384,N_29141);
nand UO_2423 (O_2423,N_29689,N_29003);
or UO_2424 (O_2424,N_29843,N_28944);
xnor UO_2425 (O_2425,N_29114,N_29521);
or UO_2426 (O_2426,N_28899,N_29353);
or UO_2427 (O_2427,N_28684,N_29766);
or UO_2428 (O_2428,N_28853,N_29371);
and UO_2429 (O_2429,N_29768,N_29911);
and UO_2430 (O_2430,N_29211,N_28527);
or UO_2431 (O_2431,N_29839,N_28837);
nor UO_2432 (O_2432,N_28696,N_29903);
or UO_2433 (O_2433,N_29777,N_28678);
xor UO_2434 (O_2434,N_28726,N_29564);
and UO_2435 (O_2435,N_29556,N_28921);
and UO_2436 (O_2436,N_29346,N_28630);
or UO_2437 (O_2437,N_29544,N_29149);
or UO_2438 (O_2438,N_29216,N_28874);
or UO_2439 (O_2439,N_29740,N_28825);
xor UO_2440 (O_2440,N_28975,N_28575);
nor UO_2441 (O_2441,N_29760,N_28953);
xor UO_2442 (O_2442,N_28721,N_29158);
nor UO_2443 (O_2443,N_29139,N_28625);
xnor UO_2444 (O_2444,N_29726,N_29002);
and UO_2445 (O_2445,N_29953,N_29430);
nor UO_2446 (O_2446,N_29426,N_29780);
xor UO_2447 (O_2447,N_29056,N_29410);
or UO_2448 (O_2448,N_28513,N_29472);
xor UO_2449 (O_2449,N_29837,N_29815);
or UO_2450 (O_2450,N_28554,N_29030);
xor UO_2451 (O_2451,N_29388,N_29916);
nor UO_2452 (O_2452,N_29764,N_29279);
and UO_2453 (O_2453,N_29984,N_29331);
xor UO_2454 (O_2454,N_29233,N_29882);
or UO_2455 (O_2455,N_28660,N_29920);
nand UO_2456 (O_2456,N_29782,N_28505);
or UO_2457 (O_2457,N_29579,N_28551);
and UO_2458 (O_2458,N_29214,N_29228);
nor UO_2459 (O_2459,N_29010,N_28601);
nor UO_2460 (O_2460,N_29226,N_29710);
or UO_2461 (O_2461,N_28768,N_29178);
or UO_2462 (O_2462,N_28985,N_29674);
and UO_2463 (O_2463,N_29126,N_28699);
nand UO_2464 (O_2464,N_28592,N_29886);
nand UO_2465 (O_2465,N_28653,N_28684);
nor UO_2466 (O_2466,N_29446,N_29746);
and UO_2467 (O_2467,N_29948,N_29130);
and UO_2468 (O_2468,N_29336,N_29824);
and UO_2469 (O_2469,N_29349,N_28566);
or UO_2470 (O_2470,N_28565,N_29945);
and UO_2471 (O_2471,N_28779,N_29831);
and UO_2472 (O_2472,N_28772,N_29677);
xnor UO_2473 (O_2473,N_28779,N_29344);
or UO_2474 (O_2474,N_28723,N_29431);
nand UO_2475 (O_2475,N_28882,N_28995);
nand UO_2476 (O_2476,N_29025,N_29762);
xor UO_2477 (O_2477,N_29843,N_28642);
and UO_2478 (O_2478,N_28981,N_29746);
or UO_2479 (O_2479,N_28522,N_29912);
and UO_2480 (O_2480,N_29848,N_29354);
or UO_2481 (O_2481,N_29344,N_29625);
and UO_2482 (O_2482,N_28587,N_29394);
and UO_2483 (O_2483,N_29367,N_29208);
xnor UO_2484 (O_2484,N_28743,N_29195);
nor UO_2485 (O_2485,N_28776,N_28733);
nor UO_2486 (O_2486,N_28954,N_29437);
or UO_2487 (O_2487,N_28658,N_29073);
or UO_2488 (O_2488,N_28877,N_29294);
xor UO_2489 (O_2489,N_28833,N_29376);
or UO_2490 (O_2490,N_29552,N_28795);
xnor UO_2491 (O_2491,N_29641,N_29072);
nand UO_2492 (O_2492,N_29630,N_29056);
xor UO_2493 (O_2493,N_28677,N_29222);
and UO_2494 (O_2494,N_29254,N_29860);
nor UO_2495 (O_2495,N_28581,N_29158);
xnor UO_2496 (O_2496,N_29697,N_28909);
nand UO_2497 (O_2497,N_29721,N_29496);
and UO_2498 (O_2498,N_29106,N_29773);
nor UO_2499 (O_2499,N_29507,N_29935);
nor UO_2500 (O_2500,N_28684,N_29973);
and UO_2501 (O_2501,N_28777,N_29725);
and UO_2502 (O_2502,N_29531,N_29249);
or UO_2503 (O_2503,N_29964,N_29450);
xnor UO_2504 (O_2504,N_29970,N_29108);
nor UO_2505 (O_2505,N_28956,N_29182);
and UO_2506 (O_2506,N_29687,N_29367);
xor UO_2507 (O_2507,N_29859,N_28522);
xnor UO_2508 (O_2508,N_28599,N_29915);
or UO_2509 (O_2509,N_29300,N_29153);
or UO_2510 (O_2510,N_28986,N_28910);
xor UO_2511 (O_2511,N_29638,N_29175);
nand UO_2512 (O_2512,N_29734,N_29796);
or UO_2513 (O_2513,N_29245,N_29124);
nor UO_2514 (O_2514,N_29098,N_29666);
nand UO_2515 (O_2515,N_29814,N_29962);
nor UO_2516 (O_2516,N_29240,N_29345);
nor UO_2517 (O_2517,N_29829,N_29595);
nor UO_2518 (O_2518,N_28535,N_29655);
or UO_2519 (O_2519,N_29367,N_29574);
and UO_2520 (O_2520,N_28627,N_29441);
nor UO_2521 (O_2521,N_28586,N_29774);
xnor UO_2522 (O_2522,N_29106,N_29506);
nand UO_2523 (O_2523,N_29490,N_29693);
xor UO_2524 (O_2524,N_29398,N_28977);
or UO_2525 (O_2525,N_28892,N_29714);
nor UO_2526 (O_2526,N_29607,N_29456);
xor UO_2527 (O_2527,N_29133,N_29780);
xnor UO_2528 (O_2528,N_29277,N_29082);
or UO_2529 (O_2529,N_28711,N_29388);
nand UO_2530 (O_2530,N_29208,N_29457);
or UO_2531 (O_2531,N_29994,N_29677);
and UO_2532 (O_2532,N_29007,N_29842);
and UO_2533 (O_2533,N_29397,N_29504);
xnor UO_2534 (O_2534,N_29986,N_29168);
or UO_2535 (O_2535,N_29012,N_29458);
nor UO_2536 (O_2536,N_28776,N_29147);
or UO_2537 (O_2537,N_29094,N_29965);
and UO_2538 (O_2538,N_29641,N_29876);
xnor UO_2539 (O_2539,N_28693,N_29802);
nand UO_2540 (O_2540,N_29919,N_29819);
nor UO_2541 (O_2541,N_29683,N_29463);
or UO_2542 (O_2542,N_29898,N_28528);
nor UO_2543 (O_2543,N_29408,N_28676);
nor UO_2544 (O_2544,N_28810,N_29697);
and UO_2545 (O_2545,N_28650,N_28830);
and UO_2546 (O_2546,N_29575,N_29724);
and UO_2547 (O_2547,N_29977,N_28969);
and UO_2548 (O_2548,N_28754,N_29242);
and UO_2549 (O_2549,N_29712,N_29458);
and UO_2550 (O_2550,N_28604,N_29758);
or UO_2551 (O_2551,N_29516,N_29761);
nand UO_2552 (O_2552,N_29922,N_29849);
nor UO_2553 (O_2553,N_29057,N_29237);
xnor UO_2554 (O_2554,N_29908,N_28993);
or UO_2555 (O_2555,N_29949,N_28646);
nand UO_2556 (O_2556,N_29296,N_28650);
and UO_2557 (O_2557,N_29734,N_29068);
nor UO_2558 (O_2558,N_29995,N_29756);
nor UO_2559 (O_2559,N_28546,N_28987);
nand UO_2560 (O_2560,N_28615,N_29203);
xnor UO_2561 (O_2561,N_28937,N_29756);
xnor UO_2562 (O_2562,N_29872,N_28596);
nor UO_2563 (O_2563,N_29695,N_28951);
and UO_2564 (O_2564,N_29971,N_29357);
nand UO_2565 (O_2565,N_29050,N_29623);
and UO_2566 (O_2566,N_28973,N_29335);
or UO_2567 (O_2567,N_29106,N_29140);
nand UO_2568 (O_2568,N_29850,N_29630);
or UO_2569 (O_2569,N_28689,N_28731);
and UO_2570 (O_2570,N_28849,N_29170);
and UO_2571 (O_2571,N_28637,N_29326);
or UO_2572 (O_2572,N_29219,N_29157);
and UO_2573 (O_2573,N_28856,N_28605);
nor UO_2574 (O_2574,N_29461,N_28536);
or UO_2575 (O_2575,N_29495,N_28937);
or UO_2576 (O_2576,N_28882,N_28538);
or UO_2577 (O_2577,N_29496,N_28987);
nor UO_2578 (O_2578,N_28948,N_29699);
xnor UO_2579 (O_2579,N_29610,N_29398);
and UO_2580 (O_2580,N_29519,N_29430);
xnor UO_2581 (O_2581,N_28763,N_29251);
or UO_2582 (O_2582,N_28856,N_28779);
or UO_2583 (O_2583,N_29161,N_28855);
nand UO_2584 (O_2584,N_28859,N_28595);
nand UO_2585 (O_2585,N_29477,N_29138);
or UO_2586 (O_2586,N_29572,N_29120);
xor UO_2587 (O_2587,N_29302,N_29897);
nor UO_2588 (O_2588,N_29575,N_29820);
or UO_2589 (O_2589,N_29332,N_29608);
nand UO_2590 (O_2590,N_28707,N_29380);
or UO_2591 (O_2591,N_29319,N_29758);
and UO_2592 (O_2592,N_29865,N_28501);
nand UO_2593 (O_2593,N_29109,N_28669);
nand UO_2594 (O_2594,N_28942,N_28778);
nand UO_2595 (O_2595,N_29737,N_28837);
xnor UO_2596 (O_2596,N_29135,N_29491);
or UO_2597 (O_2597,N_29659,N_28781);
or UO_2598 (O_2598,N_29652,N_29438);
and UO_2599 (O_2599,N_28852,N_28740);
nor UO_2600 (O_2600,N_29986,N_28784);
xnor UO_2601 (O_2601,N_29762,N_29638);
or UO_2602 (O_2602,N_29454,N_29031);
xnor UO_2603 (O_2603,N_28720,N_29938);
or UO_2604 (O_2604,N_29761,N_28946);
nor UO_2605 (O_2605,N_29956,N_29046);
xnor UO_2606 (O_2606,N_29471,N_29211);
nor UO_2607 (O_2607,N_29775,N_29464);
and UO_2608 (O_2608,N_29359,N_29037);
or UO_2609 (O_2609,N_28763,N_29846);
nor UO_2610 (O_2610,N_28851,N_29414);
nor UO_2611 (O_2611,N_29156,N_28958);
and UO_2612 (O_2612,N_29478,N_28524);
nand UO_2613 (O_2613,N_29887,N_29578);
nand UO_2614 (O_2614,N_29886,N_29339);
and UO_2615 (O_2615,N_29691,N_28868);
xnor UO_2616 (O_2616,N_29947,N_29303);
xor UO_2617 (O_2617,N_28745,N_29433);
and UO_2618 (O_2618,N_29911,N_29462);
nand UO_2619 (O_2619,N_29789,N_29459);
nand UO_2620 (O_2620,N_29619,N_29803);
and UO_2621 (O_2621,N_28886,N_29179);
nand UO_2622 (O_2622,N_29377,N_29498);
xnor UO_2623 (O_2623,N_29874,N_29551);
or UO_2624 (O_2624,N_29561,N_29567);
xnor UO_2625 (O_2625,N_28768,N_29979);
nand UO_2626 (O_2626,N_29208,N_29193);
xor UO_2627 (O_2627,N_29431,N_29458);
and UO_2628 (O_2628,N_29720,N_28789);
xor UO_2629 (O_2629,N_29755,N_28607);
nand UO_2630 (O_2630,N_28799,N_28567);
nor UO_2631 (O_2631,N_29603,N_29630);
xor UO_2632 (O_2632,N_28853,N_29811);
nand UO_2633 (O_2633,N_29734,N_29374);
xnor UO_2634 (O_2634,N_29380,N_29612);
or UO_2635 (O_2635,N_29861,N_29632);
xor UO_2636 (O_2636,N_29358,N_29150);
nand UO_2637 (O_2637,N_29834,N_29174);
nand UO_2638 (O_2638,N_29728,N_29189);
and UO_2639 (O_2639,N_28672,N_29420);
and UO_2640 (O_2640,N_29788,N_29028);
nor UO_2641 (O_2641,N_28760,N_29021);
and UO_2642 (O_2642,N_29443,N_28693);
xnor UO_2643 (O_2643,N_29588,N_29559);
nand UO_2644 (O_2644,N_29672,N_29631);
nand UO_2645 (O_2645,N_29032,N_29402);
or UO_2646 (O_2646,N_29303,N_28923);
and UO_2647 (O_2647,N_29314,N_28518);
nor UO_2648 (O_2648,N_28991,N_28977);
xor UO_2649 (O_2649,N_28529,N_28760);
and UO_2650 (O_2650,N_29058,N_29753);
and UO_2651 (O_2651,N_28933,N_28690);
or UO_2652 (O_2652,N_29725,N_29328);
nand UO_2653 (O_2653,N_28706,N_28716);
xnor UO_2654 (O_2654,N_28566,N_29900);
nor UO_2655 (O_2655,N_28933,N_28928);
nand UO_2656 (O_2656,N_28749,N_29984);
and UO_2657 (O_2657,N_28728,N_29177);
nand UO_2658 (O_2658,N_28775,N_29461);
and UO_2659 (O_2659,N_29173,N_29313);
or UO_2660 (O_2660,N_28809,N_28891);
or UO_2661 (O_2661,N_29872,N_29542);
or UO_2662 (O_2662,N_28602,N_29377);
nand UO_2663 (O_2663,N_29012,N_29488);
or UO_2664 (O_2664,N_29200,N_29619);
xnor UO_2665 (O_2665,N_28981,N_29955);
nand UO_2666 (O_2666,N_28649,N_28952);
or UO_2667 (O_2667,N_29969,N_28742);
xor UO_2668 (O_2668,N_29757,N_29233);
xnor UO_2669 (O_2669,N_29800,N_29313);
nor UO_2670 (O_2670,N_28843,N_29134);
or UO_2671 (O_2671,N_28501,N_28532);
nand UO_2672 (O_2672,N_28819,N_29498);
nor UO_2673 (O_2673,N_28964,N_28727);
and UO_2674 (O_2674,N_29668,N_28966);
nor UO_2675 (O_2675,N_29818,N_29188);
nor UO_2676 (O_2676,N_28964,N_28980);
nand UO_2677 (O_2677,N_28998,N_29778);
nor UO_2678 (O_2678,N_28889,N_29372);
nor UO_2679 (O_2679,N_28558,N_29597);
xnor UO_2680 (O_2680,N_28613,N_29988);
or UO_2681 (O_2681,N_29335,N_28638);
and UO_2682 (O_2682,N_29131,N_29319);
nand UO_2683 (O_2683,N_28982,N_29455);
nor UO_2684 (O_2684,N_29898,N_29279);
nand UO_2685 (O_2685,N_29389,N_29410);
or UO_2686 (O_2686,N_29612,N_29520);
and UO_2687 (O_2687,N_28528,N_28711);
xnor UO_2688 (O_2688,N_28600,N_29472);
nor UO_2689 (O_2689,N_29722,N_29858);
xnor UO_2690 (O_2690,N_29508,N_29454);
or UO_2691 (O_2691,N_29158,N_29602);
xor UO_2692 (O_2692,N_29889,N_28864);
xor UO_2693 (O_2693,N_28753,N_29469);
nor UO_2694 (O_2694,N_29897,N_29148);
xor UO_2695 (O_2695,N_29827,N_28796);
xor UO_2696 (O_2696,N_28822,N_28766);
or UO_2697 (O_2697,N_28696,N_29315);
and UO_2698 (O_2698,N_29497,N_28597);
xor UO_2699 (O_2699,N_29036,N_29147);
or UO_2700 (O_2700,N_29547,N_29162);
nand UO_2701 (O_2701,N_28716,N_29146);
or UO_2702 (O_2702,N_29634,N_28569);
nor UO_2703 (O_2703,N_29676,N_29845);
nand UO_2704 (O_2704,N_29937,N_28845);
and UO_2705 (O_2705,N_29404,N_28697);
and UO_2706 (O_2706,N_29011,N_29878);
nor UO_2707 (O_2707,N_29116,N_29018);
xor UO_2708 (O_2708,N_29030,N_29370);
xnor UO_2709 (O_2709,N_29948,N_28735);
or UO_2710 (O_2710,N_29415,N_29682);
and UO_2711 (O_2711,N_29115,N_28551);
or UO_2712 (O_2712,N_29007,N_28799);
and UO_2713 (O_2713,N_28988,N_29900);
nor UO_2714 (O_2714,N_29631,N_29571);
xnor UO_2715 (O_2715,N_28502,N_29035);
nand UO_2716 (O_2716,N_28889,N_29501);
nand UO_2717 (O_2717,N_29610,N_29042);
and UO_2718 (O_2718,N_29245,N_29462);
nand UO_2719 (O_2719,N_29420,N_28566);
or UO_2720 (O_2720,N_28828,N_28912);
nand UO_2721 (O_2721,N_29302,N_28664);
xnor UO_2722 (O_2722,N_28690,N_29031);
nand UO_2723 (O_2723,N_28724,N_29201);
nor UO_2724 (O_2724,N_28805,N_29527);
nor UO_2725 (O_2725,N_29196,N_29163);
nor UO_2726 (O_2726,N_29527,N_29642);
nand UO_2727 (O_2727,N_28960,N_29283);
xnor UO_2728 (O_2728,N_29344,N_29698);
nand UO_2729 (O_2729,N_29693,N_29494);
xor UO_2730 (O_2730,N_28719,N_28807);
xnor UO_2731 (O_2731,N_29484,N_29551);
or UO_2732 (O_2732,N_29860,N_29148);
xnor UO_2733 (O_2733,N_28536,N_29491);
nand UO_2734 (O_2734,N_29191,N_29155);
nor UO_2735 (O_2735,N_29064,N_28831);
and UO_2736 (O_2736,N_28938,N_29120);
xnor UO_2737 (O_2737,N_29617,N_28521);
nand UO_2738 (O_2738,N_29244,N_28909);
nand UO_2739 (O_2739,N_29398,N_29857);
nor UO_2740 (O_2740,N_29807,N_28745);
nand UO_2741 (O_2741,N_28797,N_28940);
nor UO_2742 (O_2742,N_28710,N_29291);
nand UO_2743 (O_2743,N_29287,N_29478);
and UO_2744 (O_2744,N_29221,N_29321);
or UO_2745 (O_2745,N_29276,N_29003);
nor UO_2746 (O_2746,N_29231,N_29060);
and UO_2747 (O_2747,N_28986,N_29530);
and UO_2748 (O_2748,N_28522,N_29161);
and UO_2749 (O_2749,N_29381,N_29044);
nand UO_2750 (O_2750,N_29813,N_29420);
and UO_2751 (O_2751,N_28917,N_28571);
nand UO_2752 (O_2752,N_29756,N_29776);
xor UO_2753 (O_2753,N_29803,N_29726);
xor UO_2754 (O_2754,N_29810,N_29128);
nand UO_2755 (O_2755,N_29413,N_29813);
nand UO_2756 (O_2756,N_29975,N_29593);
xor UO_2757 (O_2757,N_29032,N_29897);
and UO_2758 (O_2758,N_28643,N_29764);
and UO_2759 (O_2759,N_29905,N_28537);
nand UO_2760 (O_2760,N_28926,N_29521);
nor UO_2761 (O_2761,N_28538,N_29498);
nor UO_2762 (O_2762,N_29018,N_28772);
nor UO_2763 (O_2763,N_29042,N_29479);
or UO_2764 (O_2764,N_29003,N_28772);
nor UO_2765 (O_2765,N_29627,N_28737);
nand UO_2766 (O_2766,N_29317,N_28673);
xor UO_2767 (O_2767,N_28815,N_28717);
xnor UO_2768 (O_2768,N_28633,N_29087);
or UO_2769 (O_2769,N_28813,N_29017);
xnor UO_2770 (O_2770,N_29358,N_28642);
xor UO_2771 (O_2771,N_29155,N_28609);
and UO_2772 (O_2772,N_28715,N_29594);
xor UO_2773 (O_2773,N_28905,N_28536);
nand UO_2774 (O_2774,N_28885,N_29466);
or UO_2775 (O_2775,N_29673,N_29278);
nand UO_2776 (O_2776,N_29775,N_29360);
xor UO_2777 (O_2777,N_29608,N_29063);
and UO_2778 (O_2778,N_29418,N_28534);
and UO_2779 (O_2779,N_29644,N_29942);
and UO_2780 (O_2780,N_29963,N_29471);
nand UO_2781 (O_2781,N_29622,N_29597);
xnor UO_2782 (O_2782,N_29881,N_29852);
nand UO_2783 (O_2783,N_29053,N_29045);
nand UO_2784 (O_2784,N_28968,N_29282);
and UO_2785 (O_2785,N_28554,N_28689);
xor UO_2786 (O_2786,N_29348,N_29714);
xor UO_2787 (O_2787,N_29914,N_29495);
xnor UO_2788 (O_2788,N_29270,N_29445);
or UO_2789 (O_2789,N_29700,N_29798);
xor UO_2790 (O_2790,N_29645,N_28548);
or UO_2791 (O_2791,N_28770,N_29770);
and UO_2792 (O_2792,N_29578,N_28921);
and UO_2793 (O_2793,N_29151,N_28982);
or UO_2794 (O_2794,N_29454,N_28705);
nor UO_2795 (O_2795,N_29293,N_29876);
and UO_2796 (O_2796,N_29953,N_28886);
nor UO_2797 (O_2797,N_29821,N_29594);
xnor UO_2798 (O_2798,N_29982,N_28549);
nor UO_2799 (O_2799,N_29634,N_28632);
nor UO_2800 (O_2800,N_29438,N_29399);
or UO_2801 (O_2801,N_29919,N_28807);
and UO_2802 (O_2802,N_28740,N_28612);
or UO_2803 (O_2803,N_29921,N_29755);
xnor UO_2804 (O_2804,N_29002,N_29780);
xnor UO_2805 (O_2805,N_28751,N_29372);
nand UO_2806 (O_2806,N_28849,N_29492);
nor UO_2807 (O_2807,N_29854,N_29259);
nor UO_2808 (O_2808,N_29274,N_28504);
nand UO_2809 (O_2809,N_29154,N_29497);
nor UO_2810 (O_2810,N_28549,N_29555);
nor UO_2811 (O_2811,N_29413,N_28580);
nor UO_2812 (O_2812,N_28828,N_28653);
nor UO_2813 (O_2813,N_29612,N_29684);
or UO_2814 (O_2814,N_29779,N_29100);
nor UO_2815 (O_2815,N_28781,N_29108);
or UO_2816 (O_2816,N_29552,N_29173);
nand UO_2817 (O_2817,N_28747,N_29514);
xnor UO_2818 (O_2818,N_29398,N_28833);
xnor UO_2819 (O_2819,N_29386,N_29843);
nor UO_2820 (O_2820,N_29266,N_29070);
nor UO_2821 (O_2821,N_28571,N_28970);
or UO_2822 (O_2822,N_29917,N_28644);
nor UO_2823 (O_2823,N_29039,N_28579);
nand UO_2824 (O_2824,N_29223,N_29198);
and UO_2825 (O_2825,N_28914,N_28537);
nand UO_2826 (O_2826,N_28733,N_29110);
nand UO_2827 (O_2827,N_29779,N_29195);
xor UO_2828 (O_2828,N_29562,N_29526);
or UO_2829 (O_2829,N_29518,N_28552);
xnor UO_2830 (O_2830,N_28940,N_28884);
and UO_2831 (O_2831,N_29334,N_29895);
and UO_2832 (O_2832,N_29329,N_29966);
xor UO_2833 (O_2833,N_28834,N_29678);
or UO_2834 (O_2834,N_29461,N_29143);
or UO_2835 (O_2835,N_28875,N_29345);
and UO_2836 (O_2836,N_29435,N_29781);
xor UO_2837 (O_2837,N_29559,N_28842);
and UO_2838 (O_2838,N_28520,N_29946);
xnor UO_2839 (O_2839,N_29188,N_29216);
or UO_2840 (O_2840,N_29839,N_29120);
and UO_2841 (O_2841,N_28795,N_29089);
nand UO_2842 (O_2842,N_29378,N_29549);
xnor UO_2843 (O_2843,N_29770,N_29970);
and UO_2844 (O_2844,N_28962,N_29594);
and UO_2845 (O_2845,N_29331,N_29936);
or UO_2846 (O_2846,N_29420,N_29494);
nor UO_2847 (O_2847,N_28643,N_29164);
nand UO_2848 (O_2848,N_29259,N_28666);
or UO_2849 (O_2849,N_29945,N_29279);
xor UO_2850 (O_2850,N_29561,N_29542);
and UO_2851 (O_2851,N_28634,N_28808);
and UO_2852 (O_2852,N_28811,N_29473);
and UO_2853 (O_2853,N_28680,N_29629);
nor UO_2854 (O_2854,N_29955,N_29511);
or UO_2855 (O_2855,N_28963,N_29956);
and UO_2856 (O_2856,N_29285,N_28866);
xor UO_2857 (O_2857,N_29130,N_29531);
and UO_2858 (O_2858,N_29472,N_29922);
and UO_2859 (O_2859,N_28711,N_29765);
nor UO_2860 (O_2860,N_28780,N_29125);
nand UO_2861 (O_2861,N_29567,N_29252);
or UO_2862 (O_2862,N_28926,N_29157);
or UO_2863 (O_2863,N_29704,N_29879);
xnor UO_2864 (O_2864,N_29267,N_29278);
xnor UO_2865 (O_2865,N_28940,N_29867);
and UO_2866 (O_2866,N_28732,N_29673);
xor UO_2867 (O_2867,N_29583,N_28626);
or UO_2868 (O_2868,N_29827,N_28878);
and UO_2869 (O_2869,N_29274,N_29718);
nor UO_2870 (O_2870,N_28893,N_28655);
xor UO_2871 (O_2871,N_28859,N_28950);
xor UO_2872 (O_2872,N_29618,N_29962);
xnor UO_2873 (O_2873,N_29571,N_29171);
nand UO_2874 (O_2874,N_29892,N_29494);
or UO_2875 (O_2875,N_29006,N_28627);
nand UO_2876 (O_2876,N_29621,N_29758);
or UO_2877 (O_2877,N_29323,N_29942);
nor UO_2878 (O_2878,N_29166,N_28558);
nand UO_2879 (O_2879,N_29934,N_29263);
nand UO_2880 (O_2880,N_28598,N_29881);
or UO_2881 (O_2881,N_29207,N_29498);
nor UO_2882 (O_2882,N_29736,N_29933);
or UO_2883 (O_2883,N_28801,N_29497);
and UO_2884 (O_2884,N_29377,N_29692);
nor UO_2885 (O_2885,N_28534,N_29419);
nor UO_2886 (O_2886,N_28970,N_28602);
and UO_2887 (O_2887,N_29183,N_29064);
nor UO_2888 (O_2888,N_29377,N_28988);
and UO_2889 (O_2889,N_29734,N_28703);
nor UO_2890 (O_2890,N_29662,N_28784);
or UO_2891 (O_2891,N_29749,N_29429);
xor UO_2892 (O_2892,N_29435,N_28667);
or UO_2893 (O_2893,N_28746,N_29858);
or UO_2894 (O_2894,N_29525,N_29424);
nor UO_2895 (O_2895,N_29902,N_28649);
and UO_2896 (O_2896,N_29175,N_28989);
xnor UO_2897 (O_2897,N_29381,N_28910);
nor UO_2898 (O_2898,N_29788,N_29751);
and UO_2899 (O_2899,N_28695,N_28629);
nor UO_2900 (O_2900,N_28883,N_28746);
xor UO_2901 (O_2901,N_29884,N_29971);
and UO_2902 (O_2902,N_28984,N_29279);
nand UO_2903 (O_2903,N_29079,N_29049);
and UO_2904 (O_2904,N_28919,N_29755);
xnor UO_2905 (O_2905,N_29809,N_29146);
or UO_2906 (O_2906,N_28846,N_29873);
or UO_2907 (O_2907,N_29575,N_28665);
xnor UO_2908 (O_2908,N_29378,N_29056);
or UO_2909 (O_2909,N_28757,N_29235);
and UO_2910 (O_2910,N_29201,N_29020);
xnor UO_2911 (O_2911,N_29515,N_29767);
and UO_2912 (O_2912,N_29987,N_29976);
nand UO_2913 (O_2913,N_29516,N_29025);
nor UO_2914 (O_2914,N_29993,N_29360);
nor UO_2915 (O_2915,N_29238,N_29029);
xnor UO_2916 (O_2916,N_28773,N_29872);
nor UO_2917 (O_2917,N_29640,N_29544);
nor UO_2918 (O_2918,N_29371,N_29616);
nor UO_2919 (O_2919,N_29101,N_29537);
nor UO_2920 (O_2920,N_28601,N_28866);
nand UO_2921 (O_2921,N_28805,N_29496);
or UO_2922 (O_2922,N_29714,N_29167);
and UO_2923 (O_2923,N_29364,N_29981);
nand UO_2924 (O_2924,N_29399,N_29112);
and UO_2925 (O_2925,N_29369,N_29617);
nand UO_2926 (O_2926,N_28550,N_28877);
nand UO_2927 (O_2927,N_28793,N_29906);
xor UO_2928 (O_2928,N_29211,N_28526);
nand UO_2929 (O_2929,N_29634,N_29156);
and UO_2930 (O_2930,N_28633,N_29826);
nand UO_2931 (O_2931,N_29828,N_29699);
nand UO_2932 (O_2932,N_28970,N_28975);
and UO_2933 (O_2933,N_28878,N_29598);
xor UO_2934 (O_2934,N_29699,N_28821);
nor UO_2935 (O_2935,N_28744,N_28911);
xnor UO_2936 (O_2936,N_29512,N_29036);
or UO_2937 (O_2937,N_29546,N_29340);
and UO_2938 (O_2938,N_28846,N_29110);
nor UO_2939 (O_2939,N_29409,N_28635);
nand UO_2940 (O_2940,N_29273,N_29371);
nor UO_2941 (O_2941,N_29873,N_28714);
nor UO_2942 (O_2942,N_29297,N_29854);
or UO_2943 (O_2943,N_29273,N_28587);
nor UO_2944 (O_2944,N_28560,N_28868);
and UO_2945 (O_2945,N_29695,N_29156);
and UO_2946 (O_2946,N_29990,N_29010);
or UO_2947 (O_2947,N_29248,N_29238);
nand UO_2948 (O_2948,N_28946,N_28891);
xor UO_2949 (O_2949,N_28961,N_29213);
xor UO_2950 (O_2950,N_29815,N_28605);
and UO_2951 (O_2951,N_29872,N_28586);
nor UO_2952 (O_2952,N_29211,N_29991);
or UO_2953 (O_2953,N_28880,N_29419);
nand UO_2954 (O_2954,N_29497,N_29371);
nand UO_2955 (O_2955,N_29825,N_29577);
and UO_2956 (O_2956,N_29302,N_28693);
nand UO_2957 (O_2957,N_28534,N_29330);
and UO_2958 (O_2958,N_29093,N_29019);
xnor UO_2959 (O_2959,N_29767,N_29431);
xor UO_2960 (O_2960,N_28932,N_29284);
and UO_2961 (O_2961,N_28528,N_28609);
nand UO_2962 (O_2962,N_29960,N_29878);
nand UO_2963 (O_2963,N_29809,N_28816);
and UO_2964 (O_2964,N_29210,N_28915);
and UO_2965 (O_2965,N_28891,N_28742);
or UO_2966 (O_2966,N_29801,N_29690);
and UO_2967 (O_2967,N_29051,N_29357);
nand UO_2968 (O_2968,N_29555,N_28543);
xnor UO_2969 (O_2969,N_29958,N_29364);
or UO_2970 (O_2970,N_29173,N_29967);
xnor UO_2971 (O_2971,N_29115,N_29492);
and UO_2972 (O_2972,N_29428,N_29792);
nand UO_2973 (O_2973,N_28553,N_28911);
xor UO_2974 (O_2974,N_29692,N_29227);
and UO_2975 (O_2975,N_28559,N_28708);
nor UO_2976 (O_2976,N_28809,N_28945);
xor UO_2977 (O_2977,N_28662,N_29288);
nor UO_2978 (O_2978,N_29834,N_29112);
nand UO_2979 (O_2979,N_29468,N_29367);
and UO_2980 (O_2980,N_28643,N_29605);
nor UO_2981 (O_2981,N_29102,N_29970);
xnor UO_2982 (O_2982,N_29147,N_29677);
and UO_2983 (O_2983,N_29800,N_28784);
xor UO_2984 (O_2984,N_29147,N_29892);
nor UO_2985 (O_2985,N_29085,N_28869);
and UO_2986 (O_2986,N_29909,N_28514);
xor UO_2987 (O_2987,N_28929,N_28905);
and UO_2988 (O_2988,N_28998,N_29271);
nand UO_2989 (O_2989,N_29891,N_28935);
and UO_2990 (O_2990,N_29687,N_29773);
nand UO_2991 (O_2991,N_29488,N_28626);
nand UO_2992 (O_2992,N_28905,N_29013);
and UO_2993 (O_2993,N_28519,N_28702);
xnor UO_2994 (O_2994,N_29599,N_28714);
or UO_2995 (O_2995,N_29650,N_28924);
xor UO_2996 (O_2996,N_29559,N_28591);
and UO_2997 (O_2997,N_28947,N_28965);
xor UO_2998 (O_2998,N_29940,N_29056);
or UO_2999 (O_2999,N_29235,N_29527);
and UO_3000 (O_3000,N_29894,N_29540);
xnor UO_3001 (O_3001,N_29434,N_28709);
or UO_3002 (O_3002,N_29908,N_29159);
nand UO_3003 (O_3003,N_28975,N_29029);
or UO_3004 (O_3004,N_28946,N_29313);
nor UO_3005 (O_3005,N_29018,N_29994);
nand UO_3006 (O_3006,N_29081,N_29962);
and UO_3007 (O_3007,N_29841,N_28632);
and UO_3008 (O_3008,N_28741,N_29380);
nand UO_3009 (O_3009,N_29847,N_28937);
and UO_3010 (O_3010,N_29326,N_29743);
and UO_3011 (O_3011,N_29478,N_29300);
and UO_3012 (O_3012,N_28662,N_29664);
xor UO_3013 (O_3013,N_29781,N_29144);
and UO_3014 (O_3014,N_29844,N_28910);
nand UO_3015 (O_3015,N_29325,N_28769);
xnor UO_3016 (O_3016,N_28570,N_29380);
and UO_3017 (O_3017,N_28565,N_29973);
xnor UO_3018 (O_3018,N_29209,N_28818);
or UO_3019 (O_3019,N_29079,N_29032);
and UO_3020 (O_3020,N_29094,N_29938);
and UO_3021 (O_3021,N_28589,N_29189);
xor UO_3022 (O_3022,N_29120,N_28899);
xnor UO_3023 (O_3023,N_29130,N_28524);
and UO_3024 (O_3024,N_29364,N_29923);
nor UO_3025 (O_3025,N_29292,N_28595);
nor UO_3026 (O_3026,N_28740,N_29633);
nor UO_3027 (O_3027,N_29606,N_29620);
nor UO_3028 (O_3028,N_29750,N_28882);
nand UO_3029 (O_3029,N_29693,N_29713);
or UO_3030 (O_3030,N_28500,N_28912);
nor UO_3031 (O_3031,N_29337,N_28677);
xor UO_3032 (O_3032,N_29037,N_28877);
or UO_3033 (O_3033,N_29744,N_28511);
xnor UO_3034 (O_3034,N_29355,N_29983);
nand UO_3035 (O_3035,N_29657,N_29044);
nand UO_3036 (O_3036,N_28747,N_29424);
and UO_3037 (O_3037,N_29203,N_28537);
nand UO_3038 (O_3038,N_29690,N_29255);
and UO_3039 (O_3039,N_28510,N_29935);
and UO_3040 (O_3040,N_29529,N_28550);
nor UO_3041 (O_3041,N_28976,N_28764);
xor UO_3042 (O_3042,N_28512,N_29688);
nand UO_3043 (O_3043,N_29424,N_29321);
and UO_3044 (O_3044,N_29946,N_28719);
and UO_3045 (O_3045,N_29763,N_29892);
nand UO_3046 (O_3046,N_29179,N_29772);
nor UO_3047 (O_3047,N_29201,N_29967);
and UO_3048 (O_3048,N_28859,N_29814);
and UO_3049 (O_3049,N_29858,N_29097);
nand UO_3050 (O_3050,N_29101,N_29230);
xor UO_3051 (O_3051,N_28987,N_29739);
and UO_3052 (O_3052,N_29924,N_29124);
and UO_3053 (O_3053,N_29691,N_28904);
nand UO_3054 (O_3054,N_29516,N_29067);
nor UO_3055 (O_3055,N_28768,N_29000);
or UO_3056 (O_3056,N_29190,N_29988);
nand UO_3057 (O_3057,N_29023,N_29125);
nand UO_3058 (O_3058,N_29992,N_29723);
nor UO_3059 (O_3059,N_29270,N_29003);
or UO_3060 (O_3060,N_28612,N_28564);
nor UO_3061 (O_3061,N_28652,N_29082);
or UO_3062 (O_3062,N_29323,N_28625);
and UO_3063 (O_3063,N_28870,N_28613);
xor UO_3064 (O_3064,N_29574,N_29164);
or UO_3065 (O_3065,N_29924,N_29850);
and UO_3066 (O_3066,N_29131,N_28684);
nor UO_3067 (O_3067,N_29079,N_29921);
and UO_3068 (O_3068,N_28569,N_29871);
or UO_3069 (O_3069,N_28779,N_29380);
or UO_3070 (O_3070,N_29448,N_29713);
xor UO_3071 (O_3071,N_28624,N_28880);
xor UO_3072 (O_3072,N_29948,N_28801);
and UO_3073 (O_3073,N_28995,N_29973);
nor UO_3074 (O_3074,N_29889,N_28515);
and UO_3075 (O_3075,N_28737,N_29667);
or UO_3076 (O_3076,N_29478,N_28539);
nor UO_3077 (O_3077,N_29836,N_29448);
nor UO_3078 (O_3078,N_29913,N_29759);
xnor UO_3079 (O_3079,N_29740,N_28816);
nand UO_3080 (O_3080,N_29781,N_28505);
xor UO_3081 (O_3081,N_29412,N_28999);
and UO_3082 (O_3082,N_29323,N_29818);
or UO_3083 (O_3083,N_29401,N_29223);
nor UO_3084 (O_3084,N_29883,N_28800);
nor UO_3085 (O_3085,N_29022,N_29109);
xnor UO_3086 (O_3086,N_28629,N_28569);
nand UO_3087 (O_3087,N_28805,N_28667);
or UO_3088 (O_3088,N_29614,N_28967);
xnor UO_3089 (O_3089,N_29658,N_28518);
xor UO_3090 (O_3090,N_29710,N_29403);
nor UO_3091 (O_3091,N_29231,N_29489);
xnor UO_3092 (O_3092,N_29263,N_29025);
xor UO_3093 (O_3093,N_29081,N_28840);
or UO_3094 (O_3094,N_28805,N_28592);
nor UO_3095 (O_3095,N_29142,N_29025);
xnor UO_3096 (O_3096,N_29025,N_29757);
and UO_3097 (O_3097,N_29321,N_29278);
xor UO_3098 (O_3098,N_29991,N_29711);
nand UO_3099 (O_3099,N_29779,N_28603);
nor UO_3100 (O_3100,N_28916,N_29246);
and UO_3101 (O_3101,N_29118,N_29450);
and UO_3102 (O_3102,N_28662,N_29914);
xor UO_3103 (O_3103,N_29020,N_29941);
xnor UO_3104 (O_3104,N_28700,N_29877);
nor UO_3105 (O_3105,N_29407,N_29824);
and UO_3106 (O_3106,N_28964,N_29559);
and UO_3107 (O_3107,N_29092,N_29227);
nand UO_3108 (O_3108,N_29043,N_29958);
or UO_3109 (O_3109,N_29966,N_29302);
or UO_3110 (O_3110,N_28740,N_29484);
nand UO_3111 (O_3111,N_29670,N_29937);
nand UO_3112 (O_3112,N_29570,N_29096);
nor UO_3113 (O_3113,N_29861,N_29957);
xnor UO_3114 (O_3114,N_29292,N_29366);
nor UO_3115 (O_3115,N_28861,N_28595);
and UO_3116 (O_3116,N_29967,N_29903);
nand UO_3117 (O_3117,N_29376,N_29689);
and UO_3118 (O_3118,N_28947,N_29581);
xnor UO_3119 (O_3119,N_28854,N_29444);
and UO_3120 (O_3120,N_29631,N_28738);
or UO_3121 (O_3121,N_29754,N_29885);
or UO_3122 (O_3122,N_29170,N_29954);
nand UO_3123 (O_3123,N_28930,N_29757);
or UO_3124 (O_3124,N_28767,N_29029);
nor UO_3125 (O_3125,N_29747,N_28748);
and UO_3126 (O_3126,N_29214,N_29544);
nor UO_3127 (O_3127,N_28980,N_28740);
xor UO_3128 (O_3128,N_29119,N_28659);
nor UO_3129 (O_3129,N_29911,N_29095);
xnor UO_3130 (O_3130,N_28516,N_29422);
nor UO_3131 (O_3131,N_28875,N_29742);
and UO_3132 (O_3132,N_29185,N_29417);
nand UO_3133 (O_3133,N_28703,N_28527);
and UO_3134 (O_3134,N_29595,N_28843);
nor UO_3135 (O_3135,N_29691,N_28564);
nor UO_3136 (O_3136,N_28808,N_28990);
and UO_3137 (O_3137,N_29824,N_29006);
nand UO_3138 (O_3138,N_28574,N_29866);
xnor UO_3139 (O_3139,N_29065,N_29872);
and UO_3140 (O_3140,N_29132,N_28548);
nor UO_3141 (O_3141,N_29196,N_29029);
and UO_3142 (O_3142,N_28654,N_29360);
nand UO_3143 (O_3143,N_29803,N_29805);
and UO_3144 (O_3144,N_29325,N_29191);
or UO_3145 (O_3145,N_28803,N_29217);
or UO_3146 (O_3146,N_28727,N_29569);
xor UO_3147 (O_3147,N_29584,N_29994);
nand UO_3148 (O_3148,N_29505,N_29404);
or UO_3149 (O_3149,N_29204,N_29413);
or UO_3150 (O_3150,N_29925,N_28829);
or UO_3151 (O_3151,N_29470,N_29710);
and UO_3152 (O_3152,N_29763,N_29909);
and UO_3153 (O_3153,N_28599,N_28775);
xor UO_3154 (O_3154,N_29954,N_29599);
nand UO_3155 (O_3155,N_28954,N_29264);
and UO_3156 (O_3156,N_29481,N_28840);
and UO_3157 (O_3157,N_29303,N_29123);
xnor UO_3158 (O_3158,N_28595,N_28655);
nand UO_3159 (O_3159,N_28504,N_29908);
nand UO_3160 (O_3160,N_29593,N_29693);
or UO_3161 (O_3161,N_28896,N_28661);
xnor UO_3162 (O_3162,N_28916,N_29385);
nor UO_3163 (O_3163,N_28854,N_29863);
nand UO_3164 (O_3164,N_29803,N_29385);
xnor UO_3165 (O_3165,N_29208,N_29447);
and UO_3166 (O_3166,N_29829,N_28949);
nor UO_3167 (O_3167,N_29410,N_28796);
xor UO_3168 (O_3168,N_28811,N_28871);
and UO_3169 (O_3169,N_28619,N_29705);
nand UO_3170 (O_3170,N_29651,N_28676);
or UO_3171 (O_3171,N_28777,N_29418);
xnor UO_3172 (O_3172,N_29165,N_29719);
or UO_3173 (O_3173,N_29379,N_29558);
nor UO_3174 (O_3174,N_29369,N_29359);
and UO_3175 (O_3175,N_29237,N_29009);
nand UO_3176 (O_3176,N_29789,N_28943);
xor UO_3177 (O_3177,N_29557,N_28845);
nand UO_3178 (O_3178,N_29411,N_29603);
xnor UO_3179 (O_3179,N_28607,N_29714);
or UO_3180 (O_3180,N_28632,N_29633);
and UO_3181 (O_3181,N_29062,N_29824);
and UO_3182 (O_3182,N_28791,N_29351);
xnor UO_3183 (O_3183,N_28818,N_28620);
and UO_3184 (O_3184,N_28753,N_29690);
nand UO_3185 (O_3185,N_29000,N_28506);
nand UO_3186 (O_3186,N_29851,N_29683);
and UO_3187 (O_3187,N_29934,N_29968);
nor UO_3188 (O_3188,N_29890,N_29468);
and UO_3189 (O_3189,N_29769,N_29278);
nor UO_3190 (O_3190,N_29807,N_29855);
nand UO_3191 (O_3191,N_29228,N_29953);
or UO_3192 (O_3192,N_29831,N_29497);
or UO_3193 (O_3193,N_28969,N_29756);
xnor UO_3194 (O_3194,N_29169,N_28650);
nand UO_3195 (O_3195,N_28807,N_28815);
nand UO_3196 (O_3196,N_28602,N_28891);
nand UO_3197 (O_3197,N_29284,N_29710);
nor UO_3198 (O_3198,N_29350,N_28835);
nand UO_3199 (O_3199,N_29195,N_29411);
or UO_3200 (O_3200,N_28826,N_28712);
or UO_3201 (O_3201,N_28542,N_29037);
and UO_3202 (O_3202,N_29579,N_29747);
nand UO_3203 (O_3203,N_29534,N_29562);
or UO_3204 (O_3204,N_28921,N_28807);
and UO_3205 (O_3205,N_29998,N_29717);
or UO_3206 (O_3206,N_28562,N_29562);
or UO_3207 (O_3207,N_29240,N_29581);
xor UO_3208 (O_3208,N_29654,N_28895);
and UO_3209 (O_3209,N_29399,N_28605);
xor UO_3210 (O_3210,N_29170,N_29042);
nor UO_3211 (O_3211,N_28881,N_29254);
nand UO_3212 (O_3212,N_29943,N_28605);
nor UO_3213 (O_3213,N_28661,N_29010);
xnor UO_3214 (O_3214,N_28712,N_29093);
or UO_3215 (O_3215,N_28867,N_29022);
xor UO_3216 (O_3216,N_29083,N_29310);
or UO_3217 (O_3217,N_29789,N_28950);
xor UO_3218 (O_3218,N_29651,N_29910);
nand UO_3219 (O_3219,N_29540,N_29950);
xor UO_3220 (O_3220,N_29475,N_29301);
or UO_3221 (O_3221,N_28878,N_29500);
xnor UO_3222 (O_3222,N_28923,N_29257);
xnor UO_3223 (O_3223,N_29674,N_29477);
nor UO_3224 (O_3224,N_29450,N_29808);
nor UO_3225 (O_3225,N_28675,N_29430);
nand UO_3226 (O_3226,N_29711,N_28872);
and UO_3227 (O_3227,N_29617,N_29339);
or UO_3228 (O_3228,N_28561,N_28694);
and UO_3229 (O_3229,N_28697,N_29852);
xor UO_3230 (O_3230,N_28519,N_29545);
nor UO_3231 (O_3231,N_29763,N_28694);
or UO_3232 (O_3232,N_29568,N_29135);
xor UO_3233 (O_3233,N_28674,N_28703);
xnor UO_3234 (O_3234,N_29154,N_29106);
or UO_3235 (O_3235,N_28732,N_28702);
and UO_3236 (O_3236,N_28649,N_29553);
xor UO_3237 (O_3237,N_28767,N_29706);
nor UO_3238 (O_3238,N_28778,N_29981);
or UO_3239 (O_3239,N_29001,N_28521);
nand UO_3240 (O_3240,N_29908,N_29141);
and UO_3241 (O_3241,N_29901,N_28959);
or UO_3242 (O_3242,N_29632,N_29133);
nand UO_3243 (O_3243,N_28813,N_29828);
and UO_3244 (O_3244,N_29442,N_28502);
and UO_3245 (O_3245,N_28688,N_29259);
and UO_3246 (O_3246,N_29698,N_28804);
xnor UO_3247 (O_3247,N_29807,N_29836);
and UO_3248 (O_3248,N_28871,N_29430);
and UO_3249 (O_3249,N_28828,N_29403);
or UO_3250 (O_3250,N_28549,N_29470);
xnor UO_3251 (O_3251,N_29011,N_28633);
nand UO_3252 (O_3252,N_28573,N_29686);
or UO_3253 (O_3253,N_29569,N_29858);
and UO_3254 (O_3254,N_29773,N_29608);
xnor UO_3255 (O_3255,N_29888,N_29527);
xnor UO_3256 (O_3256,N_28544,N_29066);
or UO_3257 (O_3257,N_28917,N_28616);
nor UO_3258 (O_3258,N_29363,N_29703);
xor UO_3259 (O_3259,N_29202,N_29285);
xnor UO_3260 (O_3260,N_29800,N_29215);
or UO_3261 (O_3261,N_29116,N_29121);
nand UO_3262 (O_3262,N_28766,N_29593);
or UO_3263 (O_3263,N_29195,N_28666);
nor UO_3264 (O_3264,N_29782,N_29654);
nand UO_3265 (O_3265,N_28868,N_29826);
or UO_3266 (O_3266,N_29807,N_28744);
nand UO_3267 (O_3267,N_29252,N_29452);
and UO_3268 (O_3268,N_29374,N_28921);
or UO_3269 (O_3269,N_29249,N_28871);
and UO_3270 (O_3270,N_28508,N_28728);
and UO_3271 (O_3271,N_29447,N_29406);
and UO_3272 (O_3272,N_28895,N_28813);
xor UO_3273 (O_3273,N_29365,N_29991);
nor UO_3274 (O_3274,N_29397,N_28938);
and UO_3275 (O_3275,N_28570,N_29012);
nand UO_3276 (O_3276,N_29093,N_28592);
nand UO_3277 (O_3277,N_29250,N_28528);
xnor UO_3278 (O_3278,N_28567,N_29375);
xor UO_3279 (O_3279,N_29401,N_29354);
nor UO_3280 (O_3280,N_29144,N_28848);
or UO_3281 (O_3281,N_29650,N_28790);
nand UO_3282 (O_3282,N_29934,N_28725);
or UO_3283 (O_3283,N_29658,N_29080);
xnor UO_3284 (O_3284,N_29452,N_29259);
and UO_3285 (O_3285,N_29601,N_29091);
xor UO_3286 (O_3286,N_29831,N_29206);
nand UO_3287 (O_3287,N_29917,N_29438);
and UO_3288 (O_3288,N_28955,N_28949);
nand UO_3289 (O_3289,N_28867,N_29818);
and UO_3290 (O_3290,N_29930,N_29594);
xnor UO_3291 (O_3291,N_29508,N_29451);
nand UO_3292 (O_3292,N_29990,N_29483);
nand UO_3293 (O_3293,N_29070,N_29711);
nand UO_3294 (O_3294,N_29037,N_29432);
and UO_3295 (O_3295,N_29897,N_29078);
nand UO_3296 (O_3296,N_29330,N_28745);
nand UO_3297 (O_3297,N_29163,N_29388);
nor UO_3298 (O_3298,N_28750,N_29483);
or UO_3299 (O_3299,N_29294,N_29814);
nor UO_3300 (O_3300,N_29096,N_29270);
xnor UO_3301 (O_3301,N_29441,N_28556);
nor UO_3302 (O_3302,N_28949,N_29581);
nor UO_3303 (O_3303,N_28943,N_29154);
or UO_3304 (O_3304,N_29327,N_29405);
or UO_3305 (O_3305,N_28591,N_28622);
nor UO_3306 (O_3306,N_29202,N_29227);
or UO_3307 (O_3307,N_29454,N_29981);
nand UO_3308 (O_3308,N_29101,N_29175);
or UO_3309 (O_3309,N_29627,N_28705);
nand UO_3310 (O_3310,N_29470,N_29243);
nor UO_3311 (O_3311,N_29232,N_28922);
nand UO_3312 (O_3312,N_29995,N_28889);
nand UO_3313 (O_3313,N_29706,N_29878);
nand UO_3314 (O_3314,N_29469,N_29573);
nand UO_3315 (O_3315,N_28719,N_29737);
xnor UO_3316 (O_3316,N_29659,N_28863);
and UO_3317 (O_3317,N_28997,N_28669);
xor UO_3318 (O_3318,N_28548,N_29774);
and UO_3319 (O_3319,N_28731,N_29743);
nand UO_3320 (O_3320,N_28960,N_28964);
and UO_3321 (O_3321,N_29049,N_29177);
and UO_3322 (O_3322,N_28556,N_29249);
or UO_3323 (O_3323,N_29361,N_28921);
or UO_3324 (O_3324,N_29782,N_28585);
and UO_3325 (O_3325,N_29005,N_29935);
or UO_3326 (O_3326,N_29189,N_29628);
xor UO_3327 (O_3327,N_29623,N_28595);
nand UO_3328 (O_3328,N_29564,N_28808);
xnor UO_3329 (O_3329,N_29138,N_29287);
and UO_3330 (O_3330,N_28919,N_29351);
nand UO_3331 (O_3331,N_29092,N_29824);
nand UO_3332 (O_3332,N_28976,N_29439);
nand UO_3333 (O_3333,N_29259,N_28555);
xor UO_3334 (O_3334,N_28776,N_28636);
nor UO_3335 (O_3335,N_29963,N_29763);
nand UO_3336 (O_3336,N_28765,N_29800);
xnor UO_3337 (O_3337,N_29484,N_29355);
or UO_3338 (O_3338,N_29332,N_29800);
nand UO_3339 (O_3339,N_29765,N_29583);
and UO_3340 (O_3340,N_29065,N_28871);
xnor UO_3341 (O_3341,N_29547,N_29049);
and UO_3342 (O_3342,N_29130,N_28802);
nor UO_3343 (O_3343,N_29655,N_28645);
xnor UO_3344 (O_3344,N_29523,N_29335);
or UO_3345 (O_3345,N_29315,N_29044);
nor UO_3346 (O_3346,N_28839,N_28601);
or UO_3347 (O_3347,N_28835,N_29996);
xnor UO_3348 (O_3348,N_29253,N_28934);
nand UO_3349 (O_3349,N_29827,N_29597);
xnor UO_3350 (O_3350,N_29559,N_29644);
xor UO_3351 (O_3351,N_28985,N_29891);
nor UO_3352 (O_3352,N_28957,N_29514);
nor UO_3353 (O_3353,N_28830,N_29459);
and UO_3354 (O_3354,N_29892,N_28601);
and UO_3355 (O_3355,N_29420,N_28823);
or UO_3356 (O_3356,N_29065,N_28982);
and UO_3357 (O_3357,N_29543,N_29509);
xor UO_3358 (O_3358,N_28707,N_29833);
nor UO_3359 (O_3359,N_28728,N_28843);
xor UO_3360 (O_3360,N_29970,N_29973);
xnor UO_3361 (O_3361,N_28907,N_29314);
and UO_3362 (O_3362,N_29277,N_29147);
or UO_3363 (O_3363,N_28533,N_29724);
and UO_3364 (O_3364,N_29873,N_29077);
or UO_3365 (O_3365,N_29624,N_28897);
or UO_3366 (O_3366,N_29037,N_29194);
and UO_3367 (O_3367,N_28752,N_29791);
nor UO_3368 (O_3368,N_29420,N_29671);
and UO_3369 (O_3369,N_29239,N_28975);
or UO_3370 (O_3370,N_28756,N_28697);
xnor UO_3371 (O_3371,N_29625,N_29271);
nor UO_3372 (O_3372,N_29254,N_29413);
or UO_3373 (O_3373,N_28830,N_28721);
and UO_3374 (O_3374,N_29745,N_29292);
and UO_3375 (O_3375,N_29615,N_28802);
nand UO_3376 (O_3376,N_29459,N_28696);
or UO_3377 (O_3377,N_28987,N_28724);
nor UO_3378 (O_3378,N_28515,N_28889);
nor UO_3379 (O_3379,N_28762,N_29587);
or UO_3380 (O_3380,N_29085,N_29190);
and UO_3381 (O_3381,N_29803,N_29844);
nand UO_3382 (O_3382,N_29737,N_28642);
xor UO_3383 (O_3383,N_29212,N_28570);
and UO_3384 (O_3384,N_29805,N_29719);
or UO_3385 (O_3385,N_29197,N_29506);
or UO_3386 (O_3386,N_29934,N_29767);
or UO_3387 (O_3387,N_29617,N_29677);
xnor UO_3388 (O_3388,N_29062,N_29381);
nand UO_3389 (O_3389,N_28998,N_28871);
xor UO_3390 (O_3390,N_28636,N_29581);
nor UO_3391 (O_3391,N_29120,N_29049);
xor UO_3392 (O_3392,N_29788,N_28558);
nor UO_3393 (O_3393,N_28942,N_29349);
and UO_3394 (O_3394,N_29328,N_28885);
and UO_3395 (O_3395,N_29287,N_29274);
and UO_3396 (O_3396,N_29204,N_29313);
and UO_3397 (O_3397,N_29967,N_29652);
and UO_3398 (O_3398,N_28736,N_29165);
xor UO_3399 (O_3399,N_28768,N_29038);
xor UO_3400 (O_3400,N_28848,N_28948);
nor UO_3401 (O_3401,N_29896,N_29246);
xnor UO_3402 (O_3402,N_28628,N_29493);
and UO_3403 (O_3403,N_29742,N_29463);
xor UO_3404 (O_3404,N_29734,N_29041);
and UO_3405 (O_3405,N_28701,N_29314);
or UO_3406 (O_3406,N_28730,N_29867);
or UO_3407 (O_3407,N_29178,N_29884);
and UO_3408 (O_3408,N_29753,N_29372);
nor UO_3409 (O_3409,N_29540,N_29171);
nand UO_3410 (O_3410,N_29419,N_29331);
and UO_3411 (O_3411,N_29001,N_29249);
nor UO_3412 (O_3412,N_29356,N_28774);
and UO_3413 (O_3413,N_29883,N_29760);
or UO_3414 (O_3414,N_29926,N_28567);
nor UO_3415 (O_3415,N_28682,N_29566);
and UO_3416 (O_3416,N_29841,N_29996);
or UO_3417 (O_3417,N_28971,N_29466);
xnor UO_3418 (O_3418,N_29850,N_28930);
nand UO_3419 (O_3419,N_29060,N_28679);
xnor UO_3420 (O_3420,N_29761,N_29877);
or UO_3421 (O_3421,N_28958,N_28581);
and UO_3422 (O_3422,N_29468,N_29837);
nor UO_3423 (O_3423,N_29823,N_29518);
nand UO_3424 (O_3424,N_28507,N_28662);
or UO_3425 (O_3425,N_29884,N_29970);
nor UO_3426 (O_3426,N_29180,N_29538);
nor UO_3427 (O_3427,N_29066,N_29127);
nor UO_3428 (O_3428,N_28727,N_28629);
nor UO_3429 (O_3429,N_29944,N_29160);
nor UO_3430 (O_3430,N_29394,N_29644);
and UO_3431 (O_3431,N_29445,N_29870);
xnor UO_3432 (O_3432,N_29938,N_28569);
nor UO_3433 (O_3433,N_29274,N_28736);
or UO_3434 (O_3434,N_28641,N_28998);
and UO_3435 (O_3435,N_29733,N_29235);
xnor UO_3436 (O_3436,N_29264,N_29741);
xnor UO_3437 (O_3437,N_29311,N_28950);
xor UO_3438 (O_3438,N_29029,N_29853);
nand UO_3439 (O_3439,N_28810,N_28672);
xnor UO_3440 (O_3440,N_29637,N_29982);
nand UO_3441 (O_3441,N_29071,N_29939);
and UO_3442 (O_3442,N_29357,N_29362);
and UO_3443 (O_3443,N_29454,N_29209);
and UO_3444 (O_3444,N_28883,N_29327);
or UO_3445 (O_3445,N_29309,N_29387);
nor UO_3446 (O_3446,N_29708,N_28927);
and UO_3447 (O_3447,N_29346,N_29119);
nor UO_3448 (O_3448,N_29687,N_28850);
nor UO_3449 (O_3449,N_29301,N_28568);
or UO_3450 (O_3450,N_29780,N_29842);
nand UO_3451 (O_3451,N_28576,N_28952);
and UO_3452 (O_3452,N_29953,N_29693);
and UO_3453 (O_3453,N_29405,N_28804);
nand UO_3454 (O_3454,N_29177,N_28957);
and UO_3455 (O_3455,N_28964,N_28662);
nand UO_3456 (O_3456,N_29190,N_28508);
xnor UO_3457 (O_3457,N_28975,N_28528);
or UO_3458 (O_3458,N_29759,N_28995);
xor UO_3459 (O_3459,N_29015,N_28659);
xor UO_3460 (O_3460,N_29588,N_29603);
xor UO_3461 (O_3461,N_29356,N_29279);
nor UO_3462 (O_3462,N_28884,N_28527);
xor UO_3463 (O_3463,N_28984,N_29523);
xor UO_3464 (O_3464,N_29283,N_29445);
and UO_3465 (O_3465,N_28797,N_28724);
xor UO_3466 (O_3466,N_29685,N_28741);
or UO_3467 (O_3467,N_29281,N_29288);
xnor UO_3468 (O_3468,N_29615,N_28590);
nand UO_3469 (O_3469,N_29726,N_28955);
nor UO_3470 (O_3470,N_28618,N_29113);
and UO_3471 (O_3471,N_28959,N_28598);
and UO_3472 (O_3472,N_28986,N_29562);
or UO_3473 (O_3473,N_29155,N_29015);
or UO_3474 (O_3474,N_29237,N_28576);
nor UO_3475 (O_3475,N_29429,N_29458);
nor UO_3476 (O_3476,N_28618,N_29940);
nand UO_3477 (O_3477,N_29706,N_29132);
nor UO_3478 (O_3478,N_29705,N_29874);
and UO_3479 (O_3479,N_29049,N_29722);
or UO_3480 (O_3480,N_29612,N_29809);
nand UO_3481 (O_3481,N_28502,N_29926);
nor UO_3482 (O_3482,N_29039,N_29000);
and UO_3483 (O_3483,N_28604,N_29395);
or UO_3484 (O_3484,N_28885,N_29172);
and UO_3485 (O_3485,N_29730,N_29789);
xor UO_3486 (O_3486,N_29868,N_28526);
or UO_3487 (O_3487,N_28846,N_29719);
xor UO_3488 (O_3488,N_29878,N_28504);
nand UO_3489 (O_3489,N_28621,N_29823);
nor UO_3490 (O_3490,N_28838,N_29611);
or UO_3491 (O_3491,N_28605,N_28515);
or UO_3492 (O_3492,N_29934,N_29594);
nor UO_3493 (O_3493,N_29654,N_28887);
or UO_3494 (O_3494,N_28717,N_29962);
or UO_3495 (O_3495,N_29975,N_29793);
and UO_3496 (O_3496,N_29371,N_29820);
nand UO_3497 (O_3497,N_29366,N_28635);
nor UO_3498 (O_3498,N_29333,N_29545);
and UO_3499 (O_3499,N_29928,N_28568);
endmodule