module basic_2500_25000_3000_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1798,In_1194);
and U1 (N_1,In_394,In_2178);
nor U2 (N_2,In_1512,In_898);
xor U3 (N_3,In_2274,In_364);
or U4 (N_4,In_863,In_1635);
and U5 (N_5,In_116,In_1371);
and U6 (N_6,In_1484,In_195);
nor U7 (N_7,In_938,In_2177);
xnor U8 (N_8,In_2105,In_536);
and U9 (N_9,In_2206,In_1030);
and U10 (N_10,In_178,In_1646);
nand U11 (N_11,In_737,In_982);
xor U12 (N_12,In_1265,In_2323);
nor U13 (N_13,In_1136,In_2279);
or U14 (N_14,In_416,In_1205);
or U15 (N_15,In_2422,In_2282);
xor U16 (N_16,In_730,In_2155);
or U17 (N_17,In_872,In_1887);
and U18 (N_18,In_298,In_476);
nor U19 (N_19,In_1970,In_468);
xor U20 (N_20,In_1775,In_2065);
xor U21 (N_21,In_1153,In_1303);
and U22 (N_22,In_1425,In_135);
and U23 (N_23,In_551,In_1319);
and U24 (N_24,In_1279,In_2337);
and U25 (N_25,In_1150,In_2154);
nand U26 (N_26,In_234,In_207);
or U27 (N_27,In_1399,In_1162);
xor U28 (N_28,In_1634,In_1382);
nand U29 (N_29,In_2479,In_277);
nor U30 (N_30,In_1507,In_398);
nand U31 (N_31,In_232,In_1107);
or U32 (N_32,In_3,In_2445);
nand U33 (N_33,In_817,In_2461);
and U34 (N_34,In_179,In_1800);
nand U35 (N_35,In_875,In_169);
xor U36 (N_36,In_334,In_333);
and U37 (N_37,In_291,In_1936);
nand U38 (N_38,In_1216,In_2275);
nand U39 (N_39,In_351,In_1051);
xnor U40 (N_40,In_2372,In_2345);
or U41 (N_41,In_976,In_63);
nor U42 (N_42,In_858,In_1964);
xnor U43 (N_43,In_945,In_672);
or U44 (N_44,In_498,In_1526);
nor U45 (N_45,In_1890,In_246);
or U46 (N_46,In_1917,In_668);
nor U47 (N_47,In_1274,In_6);
nor U48 (N_48,In_735,In_1891);
or U49 (N_49,In_1055,In_430);
xor U50 (N_50,In_1294,In_1199);
nor U51 (N_51,In_2293,In_896);
xor U52 (N_52,In_2472,In_2000);
nor U53 (N_53,In_2108,In_683);
nand U54 (N_54,In_1861,In_247);
nor U55 (N_55,In_1674,In_2020);
nand U56 (N_56,In_961,In_2348);
or U57 (N_57,In_5,In_1852);
and U58 (N_58,In_1956,In_1942);
and U59 (N_59,In_332,In_537);
or U60 (N_60,In_2227,In_255);
and U61 (N_61,In_1748,In_105);
nor U62 (N_62,In_2336,In_1214);
nor U63 (N_63,In_1187,In_2078);
nand U64 (N_64,In_317,In_475);
xnor U65 (N_65,In_915,In_611);
and U66 (N_66,In_2278,In_1139);
nand U67 (N_67,In_729,In_1731);
or U68 (N_68,In_710,In_1868);
nand U69 (N_69,In_2314,In_840);
or U70 (N_70,In_1811,In_2230);
nand U71 (N_71,In_558,In_433);
or U72 (N_72,In_2368,In_702);
or U73 (N_73,In_1571,In_1928);
xor U74 (N_74,In_306,In_2437);
and U75 (N_75,In_2481,In_1448);
or U76 (N_76,In_233,In_1036);
and U77 (N_77,In_757,In_1119);
xor U78 (N_78,In_1016,In_1588);
nor U79 (N_79,In_153,In_1025);
xnor U80 (N_80,In_2001,In_309);
or U81 (N_81,In_4,In_1268);
or U82 (N_82,In_830,In_1178);
or U83 (N_83,In_2210,In_2388);
nor U84 (N_84,In_345,In_36);
or U85 (N_85,In_21,In_1329);
nor U86 (N_86,In_1832,In_1758);
or U87 (N_87,In_1113,In_1723);
nor U88 (N_88,In_194,In_1567);
and U89 (N_89,In_821,In_2387);
and U90 (N_90,In_562,In_2113);
nor U91 (N_91,In_788,In_1631);
nor U92 (N_92,In_2013,In_571);
or U93 (N_93,In_1170,In_970);
xnor U94 (N_94,In_2369,In_884);
xor U95 (N_95,In_174,In_222);
nor U96 (N_96,In_1725,In_1420);
xnor U97 (N_97,In_184,In_1152);
or U98 (N_98,In_390,In_2112);
and U99 (N_99,In_1317,In_254);
nor U100 (N_100,In_926,In_1255);
xnor U101 (N_101,In_1801,In_1378);
xor U102 (N_102,In_1632,In_663);
or U103 (N_103,In_916,In_1168);
or U104 (N_104,In_2299,In_1392);
xnor U105 (N_105,In_533,In_1383);
and U106 (N_106,In_202,In_1235);
xnor U107 (N_107,In_764,In_41);
or U108 (N_108,In_856,In_1729);
and U109 (N_109,In_2285,In_1081);
nand U110 (N_110,In_2087,In_56);
and U111 (N_111,In_446,In_2166);
and U112 (N_112,In_1285,In_2484);
and U113 (N_113,In_943,In_260);
xor U114 (N_114,In_199,In_1493);
and U115 (N_115,In_1957,In_1395);
or U116 (N_116,In_1941,In_1599);
nor U117 (N_117,In_1389,In_1892);
nand U118 (N_118,In_673,In_2332);
or U119 (N_119,In_1940,In_888);
and U120 (N_120,In_1447,In_1000);
and U121 (N_121,In_2325,In_183);
nor U122 (N_122,In_822,In_2106);
or U123 (N_123,In_708,In_977);
or U124 (N_124,In_2216,In_2208);
and U125 (N_125,In_294,In_1144);
or U126 (N_126,In_1437,In_972);
xor U127 (N_127,In_1196,In_1446);
nor U128 (N_128,In_2027,In_1760);
nor U129 (N_129,In_1562,In_2257);
and U130 (N_130,In_550,In_1580);
or U131 (N_131,In_2264,In_1440);
or U132 (N_132,In_1471,In_2362);
nand U133 (N_133,In_1985,In_559);
nor U134 (N_134,In_1829,In_1839);
nand U135 (N_135,In_805,In_1023);
nand U136 (N_136,In_2086,In_635);
and U137 (N_137,In_1988,In_2485);
nand U138 (N_138,In_1078,In_1593);
or U139 (N_139,In_1769,In_1530);
nor U140 (N_140,In_2043,In_758);
or U141 (N_141,In_2196,In_2315);
nor U142 (N_142,In_762,In_1997);
nor U143 (N_143,In_1766,In_1911);
nand U144 (N_144,In_934,In_743);
nand U145 (N_145,In_18,In_423);
and U146 (N_146,In_761,In_2344);
and U147 (N_147,In_1370,In_2410);
nor U148 (N_148,In_1648,In_1824);
and U149 (N_149,In_284,In_2417);
nor U150 (N_150,In_578,In_1394);
nand U151 (N_151,In_387,In_2);
or U152 (N_152,In_1601,In_1918);
nor U153 (N_153,In_1046,In_89);
and U154 (N_154,In_2188,In_1529);
nand U155 (N_155,In_1838,In_1578);
xnor U156 (N_156,In_2312,In_1254);
nor U157 (N_157,In_918,In_1172);
and U158 (N_158,In_2042,In_742);
nand U159 (N_159,In_2038,In_1156);
nor U160 (N_160,In_2393,In_2017);
or U161 (N_161,In_1082,In_2357);
or U162 (N_162,In_434,In_2195);
nor U163 (N_163,In_1263,In_819);
nand U164 (N_164,In_1921,In_981);
nor U165 (N_165,In_186,In_523);
nor U166 (N_166,In_1999,In_458);
xor U167 (N_167,In_1974,In_2173);
nor U168 (N_168,In_1746,In_1292);
nand U169 (N_169,In_2404,In_1304);
nand U170 (N_170,In_584,In_767);
nor U171 (N_171,In_1176,In_336);
nand U172 (N_172,In_950,In_595);
nand U173 (N_173,In_2100,In_1197);
and U174 (N_174,In_119,In_827);
or U175 (N_175,In_2254,In_1834);
nor U176 (N_176,In_958,In_1939);
xor U177 (N_177,In_1017,In_392);
nor U178 (N_178,In_1772,In_1969);
nand U179 (N_179,In_2238,In_479);
or U180 (N_180,In_1174,In_2204);
or U181 (N_181,In_1784,In_1438);
and U182 (N_182,In_964,In_1788);
and U183 (N_183,In_1905,In_1825);
nor U184 (N_184,In_642,In_2163);
xor U185 (N_185,In_1753,In_2328);
xnor U186 (N_186,In_2438,In_1923);
or U187 (N_187,In_32,In_2433);
nor U188 (N_188,In_460,In_1125);
and U189 (N_189,In_1703,In_2077);
nor U190 (N_190,In_1384,In_1109);
xor U191 (N_191,In_1871,In_660);
nor U192 (N_192,In_2449,In_1071);
nand U193 (N_193,In_2110,In_2129);
and U194 (N_194,In_2249,In_1568);
or U195 (N_195,In_955,In_1224);
or U196 (N_196,In_2489,In_1124);
or U197 (N_197,In_1540,In_1434);
nor U198 (N_198,In_1966,In_652);
nand U199 (N_199,In_513,In_303);
xor U200 (N_200,In_1551,In_581);
xor U201 (N_201,In_771,In_1426);
nand U202 (N_202,In_1642,In_1318);
nand U203 (N_203,In_753,In_615);
nor U204 (N_204,In_1850,In_70);
xnor U205 (N_205,In_2320,In_1163);
nand U206 (N_206,In_2058,In_1706);
nor U207 (N_207,In_2473,In_1714);
or U208 (N_208,In_215,In_52);
nand U209 (N_209,In_1295,In_264);
nor U210 (N_210,In_1955,In_714);
nor U211 (N_211,In_1277,In_2308);
nor U212 (N_212,In_1536,In_98);
nand U213 (N_213,In_520,In_1142);
nor U214 (N_214,In_698,In_225);
or U215 (N_215,In_488,In_1542);
or U216 (N_216,In_741,In_930);
nor U217 (N_217,In_1469,In_807);
nor U218 (N_218,In_2191,In_2174);
nand U219 (N_219,In_1417,In_1184);
or U220 (N_220,In_1091,In_644);
and U221 (N_221,In_1881,In_1090);
and U222 (N_222,In_1745,In_385);
and U223 (N_223,In_785,In_2454);
nand U224 (N_224,In_440,In_1486);
nor U225 (N_225,In_780,In_1681);
or U226 (N_226,In_573,In_1179);
nand U227 (N_227,In_2213,In_1543);
or U228 (N_228,In_2470,In_799);
and U229 (N_229,In_1620,In_342);
nand U230 (N_230,In_889,In_1198);
and U231 (N_231,In_1155,In_1203);
nand U232 (N_232,In_2132,In_1700);
nand U233 (N_233,In_1963,In_641);
nor U234 (N_234,In_833,In_1668);
nand U235 (N_235,In_1768,In_2358);
xor U236 (N_236,In_2075,In_2356);
or U237 (N_237,In_1993,In_2343);
or U238 (N_238,In_2294,In_2015);
nor U239 (N_239,In_1306,In_132);
and U240 (N_240,In_1652,In_2046);
nand U241 (N_241,In_740,In_797);
nand U242 (N_242,In_280,In_421);
xnor U243 (N_243,In_1487,In_804);
xnor U244 (N_244,In_293,In_505);
and U245 (N_245,In_1931,In_218);
and U246 (N_246,In_1146,In_667);
or U247 (N_247,In_1056,In_1579);
nor U248 (N_248,In_1611,In_828);
xor U249 (N_249,In_193,In_2403);
nor U250 (N_250,In_1009,In_794);
nor U251 (N_251,In_883,In_1926);
xnor U252 (N_252,In_902,In_599);
and U253 (N_253,In_1315,In_449);
nor U254 (N_254,In_2237,In_1151);
xor U255 (N_255,In_868,In_846);
or U256 (N_256,In_181,In_789);
xor U257 (N_257,In_1996,In_1771);
or U258 (N_258,In_590,In_2400);
and U259 (N_259,In_1754,In_473);
and U260 (N_260,In_478,In_1247);
and U261 (N_261,In_1876,In_1903);
nor U262 (N_262,In_709,In_2071);
or U263 (N_263,In_1671,In_355);
nor U264 (N_264,In_2051,In_404);
xnor U265 (N_265,In_2450,In_2491);
and U266 (N_266,In_2242,In_1385);
and U267 (N_267,In_1206,In_606);
nand U268 (N_268,In_405,In_439);
and U269 (N_269,In_880,In_1264);
xor U270 (N_270,In_75,In_665);
nand U271 (N_271,In_2447,In_1060);
xor U272 (N_272,In_912,In_1138);
xnor U273 (N_273,In_2271,In_2025);
or U274 (N_274,In_1072,In_80);
or U275 (N_275,In_1356,In_1687);
nand U276 (N_276,In_2309,In_2465);
nor U277 (N_277,In_125,In_2121);
xor U278 (N_278,In_419,In_1074);
nor U279 (N_279,In_2119,In_684);
nand U280 (N_280,In_1869,In_2424);
xnor U281 (N_281,In_1331,In_700);
nor U282 (N_282,In_678,In_674);
and U283 (N_283,In_2059,In_1504);
xor U284 (N_284,In_1882,In_2260);
nor U285 (N_285,In_834,In_1128);
or U286 (N_286,In_173,In_2091);
or U287 (N_287,In_980,In_1335);
nor U288 (N_288,In_638,In_1951);
nand U289 (N_289,In_524,In_349);
nand U290 (N_290,In_593,In_1299);
or U291 (N_291,In_1010,In_1740);
and U292 (N_292,In_1033,In_413);
nand U293 (N_293,In_1131,In_899);
nor U294 (N_294,In_576,In_495);
nand U295 (N_295,In_1597,In_216);
xnor U296 (N_296,In_2187,In_72);
nand U297 (N_297,In_453,In_50);
nor U298 (N_298,In_2427,In_464);
nand U299 (N_299,In_83,In_1482);
and U300 (N_300,In_1201,In_278);
xnor U301 (N_301,In_2167,In_1358);
nand U302 (N_302,In_438,In_29);
and U303 (N_303,In_26,In_2389);
and U304 (N_304,In_230,In_1717);
xnor U305 (N_305,In_2033,In_2109);
nand U306 (N_306,In_2240,In_1814);
xor U307 (N_307,In_242,In_2120);
nor U308 (N_308,In_93,In_1439);
or U309 (N_309,In_1860,In_1616);
and U310 (N_310,In_1689,In_1325);
and U311 (N_311,In_1792,In_397);
nor U312 (N_312,In_2317,In_1727);
nand U313 (N_313,In_1020,In_602);
xnor U314 (N_314,In_969,In_2295);
nand U315 (N_315,In_1161,In_2482);
and U316 (N_316,In_2444,In_490);
nand U317 (N_317,In_847,In_1391);
xnor U318 (N_318,In_417,In_1553);
or U319 (N_319,In_2353,In_589);
and U320 (N_320,In_258,In_1699);
nor U321 (N_321,In_67,In_909);
xnor U322 (N_322,In_2367,In_472);
nor U323 (N_323,In_2340,In_1872);
xnor U324 (N_324,In_2319,In_1961);
or U325 (N_325,In_28,In_2192);
and U326 (N_326,In_1675,In_855);
and U327 (N_327,In_925,In_2172);
nand U328 (N_328,In_1716,In_503);
nand U329 (N_329,In_1453,In_2497);
xnor U330 (N_330,In_377,In_1780);
nor U331 (N_331,In_66,In_1628);
nand U332 (N_332,In_170,In_1252);
or U333 (N_333,In_849,In_1467);
xnor U334 (N_334,In_1100,In_73);
or U335 (N_335,In_1495,In_211);
nand U336 (N_336,In_1641,In_656);
or U337 (N_337,In_983,In_1701);
nand U338 (N_338,In_2009,In_1626);
nand U339 (N_339,In_570,In_97);
nand U340 (N_340,In_2316,In_2251);
or U341 (N_341,In_2068,In_647);
xor U342 (N_342,In_1065,In_273);
and U343 (N_343,In_2492,In_565);
and U344 (N_344,In_1333,In_190);
xnor U345 (N_345,In_2239,In_738);
and U346 (N_346,In_456,In_1028);
nand U347 (N_347,In_2234,In_1857);
and U348 (N_348,In_965,In_2304);
nor U349 (N_349,In_1667,In_2217);
or U350 (N_350,In_2161,In_1708);
nand U351 (N_351,In_76,In_1045);
or U352 (N_352,In_784,In_2127);
or U353 (N_353,In_689,In_1840);
nor U354 (N_354,In_2231,In_16);
nor U355 (N_355,In_1515,In_2375);
and U356 (N_356,In_205,In_881);
xnor U357 (N_357,In_92,In_792);
xor U358 (N_358,In_1229,In_905);
or U359 (N_359,In_997,In_724);
xnor U360 (N_360,In_313,In_2480);
xor U361 (N_361,In_989,In_1544);
nor U362 (N_362,In_1980,In_1519);
and U363 (N_363,In_781,In_608);
nand U364 (N_364,In_2175,In_2256);
nor U365 (N_365,In_862,In_1411);
or U366 (N_366,In_813,In_2430);
nand U367 (N_367,In_556,In_424);
nor U368 (N_368,In_1261,In_1014);
xor U369 (N_369,In_2269,In_1272);
nand U370 (N_370,In_444,In_770);
nand U371 (N_371,In_162,In_2266);
xor U372 (N_372,In_428,In_1057);
and U373 (N_373,In_544,In_1135);
nand U374 (N_374,In_415,In_1313);
nand U375 (N_375,In_1525,In_2402);
nor U376 (N_376,In_323,In_1431);
xor U377 (N_377,In_111,In_1381);
xor U378 (N_378,In_2258,In_376);
or U379 (N_379,In_1449,In_1106);
xor U380 (N_380,In_616,In_1226);
nor U381 (N_381,In_1193,In_311);
nand U382 (N_382,In_204,In_266);
nand U383 (N_383,In_814,In_966);
nor U384 (N_384,In_2399,In_1204);
nand U385 (N_385,In_1653,In_1602);
nand U386 (N_386,In_88,In_962);
and U387 (N_387,In_370,In_1063);
nor U388 (N_388,In_2351,In_871);
and U389 (N_389,In_1837,In_425);
and U390 (N_390,In_759,In_1552);
nor U391 (N_391,In_474,In_2153);
or U392 (N_392,In_1685,In_2081);
nand U393 (N_393,In_297,In_1645);
nor U394 (N_394,In_1427,In_134);
and U395 (N_395,In_1624,In_1596);
nor U396 (N_396,In_1696,In_1141);
or U397 (N_397,In_874,In_1924);
or U398 (N_398,In_212,In_133);
or U399 (N_399,In_2494,In_777);
xor U400 (N_400,In_493,In_112);
and U401 (N_401,In_2324,In_538);
xor U402 (N_402,In_1442,In_1481);
or U403 (N_403,In_442,In_1606);
xor U404 (N_404,In_2157,In_2232);
and U405 (N_405,In_2018,In_577);
or U406 (N_406,In_1108,In_1751);
nor U407 (N_407,In_585,In_2331);
xor U408 (N_408,In_913,In_1779);
nor U409 (N_409,In_2220,In_118);
xor U410 (N_410,In_931,In_1116);
xor U411 (N_411,In_773,In_2062);
and U412 (N_412,In_1958,In_876);
or U413 (N_413,In_2276,In_1396);
or U414 (N_414,In_127,In_557);
nor U415 (N_415,In_2082,In_353);
nor U416 (N_416,In_1401,In_1367);
xnor U417 (N_417,In_869,In_1232);
nor U418 (N_418,In_60,In_1965);
or U419 (N_419,In_235,In_2211);
xor U420 (N_420,In_1586,In_1973);
and U421 (N_421,In_1669,In_1982);
or U422 (N_422,In_2434,In_1896);
xor U423 (N_423,In_1995,In_227);
xor U424 (N_424,In_406,In_588);
and U425 (N_425,In_1743,In_2198);
nand U426 (N_426,In_509,In_1804);
nor U427 (N_427,In_1305,In_383);
nor U428 (N_428,In_1910,In_2138);
nor U429 (N_429,In_2487,In_2477);
xnor U430 (N_430,In_787,In_400);
and U431 (N_431,In_942,In_1222);
xnor U432 (N_432,In_252,In_2456);
nand U433 (N_433,In_1516,In_1534);
xnor U434 (N_434,In_1339,In_928);
or U435 (N_435,In_1475,In_51);
and U436 (N_436,In_1640,In_337);
xor U437 (N_437,In_2117,In_20);
and U438 (N_438,In_734,In_2142);
nor U439 (N_439,In_82,In_19);
nor U440 (N_440,In_748,In_57);
nand U441 (N_441,In_343,In_2439);
nor U442 (N_442,In_2028,In_1465);
nor U443 (N_443,In_2074,In_713);
or U444 (N_444,In_1621,In_2248);
nand U445 (N_445,In_1585,In_511);
xnor U446 (N_446,In_285,In_219);
or U447 (N_447,In_1018,In_482);
or U448 (N_448,In_240,In_1207);
xnor U449 (N_449,In_658,In_987);
or U450 (N_450,In_572,In_2458);
nand U451 (N_451,In_2453,In_727);
nand U452 (N_452,In_1592,In_1665);
nand U453 (N_453,In_1137,In_1246);
and U454 (N_454,In_2339,In_528);
or U455 (N_455,In_2250,In_1388);
or U456 (N_456,In_2338,In_1533);
and U457 (N_457,In_282,In_640);
xor U458 (N_458,In_2286,In_330);
xnor U459 (N_459,In_717,In_1455);
nor U460 (N_460,In_136,In_1459);
nand U461 (N_461,In_391,In_1278);
nand U462 (N_462,In_1445,In_1686);
or U463 (N_463,In_826,In_1472);
or U464 (N_464,In_1796,In_2094);
xor U465 (N_465,In_2415,In_1244);
nor U466 (N_466,In_2176,In_944);
or U467 (N_467,In_2291,In_1143);
nor U468 (N_468,In_1595,In_1799);
nand U469 (N_469,In_107,In_2281);
or U470 (N_470,In_2383,In_1186);
or U471 (N_471,In_123,In_279);
xor U472 (N_472,In_2499,In_2098);
and U473 (N_473,In_1841,In_995);
and U474 (N_474,In_1826,In_1697);
nor U475 (N_475,In_2036,In_1879);
or U476 (N_476,In_1130,In_253);
or U477 (N_477,In_64,In_304);
or U478 (N_478,In_1169,In_2448);
nand U479 (N_479,In_914,In_2131);
nor U480 (N_480,In_1907,In_614);
xor U481 (N_481,In_477,In_2493);
and U482 (N_482,In_1777,In_1403);
xnor U483 (N_483,In_1524,In_1884);
nand U484 (N_484,In_1875,In_1989);
or U485 (N_485,In_2245,In_1419);
nand U486 (N_486,In_25,In_1160);
and U487 (N_487,In_1927,In_1877);
and U488 (N_488,In_643,In_403);
nand U489 (N_489,In_932,In_750);
and U490 (N_490,In_680,In_165);
nand U491 (N_491,In_163,In_160);
nand U492 (N_492,In_703,In_1791);
or U493 (N_493,In_739,In_1258);
or U494 (N_494,In_308,In_1145);
or U495 (N_495,In_2061,In_1498);
and U496 (N_496,In_1221,In_974);
or U497 (N_497,In_2305,In_2099);
and U498 (N_498,In_412,In_893);
and U499 (N_499,In_1464,In_775);
nor U500 (N_500,In_555,In_270);
or U501 (N_501,In_2310,In_1324);
nand U502 (N_502,In_1659,In_648);
xor U503 (N_503,In_1577,In_1809);
or U504 (N_504,In_1767,In_1476);
or U505 (N_505,In_1874,In_27);
or U506 (N_506,In_1070,In_1898);
and U507 (N_507,In_1177,In_2468);
nand U508 (N_508,In_1786,In_693);
and U509 (N_509,In_243,In_963);
nor U510 (N_510,In_1503,In_1615);
nand U511 (N_511,In_2052,In_1460);
nand U512 (N_512,In_43,In_1510);
or U513 (N_513,In_2236,In_2335);
xnor U514 (N_514,In_617,In_1554);
nand U515 (N_515,In_1774,In_431);
or U516 (N_516,In_37,In_1271);
or U517 (N_517,In_2149,In_801);
xnor U518 (N_518,In_100,In_650);
nand U519 (N_519,In_238,In_1240);
nand U520 (N_520,In_2021,In_1122);
xor U521 (N_521,In_592,In_621);
xnor U522 (N_522,In_568,In_979);
and U523 (N_523,In_1086,In_1564);
or U524 (N_524,In_268,In_2193);
and U525 (N_525,In_491,In_122);
xor U526 (N_526,In_329,In_583);
and U527 (N_527,In_2307,In_927);
nor U528 (N_528,In_1280,In_747);
nor U529 (N_529,In_808,In_1575);
and U530 (N_530,In_462,In_1720);
and U531 (N_531,In_1680,In_1350);
or U532 (N_532,In_953,In_686);
or U533 (N_533,In_1110,In_257);
xnor U534 (N_534,In_1104,In_481);
nand U535 (N_535,In_697,In_1302);
or U536 (N_536,In_1833,In_1239);
and U537 (N_537,In_224,In_831);
nor U538 (N_538,In_2134,In_654);
nor U539 (N_539,In_2443,In_1032);
and U540 (N_540,In_2469,In_2012);
nand U541 (N_541,In_1678,In_1807);
and U542 (N_542,In_1443,In_2341);
xnor U543 (N_543,In_1225,In_384);
nor U544 (N_544,In_755,In_2139);
and U545 (N_545,In_220,In_2390);
nor U546 (N_546,In_1468,In_2429);
and U547 (N_547,In_1165,In_489);
and U548 (N_548,In_1374,In_984);
and U549 (N_549,In_1867,In_901);
and U550 (N_550,In_2024,In_1479);
or U551 (N_551,In_679,In_587);
nand U552 (N_552,In_1015,In_2392);
xnor U553 (N_553,In_1167,In_241);
nand U554 (N_554,In_2045,In_2047);
nand U555 (N_555,In_485,In_1715);
or U556 (N_556,In_1357,In_167);
nor U557 (N_557,In_1132,In_1994);
nor U558 (N_558,In_1737,In_2118);
nand U559 (N_559,In_722,In_507);
and U560 (N_560,In_85,In_1347);
xnor U561 (N_561,In_699,In_626);
xor U562 (N_562,In_609,In_1573);
xnor U563 (N_563,In_1781,In_2203);
nor U564 (N_564,In_798,In_998);
xnor U565 (N_565,In_1912,In_1738);
xnor U566 (N_566,In_2162,In_603);
nor U567 (N_567,In_1352,In_91);
nand U568 (N_568,In_820,In_1864);
and U569 (N_569,In_180,In_633);
and U570 (N_570,In_861,In_1855);
xnor U571 (N_571,In_2003,In_772);
nor U572 (N_572,In_2288,In_138);
nand U573 (N_573,In_1022,In_237);
nor U574 (N_574,In_2426,In_1485);
nand U575 (N_575,In_466,In_2406);
and U576 (N_576,In_1808,In_923);
nand U577 (N_577,In_1050,In_749);
and U578 (N_578,In_1581,In_1296);
nor U579 (N_579,In_1096,In_1462);
nor U580 (N_580,In_1456,In_1762);
xor U581 (N_581,In_346,In_2189);
or U582 (N_582,In_1379,In_2432);
or U583 (N_583,In_373,In_988);
or U584 (N_584,In_327,In_1267);
or U585 (N_585,In_1262,In_2297);
and U586 (N_586,In_2466,In_1747);
xnor U587 (N_587,In_848,In_1932);
and U588 (N_588,In_1452,In_11);
xor U589 (N_589,In_1087,In_1330);
nand U590 (N_590,In_552,In_445);
and U591 (N_591,In_15,In_2005);
or U592 (N_592,In_903,In_1338);
nand U593 (N_593,In_522,In_1019);
or U594 (N_594,In_1251,In_2327);
nor U595 (N_595,In_1590,In_1337);
and U596 (N_596,In_1436,In_164);
xor U597 (N_597,In_1260,In_1415);
and U598 (N_598,In_341,In_1531);
xor U599 (N_599,In_1517,In_629);
nor U600 (N_600,In_2352,In_2411);
nand U601 (N_601,In_993,In_271);
nand U602 (N_602,In_1514,In_2476);
nor U603 (N_603,In_1360,In_1639);
or U604 (N_604,In_1992,In_1657);
nor U605 (N_605,In_49,In_600);
nand U606 (N_606,In_1359,In_1375);
nand U607 (N_607,In_539,In_410);
or U608 (N_608,In_1764,In_1288);
or U609 (N_609,In_1920,In_357);
xnor U610 (N_610,In_661,In_2049);
or U611 (N_611,In_371,In_322);
xnor U612 (N_612,In_2326,In_2330);
xnor U613 (N_613,In_436,In_188);
or U614 (N_614,In_887,In_2158);
or U615 (N_615,In_1854,In_1813);
nor U616 (N_616,In_175,In_746);
xnor U617 (N_617,In_1497,In_1282);
and U618 (N_618,In_201,In_929);
and U619 (N_619,In_1126,In_1906);
xnor U620 (N_620,In_2067,In_1248);
and U621 (N_621,In_1105,In_1129);
and U622 (N_622,In_379,In_1410);
nand U623 (N_623,In_1035,In_244);
nand U624 (N_624,In_569,In_815);
nand U625 (N_625,In_286,In_1351);
nand U626 (N_626,In_77,In_409);
xnor U627 (N_627,In_300,In_1750);
and U628 (N_628,In_1661,In_1865);
nand U629 (N_629,In_574,In_2200);
or U630 (N_630,In_2407,In_514);
nor U631 (N_631,In_1007,In_71);
nor U632 (N_632,In_1984,In_17);
nand U633 (N_633,In_594,In_1759);
and U634 (N_634,In_23,In_81);
nand U635 (N_635,In_356,In_1376);
and U636 (N_636,In_38,In_670);
nand U637 (N_637,In_143,In_1684);
or U638 (N_638,In_139,In_1889);
xnor U639 (N_639,In_275,In_2428);
nor U640 (N_640,In_469,In_1218);
nor U641 (N_641,In_389,In_776);
or U642 (N_642,In_1366,In_2457);
and U643 (N_643,In_1967,In_560);
or U644 (N_644,In_991,In_1817);
nor U645 (N_645,In_10,In_84);
nor U646 (N_646,In_261,In_1223);
or U647 (N_647,In_1276,In_2361);
nor U648 (N_648,In_2066,In_375);
or U649 (N_649,In_1925,In_1726);
nor U650 (N_650,In_2207,In_1763);
nand U651 (N_651,In_182,In_911);
nor U652 (N_652,In_1589,In_1068);
or U653 (N_653,In_1506,In_1622);
nor U654 (N_654,In_206,In_1843);
nor U655 (N_655,In_2329,In_1986);
or U656 (N_656,In_113,In_1114);
nand U657 (N_657,In_854,In_1237);
xnor U658 (N_658,In_809,In_676);
nand U659 (N_659,In_1823,In_1845);
nand U660 (N_660,In_1991,In_1563);
xnor U661 (N_661,In_2164,In_2011);
or U662 (N_662,In_121,In_1679);
nand U663 (N_663,In_604,In_74);
or U664 (N_664,In_1293,In_1730);
nand U665 (N_665,In_2364,In_2301);
xor U666 (N_666,In_908,In_810);
xnor U667 (N_667,In_766,In_1253);
xnor U668 (N_668,In_579,In_2354);
nand U669 (N_669,In_949,In_1242);
nor U670 (N_670,In_1698,In_2093);
xor U671 (N_671,In_1971,In_2272);
and U672 (N_672,In_2097,In_1732);
nor U673 (N_673,In_1744,In_681);
xnor U674 (N_674,In_2202,In_1692);
nor U675 (N_675,In_711,In_2014);
nor U676 (N_676,In_2079,In_22);
or U677 (N_677,In_1102,In_114);
or U678 (N_678,In_2420,In_45);
nand U679 (N_679,In_1693,In_1097);
or U680 (N_680,In_712,In_281);
and U681 (N_681,In_2471,In_1916);
nor U682 (N_682,In_1309,In_380);
xor U683 (N_683,In_1094,In_567);
nand U684 (N_684,In_2029,In_2169);
nand U685 (N_685,In_109,In_2141);
or U686 (N_686,In_2385,In_68);
xnor U687 (N_687,In_853,In_115);
and U688 (N_688,In_2321,In_429);
nand U689 (N_689,In_1943,In_471);
nand U690 (N_690,In_720,In_718);
or U691 (N_691,In_2073,In_2459);
xor U692 (N_692,In_2435,In_812);
and U693 (N_693,In_414,In_1336);
or U694 (N_694,In_2104,In_210);
nor U695 (N_695,In_1915,In_324);
and U696 (N_696,In_721,In_1572);
nand U697 (N_697,In_504,In_2222);
and U698 (N_698,In_1603,In_1546);
nand U699 (N_699,In_1883,In_1987);
or U700 (N_700,In_1950,In_939);
nor U701 (N_701,In_1728,In_1856);
and U702 (N_702,In_2379,In_2002);
nand U703 (N_703,In_484,In_857);
and U704 (N_704,In_1488,In_407);
and U705 (N_705,In_1215,In_518);
and U706 (N_706,In_1227,In_620);
nor U707 (N_707,In_941,In_907);
and U708 (N_708,In_1569,In_783);
nor U709 (N_709,In_2488,In_62);
and U710 (N_710,In_933,In_1724);
nor U711 (N_711,In_2054,In_2441);
nand U712 (N_712,In_1202,In_1195);
nor U713 (N_713,In_1217,In_2244);
nor U714 (N_714,In_836,In_1250);
nor U715 (N_715,In_1582,In_2380);
xnor U716 (N_716,In_288,In_1527);
and U717 (N_717,In_1049,In_1406);
and U718 (N_718,In_2302,In_1213);
and U719 (N_719,In_769,In_1643);
nand U720 (N_720,In_628,In_108);
and U721 (N_721,In_1409,In_515);
nor U722 (N_722,In_374,In_1080);
and U723 (N_723,In_87,In_1549);
nor U724 (N_724,In_1719,In_870);
nand U725 (N_725,In_2280,In_2463);
nor U726 (N_726,In_2475,In_187);
nor U727 (N_727,In_226,In_2255);
xor U728 (N_728,In_126,In_1576);
xnor U729 (N_729,In_1556,In_259);
nand U730 (N_730,In_104,In_2366);
or U731 (N_731,In_1900,In_1948);
xor U732 (N_732,In_1238,In_506);
nor U733 (N_733,In_2464,In_1977);
nand U734 (N_734,In_996,In_1390);
nand U735 (N_735,In_1400,In_1782);
nand U736 (N_736,In_144,In_1897);
nor U737 (N_737,In_443,In_1691);
nand U738 (N_738,In_1660,In_1828);
nor U739 (N_739,In_723,In_2373);
or U740 (N_740,In_2350,In_229);
or U741 (N_741,In_2267,In_1518);
nand U742 (N_742,In_223,In_864);
or U743 (N_743,In_1307,In_1101);
or U744 (N_744,In_2483,In_2165);
nand U745 (N_745,In_763,In_2376);
nand U746 (N_746,In_269,In_1610);
xnor U747 (N_747,In_47,In_1323);
nand U748 (N_748,In_131,In_1386);
nor U749 (N_749,In_1341,In_2026);
nor U750 (N_750,In_1998,In_365);
or U751 (N_751,In_363,In_2182);
and U752 (N_752,In_256,In_1937);
nand U753 (N_753,In_2370,In_352);
xnor U754 (N_754,In_1127,In_55);
xor U755 (N_755,In_1477,In_1904);
and U756 (N_756,In_1816,In_2284);
nand U757 (N_757,In_806,In_1757);
and U758 (N_758,In_2365,In_147);
or U759 (N_759,In_2007,In_2179);
and U760 (N_760,In_2034,In_2006);
or U761 (N_761,In_1528,In_1181);
nand U762 (N_762,In_1038,In_731);
nand U763 (N_763,In_2223,In_214);
or U764 (N_764,In_2259,In_2219);
nor U765 (N_765,In_900,In_1733);
nand U766 (N_766,In_1945,In_1600);
or U767 (N_767,In_1899,In_2270);
nand U768 (N_768,In_2311,In_957);
nor U769 (N_769,In_2486,In_1257);
xnor U770 (N_770,In_1220,In_845);
nor U771 (N_771,In_2041,In_2050);
nand U772 (N_772,In_1343,In_1818);
or U773 (N_773,In_752,In_2382);
nand U774 (N_774,In_818,In_2268);
and U775 (N_775,In_142,In_2423);
xnor U776 (N_776,In_1847,In_2072);
nor U777 (N_777,In_1345,In_732);
nand U778 (N_778,In_1059,In_8);
nor U779 (N_779,In_2490,In_99);
or U780 (N_780,In_2313,In_1848);
and U781 (N_781,In_393,In_2349);
nor U782 (N_782,In_203,In_420);
xor U783 (N_783,In_1946,In_378);
xnor U784 (N_784,In_1058,In_631);
and U785 (N_785,In_1630,In_895);
or U786 (N_786,In_760,In_885);
nand U787 (N_787,In_2333,In_580);
xnor U788 (N_788,In_1978,In_1947);
nor U789 (N_789,In_1663,In_1308);
xor U790 (N_790,In_541,In_172);
nor U791 (N_791,In_1321,In_2126);
or U792 (N_792,In_632,In_529);
nor U793 (N_793,In_2440,In_1557);
nand U794 (N_794,In_1316,In_437);
nor U795 (N_795,In_196,In_563);
nor U796 (N_796,In_890,In_1256);
or U797 (N_797,In_531,In_1054);
and U798 (N_798,In_2377,In_42);
nand U799 (N_799,In_1990,In_231);
and U800 (N_800,In_155,In_2386);
nand U801 (N_801,In_1120,In_1149);
and U802 (N_802,In_696,In_2253);
nor U803 (N_803,In_564,In_31);
nand U804 (N_804,In_1523,In_2143);
xor U805 (N_805,In_1344,In_1441);
xnor U806 (N_806,In_2168,In_110);
nand U807 (N_807,In_1422,In_312);
nand U808 (N_808,In_795,In_1066);
xnor U809 (N_809,In_46,In_649);
xor U810 (N_810,In_1397,In_1721);
or U811 (N_811,In_2460,In_2292);
and U812 (N_812,In_517,In_1789);
nand U813 (N_813,In_2235,In_48);
nor U814 (N_814,In_1694,In_1064);
nand U815 (N_815,In_1770,In_756);
or U816 (N_816,In_591,In_1322);
nand U817 (N_817,In_873,In_1702);
nand U818 (N_818,In_1778,In_1241);
or U819 (N_819,In_315,In_662);
or U820 (N_820,In_2381,In_459);
or U821 (N_821,In_53,In_586);
nand U822 (N_822,In_1053,In_128);
or U823 (N_823,In_2413,In_994);
nand U824 (N_824,In_1429,In_166);
or U825 (N_825,In_1895,In_1954);
xnor U826 (N_826,In_691,In_470);
or U827 (N_827,In_177,In_276);
xnor U828 (N_828,In_1148,In_1500);
nand U829 (N_829,In_347,In_2044);
and U830 (N_830,In_40,In_1929);
and U831 (N_831,In_1710,In_1756);
or U832 (N_832,In_1619,In_841);
and U833 (N_833,In_967,In_1121);
nand U834 (N_834,In_1583,In_1416);
nor U835 (N_835,In_1349,In_1407);
or U836 (N_836,In_975,In_239);
or U837 (N_837,In_59,In_296);
nand U838 (N_838,In_765,In_2084);
and U839 (N_839,In_2229,In_1031);
nand U840 (N_840,In_951,In_1450);
or U841 (N_841,In_1548,In_2053);
or U842 (N_842,In_1369,In_1005);
nor U843 (N_843,In_348,In_447);
nor U844 (N_844,In_1365,In_2218);
and U845 (N_845,In_1291,In_2057);
xor U846 (N_846,In_2035,In_1960);
or U847 (N_847,In_948,In_1682);
or U848 (N_848,In_623,In_497);
xor U849 (N_849,In_372,In_2360);
xor U850 (N_850,In_946,In_158);
nor U851 (N_851,In_2221,In_1189);
nor U852 (N_852,In_1099,In_1310);
xor U853 (N_853,In_140,In_1901);
xnor U854 (N_854,In_408,In_1301);
or U855 (N_855,In_1935,In_328);
nand U856 (N_856,In_2039,In_2298);
and U857 (N_857,In_1736,In_314);
xnor U858 (N_858,In_0,In_1326);
xor U859 (N_859,In_1908,In_1249);
and U860 (N_860,In_1902,In_1259);
and U861 (N_861,In_1180,In_1284);
and U862 (N_862,In_1283,In_2116);
nand U863 (N_863,In_457,In_2252);
or U864 (N_864,In_1075,In_1537);
or U865 (N_865,In_1565,In_451);
xnor U866 (N_866,In_2069,In_2419);
and U867 (N_867,In_1797,In_532);
xor U868 (N_868,In_1672,In_1034);
nand U869 (N_869,In_1270,In_2040);
and U870 (N_870,In_1062,In_596);
or U871 (N_871,In_1228,In_1157);
or U872 (N_872,In_527,In_1067);
nor U873 (N_873,In_1520,In_687);
nor U874 (N_874,In_1972,In_1734);
nand U875 (N_875,In_2425,In_290);
or U876 (N_876,In_1741,In_1803);
nor U877 (N_877,In_501,In_151);
nand U878 (N_878,In_1496,In_367);
nand U879 (N_879,In_2137,In_726);
and U880 (N_880,In_39,In_1134);
and U881 (N_881,In_1962,In_86);
or U882 (N_882,In_651,In_2303);
and U883 (N_883,In_675,In_2296);
xor U884 (N_884,In_736,In_978);
nor U885 (N_885,In_427,In_986);
nand U886 (N_886,In_886,In_1083);
nand U887 (N_887,In_338,In_1560);
nor U888 (N_888,In_1959,In_919);
or U889 (N_889,In_1790,In_321);
and U890 (N_890,In_2185,In_1851);
xnor U891 (N_891,In_54,In_2125);
and U892 (N_892,In_265,In_1666);
or U893 (N_893,In_1711,In_1089);
xor U894 (N_894,In_1354,In_685);
nand U895 (N_895,In_844,In_1041);
and U896 (N_896,In_897,In_2031);
xor U897 (N_897,In_316,In_129);
xnor U898 (N_898,In_796,In_2016);
and U899 (N_899,In_1983,In_1191);
or U900 (N_900,In_2101,In_360);
or U901 (N_901,In_1812,In_395);
nor U902 (N_902,In_145,In_2037);
nand U903 (N_903,In_267,In_2205);
and U904 (N_904,In_973,In_2378);
xor U905 (N_905,In_1432,In_999);
nand U906 (N_906,In_198,In_1594);
or U907 (N_907,In_1806,In_335);
xor U908 (N_908,In_1555,In_2090);
xnor U909 (N_909,In_1490,In_1783);
and U910 (N_910,In_1934,In_671);
nor U911 (N_911,In_1718,In_1368);
xnor U912 (N_912,In_262,In_630);
nand U913 (N_913,In_1938,In_2277);
nand U914 (N_914,In_1511,In_1236);
or U915 (N_915,In_30,In_2342);
xor U916 (N_916,In_2089,In_2115);
nand U917 (N_917,In_480,In_829);
and U918 (N_918,In_1183,In_2022);
or U919 (N_919,In_838,In_2262);
nand U920 (N_920,In_1651,In_320);
nand U921 (N_921,In_96,In_639);
xor U922 (N_922,In_2397,In_1618);
and U923 (N_923,In_688,In_35);
xnor U924 (N_924,In_1478,In_1644);
nor U925 (N_925,In_106,In_2032);
nand U926 (N_926,In_1933,In_1433);
and U927 (N_927,In_877,In_197);
nor U928 (N_928,In_1623,In_1405);
or U929 (N_929,In_299,In_1695);
xnor U930 (N_930,In_354,In_985);
and U931 (N_931,In_1739,In_455);
nand U932 (N_932,In_1171,In_865);
or U933 (N_933,In_2124,In_1598);
xor U934 (N_934,In_1968,In_2092);
nor U935 (N_935,In_754,In_1846);
xnor U936 (N_936,In_1361,In_1002);
or U937 (N_937,In_487,In_1922);
xor U938 (N_938,In_1243,In_694);
xor U939 (N_939,In_2145,In_263);
and U940 (N_940,In_1164,In_725);
and U941 (N_941,In_878,In_1412);
xor U942 (N_942,In_582,In_1794);
nand U943 (N_943,In_1853,In_1233);
nand U944 (N_944,In_751,In_1048);
nand U945 (N_945,In_1492,In_2201);
and U946 (N_946,In_1085,In_1413);
or U947 (N_947,In_1636,In_2146);
nand U948 (N_948,In_2265,In_1705);
nand U949 (N_949,In_65,In_1570);
or U950 (N_950,In_319,In_1037);
nand U951 (N_951,In_1003,In_607);
nor U952 (N_952,In_605,In_295);
and U953 (N_953,In_548,In_508);
nand U954 (N_954,In_171,In_1402);
nor U955 (N_955,In_1118,In_1269);
or U956 (N_956,In_677,In_892);
xor U957 (N_957,In_318,In_786);
nor U958 (N_958,In_2371,In_12);
nand U959 (N_959,In_2418,In_1480);
xnor U960 (N_960,In_302,In_1208);
xor U961 (N_961,In_1893,In_2008);
nand U962 (N_962,In_705,In_1830);
nand U963 (N_963,In_441,In_1047);
nor U964 (N_964,In_7,In_185);
and U965 (N_965,In_779,In_2498);
and U966 (N_966,In_1076,In_1609);
nor U967 (N_967,In_2334,In_2467);
xnor U968 (N_968,In_1541,In_1785);
xor U969 (N_969,In_1776,In_922);
nand U970 (N_970,In_2140,In_1311);
and U971 (N_971,In_1713,In_850);
and U972 (N_972,In_1173,In_891);
or U973 (N_973,In_1755,In_2363);
and U974 (N_974,In_782,In_1831);
and U975 (N_975,In_1712,In_2151);
and U976 (N_976,In_1069,In_272);
nand U977 (N_977,In_492,In_368);
nor U978 (N_978,In_1880,In_2318);
nor U979 (N_979,In_664,In_14);
nand U980 (N_980,In_778,In_1688);
nand U981 (N_981,In_2408,In_58);
nand U982 (N_982,In_1029,In_94);
nor U983 (N_983,In_510,In_1112);
or U984 (N_984,In_1377,In_1944);
and U985 (N_985,In_401,In_13);
nand U986 (N_986,In_852,In_2233);
nor U987 (N_987,In_917,In_904);
xor U988 (N_988,In_2261,In_2414);
or U989 (N_989,In_1231,In_1006);
nand U990 (N_990,In_1212,In_1676);
xor U991 (N_991,In_1836,In_2010);
nand U992 (N_992,In_1470,In_44);
nor U993 (N_993,In_1707,In_1550);
xnor U994 (N_994,In_637,In_659);
nand U995 (N_995,In_9,In_627);
nor U996 (N_996,In_1545,In_331);
and U997 (N_997,In_137,In_422);
xor U998 (N_998,In_1418,In_612);
nor U999 (N_999,In_521,In_1873);
and U1000 (N_1000,In_1835,In_2215);
nor U1001 (N_1001,In_634,In_618);
nor U1002 (N_1002,In_340,In_301);
xnor U1003 (N_1003,In_1863,In_2442);
nand U1004 (N_1004,In_657,In_719);
xnor U1005 (N_1005,In_1793,In_1428);
nor U1006 (N_1006,In_1457,In_1073);
or U1007 (N_1007,In_2056,In_465);
nand U1008 (N_1008,In_2283,In_2243);
nor U1009 (N_1009,In_1424,In_157);
nand U1010 (N_1010,In_103,In_1870);
nor U1011 (N_1011,In_152,In_2133);
xor U1012 (N_1012,In_141,In_1077);
xor U1013 (N_1013,In_2396,In_1613);
nand U1014 (N_1014,In_1662,In_1001);
nand U1015 (N_1015,In_1140,In_1658);
and U1016 (N_1016,In_34,In_2209);
or U1017 (N_1017,In_690,In_2290);
xor U1018 (N_1018,In_1334,In_1930);
or U1019 (N_1019,In_1844,In_1027);
nor U1020 (N_1020,In_519,In_388);
xor U1021 (N_1021,In_2130,In_952);
and U1022 (N_1022,In_542,In_2226);
xor U1023 (N_1023,In_1147,In_1505);
nor U1024 (N_1024,In_381,In_432);
and U1025 (N_1025,In_1532,In_1210);
xnor U1026 (N_1026,In_1052,In_811);
or U1027 (N_1027,In_1827,In_2180);
and U1028 (N_1028,In_249,In_867);
xnor U1029 (N_1029,In_1607,In_1787);
nand U1030 (N_1030,In_1454,In_307);
xor U1031 (N_1031,In_2055,In_117);
nand U1032 (N_1032,In_653,In_866);
nor U1033 (N_1033,In_463,In_168);
nor U1034 (N_1034,In_1093,In_793);
and U1035 (N_1035,In_150,In_2474);
nor U1036 (N_1036,In_1332,In_1300);
nand U1037 (N_1037,In_601,In_2096);
xor U1038 (N_1038,In_1513,In_2085);
xor U1039 (N_1039,In_2214,In_274);
xor U1040 (N_1040,In_860,In_1765);
or U1041 (N_1041,In_1752,In_2394);
and U1042 (N_1042,In_1088,In_1012);
and U1043 (N_1043,In_310,In_200);
nand U1044 (N_1044,In_192,In_1342);
and U1045 (N_1045,In_1380,In_1115);
xor U1046 (N_1046,In_2156,In_1281);
xor U1047 (N_1047,In_990,In_597);
nor U1048 (N_1048,In_1286,In_2183);
nor U1049 (N_1049,In_1404,In_1483);
and U1050 (N_1050,In_2401,In_816);
and U1051 (N_1051,In_494,In_2395);
or U1052 (N_1052,In_516,In_937);
nor U1053 (N_1053,In_411,In_1158);
xor U1054 (N_1054,In_130,In_78);
nand U1055 (N_1055,In_2095,In_1348);
xor U1056 (N_1056,In_448,In_1435);
xnor U1057 (N_1057,In_1414,In_1638);
nor U1058 (N_1058,In_1327,In_1501);
nand U1059 (N_1059,In_1894,In_669);
nor U1060 (N_1060,In_1209,In_2171);
nand U1061 (N_1061,In_1275,In_326);
nand U1062 (N_1062,In_369,In_745);
or U1063 (N_1063,In_843,In_1266);
nand U1064 (N_1064,In_1521,In_910);
nand U1065 (N_1065,In_1683,In_24);
or U1066 (N_1066,In_1364,In_622);
and U1067 (N_1067,In_1092,In_1561);
nor U1068 (N_1068,In_2048,In_1166);
nor U1069 (N_1069,In_619,In_454);
or U1070 (N_1070,In_61,In_2289);
nor U1071 (N_1071,In_1491,In_2273);
or U1072 (N_1072,In_2186,In_1608);
or U1073 (N_1073,In_1387,In_1612);
xnor U1074 (N_1074,In_1866,In_894);
nor U1075 (N_1075,In_1509,In_1182);
and U1076 (N_1076,In_960,In_1819);
and U1077 (N_1077,In_2064,In_2123);
xnor U1078 (N_1078,In_2455,In_1159);
or U1079 (N_1079,In_502,In_924);
nand U1080 (N_1080,In_2398,In_549);
and U1081 (N_1081,In_2347,In_1742);
nor U1082 (N_1082,In_1287,In_228);
nor U1083 (N_1083,In_2478,In_655);
nor U1084 (N_1084,In_2263,In_148);
or U1085 (N_1085,In_1690,In_1098);
and U1086 (N_1086,In_1393,In_189);
and U1087 (N_1087,In_2300,In_598);
xnor U1088 (N_1088,In_1061,In_2080);
nand U1089 (N_1089,In_2004,In_2103);
or U1090 (N_1090,In_350,In_1587);
or U1091 (N_1091,In_554,In_79);
and U1092 (N_1092,In_1190,In_1558);
and U1093 (N_1093,In_2019,In_1539);
and U1094 (N_1094,In_2063,In_33);
xor U1095 (N_1095,In_2355,In_366);
xor U1096 (N_1096,In_2030,In_2409);
or U1097 (N_1097,In_2412,In_120);
nand U1098 (N_1098,In_1346,In_1289);
nand U1099 (N_1099,In_1111,In_2083);
xor U1100 (N_1100,In_613,In_1320);
nand U1101 (N_1101,In_1735,In_2147);
nand U1102 (N_1102,In_2247,In_2060);
xnor U1103 (N_1103,In_1647,In_2452);
xnor U1104 (N_1104,In_1133,In_624);
or U1105 (N_1105,In_715,In_450);
xor U1106 (N_1106,In_344,In_161);
and U1107 (N_1107,In_2114,In_803);
and U1108 (N_1108,In_2374,In_486);
nand U1109 (N_1109,In_2451,In_1461);
and U1110 (N_1110,In_543,In_2190);
and U1111 (N_1111,In_217,In_1103);
or U1112 (N_1112,In_1355,In_2150);
xor U1113 (N_1113,In_2181,In_566);
nor U1114 (N_1114,In_935,In_2405);
and U1115 (N_1115,In_1858,In_824);
nor U1116 (N_1116,In_1473,In_1040);
nand U1117 (N_1117,In_1185,In_1886);
or U1118 (N_1118,In_2023,In_396);
nand U1119 (N_1119,In_1849,In_1290);
or U1120 (N_1120,In_102,In_2228);
or U1121 (N_1121,In_791,In_1117);
nor U1122 (N_1122,In_992,In_2384);
nor U1123 (N_1123,In_2446,In_728);
nand U1124 (N_1124,In_250,In_325);
and U1125 (N_1125,In_467,In_2111);
or U1126 (N_1126,In_959,In_1952);
and U1127 (N_1127,In_2359,In_2496);
nand U1128 (N_1128,In_790,In_1175);
nand U1129 (N_1129,In_561,In_1547);
and U1130 (N_1130,In_1458,In_553);
nor U1131 (N_1131,In_283,In_1042);
xnor U1132 (N_1132,In_2184,In_1909);
and U1133 (N_1133,In_832,In_1353);
nand U1134 (N_1134,In_1650,In_1);
and U1135 (N_1135,In_2148,In_213);
nor U1136 (N_1136,In_1408,In_2416);
nor U1137 (N_1137,In_1979,In_823);
nand U1138 (N_1138,In_2246,In_287);
nor U1139 (N_1139,In_2122,In_176);
or U1140 (N_1140,In_1026,In_1649);
xor U1141 (N_1141,In_1614,In_954);
nor U1142 (N_1142,In_540,In_879);
nor U1143 (N_1143,In_358,In_921);
or U1144 (N_1144,In_2107,In_1312);
and U1145 (N_1145,In_418,In_2241);
nor U1146 (N_1146,In_920,In_1914);
nand U1147 (N_1147,In_1340,In_426);
and U1148 (N_1148,In_1508,In_1474);
nand U1149 (N_1149,In_839,In_1362);
xnor U1150 (N_1150,In_1024,In_1604);
and U1151 (N_1151,In_2322,In_1043);
and U1152 (N_1152,In_2462,In_2287);
nor U1153 (N_1153,In_940,In_1913);
and U1154 (N_1154,In_1444,In_704);
xnor U1155 (N_1155,In_968,In_2152);
nand U1156 (N_1156,In_2070,In_2088);
nor U1157 (N_1157,In_535,In_512);
xor U1158 (N_1158,In_1011,In_305);
nor U1159 (N_1159,In_1981,In_534);
xnor U1160 (N_1160,In_707,In_1004);
nand U1161 (N_1161,In_500,In_2170);
and U1162 (N_1162,In_1219,In_159);
nand U1163 (N_1163,In_2421,In_1200);
nand U1164 (N_1164,In_1535,In_2197);
and U1165 (N_1165,In_156,In_1192);
nand U1166 (N_1166,In_646,In_2199);
xnor U1167 (N_1167,In_1154,In_1859);
nand U1168 (N_1168,In_251,In_1953);
xor U1169 (N_1169,In_1522,In_842);
and U1170 (N_1170,In_1976,In_744);
xnor U1171 (N_1171,In_1822,In_1123);
and U1172 (N_1172,In_768,In_1842);
xor U1173 (N_1173,In_2128,In_547);
or U1174 (N_1174,In_1654,In_859);
xnor U1175 (N_1175,In_2160,In_851);
nor U1176 (N_1176,In_1810,In_625);
nand U1177 (N_1177,In_1298,In_1821);
and U1178 (N_1178,In_90,In_435);
or U1179 (N_1179,In_1466,In_2212);
or U1180 (N_1180,In_1230,In_695);
xor U1181 (N_1181,In_2136,In_1430);
nand U1182 (N_1182,In_1749,In_1795);
or U1183 (N_1183,In_292,In_2224);
and U1184 (N_1184,In_956,In_69);
nor U1185 (N_1185,In_1664,In_1451);
xor U1186 (N_1186,In_452,In_221);
or U1187 (N_1187,In_1373,In_245);
nand U1188 (N_1188,In_575,In_1805);
and U1189 (N_1189,In_971,In_248);
and U1190 (N_1190,In_1363,In_1591);
and U1191 (N_1191,In_1633,In_706);
nor U1192 (N_1192,In_483,In_936);
nand U1193 (N_1193,In_526,In_545);
or U1194 (N_1194,In_701,In_399);
xor U1195 (N_1195,In_1328,In_1273);
and U1196 (N_1196,In_1297,In_362);
and U1197 (N_1197,In_947,In_835);
xnor U1198 (N_1198,In_1627,In_1637);
nand U1199 (N_1199,In_802,In_682);
xnor U1200 (N_1200,In_1044,In_1722);
xnor U1201 (N_1201,In_636,In_1489);
nor U1202 (N_1202,In_1949,In_1566);
nor U1203 (N_1203,In_825,In_2144);
or U1204 (N_1204,In_2135,In_1234);
nor U1205 (N_1205,In_1704,In_361);
xor U1206 (N_1206,In_716,In_124);
xnor U1207 (N_1207,In_1574,In_666);
xor U1208 (N_1208,In_154,In_882);
and U1209 (N_1209,In_1463,In_1655);
or U1210 (N_1210,In_209,In_2431);
xnor U1211 (N_1211,In_733,In_2225);
and U1212 (N_1212,In_499,In_2306);
nand U1213 (N_1213,In_1656,In_2159);
or U1214 (N_1214,In_1211,In_496);
nor U1215 (N_1215,In_1975,In_525);
xnor U1216 (N_1216,In_530,In_1673);
xnor U1217 (N_1217,In_1584,In_2076);
or U1218 (N_1218,In_1605,In_1095);
and U1219 (N_1219,In_1559,In_1625);
or U1220 (N_1220,In_1670,In_546);
xor U1221 (N_1221,In_461,In_146);
and U1222 (N_1222,In_2194,In_1862);
or U1223 (N_1223,In_339,In_1878);
and U1224 (N_1224,In_1677,In_1398);
xnor U1225 (N_1225,In_774,In_95);
and U1226 (N_1226,In_1885,In_1773);
nand U1227 (N_1227,In_1245,In_906);
or U1228 (N_1228,In_645,In_2391);
xor U1229 (N_1229,In_1617,In_1815);
and U1230 (N_1230,In_1372,In_382);
and U1231 (N_1231,In_610,In_402);
nand U1232 (N_1232,In_386,In_1008);
xor U1233 (N_1233,In_359,In_1629);
nand U1234 (N_1234,In_1421,In_1188);
nand U1235 (N_1235,In_800,In_2102);
nand U1236 (N_1236,In_1502,In_208);
nand U1237 (N_1237,In_1538,In_692);
nand U1238 (N_1238,In_1494,In_1919);
nand U1239 (N_1239,In_191,In_1499);
nor U1240 (N_1240,In_101,In_236);
xnor U1241 (N_1241,In_1802,In_1039);
nor U1242 (N_1242,In_1079,In_1021);
nand U1243 (N_1243,In_149,In_2436);
and U1244 (N_1244,In_1820,In_1314);
nand U1245 (N_1245,In_1013,In_837);
and U1246 (N_1246,In_2495,In_2346);
nand U1247 (N_1247,In_1888,In_1709);
xor U1248 (N_1248,In_1084,In_1423);
xnor U1249 (N_1249,In_1761,In_289);
nand U1250 (N_1250,In_1123,In_101);
xnor U1251 (N_1251,In_306,In_2433);
nand U1252 (N_1252,In_450,In_495);
nor U1253 (N_1253,In_2332,In_563);
xor U1254 (N_1254,In_1453,In_2344);
xor U1255 (N_1255,In_478,In_2033);
xnor U1256 (N_1256,In_12,In_117);
nand U1257 (N_1257,In_1198,In_418);
xor U1258 (N_1258,In_608,In_729);
xor U1259 (N_1259,In_1794,In_714);
or U1260 (N_1260,In_384,In_515);
xnor U1261 (N_1261,In_2320,In_2103);
xnor U1262 (N_1262,In_479,In_1119);
xor U1263 (N_1263,In_671,In_1826);
or U1264 (N_1264,In_710,In_542);
xor U1265 (N_1265,In_171,In_1837);
or U1266 (N_1266,In_1662,In_1231);
or U1267 (N_1267,In_1164,In_2446);
and U1268 (N_1268,In_646,In_544);
xor U1269 (N_1269,In_728,In_762);
xnor U1270 (N_1270,In_1069,In_718);
nand U1271 (N_1271,In_1765,In_1088);
nand U1272 (N_1272,In_2125,In_818);
or U1273 (N_1273,In_388,In_725);
nor U1274 (N_1274,In_487,In_253);
xnor U1275 (N_1275,In_1158,In_1678);
nor U1276 (N_1276,In_1921,In_2417);
nor U1277 (N_1277,In_1993,In_722);
nor U1278 (N_1278,In_327,In_1195);
xnor U1279 (N_1279,In_1249,In_836);
xnor U1280 (N_1280,In_1036,In_1292);
xnor U1281 (N_1281,In_471,In_2312);
nand U1282 (N_1282,In_85,In_1604);
or U1283 (N_1283,In_742,In_708);
nor U1284 (N_1284,In_1161,In_960);
xnor U1285 (N_1285,In_2003,In_1880);
xnor U1286 (N_1286,In_736,In_1379);
nand U1287 (N_1287,In_1745,In_1060);
xor U1288 (N_1288,In_289,In_1374);
or U1289 (N_1289,In_1409,In_340);
nor U1290 (N_1290,In_1580,In_2305);
and U1291 (N_1291,In_1687,In_666);
or U1292 (N_1292,In_1770,In_1404);
xor U1293 (N_1293,In_573,In_1964);
nand U1294 (N_1294,In_1589,In_166);
and U1295 (N_1295,In_869,In_2175);
or U1296 (N_1296,In_826,In_798);
nor U1297 (N_1297,In_239,In_1142);
xor U1298 (N_1298,In_557,In_1431);
and U1299 (N_1299,In_2003,In_1131);
xnor U1300 (N_1300,In_720,In_1938);
nand U1301 (N_1301,In_757,In_411);
nor U1302 (N_1302,In_1511,In_1476);
and U1303 (N_1303,In_996,In_1315);
nand U1304 (N_1304,In_1406,In_1039);
nor U1305 (N_1305,In_906,In_395);
nor U1306 (N_1306,In_1998,In_185);
xnor U1307 (N_1307,In_1405,In_941);
nor U1308 (N_1308,In_1022,In_11);
nor U1309 (N_1309,In_2158,In_389);
nand U1310 (N_1310,In_765,In_1482);
and U1311 (N_1311,In_380,In_19);
nor U1312 (N_1312,In_746,In_325);
and U1313 (N_1313,In_899,In_1884);
nand U1314 (N_1314,In_604,In_2429);
or U1315 (N_1315,In_1915,In_932);
nand U1316 (N_1316,In_2379,In_1065);
or U1317 (N_1317,In_2237,In_540);
nor U1318 (N_1318,In_2118,In_1952);
xnor U1319 (N_1319,In_570,In_1680);
xnor U1320 (N_1320,In_763,In_740);
nor U1321 (N_1321,In_562,In_1527);
or U1322 (N_1322,In_718,In_1723);
and U1323 (N_1323,In_1235,In_2284);
xnor U1324 (N_1324,In_1129,In_515);
xor U1325 (N_1325,In_1963,In_1406);
and U1326 (N_1326,In_949,In_1731);
xor U1327 (N_1327,In_98,In_2085);
nand U1328 (N_1328,In_2475,In_139);
nor U1329 (N_1329,In_2115,In_1003);
or U1330 (N_1330,In_219,In_354);
or U1331 (N_1331,In_549,In_336);
nand U1332 (N_1332,In_1833,In_121);
xnor U1333 (N_1333,In_374,In_1832);
and U1334 (N_1334,In_436,In_677);
nand U1335 (N_1335,In_1471,In_1061);
and U1336 (N_1336,In_1870,In_18);
nand U1337 (N_1337,In_2239,In_410);
xnor U1338 (N_1338,In_2481,In_1801);
and U1339 (N_1339,In_1346,In_2491);
xor U1340 (N_1340,In_1536,In_1976);
nand U1341 (N_1341,In_1475,In_561);
nor U1342 (N_1342,In_547,In_421);
and U1343 (N_1343,In_2205,In_208);
and U1344 (N_1344,In_550,In_2451);
nand U1345 (N_1345,In_2354,In_2416);
nor U1346 (N_1346,In_268,In_975);
xor U1347 (N_1347,In_2238,In_1693);
and U1348 (N_1348,In_1048,In_1513);
and U1349 (N_1349,In_233,In_458);
nand U1350 (N_1350,In_1807,In_988);
nand U1351 (N_1351,In_930,In_871);
or U1352 (N_1352,In_73,In_724);
xnor U1353 (N_1353,In_34,In_2478);
nand U1354 (N_1354,In_2417,In_324);
nand U1355 (N_1355,In_874,In_1294);
nor U1356 (N_1356,In_729,In_1462);
nor U1357 (N_1357,In_469,In_1776);
nand U1358 (N_1358,In_1762,In_172);
xor U1359 (N_1359,In_412,In_1559);
nor U1360 (N_1360,In_2383,In_207);
xor U1361 (N_1361,In_1014,In_92);
and U1362 (N_1362,In_1656,In_1057);
nand U1363 (N_1363,In_1762,In_514);
xor U1364 (N_1364,In_414,In_1254);
and U1365 (N_1365,In_2082,In_2196);
nand U1366 (N_1366,In_472,In_2179);
xnor U1367 (N_1367,In_2137,In_466);
nor U1368 (N_1368,In_1027,In_1415);
nor U1369 (N_1369,In_1038,In_1950);
nand U1370 (N_1370,In_307,In_2116);
xnor U1371 (N_1371,In_507,In_1827);
nand U1372 (N_1372,In_2287,In_2466);
nor U1373 (N_1373,In_2403,In_2115);
nor U1374 (N_1374,In_349,In_1291);
xnor U1375 (N_1375,In_1689,In_402);
or U1376 (N_1376,In_809,In_1529);
nor U1377 (N_1377,In_727,In_614);
nor U1378 (N_1378,In_379,In_1418);
nand U1379 (N_1379,In_986,In_553);
and U1380 (N_1380,In_1464,In_1946);
nand U1381 (N_1381,In_856,In_1196);
nor U1382 (N_1382,In_1083,In_1542);
nand U1383 (N_1383,In_661,In_2487);
or U1384 (N_1384,In_471,In_862);
xnor U1385 (N_1385,In_2171,In_667);
xor U1386 (N_1386,In_2144,In_1458);
xnor U1387 (N_1387,In_1782,In_455);
xnor U1388 (N_1388,In_1066,In_1893);
or U1389 (N_1389,In_1272,In_1325);
nor U1390 (N_1390,In_729,In_808);
and U1391 (N_1391,In_2360,In_160);
and U1392 (N_1392,In_509,In_2195);
nor U1393 (N_1393,In_244,In_2024);
nand U1394 (N_1394,In_79,In_1957);
nand U1395 (N_1395,In_1619,In_1223);
xor U1396 (N_1396,In_904,In_472);
and U1397 (N_1397,In_1336,In_1271);
or U1398 (N_1398,In_2171,In_2162);
nor U1399 (N_1399,In_2111,In_2061);
nand U1400 (N_1400,In_2032,In_1433);
xor U1401 (N_1401,In_1532,In_655);
or U1402 (N_1402,In_297,In_869);
nand U1403 (N_1403,In_1090,In_1850);
and U1404 (N_1404,In_85,In_714);
nor U1405 (N_1405,In_1844,In_1905);
and U1406 (N_1406,In_1466,In_1792);
nor U1407 (N_1407,In_2300,In_438);
xnor U1408 (N_1408,In_1990,In_2454);
xor U1409 (N_1409,In_1643,In_2039);
or U1410 (N_1410,In_353,In_907);
xnor U1411 (N_1411,In_2251,In_791);
or U1412 (N_1412,In_1546,In_1517);
nor U1413 (N_1413,In_1418,In_435);
and U1414 (N_1414,In_2111,In_2366);
nand U1415 (N_1415,In_1014,In_1378);
xnor U1416 (N_1416,In_309,In_2060);
nand U1417 (N_1417,In_2386,In_1815);
and U1418 (N_1418,In_671,In_1493);
or U1419 (N_1419,In_1506,In_1427);
nor U1420 (N_1420,In_716,In_374);
and U1421 (N_1421,In_2441,In_2031);
and U1422 (N_1422,In_287,In_676);
xor U1423 (N_1423,In_1925,In_1958);
nand U1424 (N_1424,In_1436,In_1828);
or U1425 (N_1425,In_2130,In_798);
xor U1426 (N_1426,In_1295,In_218);
nor U1427 (N_1427,In_2414,In_1196);
and U1428 (N_1428,In_1042,In_2225);
nand U1429 (N_1429,In_648,In_219);
and U1430 (N_1430,In_245,In_1945);
and U1431 (N_1431,In_1778,In_1921);
nor U1432 (N_1432,In_1259,In_887);
xor U1433 (N_1433,In_1261,In_1682);
xnor U1434 (N_1434,In_1034,In_1079);
or U1435 (N_1435,In_1798,In_1150);
nor U1436 (N_1436,In_328,In_649);
or U1437 (N_1437,In_1102,In_510);
xnor U1438 (N_1438,In_1540,In_1788);
nand U1439 (N_1439,In_2378,In_492);
xor U1440 (N_1440,In_359,In_920);
xnor U1441 (N_1441,In_796,In_778);
or U1442 (N_1442,In_1509,In_67);
and U1443 (N_1443,In_1166,In_2300);
nand U1444 (N_1444,In_2372,In_2072);
nand U1445 (N_1445,In_2057,In_107);
nor U1446 (N_1446,In_336,In_1145);
and U1447 (N_1447,In_945,In_2471);
and U1448 (N_1448,In_306,In_286);
or U1449 (N_1449,In_2062,In_1343);
and U1450 (N_1450,In_1915,In_2083);
xnor U1451 (N_1451,In_1701,In_2047);
xnor U1452 (N_1452,In_941,In_330);
nand U1453 (N_1453,In_1734,In_1313);
nand U1454 (N_1454,In_1626,In_1221);
and U1455 (N_1455,In_822,In_410);
or U1456 (N_1456,In_1940,In_1858);
nor U1457 (N_1457,In_1559,In_173);
nand U1458 (N_1458,In_2191,In_1464);
nor U1459 (N_1459,In_187,In_1409);
nor U1460 (N_1460,In_1927,In_201);
nand U1461 (N_1461,In_403,In_2412);
or U1462 (N_1462,In_1363,In_1349);
and U1463 (N_1463,In_2148,In_797);
nor U1464 (N_1464,In_384,In_2362);
nand U1465 (N_1465,In_480,In_766);
nor U1466 (N_1466,In_2366,In_2162);
nand U1467 (N_1467,In_256,In_1191);
and U1468 (N_1468,In_627,In_1867);
and U1469 (N_1469,In_1492,In_311);
nand U1470 (N_1470,In_458,In_1705);
nand U1471 (N_1471,In_422,In_467);
or U1472 (N_1472,In_2129,In_2101);
xor U1473 (N_1473,In_1781,In_1686);
nor U1474 (N_1474,In_1945,In_1346);
xor U1475 (N_1475,In_1860,In_251);
nand U1476 (N_1476,In_781,In_940);
nor U1477 (N_1477,In_1363,In_2388);
xor U1478 (N_1478,In_816,In_1473);
nand U1479 (N_1479,In_2355,In_1036);
nor U1480 (N_1480,In_2428,In_490);
nand U1481 (N_1481,In_679,In_1340);
or U1482 (N_1482,In_2016,In_2093);
nor U1483 (N_1483,In_236,In_154);
nand U1484 (N_1484,In_1974,In_444);
nor U1485 (N_1485,In_264,In_1373);
nand U1486 (N_1486,In_2325,In_370);
nor U1487 (N_1487,In_1806,In_767);
xor U1488 (N_1488,In_2449,In_2165);
nand U1489 (N_1489,In_995,In_2086);
xnor U1490 (N_1490,In_2470,In_1898);
and U1491 (N_1491,In_1891,In_2464);
or U1492 (N_1492,In_2212,In_2110);
nor U1493 (N_1493,In_1250,In_1559);
xnor U1494 (N_1494,In_2067,In_2165);
xnor U1495 (N_1495,In_118,In_1568);
nor U1496 (N_1496,In_506,In_361);
and U1497 (N_1497,In_716,In_1570);
xor U1498 (N_1498,In_1146,In_2225);
xnor U1499 (N_1499,In_831,In_364);
nand U1500 (N_1500,In_718,In_822);
nand U1501 (N_1501,In_972,In_1390);
or U1502 (N_1502,In_2373,In_1826);
nor U1503 (N_1503,In_266,In_2126);
or U1504 (N_1504,In_1856,In_569);
nand U1505 (N_1505,In_1217,In_1076);
xnor U1506 (N_1506,In_1793,In_1651);
xnor U1507 (N_1507,In_1533,In_865);
and U1508 (N_1508,In_2047,In_84);
and U1509 (N_1509,In_113,In_1197);
or U1510 (N_1510,In_1082,In_925);
nor U1511 (N_1511,In_2001,In_486);
xor U1512 (N_1512,In_549,In_538);
or U1513 (N_1513,In_1876,In_642);
xor U1514 (N_1514,In_673,In_1979);
and U1515 (N_1515,In_1846,In_1580);
or U1516 (N_1516,In_189,In_1987);
xor U1517 (N_1517,In_283,In_1815);
xor U1518 (N_1518,In_2160,In_1684);
and U1519 (N_1519,In_977,In_1077);
and U1520 (N_1520,In_489,In_802);
nor U1521 (N_1521,In_1494,In_288);
or U1522 (N_1522,In_540,In_1293);
or U1523 (N_1523,In_1102,In_720);
nand U1524 (N_1524,In_687,In_1708);
nand U1525 (N_1525,In_160,In_1306);
nor U1526 (N_1526,In_37,In_402);
nand U1527 (N_1527,In_908,In_1283);
or U1528 (N_1528,In_23,In_1929);
and U1529 (N_1529,In_2366,In_2484);
nor U1530 (N_1530,In_1205,In_1735);
or U1531 (N_1531,In_1484,In_2168);
and U1532 (N_1532,In_675,In_776);
nor U1533 (N_1533,In_142,In_2307);
xnor U1534 (N_1534,In_1162,In_67);
nand U1535 (N_1535,In_1938,In_2427);
nand U1536 (N_1536,In_761,In_578);
or U1537 (N_1537,In_1760,In_1014);
nand U1538 (N_1538,In_2432,In_1554);
xor U1539 (N_1539,In_1161,In_2133);
xnor U1540 (N_1540,In_1681,In_1520);
nand U1541 (N_1541,In_612,In_1041);
or U1542 (N_1542,In_2183,In_451);
nand U1543 (N_1543,In_326,In_2128);
or U1544 (N_1544,In_1189,In_82);
and U1545 (N_1545,In_1488,In_943);
and U1546 (N_1546,In_1610,In_1651);
nand U1547 (N_1547,In_987,In_673);
nor U1548 (N_1548,In_686,In_1714);
and U1549 (N_1549,In_1362,In_1722);
nor U1550 (N_1550,In_2242,In_551);
xnor U1551 (N_1551,In_2070,In_1314);
nor U1552 (N_1552,In_549,In_320);
and U1553 (N_1553,In_587,In_2024);
nor U1554 (N_1554,In_2338,In_2375);
and U1555 (N_1555,In_112,In_1912);
or U1556 (N_1556,In_1895,In_500);
and U1557 (N_1557,In_1375,In_292);
xor U1558 (N_1558,In_1894,In_2385);
and U1559 (N_1559,In_2318,In_962);
xor U1560 (N_1560,In_1283,In_2242);
xor U1561 (N_1561,In_2210,In_1768);
xor U1562 (N_1562,In_922,In_771);
and U1563 (N_1563,In_2007,In_43);
and U1564 (N_1564,In_2266,In_1141);
and U1565 (N_1565,In_2024,In_1381);
nand U1566 (N_1566,In_2283,In_380);
or U1567 (N_1567,In_1350,In_76);
and U1568 (N_1568,In_185,In_1280);
nor U1569 (N_1569,In_1051,In_2055);
nor U1570 (N_1570,In_1673,In_2028);
or U1571 (N_1571,In_1000,In_2104);
nor U1572 (N_1572,In_571,In_2349);
nor U1573 (N_1573,In_170,In_657);
nand U1574 (N_1574,In_1381,In_116);
or U1575 (N_1575,In_790,In_169);
or U1576 (N_1576,In_699,In_724);
nor U1577 (N_1577,In_820,In_84);
nand U1578 (N_1578,In_1058,In_1824);
nand U1579 (N_1579,In_2073,In_700);
nand U1580 (N_1580,In_627,In_2498);
nand U1581 (N_1581,In_85,In_1046);
xor U1582 (N_1582,In_655,In_942);
or U1583 (N_1583,In_1378,In_2280);
xor U1584 (N_1584,In_1363,In_2068);
or U1585 (N_1585,In_1078,In_2323);
xnor U1586 (N_1586,In_828,In_2094);
nand U1587 (N_1587,In_726,In_558);
nor U1588 (N_1588,In_1266,In_2144);
nand U1589 (N_1589,In_1363,In_1737);
or U1590 (N_1590,In_2060,In_894);
xnor U1591 (N_1591,In_94,In_1818);
and U1592 (N_1592,In_732,In_2497);
nor U1593 (N_1593,In_711,In_1823);
or U1594 (N_1594,In_1777,In_1515);
xor U1595 (N_1595,In_2221,In_1205);
nand U1596 (N_1596,In_2106,In_509);
nor U1597 (N_1597,In_1300,In_1973);
nor U1598 (N_1598,In_2342,In_2421);
nor U1599 (N_1599,In_1149,In_664);
nand U1600 (N_1600,In_1842,In_1890);
or U1601 (N_1601,In_2350,In_1462);
nor U1602 (N_1602,In_1248,In_1956);
or U1603 (N_1603,In_318,In_423);
xor U1604 (N_1604,In_613,In_381);
nand U1605 (N_1605,In_1375,In_1807);
nor U1606 (N_1606,In_151,In_359);
xor U1607 (N_1607,In_2498,In_92);
nor U1608 (N_1608,In_1513,In_1218);
or U1609 (N_1609,In_196,In_1804);
or U1610 (N_1610,In_334,In_1890);
and U1611 (N_1611,In_1817,In_216);
and U1612 (N_1612,In_727,In_2426);
or U1613 (N_1613,In_1230,In_1876);
nand U1614 (N_1614,In_908,In_2280);
nand U1615 (N_1615,In_1394,In_365);
nand U1616 (N_1616,In_1403,In_2429);
xor U1617 (N_1617,In_1677,In_286);
and U1618 (N_1618,In_680,In_1490);
nor U1619 (N_1619,In_458,In_651);
nand U1620 (N_1620,In_1495,In_1009);
nand U1621 (N_1621,In_637,In_1640);
nor U1622 (N_1622,In_1986,In_1740);
and U1623 (N_1623,In_2079,In_1538);
nand U1624 (N_1624,In_95,In_607);
and U1625 (N_1625,In_1997,In_331);
nand U1626 (N_1626,In_1687,In_1998);
nor U1627 (N_1627,In_231,In_1810);
or U1628 (N_1628,In_1113,In_2313);
xor U1629 (N_1629,In_56,In_1496);
or U1630 (N_1630,In_276,In_2279);
nor U1631 (N_1631,In_1565,In_1455);
nand U1632 (N_1632,In_893,In_211);
nor U1633 (N_1633,In_510,In_373);
nor U1634 (N_1634,In_1977,In_1449);
xor U1635 (N_1635,In_842,In_827);
xor U1636 (N_1636,In_1461,In_1994);
or U1637 (N_1637,In_1707,In_1939);
or U1638 (N_1638,In_2407,In_2435);
nand U1639 (N_1639,In_1762,In_1183);
nor U1640 (N_1640,In_1942,In_1806);
nor U1641 (N_1641,In_2387,In_2109);
or U1642 (N_1642,In_101,In_1041);
nand U1643 (N_1643,In_185,In_1783);
and U1644 (N_1644,In_1459,In_1235);
nand U1645 (N_1645,In_1250,In_1847);
and U1646 (N_1646,In_221,In_252);
xnor U1647 (N_1647,In_1843,In_884);
xor U1648 (N_1648,In_2278,In_976);
or U1649 (N_1649,In_1484,In_407);
or U1650 (N_1650,In_1216,In_2068);
and U1651 (N_1651,In_1977,In_1831);
xor U1652 (N_1652,In_1191,In_751);
xor U1653 (N_1653,In_1079,In_2289);
or U1654 (N_1654,In_516,In_1891);
or U1655 (N_1655,In_2314,In_839);
xnor U1656 (N_1656,In_271,In_2108);
or U1657 (N_1657,In_641,In_870);
xnor U1658 (N_1658,In_1900,In_895);
xor U1659 (N_1659,In_30,In_581);
or U1660 (N_1660,In_2358,In_1648);
and U1661 (N_1661,In_1196,In_1771);
and U1662 (N_1662,In_28,In_919);
nor U1663 (N_1663,In_1202,In_368);
and U1664 (N_1664,In_1038,In_1520);
nand U1665 (N_1665,In_405,In_483);
nand U1666 (N_1666,In_1815,In_2004);
nor U1667 (N_1667,In_1136,In_701);
nand U1668 (N_1668,In_763,In_752);
nand U1669 (N_1669,In_1817,In_1050);
and U1670 (N_1670,In_1370,In_1271);
nor U1671 (N_1671,In_2016,In_588);
nand U1672 (N_1672,In_26,In_1225);
nand U1673 (N_1673,In_512,In_1938);
or U1674 (N_1674,In_1443,In_37);
nand U1675 (N_1675,In_11,In_149);
or U1676 (N_1676,In_968,In_1505);
nand U1677 (N_1677,In_2070,In_275);
nand U1678 (N_1678,In_306,In_1019);
and U1679 (N_1679,In_1540,In_544);
or U1680 (N_1680,In_2394,In_1461);
or U1681 (N_1681,In_733,In_1818);
xnor U1682 (N_1682,In_1965,In_844);
or U1683 (N_1683,In_789,In_899);
nor U1684 (N_1684,In_2066,In_2003);
nor U1685 (N_1685,In_1383,In_389);
or U1686 (N_1686,In_921,In_353);
nor U1687 (N_1687,In_1376,In_691);
nor U1688 (N_1688,In_1270,In_1758);
and U1689 (N_1689,In_2223,In_1281);
nand U1690 (N_1690,In_1603,In_1776);
xnor U1691 (N_1691,In_861,In_2129);
or U1692 (N_1692,In_2223,In_1637);
and U1693 (N_1693,In_2244,In_1671);
xnor U1694 (N_1694,In_814,In_2485);
and U1695 (N_1695,In_377,In_1468);
or U1696 (N_1696,In_2361,In_574);
and U1697 (N_1697,In_384,In_1659);
nand U1698 (N_1698,In_73,In_1303);
or U1699 (N_1699,In_1999,In_1946);
or U1700 (N_1700,In_1418,In_1627);
and U1701 (N_1701,In_2118,In_2419);
xor U1702 (N_1702,In_1834,In_1589);
or U1703 (N_1703,In_347,In_795);
nor U1704 (N_1704,In_989,In_2359);
or U1705 (N_1705,In_838,In_1051);
and U1706 (N_1706,In_108,In_2205);
nor U1707 (N_1707,In_2131,In_1500);
and U1708 (N_1708,In_1258,In_1864);
xnor U1709 (N_1709,In_2085,In_1180);
nand U1710 (N_1710,In_869,In_140);
nand U1711 (N_1711,In_263,In_1570);
xor U1712 (N_1712,In_1579,In_1167);
and U1713 (N_1713,In_2289,In_271);
or U1714 (N_1714,In_1292,In_500);
nand U1715 (N_1715,In_211,In_1889);
and U1716 (N_1716,In_2237,In_881);
xor U1717 (N_1717,In_262,In_848);
or U1718 (N_1718,In_2013,In_1696);
or U1719 (N_1719,In_142,In_37);
xor U1720 (N_1720,In_406,In_801);
nand U1721 (N_1721,In_918,In_1570);
and U1722 (N_1722,In_912,In_1472);
nand U1723 (N_1723,In_529,In_288);
nor U1724 (N_1724,In_967,In_1975);
or U1725 (N_1725,In_1154,In_1042);
and U1726 (N_1726,In_981,In_182);
nor U1727 (N_1727,In_77,In_539);
or U1728 (N_1728,In_389,In_1606);
nand U1729 (N_1729,In_1451,In_824);
or U1730 (N_1730,In_1934,In_1314);
nor U1731 (N_1731,In_2217,In_2058);
or U1732 (N_1732,In_2317,In_1336);
and U1733 (N_1733,In_381,In_2373);
nand U1734 (N_1734,In_911,In_1461);
nor U1735 (N_1735,In_203,In_55);
nand U1736 (N_1736,In_794,In_2393);
nand U1737 (N_1737,In_275,In_2037);
nand U1738 (N_1738,In_1794,In_340);
or U1739 (N_1739,In_1530,In_1293);
nor U1740 (N_1740,In_1718,In_1131);
nand U1741 (N_1741,In_321,In_273);
and U1742 (N_1742,In_2130,In_1048);
or U1743 (N_1743,In_1474,In_1381);
nand U1744 (N_1744,In_1523,In_2155);
or U1745 (N_1745,In_953,In_1395);
nor U1746 (N_1746,In_1291,In_736);
nand U1747 (N_1747,In_1748,In_664);
and U1748 (N_1748,In_2150,In_2193);
and U1749 (N_1749,In_585,In_1280);
and U1750 (N_1750,In_1915,In_1494);
xor U1751 (N_1751,In_1497,In_33);
and U1752 (N_1752,In_2359,In_1280);
and U1753 (N_1753,In_2167,In_1440);
or U1754 (N_1754,In_2229,In_2374);
nor U1755 (N_1755,In_528,In_2269);
and U1756 (N_1756,In_400,In_2280);
and U1757 (N_1757,In_1634,In_380);
nor U1758 (N_1758,In_489,In_223);
nor U1759 (N_1759,In_724,In_1064);
and U1760 (N_1760,In_763,In_1731);
xor U1761 (N_1761,In_21,In_755);
or U1762 (N_1762,In_46,In_937);
or U1763 (N_1763,In_988,In_348);
or U1764 (N_1764,In_1866,In_149);
xor U1765 (N_1765,In_607,In_1543);
xnor U1766 (N_1766,In_2349,In_2021);
nand U1767 (N_1767,In_2393,In_1227);
xor U1768 (N_1768,In_2054,In_2208);
and U1769 (N_1769,In_254,In_284);
nand U1770 (N_1770,In_1635,In_2286);
and U1771 (N_1771,In_1272,In_1459);
xor U1772 (N_1772,In_866,In_234);
nor U1773 (N_1773,In_2011,In_2340);
and U1774 (N_1774,In_1394,In_1670);
xnor U1775 (N_1775,In_1110,In_1523);
xnor U1776 (N_1776,In_1499,In_215);
xor U1777 (N_1777,In_727,In_631);
xor U1778 (N_1778,In_1333,In_1790);
or U1779 (N_1779,In_1653,In_1654);
or U1780 (N_1780,In_890,In_563);
nor U1781 (N_1781,In_2100,In_302);
nor U1782 (N_1782,In_1092,In_413);
and U1783 (N_1783,In_1641,In_575);
nand U1784 (N_1784,In_1610,In_1784);
nand U1785 (N_1785,In_1277,In_1004);
xnor U1786 (N_1786,In_534,In_221);
nand U1787 (N_1787,In_1506,In_1255);
and U1788 (N_1788,In_1138,In_1105);
xnor U1789 (N_1789,In_3,In_349);
nor U1790 (N_1790,In_1973,In_898);
nor U1791 (N_1791,In_700,In_1022);
or U1792 (N_1792,In_1942,In_2178);
xor U1793 (N_1793,In_1374,In_2028);
nor U1794 (N_1794,In_2262,In_1315);
and U1795 (N_1795,In_2423,In_1137);
nand U1796 (N_1796,In_988,In_1109);
or U1797 (N_1797,In_382,In_424);
nand U1798 (N_1798,In_977,In_2065);
nand U1799 (N_1799,In_343,In_648);
and U1800 (N_1800,In_1869,In_892);
nand U1801 (N_1801,In_1468,In_2392);
xnor U1802 (N_1802,In_496,In_483);
and U1803 (N_1803,In_1123,In_1441);
nand U1804 (N_1804,In_1081,In_412);
nand U1805 (N_1805,In_535,In_2122);
xnor U1806 (N_1806,In_2025,In_2493);
or U1807 (N_1807,In_2437,In_2361);
or U1808 (N_1808,In_2282,In_1286);
and U1809 (N_1809,In_2258,In_714);
nand U1810 (N_1810,In_383,In_780);
and U1811 (N_1811,In_1288,In_482);
nor U1812 (N_1812,In_763,In_675);
nand U1813 (N_1813,In_2080,In_2260);
and U1814 (N_1814,In_727,In_2265);
and U1815 (N_1815,In_2144,In_440);
or U1816 (N_1816,In_640,In_321);
and U1817 (N_1817,In_1297,In_753);
nand U1818 (N_1818,In_287,In_1152);
and U1819 (N_1819,In_957,In_1977);
and U1820 (N_1820,In_748,In_627);
and U1821 (N_1821,In_1099,In_1488);
nor U1822 (N_1822,In_1846,In_1095);
xor U1823 (N_1823,In_2465,In_205);
nor U1824 (N_1824,In_2435,In_2486);
nand U1825 (N_1825,In_1281,In_1998);
and U1826 (N_1826,In_1729,In_941);
nor U1827 (N_1827,In_190,In_1627);
xnor U1828 (N_1828,In_1078,In_1570);
nor U1829 (N_1829,In_538,In_1278);
xor U1830 (N_1830,In_1696,In_523);
and U1831 (N_1831,In_1459,In_138);
xor U1832 (N_1832,In_1022,In_1507);
nand U1833 (N_1833,In_574,In_2462);
nand U1834 (N_1834,In_1914,In_212);
nand U1835 (N_1835,In_1177,In_1268);
xnor U1836 (N_1836,In_1457,In_1653);
or U1837 (N_1837,In_490,In_33);
nand U1838 (N_1838,In_2467,In_2275);
nor U1839 (N_1839,In_2410,In_2170);
nor U1840 (N_1840,In_625,In_1603);
nor U1841 (N_1841,In_1782,In_1423);
nand U1842 (N_1842,In_94,In_2469);
xor U1843 (N_1843,In_1952,In_153);
xor U1844 (N_1844,In_939,In_897);
nor U1845 (N_1845,In_1394,In_951);
nand U1846 (N_1846,In_2442,In_908);
xnor U1847 (N_1847,In_1187,In_1136);
and U1848 (N_1848,In_1465,In_949);
xor U1849 (N_1849,In_79,In_2457);
xor U1850 (N_1850,In_615,In_1503);
nand U1851 (N_1851,In_637,In_1109);
nand U1852 (N_1852,In_2071,In_1442);
nand U1853 (N_1853,In_1491,In_1311);
or U1854 (N_1854,In_1329,In_433);
nor U1855 (N_1855,In_1643,In_136);
xor U1856 (N_1856,In_557,In_2443);
nor U1857 (N_1857,In_202,In_755);
xor U1858 (N_1858,In_574,In_357);
or U1859 (N_1859,In_351,In_1619);
xor U1860 (N_1860,In_1472,In_2051);
and U1861 (N_1861,In_1161,In_2249);
and U1862 (N_1862,In_1088,In_1453);
nand U1863 (N_1863,In_880,In_105);
nor U1864 (N_1864,In_777,In_369);
nor U1865 (N_1865,In_1159,In_748);
nor U1866 (N_1866,In_433,In_265);
or U1867 (N_1867,In_1835,In_1857);
nor U1868 (N_1868,In_1529,In_409);
nand U1869 (N_1869,In_929,In_2124);
nand U1870 (N_1870,In_1363,In_1015);
nand U1871 (N_1871,In_572,In_165);
or U1872 (N_1872,In_2376,In_2006);
and U1873 (N_1873,In_1601,In_302);
and U1874 (N_1874,In_520,In_689);
xnor U1875 (N_1875,In_1222,In_1008);
xnor U1876 (N_1876,In_1654,In_1046);
nand U1877 (N_1877,In_1928,In_1403);
nor U1878 (N_1878,In_1571,In_612);
nand U1879 (N_1879,In_2408,In_2005);
nand U1880 (N_1880,In_1163,In_2400);
nor U1881 (N_1881,In_1002,In_15);
nor U1882 (N_1882,In_1872,In_1971);
nand U1883 (N_1883,In_1124,In_1766);
nand U1884 (N_1884,In_2216,In_754);
and U1885 (N_1885,In_1842,In_12);
nand U1886 (N_1886,In_1139,In_1424);
nand U1887 (N_1887,In_361,In_2329);
or U1888 (N_1888,In_2142,In_173);
or U1889 (N_1889,In_218,In_1880);
or U1890 (N_1890,In_1558,In_2482);
or U1891 (N_1891,In_1888,In_548);
xnor U1892 (N_1892,In_2344,In_2419);
nor U1893 (N_1893,In_1966,In_1822);
nor U1894 (N_1894,In_112,In_215);
xor U1895 (N_1895,In_1523,In_955);
and U1896 (N_1896,In_123,In_776);
nand U1897 (N_1897,In_787,In_1668);
nand U1898 (N_1898,In_577,In_306);
nand U1899 (N_1899,In_1596,In_32);
or U1900 (N_1900,In_2314,In_1822);
xor U1901 (N_1901,In_1871,In_1530);
nor U1902 (N_1902,In_2331,In_1141);
and U1903 (N_1903,In_756,In_121);
and U1904 (N_1904,In_1851,In_123);
or U1905 (N_1905,In_1299,In_605);
nand U1906 (N_1906,In_540,In_846);
or U1907 (N_1907,In_1293,In_565);
nand U1908 (N_1908,In_283,In_2153);
or U1909 (N_1909,In_1423,In_880);
xnor U1910 (N_1910,In_1332,In_2394);
xnor U1911 (N_1911,In_1728,In_652);
nor U1912 (N_1912,In_1493,In_281);
and U1913 (N_1913,In_879,In_1554);
or U1914 (N_1914,In_1275,In_2400);
nor U1915 (N_1915,In_336,In_1719);
xnor U1916 (N_1916,In_198,In_214);
nand U1917 (N_1917,In_1114,In_1643);
or U1918 (N_1918,In_2074,In_2122);
and U1919 (N_1919,In_662,In_1248);
xor U1920 (N_1920,In_938,In_506);
and U1921 (N_1921,In_65,In_783);
xnor U1922 (N_1922,In_1977,In_1127);
nand U1923 (N_1923,In_208,In_2473);
nand U1924 (N_1924,In_1678,In_392);
and U1925 (N_1925,In_1721,In_688);
xor U1926 (N_1926,In_161,In_1748);
nand U1927 (N_1927,In_1439,In_1700);
nand U1928 (N_1928,In_878,In_751);
nand U1929 (N_1929,In_1546,In_2412);
nand U1930 (N_1930,In_2351,In_1503);
or U1931 (N_1931,In_1732,In_1157);
and U1932 (N_1932,In_89,In_276);
and U1933 (N_1933,In_1908,In_580);
nand U1934 (N_1934,In_1454,In_1528);
nand U1935 (N_1935,In_1488,In_1992);
or U1936 (N_1936,In_2237,In_258);
nor U1937 (N_1937,In_666,In_1819);
and U1938 (N_1938,In_2222,In_1613);
or U1939 (N_1939,In_1001,In_2116);
and U1940 (N_1940,In_187,In_2443);
nor U1941 (N_1941,In_2193,In_2342);
nand U1942 (N_1942,In_1652,In_378);
and U1943 (N_1943,In_1011,In_1053);
and U1944 (N_1944,In_34,In_720);
or U1945 (N_1945,In_818,In_391);
xnor U1946 (N_1946,In_2122,In_2024);
or U1947 (N_1947,In_2144,In_2196);
and U1948 (N_1948,In_1787,In_731);
and U1949 (N_1949,In_384,In_1475);
or U1950 (N_1950,In_2147,In_103);
or U1951 (N_1951,In_1415,In_1280);
nor U1952 (N_1952,In_104,In_950);
or U1953 (N_1953,In_2015,In_1446);
xor U1954 (N_1954,In_1905,In_2229);
nor U1955 (N_1955,In_26,In_1857);
or U1956 (N_1956,In_2046,In_2470);
xnor U1957 (N_1957,In_329,In_1757);
xnor U1958 (N_1958,In_1297,In_1356);
nand U1959 (N_1959,In_742,In_551);
or U1960 (N_1960,In_249,In_1084);
and U1961 (N_1961,In_610,In_2471);
nand U1962 (N_1962,In_1835,In_274);
nor U1963 (N_1963,In_1092,In_173);
xnor U1964 (N_1964,In_1629,In_1768);
nand U1965 (N_1965,In_746,In_1688);
and U1966 (N_1966,In_1990,In_264);
nor U1967 (N_1967,In_1544,In_717);
and U1968 (N_1968,In_1222,In_1957);
and U1969 (N_1969,In_1615,In_2032);
nand U1970 (N_1970,In_1349,In_2477);
nor U1971 (N_1971,In_1945,In_1751);
xor U1972 (N_1972,In_1946,In_736);
nor U1973 (N_1973,In_1192,In_227);
or U1974 (N_1974,In_1916,In_2456);
xnor U1975 (N_1975,In_2102,In_1244);
nand U1976 (N_1976,In_12,In_1715);
nor U1977 (N_1977,In_542,In_2180);
or U1978 (N_1978,In_879,In_30);
or U1979 (N_1979,In_2297,In_1369);
or U1980 (N_1980,In_1206,In_2243);
xnor U1981 (N_1981,In_248,In_37);
nand U1982 (N_1982,In_104,In_733);
nand U1983 (N_1983,In_999,In_926);
and U1984 (N_1984,In_1723,In_1802);
xnor U1985 (N_1985,In_108,In_16);
xnor U1986 (N_1986,In_1279,In_1821);
or U1987 (N_1987,In_1889,In_1424);
or U1988 (N_1988,In_102,In_1767);
nor U1989 (N_1989,In_1719,In_295);
or U1990 (N_1990,In_281,In_1582);
xnor U1991 (N_1991,In_336,In_2252);
nand U1992 (N_1992,In_1377,In_574);
or U1993 (N_1993,In_1401,In_2146);
or U1994 (N_1994,In_1654,In_2396);
or U1995 (N_1995,In_2015,In_1906);
or U1996 (N_1996,In_145,In_216);
or U1997 (N_1997,In_1321,In_70);
xor U1998 (N_1998,In_1376,In_454);
nor U1999 (N_1999,In_1256,In_2171);
nor U2000 (N_2000,In_1223,In_1003);
nand U2001 (N_2001,In_54,In_1488);
nand U2002 (N_2002,In_681,In_913);
or U2003 (N_2003,In_112,In_364);
xor U2004 (N_2004,In_66,In_2310);
nor U2005 (N_2005,In_1969,In_1477);
or U2006 (N_2006,In_57,In_417);
nor U2007 (N_2007,In_109,In_257);
and U2008 (N_2008,In_1088,In_1222);
and U2009 (N_2009,In_290,In_750);
nor U2010 (N_2010,In_429,In_1600);
or U2011 (N_2011,In_1291,In_1865);
nor U2012 (N_2012,In_998,In_1754);
nand U2013 (N_2013,In_1721,In_1096);
xnor U2014 (N_2014,In_1611,In_2111);
xnor U2015 (N_2015,In_2228,In_1995);
nand U2016 (N_2016,In_2105,In_2474);
nand U2017 (N_2017,In_365,In_1592);
nand U2018 (N_2018,In_798,In_2249);
nand U2019 (N_2019,In_931,In_2062);
and U2020 (N_2020,In_1712,In_1856);
xnor U2021 (N_2021,In_1039,In_1680);
and U2022 (N_2022,In_882,In_1750);
and U2023 (N_2023,In_936,In_8);
and U2024 (N_2024,In_1996,In_159);
xor U2025 (N_2025,In_1589,In_2277);
xnor U2026 (N_2026,In_1803,In_1094);
xor U2027 (N_2027,In_198,In_1245);
nand U2028 (N_2028,In_1387,In_2095);
nand U2029 (N_2029,In_1574,In_152);
nand U2030 (N_2030,In_1632,In_1769);
or U2031 (N_2031,In_269,In_1059);
or U2032 (N_2032,In_1263,In_1332);
xor U2033 (N_2033,In_1369,In_2325);
and U2034 (N_2034,In_841,In_1087);
nor U2035 (N_2035,In_1768,In_1089);
or U2036 (N_2036,In_1274,In_1684);
nor U2037 (N_2037,In_2086,In_2475);
and U2038 (N_2038,In_463,In_504);
nand U2039 (N_2039,In_477,In_2035);
or U2040 (N_2040,In_1824,In_2107);
xor U2041 (N_2041,In_1371,In_1811);
nor U2042 (N_2042,In_106,In_843);
xor U2043 (N_2043,In_166,In_707);
and U2044 (N_2044,In_237,In_909);
nand U2045 (N_2045,In_2380,In_2462);
nand U2046 (N_2046,In_2440,In_40);
nor U2047 (N_2047,In_312,In_2095);
or U2048 (N_2048,In_115,In_1091);
nor U2049 (N_2049,In_1964,In_1872);
nand U2050 (N_2050,In_305,In_140);
or U2051 (N_2051,In_872,In_13);
and U2052 (N_2052,In_1824,In_1961);
or U2053 (N_2053,In_504,In_1193);
nor U2054 (N_2054,In_1832,In_1959);
nand U2055 (N_2055,In_194,In_290);
xor U2056 (N_2056,In_73,In_161);
and U2057 (N_2057,In_1622,In_1957);
xor U2058 (N_2058,In_308,In_2091);
or U2059 (N_2059,In_1232,In_1500);
nand U2060 (N_2060,In_2079,In_2088);
xnor U2061 (N_2061,In_224,In_1357);
nand U2062 (N_2062,In_2450,In_25);
nand U2063 (N_2063,In_1090,In_2119);
nor U2064 (N_2064,In_589,In_1820);
and U2065 (N_2065,In_1907,In_487);
xor U2066 (N_2066,In_2131,In_1350);
nand U2067 (N_2067,In_697,In_2150);
or U2068 (N_2068,In_528,In_1678);
xnor U2069 (N_2069,In_1572,In_518);
nor U2070 (N_2070,In_2166,In_2029);
and U2071 (N_2071,In_312,In_2177);
and U2072 (N_2072,In_33,In_1383);
xor U2073 (N_2073,In_1628,In_2463);
nor U2074 (N_2074,In_2082,In_1680);
nand U2075 (N_2075,In_286,In_882);
xnor U2076 (N_2076,In_2450,In_1273);
nand U2077 (N_2077,In_161,In_616);
xnor U2078 (N_2078,In_2485,In_661);
nor U2079 (N_2079,In_2125,In_252);
and U2080 (N_2080,In_2092,In_1451);
nand U2081 (N_2081,In_997,In_1892);
nor U2082 (N_2082,In_895,In_1907);
xor U2083 (N_2083,In_1660,In_1380);
nor U2084 (N_2084,In_1715,In_92);
and U2085 (N_2085,In_181,In_2109);
nor U2086 (N_2086,In_4,In_1199);
xor U2087 (N_2087,In_1381,In_2060);
nor U2088 (N_2088,In_959,In_525);
and U2089 (N_2089,In_2072,In_2452);
xnor U2090 (N_2090,In_1841,In_1964);
xnor U2091 (N_2091,In_2486,In_475);
nor U2092 (N_2092,In_2343,In_912);
nand U2093 (N_2093,In_335,In_1757);
nand U2094 (N_2094,In_717,In_1811);
nand U2095 (N_2095,In_2174,In_1663);
or U2096 (N_2096,In_1773,In_1440);
xor U2097 (N_2097,In_323,In_632);
xnor U2098 (N_2098,In_1241,In_1614);
xor U2099 (N_2099,In_698,In_1972);
or U2100 (N_2100,In_1256,In_82);
nor U2101 (N_2101,In_1052,In_593);
nor U2102 (N_2102,In_111,In_1462);
nor U2103 (N_2103,In_1269,In_1499);
or U2104 (N_2104,In_1147,In_861);
nor U2105 (N_2105,In_2308,In_1093);
or U2106 (N_2106,In_1462,In_1570);
nor U2107 (N_2107,In_730,In_1240);
xnor U2108 (N_2108,In_2325,In_533);
or U2109 (N_2109,In_814,In_197);
or U2110 (N_2110,In_1133,In_2479);
nor U2111 (N_2111,In_2175,In_2335);
xor U2112 (N_2112,In_1448,In_1678);
xnor U2113 (N_2113,In_114,In_2309);
nand U2114 (N_2114,In_496,In_926);
nand U2115 (N_2115,In_1373,In_841);
xnor U2116 (N_2116,In_1507,In_1308);
xor U2117 (N_2117,In_1434,In_1139);
xor U2118 (N_2118,In_702,In_1594);
nand U2119 (N_2119,In_1335,In_1775);
or U2120 (N_2120,In_2272,In_2088);
or U2121 (N_2121,In_328,In_1015);
xnor U2122 (N_2122,In_2415,In_1669);
and U2123 (N_2123,In_1952,In_50);
and U2124 (N_2124,In_56,In_267);
and U2125 (N_2125,In_691,In_1464);
xnor U2126 (N_2126,In_564,In_254);
nand U2127 (N_2127,In_502,In_227);
nor U2128 (N_2128,In_782,In_2363);
xor U2129 (N_2129,In_100,In_1420);
nand U2130 (N_2130,In_757,In_1103);
or U2131 (N_2131,In_356,In_837);
or U2132 (N_2132,In_793,In_495);
nand U2133 (N_2133,In_2104,In_910);
nor U2134 (N_2134,In_809,In_1072);
nor U2135 (N_2135,In_2325,In_230);
nand U2136 (N_2136,In_830,In_400);
and U2137 (N_2137,In_417,In_192);
xor U2138 (N_2138,In_2283,In_1178);
or U2139 (N_2139,In_292,In_532);
and U2140 (N_2140,In_95,In_364);
and U2141 (N_2141,In_1588,In_602);
nor U2142 (N_2142,In_1672,In_371);
or U2143 (N_2143,In_1532,In_2436);
or U2144 (N_2144,In_757,In_879);
nand U2145 (N_2145,In_1989,In_547);
nor U2146 (N_2146,In_1869,In_2193);
nor U2147 (N_2147,In_528,In_946);
and U2148 (N_2148,In_2255,In_2207);
nand U2149 (N_2149,In_2335,In_906);
or U2150 (N_2150,In_1225,In_1553);
and U2151 (N_2151,In_1417,In_790);
xor U2152 (N_2152,In_1980,In_1424);
or U2153 (N_2153,In_2346,In_814);
xor U2154 (N_2154,In_694,In_120);
nand U2155 (N_2155,In_2407,In_2276);
and U2156 (N_2156,In_756,In_1111);
nand U2157 (N_2157,In_451,In_463);
nor U2158 (N_2158,In_1587,In_1657);
nand U2159 (N_2159,In_2356,In_1922);
nor U2160 (N_2160,In_920,In_1960);
xor U2161 (N_2161,In_29,In_2101);
xnor U2162 (N_2162,In_1855,In_682);
or U2163 (N_2163,In_1440,In_1591);
and U2164 (N_2164,In_557,In_190);
or U2165 (N_2165,In_1772,In_1193);
xor U2166 (N_2166,In_1387,In_111);
or U2167 (N_2167,In_1183,In_182);
and U2168 (N_2168,In_922,In_834);
xnor U2169 (N_2169,In_1989,In_2191);
and U2170 (N_2170,In_1123,In_2443);
nor U2171 (N_2171,In_49,In_1686);
nand U2172 (N_2172,In_830,In_488);
nor U2173 (N_2173,In_1445,In_763);
nor U2174 (N_2174,In_1214,In_2067);
nor U2175 (N_2175,In_2095,In_580);
and U2176 (N_2176,In_1213,In_2202);
nand U2177 (N_2177,In_451,In_1911);
xor U2178 (N_2178,In_566,In_1931);
or U2179 (N_2179,In_8,In_962);
nand U2180 (N_2180,In_2357,In_949);
and U2181 (N_2181,In_221,In_1838);
nor U2182 (N_2182,In_666,In_818);
or U2183 (N_2183,In_1447,In_2323);
or U2184 (N_2184,In_970,In_1367);
and U2185 (N_2185,In_498,In_1514);
xor U2186 (N_2186,In_1330,In_758);
nor U2187 (N_2187,In_317,In_1731);
nand U2188 (N_2188,In_1578,In_1628);
nand U2189 (N_2189,In_538,In_219);
and U2190 (N_2190,In_1420,In_1294);
xor U2191 (N_2191,In_1978,In_1293);
nand U2192 (N_2192,In_2367,In_1588);
or U2193 (N_2193,In_284,In_1406);
or U2194 (N_2194,In_1009,In_1723);
nor U2195 (N_2195,In_400,In_502);
and U2196 (N_2196,In_2298,In_353);
nand U2197 (N_2197,In_637,In_302);
nand U2198 (N_2198,In_1808,In_1167);
nor U2199 (N_2199,In_39,In_1319);
nor U2200 (N_2200,In_1204,In_1138);
xor U2201 (N_2201,In_1053,In_338);
xnor U2202 (N_2202,In_1074,In_1097);
nand U2203 (N_2203,In_1779,In_1274);
nor U2204 (N_2204,In_1882,In_52);
nand U2205 (N_2205,In_1628,In_1228);
and U2206 (N_2206,In_2154,In_323);
and U2207 (N_2207,In_123,In_2074);
nand U2208 (N_2208,In_679,In_282);
xnor U2209 (N_2209,In_1676,In_1331);
nor U2210 (N_2210,In_511,In_1770);
nand U2211 (N_2211,In_1077,In_20);
or U2212 (N_2212,In_848,In_1234);
or U2213 (N_2213,In_1784,In_2212);
nand U2214 (N_2214,In_442,In_998);
and U2215 (N_2215,In_1779,In_843);
nand U2216 (N_2216,In_1378,In_693);
nor U2217 (N_2217,In_23,In_1664);
xor U2218 (N_2218,In_1937,In_1481);
nand U2219 (N_2219,In_1412,In_643);
xor U2220 (N_2220,In_1975,In_2052);
or U2221 (N_2221,In_1009,In_1280);
xnor U2222 (N_2222,In_1828,In_2281);
and U2223 (N_2223,In_1772,In_638);
and U2224 (N_2224,In_228,In_1114);
and U2225 (N_2225,In_1250,In_1562);
xnor U2226 (N_2226,In_2115,In_1045);
or U2227 (N_2227,In_1660,In_1302);
or U2228 (N_2228,In_288,In_1973);
xnor U2229 (N_2229,In_808,In_2220);
nand U2230 (N_2230,In_1401,In_1764);
nand U2231 (N_2231,In_102,In_1148);
and U2232 (N_2232,In_1560,In_1295);
or U2233 (N_2233,In_2311,In_1345);
xor U2234 (N_2234,In_2081,In_607);
xnor U2235 (N_2235,In_698,In_1694);
xor U2236 (N_2236,In_844,In_1009);
or U2237 (N_2237,In_1791,In_1043);
xnor U2238 (N_2238,In_1659,In_2323);
nand U2239 (N_2239,In_806,In_931);
nor U2240 (N_2240,In_1259,In_1785);
nand U2241 (N_2241,In_2496,In_2265);
xor U2242 (N_2242,In_27,In_1523);
xor U2243 (N_2243,In_750,In_2140);
nand U2244 (N_2244,In_765,In_599);
xnor U2245 (N_2245,In_904,In_1208);
nor U2246 (N_2246,In_131,In_149);
nor U2247 (N_2247,In_2358,In_1187);
xor U2248 (N_2248,In_1048,In_808);
nand U2249 (N_2249,In_1898,In_1647);
and U2250 (N_2250,In_1381,In_1868);
nand U2251 (N_2251,In_1566,In_1846);
xnor U2252 (N_2252,In_1651,In_1283);
or U2253 (N_2253,In_1116,In_1054);
nor U2254 (N_2254,In_2059,In_883);
or U2255 (N_2255,In_1344,In_1297);
nand U2256 (N_2256,In_1423,In_1780);
xor U2257 (N_2257,In_1562,In_993);
nor U2258 (N_2258,In_1156,In_1401);
or U2259 (N_2259,In_519,In_2058);
nor U2260 (N_2260,In_1854,In_2486);
xor U2261 (N_2261,In_1174,In_1532);
nor U2262 (N_2262,In_2213,In_688);
xor U2263 (N_2263,In_2375,In_756);
and U2264 (N_2264,In_1972,In_1837);
nand U2265 (N_2265,In_1098,In_2100);
or U2266 (N_2266,In_1111,In_1008);
nor U2267 (N_2267,In_1436,In_1571);
nor U2268 (N_2268,In_2227,In_2172);
or U2269 (N_2269,In_1349,In_598);
or U2270 (N_2270,In_454,In_778);
nand U2271 (N_2271,In_1024,In_1773);
nand U2272 (N_2272,In_1764,In_2235);
nand U2273 (N_2273,In_1657,In_1530);
nand U2274 (N_2274,In_2262,In_2467);
or U2275 (N_2275,In_683,In_698);
nand U2276 (N_2276,In_2075,In_1069);
nor U2277 (N_2277,In_2460,In_2187);
xnor U2278 (N_2278,In_1033,In_1569);
nor U2279 (N_2279,In_2217,In_1017);
nand U2280 (N_2280,In_693,In_2144);
and U2281 (N_2281,In_138,In_1741);
or U2282 (N_2282,In_1994,In_542);
nor U2283 (N_2283,In_445,In_167);
and U2284 (N_2284,In_193,In_1916);
and U2285 (N_2285,In_79,In_1343);
or U2286 (N_2286,In_433,In_1419);
nand U2287 (N_2287,In_817,In_647);
and U2288 (N_2288,In_2170,In_1326);
xnor U2289 (N_2289,In_1900,In_2462);
or U2290 (N_2290,In_954,In_218);
nand U2291 (N_2291,In_2292,In_2128);
nand U2292 (N_2292,In_433,In_2148);
xor U2293 (N_2293,In_947,In_572);
or U2294 (N_2294,In_603,In_643);
or U2295 (N_2295,In_1534,In_2432);
nor U2296 (N_2296,In_1728,In_823);
nor U2297 (N_2297,In_1743,In_1572);
xor U2298 (N_2298,In_1689,In_6);
xor U2299 (N_2299,In_2006,In_2164);
or U2300 (N_2300,In_2417,In_17);
or U2301 (N_2301,In_808,In_735);
nand U2302 (N_2302,In_2340,In_2262);
nand U2303 (N_2303,In_616,In_1858);
xnor U2304 (N_2304,In_2425,In_2248);
xnor U2305 (N_2305,In_1547,In_732);
xor U2306 (N_2306,In_1103,In_1020);
xnor U2307 (N_2307,In_907,In_2266);
or U2308 (N_2308,In_265,In_1561);
and U2309 (N_2309,In_347,In_2167);
nor U2310 (N_2310,In_384,In_392);
and U2311 (N_2311,In_450,In_2451);
or U2312 (N_2312,In_89,In_1217);
nand U2313 (N_2313,In_186,In_664);
nand U2314 (N_2314,In_552,In_1621);
and U2315 (N_2315,In_1711,In_1753);
nor U2316 (N_2316,In_1353,In_884);
or U2317 (N_2317,In_1293,In_703);
nand U2318 (N_2318,In_1271,In_1766);
nand U2319 (N_2319,In_350,In_1026);
nand U2320 (N_2320,In_1206,In_1369);
and U2321 (N_2321,In_1614,In_772);
xnor U2322 (N_2322,In_2140,In_1025);
and U2323 (N_2323,In_2032,In_715);
nand U2324 (N_2324,In_55,In_83);
nor U2325 (N_2325,In_1783,In_1142);
nor U2326 (N_2326,In_708,In_1026);
nor U2327 (N_2327,In_982,In_1802);
xnor U2328 (N_2328,In_185,In_2427);
xnor U2329 (N_2329,In_232,In_2071);
xnor U2330 (N_2330,In_1725,In_616);
nor U2331 (N_2331,In_521,In_628);
xor U2332 (N_2332,In_615,In_1283);
xnor U2333 (N_2333,In_1477,In_1204);
and U2334 (N_2334,In_1781,In_1438);
or U2335 (N_2335,In_92,In_1945);
and U2336 (N_2336,In_554,In_1835);
xnor U2337 (N_2337,In_1189,In_2468);
xnor U2338 (N_2338,In_768,In_896);
or U2339 (N_2339,In_5,In_1116);
or U2340 (N_2340,In_1330,In_1777);
nand U2341 (N_2341,In_427,In_1143);
and U2342 (N_2342,In_1811,In_1557);
nor U2343 (N_2343,In_1811,In_1947);
and U2344 (N_2344,In_2052,In_1715);
xor U2345 (N_2345,In_1439,In_1051);
or U2346 (N_2346,In_841,In_687);
and U2347 (N_2347,In_1236,In_1306);
nor U2348 (N_2348,In_309,In_2295);
xnor U2349 (N_2349,In_1224,In_1407);
xnor U2350 (N_2350,In_691,In_161);
xor U2351 (N_2351,In_634,In_1023);
and U2352 (N_2352,In_1137,In_335);
or U2353 (N_2353,In_2340,In_1486);
xor U2354 (N_2354,In_65,In_1464);
nand U2355 (N_2355,In_601,In_2193);
and U2356 (N_2356,In_1556,In_1808);
xor U2357 (N_2357,In_2414,In_1302);
nor U2358 (N_2358,In_541,In_212);
or U2359 (N_2359,In_2368,In_985);
nor U2360 (N_2360,In_730,In_111);
nor U2361 (N_2361,In_2348,In_1564);
and U2362 (N_2362,In_825,In_1464);
or U2363 (N_2363,In_795,In_2057);
and U2364 (N_2364,In_1042,In_1393);
xnor U2365 (N_2365,In_1705,In_1220);
nand U2366 (N_2366,In_1490,In_2262);
and U2367 (N_2367,In_21,In_78);
xnor U2368 (N_2368,In_868,In_1937);
and U2369 (N_2369,In_1213,In_1407);
nor U2370 (N_2370,In_429,In_1801);
nand U2371 (N_2371,In_2030,In_1370);
nand U2372 (N_2372,In_654,In_1340);
nand U2373 (N_2373,In_1269,In_623);
nand U2374 (N_2374,In_1254,In_2293);
or U2375 (N_2375,In_2152,In_41);
nand U2376 (N_2376,In_1021,In_2337);
xnor U2377 (N_2377,In_2065,In_1479);
or U2378 (N_2378,In_819,In_1215);
and U2379 (N_2379,In_1003,In_112);
nand U2380 (N_2380,In_1041,In_2436);
or U2381 (N_2381,In_1432,In_1313);
or U2382 (N_2382,In_1879,In_2165);
nor U2383 (N_2383,In_902,In_1007);
xnor U2384 (N_2384,In_1317,In_2314);
nor U2385 (N_2385,In_2057,In_1925);
xor U2386 (N_2386,In_1407,In_204);
nor U2387 (N_2387,In_224,In_832);
nor U2388 (N_2388,In_1351,In_1897);
nor U2389 (N_2389,In_2118,In_322);
and U2390 (N_2390,In_2285,In_2362);
nor U2391 (N_2391,In_1738,In_1694);
xor U2392 (N_2392,In_1918,In_1885);
and U2393 (N_2393,In_1493,In_1695);
nand U2394 (N_2394,In_1858,In_165);
xor U2395 (N_2395,In_68,In_1130);
xor U2396 (N_2396,In_98,In_544);
and U2397 (N_2397,In_774,In_1565);
and U2398 (N_2398,In_149,In_1975);
xnor U2399 (N_2399,In_2097,In_328);
or U2400 (N_2400,In_177,In_1049);
nand U2401 (N_2401,In_24,In_456);
nand U2402 (N_2402,In_969,In_1256);
nor U2403 (N_2403,In_392,In_2238);
nor U2404 (N_2404,In_702,In_2415);
and U2405 (N_2405,In_2263,In_1366);
nor U2406 (N_2406,In_559,In_1524);
nand U2407 (N_2407,In_1775,In_1423);
nand U2408 (N_2408,In_579,In_2281);
or U2409 (N_2409,In_1354,In_1577);
and U2410 (N_2410,In_2051,In_2286);
or U2411 (N_2411,In_2095,In_287);
nor U2412 (N_2412,In_2205,In_844);
xnor U2413 (N_2413,In_1888,In_1487);
or U2414 (N_2414,In_161,In_739);
xnor U2415 (N_2415,In_1921,In_705);
nand U2416 (N_2416,In_2026,In_1390);
xor U2417 (N_2417,In_2395,In_983);
xnor U2418 (N_2418,In_411,In_125);
or U2419 (N_2419,In_1323,In_773);
nor U2420 (N_2420,In_728,In_884);
or U2421 (N_2421,In_1711,In_1503);
xor U2422 (N_2422,In_1054,In_2146);
xnor U2423 (N_2423,In_123,In_565);
nand U2424 (N_2424,In_1457,In_1197);
nand U2425 (N_2425,In_365,In_2389);
or U2426 (N_2426,In_425,In_870);
and U2427 (N_2427,In_2475,In_2018);
nand U2428 (N_2428,In_687,In_399);
nand U2429 (N_2429,In_2373,In_97);
nand U2430 (N_2430,In_229,In_2399);
xor U2431 (N_2431,In_1163,In_533);
xnor U2432 (N_2432,In_1776,In_2260);
xor U2433 (N_2433,In_694,In_1955);
nor U2434 (N_2434,In_1673,In_1679);
nand U2435 (N_2435,In_2135,In_180);
xnor U2436 (N_2436,In_548,In_1829);
or U2437 (N_2437,In_18,In_2317);
nor U2438 (N_2438,In_1786,In_861);
xor U2439 (N_2439,In_749,In_2083);
and U2440 (N_2440,In_739,In_564);
and U2441 (N_2441,In_1639,In_395);
and U2442 (N_2442,In_1174,In_1023);
or U2443 (N_2443,In_666,In_376);
or U2444 (N_2444,In_771,In_402);
and U2445 (N_2445,In_25,In_2110);
xor U2446 (N_2446,In_178,In_2130);
or U2447 (N_2447,In_1324,In_1243);
and U2448 (N_2448,In_361,In_1078);
nand U2449 (N_2449,In_1982,In_660);
xnor U2450 (N_2450,In_731,In_1640);
nand U2451 (N_2451,In_607,In_2486);
and U2452 (N_2452,In_1425,In_1022);
nand U2453 (N_2453,In_56,In_1021);
or U2454 (N_2454,In_326,In_1173);
nand U2455 (N_2455,In_910,In_343);
nor U2456 (N_2456,In_1021,In_710);
nand U2457 (N_2457,In_550,In_1630);
or U2458 (N_2458,In_1082,In_2156);
nor U2459 (N_2459,In_1973,In_1152);
or U2460 (N_2460,In_440,In_1310);
xor U2461 (N_2461,In_2116,In_2204);
and U2462 (N_2462,In_905,In_37);
nand U2463 (N_2463,In_852,In_2419);
nor U2464 (N_2464,In_270,In_85);
nand U2465 (N_2465,In_370,In_1127);
nor U2466 (N_2466,In_679,In_809);
or U2467 (N_2467,In_543,In_325);
xnor U2468 (N_2468,In_411,In_288);
nor U2469 (N_2469,In_2345,In_566);
nand U2470 (N_2470,In_133,In_254);
nor U2471 (N_2471,In_2467,In_1155);
or U2472 (N_2472,In_306,In_1185);
xor U2473 (N_2473,In_1405,In_2401);
xnor U2474 (N_2474,In_42,In_370);
and U2475 (N_2475,In_1622,In_590);
and U2476 (N_2476,In_939,In_1124);
nand U2477 (N_2477,In_814,In_1430);
nor U2478 (N_2478,In_1683,In_1980);
nand U2479 (N_2479,In_2159,In_234);
and U2480 (N_2480,In_2294,In_64);
and U2481 (N_2481,In_2131,In_1748);
xnor U2482 (N_2482,In_1143,In_1047);
nor U2483 (N_2483,In_1415,In_1992);
or U2484 (N_2484,In_1624,In_129);
or U2485 (N_2485,In_850,In_2070);
nand U2486 (N_2486,In_1422,In_1188);
xnor U2487 (N_2487,In_844,In_558);
and U2488 (N_2488,In_434,In_415);
and U2489 (N_2489,In_1963,In_2353);
xor U2490 (N_2490,In_1769,In_866);
and U2491 (N_2491,In_130,In_944);
or U2492 (N_2492,In_1646,In_1294);
nand U2493 (N_2493,In_1906,In_936);
and U2494 (N_2494,In_18,In_2027);
or U2495 (N_2495,In_2115,In_2076);
nor U2496 (N_2496,In_1249,In_1532);
and U2497 (N_2497,In_2339,In_1553);
xnor U2498 (N_2498,In_830,In_391);
nor U2499 (N_2499,In_601,In_1789);
and U2500 (N_2500,In_695,In_303);
or U2501 (N_2501,In_2421,In_1397);
nor U2502 (N_2502,In_127,In_164);
xor U2503 (N_2503,In_1117,In_2023);
xor U2504 (N_2504,In_2090,In_1829);
or U2505 (N_2505,In_2362,In_1319);
or U2506 (N_2506,In_1822,In_1444);
or U2507 (N_2507,In_932,In_2251);
or U2508 (N_2508,In_1756,In_1108);
xor U2509 (N_2509,In_750,In_2169);
and U2510 (N_2510,In_297,In_1305);
and U2511 (N_2511,In_1592,In_595);
xnor U2512 (N_2512,In_1773,In_114);
xnor U2513 (N_2513,In_365,In_1355);
or U2514 (N_2514,In_1027,In_1456);
or U2515 (N_2515,In_968,In_597);
xor U2516 (N_2516,In_2071,In_1814);
nor U2517 (N_2517,In_696,In_241);
or U2518 (N_2518,In_1228,In_2147);
or U2519 (N_2519,In_829,In_585);
and U2520 (N_2520,In_587,In_2091);
and U2521 (N_2521,In_115,In_1043);
and U2522 (N_2522,In_1206,In_1848);
or U2523 (N_2523,In_1124,In_2312);
xnor U2524 (N_2524,In_1056,In_2257);
xor U2525 (N_2525,In_1808,In_2453);
or U2526 (N_2526,In_2430,In_489);
xnor U2527 (N_2527,In_2378,In_1102);
or U2528 (N_2528,In_475,In_2411);
and U2529 (N_2529,In_170,In_1738);
nor U2530 (N_2530,In_110,In_854);
xor U2531 (N_2531,In_1198,In_2140);
xor U2532 (N_2532,In_1557,In_2001);
nor U2533 (N_2533,In_1084,In_1065);
nand U2534 (N_2534,In_259,In_1412);
or U2535 (N_2535,In_1553,In_2470);
xor U2536 (N_2536,In_1547,In_1166);
xnor U2537 (N_2537,In_1960,In_2285);
xor U2538 (N_2538,In_1772,In_1204);
nor U2539 (N_2539,In_185,In_573);
or U2540 (N_2540,In_522,In_2306);
nor U2541 (N_2541,In_1509,In_1008);
or U2542 (N_2542,In_2479,In_77);
nor U2543 (N_2543,In_271,In_1019);
nand U2544 (N_2544,In_554,In_550);
and U2545 (N_2545,In_2315,In_758);
and U2546 (N_2546,In_1691,In_2103);
nor U2547 (N_2547,In_693,In_1766);
or U2548 (N_2548,In_353,In_1951);
nor U2549 (N_2549,In_1796,In_147);
nand U2550 (N_2550,In_2028,In_762);
nor U2551 (N_2551,In_584,In_2122);
nor U2552 (N_2552,In_136,In_780);
and U2553 (N_2553,In_1816,In_2222);
and U2554 (N_2554,In_1822,In_2353);
nand U2555 (N_2555,In_2386,In_2415);
xor U2556 (N_2556,In_418,In_832);
xor U2557 (N_2557,In_692,In_2037);
nand U2558 (N_2558,In_656,In_2342);
nand U2559 (N_2559,In_1049,In_676);
or U2560 (N_2560,In_2422,In_0);
xnor U2561 (N_2561,In_2365,In_1219);
nand U2562 (N_2562,In_1516,In_1161);
or U2563 (N_2563,In_608,In_726);
nor U2564 (N_2564,In_1551,In_2116);
and U2565 (N_2565,In_452,In_1952);
xnor U2566 (N_2566,In_1732,In_1609);
and U2567 (N_2567,In_1948,In_1114);
nand U2568 (N_2568,In_960,In_2434);
or U2569 (N_2569,In_1003,In_379);
and U2570 (N_2570,In_1857,In_370);
xor U2571 (N_2571,In_769,In_1972);
xor U2572 (N_2572,In_2200,In_1058);
or U2573 (N_2573,In_623,In_157);
nor U2574 (N_2574,In_639,In_184);
xnor U2575 (N_2575,In_1301,In_1460);
nor U2576 (N_2576,In_2376,In_1887);
or U2577 (N_2577,In_592,In_2277);
nor U2578 (N_2578,In_209,In_1481);
nor U2579 (N_2579,In_76,In_317);
and U2580 (N_2580,In_1655,In_2343);
nand U2581 (N_2581,In_365,In_377);
or U2582 (N_2582,In_1865,In_1528);
or U2583 (N_2583,In_1746,In_255);
and U2584 (N_2584,In_935,In_145);
xor U2585 (N_2585,In_851,In_1572);
xnor U2586 (N_2586,In_1938,In_74);
nand U2587 (N_2587,In_919,In_937);
or U2588 (N_2588,In_1679,In_1989);
nand U2589 (N_2589,In_2404,In_664);
nor U2590 (N_2590,In_55,In_831);
nand U2591 (N_2591,In_2037,In_2012);
or U2592 (N_2592,In_348,In_1480);
xnor U2593 (N_2593,In_2417,In_2211);
nor U2594 (N_2594,In_640,In_828);
nand U2595 (N_2595,In_1536,In_2132);
nor U2596 (N_2596,In_910,In_1409);
xor U2597 (N_2597,In_79,In_859);
nor U2598 (N_2598,In_1369,In_530);
and U2599 (N_2599,In_1088,In_1991);
and U2600 (N_2600,In_1644,In_64);
and U2601 (N_2601,In_644,In_1813);
and U2602 (N_2602,In_1240,In_3);
xnor U2603 (N_2603,In_1654,In_2349);
xnor U2604 (N_2604,In_1504,In_59);
xnor U2605 (N_2605,In_2119,In_1945);
nor U2606 (N_2606,In_698,In_13);
xnor U2607 (N_2607,In_1117,In_157);
and U2608 (N_2608,In_1408,In_1457);
or U2609 (N_2609,In_2446,In_1126);
and U2610 (N_2610,In_1330,In_428);
nor U2611 (N_2611,In_1876,In_697);
or U2612 (N_2612,In_2333,In_2030);
or U2613 (N_2613,In_1585,In_1060);
nor U2614 (N_2614,In_1616,In_1087);
or U2615 (N_2615,In_1025,In_1175);
or U2616 (N_2616,In_2122,In_1022);
nor U2617 (N_2617,In_667,In_1473);
or U2618 (N_2618,In_2117,In_2138);
nand U2619 (N_2619,In_1303,In_1099);
and U2620 (N_2620,In_1238,In_2146);
nand U2621 (N_2621,In_673,In_2195);
nor U2622 (N_2622,In_533,In_2363);
nor U2623 (N_2623,In_1378,In_1031);
or U2624 (N_2624,In_1471,In_2263);
or U2625 (N_2625,In_597,In_337);
xnor U2626 (N_2626,In_1700,In_450);
nand U2627 (N_2627,In_391,In_41);
nand U2628 (N_2628,In_1088,In_443);
xor U2629 (N_2629,In_84,In_2043);
xnor U2630 (N_2630,In_1568,In_459);
nor U2631 (N_2631,In_489,In_944);
nand U2632 (N_2632,In_1083,In_1545);
nor U2633 (N_2633,In_489,In_1210);
nor U2634 (N_2634,In_363,In_779);
xor U2635 (N_2635,In_616,In_1327);
nor U2636 (N_2636,In_1820,In_184);
xor U2637 (N_2637,In_3,In_474);
or U2638 (N_2638,In_811,In_1153);
nor U2639 (N_2639,In_752,In_1350);
nand U2640 (N_2640,In_524,In_2167);
nand U2641 (N_2641,In_162,In_1377);
nand U2642 (N_2642,In_719,In_1278);
xnor U2643 (N_2643,In_2024,In_934);
nor U2644 (N_2644,In_1825,In_873);
and U2645 (N_2645,In_1640,In_1600);
and U2646 (N_2646,In_1166,In_2324);
and U2647 (N_2647,In_1977,In_2475);
nand U2648 (N_2648,In_843,In_274);
xor U2649 (N_2649,In_223,In_2243);
nor U2650 (N_2650,In_2020,In_1040);
xor U2651 (N_2651,In_531,In_103);
nor U2652 (N_2652,In_491,In_329);
nand U2653 (N_2653,In_2000,In_1945);
nor U2654 (N_2654,In_371,In_1418);
xor U2655 (N_2655,In_1291,In_2244);
xnor U2656 (N_2656,In_154,In_2014);
and U2657 (N_2657,In_1543,In_1782);
nor U2658 (N_2658,In_2233,In_340);
xor U2659 (N_2659,In_342,In_363);
nand U2660 (N_2660,In_1105,In_2035);
nand U2661 (N_2661,In_2075,In_266);
nor U2662 (N_2662,In_767,In_2392);
nor U2663 (N_2663,In_2145,In_2284);
nand U2664 (N_2664,In_1321,In_1661);
nor U2665 (N_2665,In_2442,In_491);
or U2666 (N_2666,In_2272,In_1426);
and U2667 (N_2667,In_1157,In_702);
and U2668 (N_2668,In_1185,In_1474);
or U2669 (N_2669,In_2127,In_1461);
or U2670 (N_2670,In_1029,In_1744);
xor U2671 (N_2671,In_1137,In_585);
nand U2672 (N_2672,In_1275,In_1024);
nand U2673 (N_2673,In_2239,In_801);
nand U2674 (N_2674,In_2363,In_2435);
nand U2675 (N_2675,In_534,In_2047);
and U2676 (N_2676,In_2166,In_1675);
nand U2677 (N_2677,In_2016,In_1574);
and U2678 (N_2678,In_1842,In_247);
nor U2679 (N_2679,In_2410,In_464);
and U2680 (N_2680,In_1640,In_1967);
xor U2681 (N_2681,In_367,In_499);
or U2682 (N_2682,In_913,In_1393);
nand U2683 (N_2683,In_2195,In_312);
nor U2684 (N_2684,In_67,In_1422);
or U2685 (N_2685,In_1018,In_1633);
or U2686 (N_2686,In_2258,In_1503);
and U2687 (N_2687,In_635,In_1615);
and U2688 (N_2688,In_775,In_773);
or U2689 (N_2689,In_1538,In_304);
and U2690 (N_2690,In_1628,In_692);
xor U2691 (N_2691,In_2333,In_1135);
nor U2692 (N_2692,In_1094,In_1293);
and U2693 (N_2693,In_1175,In_819);
and U2694 (N_2694,In_264,In_565);
and U2695 (N_2695,In_1679,In_1295);
nand U2696 (N_2696,In_79,In_468);
nor U2697 (N_2697,In_849,In_1076);
and U2698 (N_2698,In_7,In_2354);
xnor U2699 (N_2699,In_402,In_2231);
xnor U2700 (N_2700,In_858,In_1045);
and U2701 (N_2701,In_147,In_2359);
nor U2702 (N_2702,In_866,In_1174);
xnor U2703 (N_2703,In_436,In_2484);
and U2704 (N_2704,In_2132,In_427);
nand U2705 (N_2705,In_1139,In_817);
xor U2706 (N_2706,In_1347,In_658);
or U2707 (N_2707,In_2448,In_1785);
xor U2708 (N_2708,In_2119,In_497);
nor U2709 (N_2709,In_2185,In_972);
and U2710 (N_2710,In_428,In_2311);
and U2711 (N_2711,In_1915,In_1945);
nor U2712 (N_2712,In_2022,In_2225);
xor U2713 (N_2713,In_2259,In_2472);
and U2714 (N_2714,In_1575,In_362);
or U2715 (N_2715,In_1135,In_317);
nor U2716 (N_2716,In_1130,In_1844);
xor U2717 (N_2717,In_476,In_2177);
nor U2718 (N_2718,In_264,In_2200);
nand U2719 (N_2719,In_1167,In_1745);
and U2720 (N_2720,In_1554,In_1965);
or U2721 (N_2721,In_1496,In_1071);
or U2722 (N_2722,In_1353,In_560);
nand U2723 (N_2723,In_1308,In_113);
xor U2724 (N_2724,In_353,In_1077);
nor U2725 (N_2725,In_1489,In_316);
or U2726 (N_2726,In_2477,In_1598);
or U2727 (N_2727,In_2113,In_25);
and U2728 (N_2728,In_1620,In_310);
nor U2729 (N_2729,In_540,In_1482);
nand U2730 (N_2730,In_1189,In_210);
or U2731 (N_2731,In_1989,In_2027);
and U2732 (N_2732,In_2278,In_406);
xor U2733 (N_2733,In_2028,In_2402);
nor U2734 (N_2734,In_1524,In_747);
xnor U2735 (N_2735,In_682,In_122);
xnor U2736 (N_2736,In_1027,In_1689);
and U2737 (N_2737,In_1167,In_2434);
nand U2738 (N_2738,In_247,In_2461);
nand U2739 (N_2739,In_679,In_1198);
nor U2740 (N_2740,In_649,In_1937);
and U2741 (N_2741,In_2253,In_1093);
or U2742 (N_2742,In_2191,In_2329);
nor U2743 (N_2743,In_1681,In_974);
xnor U2744 (N_2744,In_1594,In_1602);
and U2745 (N_2745,In_1071,In_2241);
xor U2746 (N_2746,In_2065,In_5);
nor U2747 (N_2747,In_1621,In_85);
or U2748 (N_2748,In_1845,In_787);
xor U2749 (N_2749,In_350,In_293);
nor U2750 (N_2750,In_465,In_295);
xor U2751 (N_2751,In_490,In_1048);
xnor U2752 (N_2752,In_1086,In_1174);
and U2753 (N_2753,In_826,In_947);
nand U2754 (N_2754,In_934,In_2093);
nor U2755 (N_2755,In_610,In_112);
and U2756 (N_2756,In_381,In_330);
nand U2757 (N_2757,In_1723,In_1485);
and U2758 (N_2758,In_2158,In_1020);
xor U2759 (N_2759,In_885,In_1892);
xor U2760 (N_2760,In_1919,In_1369);
xnor U2761 (N_2761,In_292,In_1974);
and U2762 (N_2762,In_354,In_1281);
xnor U2763 (N_2763,In_1111,In_1026);
and U2764 (N_2764,In_1112,In_1505);
and U2765 (N_2765,In_973,In_2222);
nor U2766 (N_2766,In_1024,In_236);
xnor U2767 (N_2767,In_1383,In_893);
nor U2768 (N_2768,In_1147,In_2008);
or U2769 (N_2769,In_1450,In_1934);
xnor U2770 (N_2770,In_2370,In_1155);
xor U2771 (N_2771,In_1624,In_1211);
and U2772 (N_2772,In_869,In_1003);
nand U2773 (N_2773,In_2363,In_2307);
nor U2774 (N_2774,In_2232,In_801);
or U2775 (N_2775,In_618,In_2085);
nor U2776 (N_2776,In_2492,In_1330);
nor U2777 (N_2777,In_876,In_1938);
xor U2778 (N_2778,In_807,In_177);
nor U2779 (N_2779,In_991,In_805);
nor U2780 (N_2780,In_2148,In_677);
xnor U2781 (N_2781,In_1393,In_1003);
xnor U2782 (N_2782,In_2457,In_1604);
nand U2783 (N_2783,In_2221,In_2425);
or U2784 (N_2784,In_506,In_1496);
xor U2785 (N_2785,In_1530,In_1851);
xnor U2786 (N_2786,In_1075,In_2369);
nor U2787 (N_2787,In_572,In_479);
nor U2788 (N_2788,In_358,In_825);
and U2789 (N_2789,In_2018,In_386);
nor U2790 (N_2790,In_565,In_580);
xor U2791 (N_2791,In_1744,In_456);
or U2792 (N_2792,In_1130,In_2351);
nand U2793 (N_2793,In_2217,In_1088);
xor U2794 (N_2794,In_1324,In_1515);
and U2795 (N_2795,In_53,In_750);
nand U2796 (N_2796,In_1579,In_1158);
nor U2797 (N_2797,In_554,In_72);
nand U2798 (N_2798,In_1165,In_1413);
or U2799 (N_2799,In_2006,In_1685);
and U2800 (N_2800,In_847,In_315);
or U2801 (N_2801,In_651,In_1292);
nand U2802 (N_2802,In_1706,In_762);
or U2803 (N_2803,In_76,In_1370);
nand U2804 (N_2804,In_1089,In_1476);
nand U2805 (N_2805,In_874,In_1560);
nand U2806 (N_2806,In_553,In_2035);
xor U2807 (N_2807,In_1791,In_862);
or U2808 (N_2808,In_1550,In_2051);
xor U2809 (N_2809,In_1542,In_951);
and U2810 (N_2810,In_1364,In_2015);
and U2811 (N_2811,In_1436,In_659);
nor U2812 (N_2812,In_2418,In_1983);
and U2813 (N_2813,In_182,In_447);
or U2814 (N_2814,In_1188,In_1211);
xnor U2815 (N_2815,In_1642,In_1348);
or U2816 (N_2816,In_1445,In_1646);
nor U2817 (N_2817,In_2344,In_688);
nand U2818 (N_2818,In_2393,In_414);
xor U2819 (N_2819,In_2143,In_448);
and U2820 (N_2820,In_1489,In_329);
nor U2821 (N_2821,In_1661,In_1711);
nor U2822 (N_2822,In_241,In_1651);
or U2823 (N_2823,In_1754,In_1842);
nand U2824 (N_2824,In_1770,In_2017);
nand U2825 (N_2825,In_1852,In_1750);
or U2826 (N_2826,In_1655,In_1487);
or U2827 (N_2827,In_2114,In_714);
or U2828 (N_2828,In_1793,In_994);
nand U2829 (N_2829,In_211,In_1790);
or U2830 (N_2830,In_2083,In_811);
nand U2831 (N_2831,In_1861,In_2362);
nand U2832 (N_2832,In_1433,In_200);
nor U2833 (N_2833,In_1353,In_626);
nand U2834 (N_2834,In_2412,In_1555);
xor U2835 (N_2835,In_312,In_1620);
nand U2836 (N_2836,In_1823,In_310);
nor U2837 (N_2837,In_1481,In_1325);
and U2838 (N_2838,In_465,In_1602);
nand U2839 (N_2839,In_538,In_2341);
and U2840 (N_2840,In_267,In_237);
nor U2841 (N_2841,In_2208,In_2003);
nand U2842 (N_2842,In_2228,In_218);
and U2843 (N_2843,In_683,In_2406);
or U2844 (N_2844,In_1910,In_2216);
xor U2845 (N_2845,In_900,In_1765);
and U2846 (N_2846,In_1478,In_383);
nor U2847 (N_2847,In_2093,In_871);
nor U2848 (N_2848,In_162,In_571);
or U2849 (N_2849,In_305,In_1694);
or U2850 (N_2850,In_409,In_677);
nor U2851 (N_2851,In_2054,In_1838);
or U2852 (N_2852,In_1414,In_1219);
and U2853 (N_2853,In_2033,In_2095);
nand U2854 (N_2854,In_116,In_1652);
and U2855 (N_2855,In_1244,In_681);
xor U2856 (N_2856,In_608,In_2192);
xor U2857 (N_2857,In_1652,In_1145);
and U2858 (N_2858,In_1951,In_327);
or U2859 (N_2859,In_279,In_2342);
nand U2860 (N_2860,In_314,In_2169);
xor U2861 (N_2861,In_1079,In_2127);
nand U2862 (N_2862,In_2260,In_1111);
and U2863 (N_2863,In_1652,In_2462);
nor U2864 (N_2864,In_1813,In_277);
xor U2865 (N_2865,In_368,In_995);
nor U2866 (N_2866,In_2421,In_2433);
xor U2867 (N_2867,In_108,In_2027);
and U2868 (N_2868,In_2419,In_965);
xor U2869 (N_2869,In_2436,In_1672);
nand U2870 (N_2870,In_823,In_2166);
nand U2871 (N_2871,In_988,In_1282);
or U2872 (N_2872,In_599,In_1943);
xnor U2873 (N_2873,In_94,In_2323);
nand U2874 (N_2874,In_329,In_859);
or U2875 (N_2875,In_927,In_2057);
xnor U2876 (N_2876,In_1417,In_422);
nand U2877 (N_2877,In_1702,In_1260);
and U2878 (N_2878,In_1365,In_1064);
and U2879 (N_2879,In_549,In_1794);
nor U2880 (N_2880,In_363,In_1718);
or U2881 (N_2881,In_2382,In_1093);
and U2882 (N_2882,In_2228,In_2105);
nand U2883 (N_2883,In_806,In_2222);
or U2884 (N_2884,In_1577,In_1277);
nor U2885 (N_2885,In_1395,In_572);
xor U2886 (N_2886,In_288,In_1035);
or U2887 (N_2887,In_801,In_2474);
nand U2888 (N_2888,In_1721,In_2185);
and U2889 (N_2889,In_2472,In_245);
or U2890 (N_2890,In_626,In_2311);
xnor U2891 (N_2891,In_1583,In_625);
or U2892 (N_2892,In_328,In_1237);
nor U2893 (N_2893,In_1962,In_948);
nand U2894 (N_2894,In_1414,In_1168);
nor U2895 (N_2895,In_1696,In_1213);
xnor U2896 (N_2896,In_438,In_1174);
or U2897 (N_2897,In_947,In_1438);
xor U2898 (N_2898,In_608,In_125);
and U2899 (N_2899,In_1337,In_2094);
nor U2900 (N_2900,In_1497,In_1506);
xnor U2901 (N_2901,In_846,In_167);
nor U2902 (N_2902,In_653,In_1814);
nor U2903 (N_2903,In_254,In_1512);
and U2904 (N_2904,In_1481,In_611);
and U2905 (N_2905,In_600,In_2128);
or U2906 (N_2906,In_984,In_2141);
and U2907 (N_2907,In_1731,In_1821);
and U2908 (N_2908,In_1681,In_1769);
nand U2909 (N_2909,In_93,In_345);
xnor U2910 (N_2910,In_41,In_701);
xor U2911 (N_2911,In_1808,In_270);
or U2912 (N_2912,In_116,In_796);
nor U2913 (N_2913,In_1644,In_890);
or U2914 (N_2914,In_866,In_1128);
nor U2915 (N_2915,In_329,In_1163);
nand U2916 (N_2916,In_383,In_360);
xor U2917 (N_2917,In_1856,In_1022);
nand U2918 (N_2918,In_2102,In_1987);
xnor U2919 (N_2919,In_975,In_2135);
nand U2920 (N_2920,In_2474,In_1437);
nor U2921 (N_2921,In_120,In_1088);
and U2922 (N_2922,In_1199,In_370);
and U2923 (N_2923,In_2079,In_214);
or U2924 (N_2924,In_366,In_1344);
and U2925 (N_2925,In_761,In_448);
and U2926 (N_2926,In_995,In_565);
xnor U2927 (N_2927,In_1644,In_2489);
nor U2928 (N_2928,In_1064,In_1871);
nand U2929 (N_2929,In_1962,In_1850);
nand U2930 (N_2930,In_724,In_1173);
and U2931 (N_2931,In_1867,In_1984);
and U2932 (N_2932,In_2408,In_1610);
nor U2933 (N_2933,In_1717,In_302);
nor U2934 (N_2934,In_738,In_1996);
and U2935 (N_2935,In_32,In_1920);
nor U2936 (N_2936,In_307,In_2395);
or U2937 (N_2937,In_1160,In_2337);
or U2938 (N_2938,In_755,In_284);
xnor U2939 (N_2939,In_140,In_2463);
and U2940 (N_2940,In_198,In_1448);
xnor U2941 (N_2941,In_2483,In_1278);
nor U2942 (N_2942,In_1512,In_1499);
or U2943 (N_2943,In_1610,In_1292);
or U2944 (N_2944,In_2021,In_652);
nor U2945 (N_2945,In_1566,In_1717);
nand U2946 (N_2946,In_1000,In_413);
nor U2947 (N_2947,In_1925,In_977);
nand U2948 (N_2948,In_72,In_2421);
and U2949 (N_2949,In_616,In_575);
xor U2950 (N_2950,In_1035,In_1488);
and U2951 (N_2951,In_503,In_2468);
xor U2952 (N_2952,In_451,In_1774);
and U2953 (N_2953,In_2444,In_1195);
or U2954 (N_2954,In_659,In_808);
nand U2955 (N_2955,In_1286,In_1540);
nand U2956 (N_2956,In_866,In_621);
xnor U2957 (N_2957,In_2148,In_227);
nor U2958 (N_2958,In_2436,In_1360);
nor U2959 (N_2959,In_1608,In_816);
nor U2960 (N_2960,In_1230,In_1642);
xnor U2961 (N_2961,In_1677,In_298);
nand U2962 (N_2962,In_649,In_335);
nand U2963 (N_2963,In_856,In_2183);
xor U2964 (N_2964,In_2336,In_470);
or U2965 (N_2965,In_2462,In_969);
nand U2966 (N_2966,In_2265,In_1349);
or U2967 (N_2967,In_1142,In_2021);
nand U2968 (N_2968,In_2311,In_987);
or U2969 (N_2969,In_2066,In_384);
xor U2970 (N_2970,In_699,In_2318);
nor U2971 (N_2971,In_1159,In_1248);
or U2972 (N_2972,In_1855,In_2161);
or U2973 (N_2973,In_2151,In_1311);
xor U2974 (N_2974,In_118,In_2417);
xor U2975 (N_2975,In_272,In_1141);
xor U2976 (N_2976,In_2408,In_253);
nor U2977 (N_2977,In_470,In_421);
nand U2978 (N_2978,In_1663,In_512);
and U2979 (N_2979,In_1279,In_2332);
and U2980 (N_2980,In_956,In_685);
nand U2981 (N_2981,In_1938,In_1255);
or U2982 (N_2982,In_1378,In_299);
nor U2983 (N_2983,In_75,In_456);
nor U2984 (N_2984,In_1485,In_1487);
xnor U2985 (N_2985,In_1490,In_569);
or U2986 (N_2986,In_345,In_1486);
and U2987 (N_2987,In_2161,In_570);
xnor U2988 (N_2988,In_1461,In_1753);
or U2989 (N_2989,In_337,In_153);
or U2990 (N_2990,In_2279,In_2471);
or U2991 (N_2991,In_1031,In_1929);
or U2992 (N_2992,In_1097,In_1999);
and U2993 (N_2993,In_711,In_6);
xnor U2994 (N_2994,In_1240,In_775);
nor U2995 (N_2995,In_2071,In_138);
nor U2996 (N_2996,In_197,In_1127);
and U2997 (N_2997,In_1732,In_1452);
xor U2998 (N_2998,In_707,In_437);
and U2999 (N_2999,In_1355,In_952);
nor U3000 (N_3000,In_502,In_2209);
nand U3001 (N_3001,In_476,In_734);
xnor U3002 (N_3002,In_167,In_314);
nand U3003 (N_3003,In_1415,In_1238);
xnor U3004 (N_3004,In_637,In_746);
nor U3005 (N_3005,In_975,In_1524);
nand U3006 (N_3006,In_1243,In_1924);
or U3007 (N_3007,In_1703,In_1036);
xnor U3008 (N_3008,In_999,In_1021);
nand U3009 (N_3009,In_168,In_1311);
nand U3010 (N_3010,In_1064,In_1156);
nand U3011 (N_3011,In_1862,In_2236);
nor U3012 (N_3012,In_1280,In_241);
or U3013 (N_3013,In_1579,In_1825);
xnor U3014 (N_3014,In_1454,In_197);
xor U3015 (N_3015,In_892,In_2299);
nand U3016 (N_3016,In_1930,In_1822);
nor U3017 (N_3017,In_1883,In_2166);
or U3018 (N_3018,In_1326,In_2267);
nand U3019 (N_3019,In_1847,In_1752);
nor U3020 (N_3020,In_1965,In_192);
nand U3021 (N_3021,In_930,In_146);
and U3022 (N_3022,In_1646,In_242);
nand U3023 (N_3023,In_1161,In_1266);
or U3024 (N_3024,In_1536,In_1992);
and U3025 (N_3025,In_1903,In_2353);
xor U3026 (N_3026,In_1644,In_1963);
or U3027 (N_3027,In_1603,In_2154);
and U3028 (N_3028,In_2047,In_48);
xor U3029 (N_3029,In_1563,In_122);
nand U3030 (N_3030,In_591,In_2227);
or U3031 (N_3031,In_1954,In_9);
or U3032 (N_3032,In_862,In_1032);
or U3033 (N_3033,In_1954,In_1436);
or U3034 (N_3034,In_955,In_1529);
nand U3035 (N_3035,In_1145,In_389);
or U3036 (N_3036,In_1100,In_9);
nor U3037 (N_3037,In_595,In_1731);
xnor U3038 (N_3038,In_810,In_364);
and U3039 (N_3039,In_1991,In_1769);
nor U3040 (N_3040,In_1603,In_2070);
and U3041 (N_3041,In_2455,In_638);
nor U3042 (N_3042,In_597,In_2403);
and U3043 (N_3043,In_1216,In_1970);
and U3044 (N_3044,In_2407,In_1591);
or U3045 (N_3045,In_2361,In_1215);
and U3046 (N_3046,In_1272,In_273);
or U3047 (N_3047,In_2370,In_971);
xor U3048 (N_3048,In_1948,In_296);
nand U3049 (N_3049,In_1478,In_902);
nand U3050 (N_3050,In_2009,In_1850);
xnor U3051 (N_3051,In_1109,In_2297);
or U3052 (N_3052,In_208,In_244);
or U3053 (N_3053,In_375,In_1832);
nor U3054 (N_3054,In_110,In_1120);
nor U3055 (N_3055,In_2077,In_747);
and U3056 (N_3056,In_1205,In_1126);
and U3057 (N_3057,In_2454,In_1576);
and U3058 (N_3058,In_686,In_129);
and U3059 (N_3059,In_2294,In_2014);
nor U3060 (N_3060,In_73,In_2319);
and U3061 (N_3061,In_577,In_468);
nor U3062 (N_3062,In_456,In_2121);
nor U3063 (N_3063,In_348,In_2007);
nand U3064 (N_3064,In_1357,In_2320);
nand U3065 (N_3065,In_1004,In_2321);
and U3066 (N_3066,In_1329,In_700);
or U3067 (N_3067,In_2078,In_275);
nor U3068 (N_3068,In_2092,In_838);
nand U3069 (N_3069,In_806,In_2251);
and U3070 (N_3070,In_817,In_1881);
xor U3071 (N_3071,In_1890,In_2037);
nand U3072 (N_3072,In_279,In_1186);
and U3073 (N_3073,In_613,In_1221);
nand U3074 (N_3074,In_1217,In_1988);
xnor U3075 (N_3075,In_1123,In_104);
or U3076 (N_3076,In_275,In_407);
nand U3077 (N_3077,In_196,In_376);
xor U3078 (N_3078,In_686,In_1013);
xnor U3079 (N_3079,In_749,In_442);
nor U3080 (N_3080,In_2182,In_1249);
xor U3081 (N_3081,In_1145,In_849);
xnor U3082 (N_3082,In_1081,In_973);
nor U3083 (N_3083,In_2345,In_364);
and U3084 (N_3084,In_160,In_1570);
nand U3085 (N_3085,In_572,In_1839);
and U3086 (N_3086,In_2212,In_2267);
xnor U3087 (N_3087,In_1905,In_1622);
xnor U3088 (N_3088,In_346,In_1259);
nand U3089 (N_3089,In_2257,In_522);
or U3090 (N_3090,In_517,In_1406);
xnor U3091 (N_3091,In_304,In_1195);
and U3092 (N_3092,In_625,In_740);
and U3093 (N_3093,In_1856,In_670);
or U3094 (N_3094,In_1392,In_951);
or U3095 (N_3095,In_898,In_980);
and U3096 (N_3096,In_466,In_415);
nand U3097 (N_3097,In_423,In_614);
nor U3098 (N_3098,In_103,In_1839);
or U3099 (N_3099,In_2064,In_301);
or U3100 (N_3100,In_200,In_901);
and U3101 (N_3101,In_1579,In_1558);
xor U3102 (N_3102,In_1625,In_902);
xor U3103 (N_3103,In_1768,In_1851);
or U3104 (N_3104,In_2213,In_1191);
or U3105 (N_3105,In_767,In_2365);
xor U3106 (N_3106,In_174,In_906);
xor U3107 (N_3107,In_1997,In_1114);
nand U3108 (N_3108,In_95,In_2116);
nand U3109 (N_3109,In_565,In_2255);
and U3110 (N_3110,In_1675,In_2259);
and U3111 (N_3111,In_502,In_949);
xor U3112 (N_3112,In_1569,In_564);
xnor U3113 (N_3113,In_548,In_581);
or U3114 (N_3114,In_2069,In_285);
and U3115 (N_3115,In_1180,In_64);
nand U3116 (N_3116,In_171,In_796);
or U3117 (N_3117,In_1885,In_1692);
and U3118 (N_3118,In_946,In_589);
nand U3119 (N_3119,In_2373,In_1916);
nor U3120 (N_3120,In_1590,In_903);
nor U3121 (N_3121,In_1902,In_171);
nand U3122 (N_3122,In_714,In_96);
and U3123 (N_3123,In_207,In_1273);
xor U3124 (N_3124,In_1409,In_2012);
nand U3125 (N_3125,In_2269,In_621);
xnor U3126 (N_3126,In_1892,In_1179);
xor U3127 (N_3127,In_1628,In_2017);
and U3128 (N_3128,In_2001,In_2387);
and U3129 (N_3129,In_428,In_1341);
nand U3130 (N_3130,In_717,In_614);
nand U3131 (N_3131,In_26,In_2447);
xor U3132 (N_3132,In_2324,In_1077);
or U3133 (N_3133,In_1856,In_402);
and U3134 (N_3134,In_124,In_1508);
nor U3135 (N_3135,In_699,In_2471);
or U3136 (N_3136,In_973,In_439);
nor U3137 (N_3137,In_2300,In_676);
or U3138 (N_3138,In_493,In_2440);
nor U3139 (N_3139,In_97,In_800);
nor U3140 (N_3140,In_218,In_2421);
and U3141 (N_3141,In_1841,In_90);
nand U3142 (N_3142,In_1721,In_1601);
nand U3143 (N_3143,In_2153,In_218);
nand U3144 (N_3144,In_1547,In_1516);
xnor U3145 (N_3145,In_869,In_188);
nor U3146 (N_3146,In_1052,In_308);
xor U3147 (N_3147,In_1629,In_2013);
or U3148 (N_3148,In_118,In_1086);
and U3149 (N_3149,In_1639,In_306);
nand U3150 (N_3150,In_2045,In_1856);
xnor U3151 (N_3151,In_1232,In_1267);
and U3152 (N_3152,In_528,In_1632);
nor U3153 (N_3153,In_234,In_1122);
xor U3154 (N_3154,In_1690,In_1110);
and U3155 (N_3155,In_1269,In_1388);
xnor U3156 (N_3156,In_2006,In_1069);
and U3157 (N_3157,In_2474,In_1436);
and U3158 (N_3158,In_1888,In_2334);
or U3159 (N_3159,In_840,In_1122);
nor U3160 (N_3160,In_453,In_2123);
nor U3161 (N_3161,In_250,In_1346);
or U3162 (N_3162,In_374,In_877);
nand U3163 (N_3163,In_1521,In_463);
and U3164 (N_3164,In_1903,In_2318);
nor U3165 (N_3165,In_1721,In_2192);
and U3166 (N_3166,In_2037,In_467);
and U3167 (N_3167,In_1446,In_1111);
nand U3168 (N_3168,In_564,In_2483);
or U3169 (N_3169,In_2350,In_862);
nor U3170 (N_3170,In_2024,In_883);
nand U3171 (N_3171,In_2086,In_1130);
nand U3172 (N_3172,In_1518,In_621);
nor U3173 (N_3173,In_753,In_671);
nor U3174 (N_3174,In_1621,In_867);
xor U3175 (N_3175,In_1471,In_2114);
nand U3176 (N_3176,In_1037,In_626);
nand U3177 (N_3177,In_2191,In_387);
nor U3178 (N_3178,In_381,In_793);
xor U3179 (N_3179,In_234,In_2029);
nand U3180 (N_3180,In_2178,In_726);
nor U3181 (N_3181,In_142,In_657);
nand U3182 (N_3182,In_2330,In_1179);
or U3183 (N_3183,In_165,In_1426);
nor U3184 (N_3184,In_1566,In_1477);
xor U3185 (N_3185,In_1148,In_2058);
xor U3186 (N_3186,In_1161,In_2109);
xnor U3187 (N_3187,In_1600,In_2101);
nor U3188 (N_3188,In_2005,In_99);
nand U3189 (N_3189,In_953,In_304);
xor U3190 (N_3190,In_2204,In_2198);
and U3191 (N_3191,In_2338,In_887);
nand U3192 (N_3192,In_2185,In_963);
or U3193 (N_3193,In_1408,In_1814);
xor U3194 (N_3194,In_627,In_1798);
nand U3195 (N_3195,In_2296,In_413);
or U3196 (N_3196,In_553,In_964);
xor U3197 (N_3197,In_117,In_632);
nor U3198 (N_3198,In_1911,In_2143);
or U3199 (N_3199,In_1437,In_2206);
xnor U3200 (N_3200,In_2227,In_647);
or U3201 (N_3201,In_2321,In_401);
nand U3202 (N_3202,In_1882,In_1714);
and U3203 (N_3203,In_2187,In_443);
or U3204 (N_3204,In_1885,In_628);
or U3205 (N_3205,In_2498,In_535);
xor U3206 (N_3206,In_2350,In_728);
nand U3207 (N_3207,In_1390,In_2215);
and U3208 (N_3208,In_375,In_1278);
xor U3209 (N_3209,In_1772,In_662);
nand U3210 (N_3210,In_1371,In_1261);
or U3211 (N_3211,In_1973,In_1827);
nand U3212 (N_3212,In_72,In_1852);
nor U3213 (N_3213,In_548,In_2172);
or U3214 (N_3214,In_1948,In_2282);
xnor U3215 (N_3215,In_1924,In_1372);
nand U3216 (N_3216,In_809,In_653);
or U3217 (N_3217,In_105,In_2076);
nor U3218 (N_3218,In_1196,In_1383);
nand U3219 (N_3219,In_1483,In_1609);
and U3220 (N_3220,In_2405,In_1470);
xor U3221 (N_3221,In_1881,In_2151);
nand U3222 (N_3222,In_284,In_2114);
nor U3223 (N_3223,In_1365,In_1659);
and U3224 (N_3224,In_2315,In_216);
nand U3225 (N_3225,In_2132,In_1363);
and U3226 (N_3226,In_904,In_2201);
nand U3227 (N_3227,In_142,In_1943);
nor U3228 (N_3228,In_776,In_1860);
and U3229 (N_3229,In_1048,In_1946);
nor U3230 (N_3230,In_487,In_733);
nand U3231 (N_3231,In_792,In_2167);
xnor U3232 (N_3232,In_1572,In_2437);
xor U3233 (N_3233,In_1376,In_1015);
and U3234 (N_3234,In_1677,In_326);
or U3235 (N_3235,In_1294,In_743);
nor U3236 (N_3236,In_1417,In_32);
or U3237 (N_3237,In_2354,In_2322);
and U3238 (N_3238,In_1621,In_2176);
and U3239 (N_3239,In_1377,In_1995);
nand U3240 (N_3240,In_653,In_2282);
and U3241 (N_3241,In_34,In_1942);
nand U3242 (N_3242,In_1316,In_1842);
xnor U3243 (N_3243,In_1722,In_1579);
nand U3244 (N_3244,In_1648,In_86);
xor U3245 (N_3245,In_63,In_659);
xor U3246 (N_3246,In_2149,In_819);
and U3247 (N_3247,In_834,In_886);
nor U3248 (N_3248,In_2355,In_2378);
nor U3249 (N_3249,In_120,In_1295);
nor U3250 (N_3250,In_519,In_2128);
xnor U3251 (N_3251,In_1718,In_729);
nand U3252 (N_3252,In_1860,In_1845);
nor U3253 (N_3253,In_244,In_46);
or U3254 (N_3254,In_586,In_1493);
xor U3255 (N_3255,In_193,In_1811);
nor U3256 (N_3256,In_611,In_2312);
or U3257 (N_3257,In_1140,In_1300);
nand U3258 (N_3258,In_895,In_2257);
and U3259 (N_3259,In_4,In_592);
and U3260 (N_3260,In_1573,In_2319);
xnor U3261 (N_3261,In_339,In_404);
nor U3262 (N_3262,In_1202,In_913);
xor U3263 (N_3263,In_1567,In_1661);
or U3264 (N_3264,In_522,In_0);
or U3265 (N_3265,In_1213,In_1292);
or U3266 (N_3266,In_1946,In_999);
and U3267 (N_3267,In_2440,In_2407);
and U3268 (N_3268,In_948,In_1941);
xnor U3269 (N_3269,In_1569,In_423);
nor U3270 (N_3270,In_2272,In_1318);
or U3271 (N_3271,In_980,In_38);
or U3272 (N_3272,In_1506,In_1395);
xor U3273 (N_3273,In_534,In_2203);
nand U3274 (N_3274,In_786,In_736);
or U3275 (N_3275,In_1636,In_2387);
or U3276 (N_3276,In_498,In_360);
nand U3277 (N_3277,In_2142,In_1684);
nor U3278 (N_3278,In_453,In_1619);
and U3279 (N_3279,In_442,In_1561);
and U3280 (N_3280,In_1038,In_1218);
nand U3281 (N_3281,In_1306,In_1421);
nand U3282 (N_3282,In_1103,In_1084);
xor U3283 (N_3283,In_98,In_969);
nand U3284 (N_3284,In_1531,In_2475);
nor U3285 (N_3285,In_1156,In_1386);
xor U3286 (N_3286,In_748,In_1493);
nand U3287 (N_3287,In_1643,In_2111);
or U3288 (N_3288,In_2061,In_35);
and U3289 (N_3289,In_1158,In_2465);
nor U3290 (N_3290,In_1060,In_597);
nor U3291 (N_3291,In_1480,In_969);
nand U3292 (N_3292,In_1302,In_2049);
or U3293 (N_3293,In_1439,In_2238);
xnor U3294 (N_3294,In_1455,In_1795);
or U3295 (N_3295,In_2418,In_1771);
nand U3296 (N_3296,In_1635,In_2308);
or U3297 (N_3297,In_1353,In_1578);
and U3298 (N_3298,In_557,In_520);
and U3299 (N_3299,In_277,In_366);
or U3300 (N_3300,In_1647,In_1053);
nand U3301 (N_3301,In_1918,In_2489);
or U3302 (N_3302,In_61,In_2195);
nor U3303 (N_3303,In_2232,In_258);
nor U3304 (N_3304,In_302,In_2351);
nor U3305 (N_3305,In_318,In_1094);
nand U3306 (N_3306,In_2378,In_1896);
and U3307 (N_3307,In_1473,In_1436);
nand U3308 (N_3308,In_322,In_134);
or U3309 (N_3309,In_1824,In_210);
and U3310 (N_3310,In_1382,In_2265);
nand U3311 (N_3311,In_2132,In_134);
nor U3312 (N_3312,In_247,In_1060);
and U3313 (N_3313,In_1010,In_1409);
nand U3314 (N_3314,In_1520,In_1127);
nand U3315 (N_3315,In_1349,In_806);
nor U3316 (N_3316,In_139,In_583);
and U3317 (N_3317,In_1664,In_1623);
and U3318 (N_3318,In_1204,In_1050);
or U3319 (N_3319,In_40,In_1453);
or U3320 (N_3320,In_1455,In_936);
nor U3321 (N_3321,In_1940,In_1094);
nor U3322 (N_3322,In_707,In_546);
or U3323 (N_3323,In_655,In_2326);
nor U3324 (N_3324,In_204,In_373);
and U3325 (N_3325,In_1042,In_201);
or U3326 (N_3326,In_413,In_88);
and U3327 (N_3327,In_647,In_2206);
or U3328 (N_3328,In_1361,In_340);
nor U3329 (N_3329,In_2013,In_1892);
and U3330 (N_3330,In_1625,In_76);
or U3331 (N_3331,In_1972,In_380);
and U3332 (N_3332,In_1577,In_1154);
xnor U3333 (N_3333,In_1220,In_1035);
or U3334 (N_3334,In_2340,In_1646);
nand U3335 (N_3335,In_344,In_953);
nand U3336 (N_3336,In_157,In_824);
and U3337 (N_3337,In_1425,In_557);
and U3338 (N_3338,In_867,In_451);
xnor U3339 (N_3339,In_1637,In_35);
and U3340 (N_3340,In_1001,In_2307);
xor U3341 (N_3341,In_2379,In_773);
or U3342 (N_3342,In_1516,In_361);
and U3343 (N_3343,In_1187,In_2185);
nand U3344 (N_3344,In_95,In_1019);
xor U3345 (N_3345,In_375,In_918);
and U3346 (N_3346,In_68,In_1728);
and U3347 (N_3347,In_1323,In_1434);
and U3348 (N_3348,In_939,In_1891);
and U3349 (N_3349,In_1516,In_286);
nand U3350 (N_3350,In_534,In_322);
xnor U3351 (N_3351,In_372,In_61);
xnor U3352 (N_3352,In_2477,In_1755);
xor U3353 (N_3353,In_591,In_1663);
xor U3354 (N_3354,In_1709,In_575);
xnor U3355 (N_3355,In_1808,In_1944);
or U3356 (N_3356,In_1793,In_2470);
nor U3357 (N_3357,In_1263,In_2023);
and U3358 (N_3358,In_2333,In_1042);
or U3359 (N_3359,In_1901,In_521);
and U3360 (N_3360,In_243,In_62);
and U3361 (N_3361,In_367,In_1347);
xor U3362 (N_3362,In_1003,In_1028);
or U3363 (N_3363,In_148,In_254);
or U3364 (N_3364,In_1292,In_1252);
or U3365 (N_3365,In_1210,In_2079);
xnor U3366 (N_3366,In_1676,In_1005);
and U3367 (N_3367,In_1943,In_2467);
xor U3368 (N_3368,In_2128,In_940);
xnor U3369 (N_3369,In_2121,In_370);
xnor U3370 (N_3370,In_901,In_1099);
nand U3371 (N_3371,In_1882,In_2140);
xnor U3372 (N_3372,In_780,In_1399);
nor U3373 (N_3373,In_990,In_1166);
xor U3374 (N_3374,In_2232,In_580);
and U3375 (N_3375,In_998,In_2470);
and U3376 (N_3376,In_1663,In_701);
nor U3377 (N_3377,In_1851,In_653);
nand U3378 (N_3378,In_1339,In_1844);
or U3379 (N_3379,In_1991,In_1779);
nor U3380 (N_3380,In_2388,In_287);
nand U3381 (N_3381,In_1069,In_2297);
nand U3382 (N_3382,In_305,In_69);
or U3383 (N_3383,In_1378,In_1883);
nand U3384 (N_3384,In_2353,In_440);
or U3385 (N_3385,In_542,In_894);
nor U3386 (N_3386,In_843,In_2183);
or U3387 (N_3387,In_471,In_14);
nor U3388 (N_3388,In_1335,In_1408);
nand U3389 (N_3389,In_2200,In_1188);
or U3390 (N_3390,In_2479,In_2295);
and U3391 (N_3391,In_1777,In_315);
and U3392 (N_3392,In_247,In_467);
nor U3393 (N_3393,In_2258,In_1634);
or U3394 (N_3394,In_1376,In_2475);
or U3395 (N_3395,In_1106,In_404);
or U3396 (N_3396,In_541,In_2229);
and U3397 (N_3397,In_2375,In_853);
nand U3398 (N_3398,In_2229,In_699);
nor U3399 (N_3399,In_1995,In_2475);
or U3400 (N_3400,In_146,In_2056);
nor U3401 (N_3401,In_1078,In_2015);
and U3402 (N_3402,In_2376,In_2131);
nand U3403 (N_3403,In_1363,In_950);
nand U3404 (N_3404,In_2456,In_1709);
and U3405 (N_3405,In_1559,In_1092);
nor U3406 (N_3406,In_2093,In_2156);
or U3407 (N_3407,In_1076,In_362);
nand U3408 (N_3408,In_1632,In_1609);
or U3409 (N_3409,In_965,In_2141);
or U3410 (N_3410,In_1313,In_1315);
nor U3411 (N_3411,In_2244,In_1567);
and U3412 (N_3412,In_556,In_2058);
nand U3413 (N_3413,In_716,In_725);
and U3414 (N_3414,In_974,In_1045);
xnor U3415 (N_3415,In_1827,In_203);
or U3416 (N_3416,In_863,In_1622);
or U3417 (N_3417,In_130,In_1095);
nor U3418 (N_3418,In_1016,In_2305);
or U3419 (N_3419,In_2251,In_2382);
nor U3420 (N_3420,In_1954,In_1114);
or U3421 (N_3421,In_13,In_1320);
nor U3422 (N_3422,In_1434,In_2403);
and U3423 (N_3423,In_967,In_893);
nand U3424 (N_3424,In_1261,In_248);
and U3425 (N_3425,In_2354,In_403);
nor U3426 (N_3426,In_234,In_1754);
xnor U3427 (N_3427,In_563,In_1531);
nand U3428 (N_3428,In_15,In_1685);
nand U3429 (N_3429,In_1507,In_1421);
or U3430 (N_3430,In_2340,In_2077);
or U3431 (N_3431,In_1384,In_2161);
nand U3432 (N_3432,In_2264,In_1809);
and U3433 (N_3433,In_1601,In_1605);
xor U3434 (N_3434,In_609,In_1503);
nor U3435 (N_3435,In_1244,In_2365);
xnor U3436 (N_3436,In_827,In_2432);
xor U3437 (N_3437,In_939,In_836);
nor U3438 (N_3438,In_1561,In_935);
nor U3439 (N_3439,In_443,In_186);
xor U3440 (N_3440,In_24,In_1412);
or U3441 (N_3441,In_994,In_1569);
or U3442 (N_3442,In_2036,In_1237);
or U3443 (N_3443,In_2457,In_1528);
nand U3444 (N_3444,In_1157,In_1751);
nand U3445 (N_3445,In_468,In_1305);
or U3446 (N_3446,In_839,In_640);
nor U3447 (N_3447,In_1743,In_2185);
or U3448 (N_3448,In_1289,In_1693);
nor U3449 (N_3449,In_2358,In_1091);
xnor U3450 (N_3450,In_694,In_1189);
xor U3451 (N_3451,In_2399,In_2236);
nor U3452 (N_3452,In_1219,In_2002);
nand U3453 (N_3453,In_72,In_408);
and U3454 (N_3454,In_74,In_1274);
or U3455 (N_3455,In_2466,In_1516);
xor U3456 (N_3456,In_1823,In_1125);
nand U3457 (N_3457,In_1953,In_1914);
nand U3458 (N_3458,In_1031,In_412);
nor U3459 (N_3459,In_1575,In_194);
or U3460 (N_3460,In_244,In_2322);
nor U3461 (N_3461,In_2395,In_501);
and U3462 (N_3462,In_2301,In_1956);
or U3463 (N_3463,In_688,In_2165);
nor U3464 (N_3464,In_870,In_595);
nand U3465 (N_3465,In_812,In_244);
nand U3466 (N_3466,In_1977,In_1752);
or U3467 (N_3467,In_676,In_995);
and U3468 (N_3468,In_1267,In_1070);
and U3469 (N_3469,In_945,In_491);
xor U3470 (N_3470,In_962,In_420);
and U3471 (N_3471,In_1265,In_1586);
nor U3472 (N_3472,In_1447,In_1934);
or U3473 (N_3473,In_2315,In_1276);
nand U3474 (N_3474,In_2109,In_1945);
nand U3475 (N_3475,In_530,In_1990);
or U3476 (N_3476,In_1312,In_1146);
nor U3477 (N_3477,In_1177,In_2224);
nor U3478 (N_3478,In_1172,In_1921);
nand U3479 (N_3479,In_873,In_1664);
nor U3480 (N_3480,In_137,In_2228);
nor U3481 (N_3481,In_226,In_896);
nor U3482 (N_3482,In_2077,In_314);
and U3483 (N_3483,In_187,In_653);
nand U3484 (N_3484,In_699,In_1508);
and U3485 (N_3485,In_440,In_2346);
nand U3486 (N_3486,In_2495,In_901);
nor U3487 (N_3487,In_1988,In_554);
nor U3488 (N_3488,In_2252,In_1888);
xnor U3489 (N_3489,In_775,In_208);
and U3490 (N_3490,In_2289,In_1980);
or U3491 (N_3491,In_1120,In_1653);
nand U3492 (N_3492,In_1287,In_411);
or U3493 (N_3493,In_1844,In_1322);
nor U3494 (N_3494,In_1545,In_2216);
nor U3495 (N_3495,In_1295,In_1931);
xnor U3496 (N_3496,In_153,In_1546);
nor U3497 (N_3497,In_23,In_2193);
or U3498 (N_3498,In_821,In_1853);
nand U3499 (N_3499,In_145,In_1454);
or U3500 (N_3500,In_523,In_2073);
or U3501 (N_3501,In_2050,In_1185);
nor U3502 (N_3502,In_1382,In_2361);
nor U3503 (N_3503,In_1617,In_1337);
or U3504 (N_3504,In_908,In_2281);
xnor U3505 (N_3505,In_758,In_1368);
xnor U3506 (N_3506,In_1356,In_2085);
nand U3507 (N_3507,In_1846,In_1105);
or U3508 (N_3508,In_2283,In_2493);
and U3509 (N_3509,In_903,In_1943);
nand U3510 (N_3510,In_1040,In_801);
xnor U3511 (N_3511,In_2242,In_1983);
and U3512 (N_3512,In_1843,In_523);
xor U3513 (N_3513,In_663,In_671);
xor U3514 (N_3514,In_1150,In_56);
or U3515 (N_3515,In_1560,In_1060);
nand U3516 (N_3516,In_123,In_802);
nor U3517 (N_3517,In_2148,In_1175);
nand U3518 (N_3518,In_2468,In_1351);
and U3519 (N_3519,In_1875,In_615);
nand U3520 (N_3520,In_922,In_1026);
nor U3521 (N_3521,In_525,In_2206);
nor U3522 (N_3522,In_2101,In_174);
or U3523 (N_3523,In_766,In_1000);
and U3524 (N_3524,In_1596,In_79);
or U3525 (N_3525,In_183,In_1156);
or U3526 (N_3526,In_253,In_1476);
nor U3527 (N_3527,In_882,In_1230);
nor U3528 (N_3528,In_1388,In_1079);
and U3529 (N_3529,In_294,In_2345);
and U3530 (N_3530,In_1001,In_382);
nand U3531 (N_3531,In_659,In_2069);
and U3532 (N_3532,In_869,In_2344);
xnor U3533 (N_3533,In_1409,In_77);
and U3534 (N_3534,In_80,In_2038);
nand U3535 (N_3535,In_136,In_644);
or U3536 (N_3536,In_530,In_2414);
and U3537 (N_3537,In_1657,In_290);
or U3538 (N_3538,In_519,In_482);
nor U3539 (N_3539,In_3,In_1740);
xor U3540 (N_3540,In_1671,In_1142);
and U3541 (N_3541,In_1434,In_87);
or U3542 (N_3542,In_1311,In_2194);
nand U3543 (N_3543,In_2242,In_1964);
or U3544 (N_3544,In_463,In_136);
or U3545 (N_3545,In_1470,In_686);
or U3546 (N_3546,In_1914,In_514);
nor U3547 (N_3547,In_1328,In_364);
xnor U3548 (N_3548,In_604,In_1317);
xnor U3549 (N_3549,In_950,In_262);
or U3550 (N_3550,In_779,In_685);
or U3551 (N_3551,In_871,In_2284);
nor U3552 (N_3552,In_625,In_2202);
nand U3553 (N_3553,In_2075,In_50);
or U3554 (N_3554,In_1570,In_107);
and U3555 (N_3555,In_1419,In_662);
xnor U3556 (N_3556,In_2343,In_1135);
nand U3557 (N_3557,In_2204,In_573);
or U3558 (N_3558,In_225,In_167);
and U3559 (N_3559,In_225,In_2378);
xnor U3560 (N_3560,In_584,In_319);
or U3561 (N_3561,In_2125,In_1052);
nand U3562 (N_3562,In_1013,In_1101);
nand U3563 (N_3563,In_2473,In_1366);
nand U3564 (N_3564,In_1181,In_1649);
nor U3565 (N_3565,In_1024,In_2037);
xor U3566 (N_3566,In_1970,In_2418);
xnor U3567 (N_3567,In_2235,In_1873);
nand U3568 (N_3568,In_1261,In_1962);
or U3569 (N_3569,In_809,In_16);
nand U3570 (N_3570,In_1888,In_1356);
or U3571 (N_3571,In_904,In_96);
xnor U3572 (N_3572,In_235,In_2407);
and U3573 (N_3573,In_2097,In_574);
xor U3574 (N_3574,In_368,In_1573);
or U3575 (N_3575,In_110,In_1848);
xor U3576 (N_3576,In_2442,In_513);
nand U3577 (N_3577,In_551,In_1492);
or U3578 (N_3578,In_87,In_676);
or U3579 (N_3579,In_1380,In_2357);
or U3580 (N_3580,In_2323,In_606);
nand U3581 (N_3581,In_720,In_781);
xor U3582 (N_3582,In_628,In_757);
and U3583 (N_3583,In_156,In_528);
nand U3584 (N_3584,In_263,In_261);
nor U3585 (N_3585,In_1256,In_1847);
nand U3586 (N_3586,In_1023,In_1209);
or U3587 (N_3587,In_2483,In_459);
xor U3588 (N_3588,In_842,In_2104);
xnor U3589 (N_3589,In_940,In_2288);
nor U3590 (N_3590,In_176,In_1776);
and U3591 (N_3591,In_841,In_410);
or U3592 (N_3592,In_1242,In_1565);
nor U3593 (N_3593,In_614,In_2091);
and U3594 (N_3594,In_1531,In_1545);
and U3595 (N_3595,In_2132,In_1853);
xnor U3596 (N_3596,In_1808,In_1794);
nor U3597 (N_3597,In_830,In_2381);
and U3598 (N_3598,In_413,In_2103);
and U3599 (N_3599,In_84,In_938);
xnor U3600 (N_3600,In_1887,In_494);
and U3601 (N_3601,In_936,In_1608);
nand U3602 (N_3602,In_2197,In_1590);
xor U3603 (N_3603,In_1862,In_2038);
and U3604 (N_3604,In_723,In_91);
xnor U3605 (N_3605,In_493,In_175);
or U3606 (N_3606,In_1797,In_743);
nor U3607 (N_3607,In_1771,In_930);
and U3608 (N_3608,In_2018,In_937);
xnor U3609 (N_3609,In_1614,In_2425);
xor U3610 (N_3610,In_1386,In_1634);
or U3611 (N_3611,In_1609,In_2214);
and U3612 (N_3612,In_2431,In_924);
nand U3613 (N_3613,In_1444,In_292);
nor U3614 (N_3614,In_700,In_1645);
xor U3615 (N_3615,In_1303,In_1942);
and U3616 (N_3616,In_534,In_1318);
nor U3617 (N_3617,In_2136,In_1586);
xor U3618 (N_3618,In_730,In_1750);
and U3619 (N_3619,In_1922,In_2081);
nor U3620 (N_3620,In_651,In_346);
xor U3621 (N_3621,In_1712,In_2114);
xnor U3622 (N_3622,In_1309,In_1943);
nand U3623 (N_3623,In_2061,In_889);
xor U3624 (N_3624,In_636,In_1525);
nor U3625 (N_3625,In_2241,In_634);
and U3626 (N_3626,In_100,In_1377);
or U3627 (N_3627,In_1086,In_2494);
nor U3628 (N_3628,In_2060,In_561);
nand U3629 (N_3629,In_1135,In_1737);
nor U3630 (N_3630,In_1209,In_225);
xor U3631 (N_3631,In_92,In_1110);
nor U3632 (N_3632,In_18,In_223);
and U3633 (N_3633,In_1129,In_1368);
and U3634 (N_3634,In_2219,In_291);
nand U3635 (N_3635,In_288,In_415);
nand U3636 (N_3636,In_1931,In_1511);
nand U3637 (N_3637,In_1625,In_137);
xor U3638 (N_3638,In_2455,In_1593);
nor U3639 (N_3639,In_1593,In_111);
xor U3640 (N_3640,In_884,In_657);
or U3641 (N_3641,In_1520,In_2276);
xnor U3642 (N_3642,In_514,In_629);
nand U3643 (N_3643,In_1709,In_2146);
and U3644 (N_3644,In_2076,In_1963);
nand U3645 (N_3645,In_1084,In_1080);
or U3646 (N_3646,In_2358,In_1736);
nor U3647 (N_3647,In_2196,In_1427);
nand U3648 (N_3648,In_1562,In_2123);
or U3649 (N_3649,In_264,In_2210);
nor U3650 (N_3650,In_674,In_1851);
nand U3651 (N_3651,In_1180,In_73);
and U3652 (N_3652,In_2184,In_579);
and U3653 (N_3653,In_1143,In_1561);
or U3654 (N_3654,In_1653,In_2497);
xor U3655 (N_3655,In_290,In_918);
nand U3656 (N_3656,In_1971,In_816);
nor U3657 (N_3657,In_467,In_1822);
or U3658 (N_3658,In_732,In_2377);
nand U3659 (N_3659,In_2408,In_875);
nor U3660 (N_3660,In_2445,In_223);
xnor U3661 (N_3661,In_1231,In_185);
xor U3662 (N_3662,In_826,In_914);
or U3663 (N_3663,In_711,In_1299);
nor U3664 (N_3664,In_52,In_1667);
nand U3665 (N_3665,In_764,In_2234);
nand U3666 (N_3666,In_1297,In_1850);
nor U3667 (N_3667,In_1749,In_604);
and U3668 (N_3668,In_876,In_1970);
or U3669 (N_3669,In_2139,In_1986);
nand U3670 (N_3670,In_44,In_1464);
or U3671 (N_3671,In_1921,In_836);
nor U3672 (N_3672,In_184,In_238);
nor U3673 (N_3673,In_1167,In_644);
nor U3674 (N_3674,In_1166,In_790);
and U3675 (N_3675,In_582,In_2330);
nand U3676 (N_3676,In_1855,In_80);
nand U3677 (N_3677,In_410,In_1413);
nor U3678 (N_3678,In_524,In_33);
and U3679 (N_3679,In_811,In_1552);
nand U3680 (N_3680,In_2201,In_1764);
and U3681 (N_3681,In_1229,In_952);
xnor U3682 (N_3682,In_2382,In_2106);
nor U3683 (N_3683,In_1566,In_820);
xor U3684 (N_3684,In_1756,In_927);
xor U3685 (N_3685,In_2256,In_1549);
or U3686 (N_3686,In_1637,In_1663);
xnor U3687 (N_3687,In_1864,In_1154);
nor U3688 (N_3688,In_917,In_2469);
and U3689 (N_3689,In_2123,In_2470);
xor U3690 (N_3690,In_696,In_1943);
xnor U3691 (N_3691,In_1241,In_629);
nand U3692 (N_3692,In_10,In_1506);
and U3693 (N_3693,In_384,In_2005);
nor U3694 (N_3694,In_684,In_536);
nor U3695 (N_3695,In_704,In_1602);
and U3696 (N_3696,In_2367,In_866);
nor U3697 (N_3697,In_454,In_1902);
xor U3698 (N_3698,In_383,In_2355);
xnor U3699 (N_3699,In_2210,In_1528);
and U3700 (N_3700,In_588,In_2069);
xnor U3701 (N_3701,In_811,In_1827);
nor U3702 (N_3702,In_190,In_1513);
or U3703 (N_3703,In_1927,In_1692);
or U3704 (N_3704,In_929,In_1700);
and U3705 (N_3705,In_254,In_931);
xor U3706 (N_3706,In_1240,In_2282);
nand U3707 (N_3707,In_637,In_2336);
xnor U3708 (N_3708,In_1784,In_753);
nand U3709 (N_3709,In_2180,In_1393);
nand U3710 (N_3710,In_1771,In_1684);
or U3711 (N_3711,In_304,In_1896);
nand U3712 (N_3712,In_1637,In_157);
or U3713 (N_3713,In_419,In_1456);
or U3714 (N_3714,In_260,In_505);
nor U3715 (N_3715,In_275,In_1802);
nor U3716 (N_3716,In_129,In_2214);
nor U3717 (N_3717,In_554,In_2213);
and U3718 (N_3718,In_1230,In_2105);
nand U3719 (N_3719,In_60,In_2153);
nand U3720 (N_3720,In_186,In_1455);
xor U3721 (N_3721,In_155,In_759);
nand U3722 (N_3722,In_293,In_1263);
nor U3723 (N_3723,In_2065,In_1690);
xor U3724 (N_3724,In_1178,In_2038);
and U3725 (N_3725,In_1533,In_797);
or U3726 (N_3726,In_1054,In_1644);
and U3727 (N_3727,In_1082,In_70);
and U3728 (N_3728,In_2193,In_1881);
or U3729 (N_3729,In_1071,In_2261);
or U3730 (N_3730,In_1881,In_2246);
nand U3731 (N_3731,In_629,In_735);
and U3732 (N_3732,In_957,In_36);
and U3733 (N_3733,In_290,In_248);
and U3734 (N_3734,In_1904,In_1849);
nand U3735 (N_3735,In_1839,In_744);
xnor U3736 (N_3736,In_364,In_2255);
nor U3737 (N_3737,In_1650,In_2295);
and U3738 (N_3738,In_1148,In_2421);
nor U3739 (N_3739,In_1323,In_841);
or U3740 (N_3740,In_54,In_1911);
nor U3741 (N_3741,In_2435,In_1283);
or U3742 (N_3742,In_2174,In_939);
or U3743 (N_3743,In_1686,In_1097);
xor U3744 (N_3744,In_485,In_1364);
and U3745 (N_3745,In_420,In_2201);
xnor U3746 (N_3746,In_1042,In_442);
xor U3747 (N_3747,In_1589,In_1127);
and U3748 (N_3748,In_122,In_161);
nand U3749 (N_3749,In_1865,In_2118);
or U3750 (N_3750,In_196,In_604);
nor U3751 (N_3751,In_1181,In_1503);
or U3752 (N_3752,In_1073,In_116);
nor U3753 (N_3753,In_1107,In_117);
nor U3754 (N_3754,In_138,In_1153);
or U3755 (N_3755,In_1893,In_2045);
xor U3756 (N_3756,In_1967,In_253);
or U3757 (N_3757,In_1003,In_1317);
nand U3758 (N_3758,In_1797,In_2169);
nor U3759 (N_3759,In_2381,In_1951);
nand U3760 (N_3760,In_1734,In_2377);
and U3761 (N_3761,In_893,In_776);
and U3762 (N_3762,In_2248,In_1468);
nor U3763 (N_3763,In_2199,In_827);
nand U3764 (N_3764,In_1912,In_1654);
and U3765 (N_3765,In_847,In_2446);
nand U3766 (N_3766,In_196,In_194);
xor U3767 (N_3767,In_562,In_1363);
nor U3768 (N_3768,In_1594,In_1121);
or U3769 (N_3769,In_625,In_1585);
or U3770 (N_3770,In_1670,In_2);
and U3771 (N_3771,In_1791,In_1283);
nor U3772 (N_3772,In_1240,In_2133);
nor U3773 (N_3773,In_2315,In_319);
nor U3774 (N_3774,In_2269,In_851);
nand U3775 (N_3775,In_852,In_935);
nand U3776 (N_3776,In_1534,In_2420);
nor U3777 (N_3777,In_254,In_1133);
nand U3778 (N_3778,In_422,In_1361);
xor U3779 (N_3779,In_1494,In_1999);
or U3780 (N_3780,In_628,In_2349);
and U3781 (N_3781,In_1821,In_2147);
or U3782 (N_3782,In_1972,In_386);
nor U3783 (N_3783,In_1987,In_886);
nand U3784 (N_3784,In_608,In_1869);
and U3785 (N_3785,In_41,In_628);
or U3786 (N_3786,In_589,In_1750);
or U3787 (N_3787,In_28,In_1566);
nand U3788 (N_3788,In_1217,In_1954);
nand U3789 (N_3789,In_869,In_1006);
nand U3790 (N_3790,In_579,In_712);
nand U3791 (N_3791,In_1721,In_711);
or U3792 (N_3792,In_1029,In_1355);
xnor U3793 (N_3793,In_2054,In_2045);
nor U3794 (N_3794,In_1595,In_22);
nand U3795 (N_3795,In_1888,In_2300);
xnor U3796 (N_3796,In_718,In_11);
or U3797 (N_3797,In_1197,In_1595);
xnor U3798 (N_3798,In_809,In_1118);
nor U3799 (N_3799,In_2331,In_272);
nand U3800 (N_3800,In_955,In_766);
xor U3801 (N_3801,In_2007,In_2461);
xnor U3802 (N_3802,In_1836,In_2100);
nand U3803 (N_3803,In_1735,In_673);
and U3804 (N_3804,In_1556,In_360);
nor U3805 (N_3805,In_46,In_345);
or U3806 (N_3806,In_412,In_582);
and U3807 (N_3807,In_50,In_498);
nor U3808 (N_3808,In_1516,In_2369);
or U3809 (N_3809,In_690,In_1220);
xor U3810 (N_3810,In_2035,In_1936);
and U3811 (N_3811,In_780,In_1672);
and U3812 (N_3812,In_1628,In_1088);
and U3813 (N_3813,In_2170,In_1419);
or U3814 (N_3814,In_1574,In_1979);
nand U3815 (N_3815,In_1446,In_2412);
nor U3816 (N_3816,In_1247,In_1345);
nand U3817 (N_3817,In_913,In_1843);
nor U3818 (N_3818,In_1376,In_1681);
nor U3819 (N_3819,In_237,In_1208);
nand U3820 (N_3820,In_743,In_838);
nand U3821 (N_3821,In_22,In_999);
xor U3822 (N_3822,In_2080,In_1250);
xnor U3823 (N_3823,In_2085,In_1667);
xor U3824 (N_3824,In_647,In_843);
nand U3825 (N_3825,In_844,In_1450);
and U3826 (N_3826,In_2416,In_1088);
and U3827 (N_3827,In_106,In_1021);
or U3828 (N_3828,In_1975,In_2060);
nand U3829 (N_3829,In_424,In_1344);
nand U3830 (N_3830,In_2082,In_1161);
xor U3831 (N_3831,In_139,In_1382);
or U3832 (N_3832,In_310,In_1553);
and U3833 (N_3833,In_1048,In_673);
nor U3834 (N_3834,In_1167,In_1764);
or U3835 (N_3835,In_2129,In_553);
nor U3836 (N_3836,In_1013,In_1823);
or U3837 (N_3837,In_368,In_1233);
or U3838 (N_3838,In_430,In_350);
nand U3839 (N_3839,In_1293,In_1220);
and U3840 (N_3840,In_1151,In_1984);
nor U3841 (N_3841,In_2069,In_747);
and U3842 (N_3842,In_168,In_1052);
or U3843 (N_3843,In_1822,In_1596);
and U3844 (N_3844,In_2418,In_1888);
nor U3845 (N_3845,In_1786,In_1066);
and U3846 (N_3846,In_1417,In_85);
and U3847 (N_3847,In_1933,In_1997);
nor U3848 (N_3848,In_505,In_278);
xnor U3849 (N_3849,In_2080,In_1073);
or U3850 (N_3850,In_1019,In_1385);
nor U3851 (N_3851,In_701,In_2184);
and U3852 (N_3852,In_10,In_1077);
or U3853 (N_3853,In_2354,In_1965);
or U3854 (N_3854,In_2407,In_445);
and U3855 (N_3855,In_793,In_398);
or U3856 (N_3856,In_2158,In_1629);
and U3857 (N_3857,In_2462,In_1723);
and U3858 (N_3858,In_2277,In_2272);
nor U3859 (N_3859,In_322,In_1889);
or U3860 (N_3860,In_483,In_1033);
or U3861 (N_3861,In_1917,In_1508);
nor U3862 (N_3862,In_411,In_1153);
nand U3863 (N_3863,In_1166,In_522);
or U3864 (N_3864,In_758,In_333);
nand U3865 (N_3865,In_1251,In_189);
xor U3866 (N_3866,In_632,In_1511);
and U3867 (N_3867,In_914,In_1756);
or U3868 (N_3868,In_2033,In_735);
and U3869 (N_3869,In_441,In_1681);
or U3870 (N_3870,In_658,In_1489);
nor U3871 (N_3871,In_1931,In_1465);
xnor U3872 (N_3872,In_1361,In_1805);
and U3873 (N_3873,In_1147,In_1409);
xor U3874 (N_3874,In_458,In_645);
xor U3875 (N_3875,In_2211,In_1978);
xor U3876 (N_3876,In_2068,In_292);
or U3877 (N_3877,In_1641,In_756);
or U3878 (N_3878,In_202,In_1947);
or U3879 (N_3879,In_79,In_1168);
xnor U3880 (N_3880,In_1203,In_2350);
xor U3881 (N_3881,In_2267,In_53);
or U3882 (N_3882,In_882,In_2285);
or U3883 (N_3883,In_2352,In_2164);
nor U3884 (N_3884,In_1184,In_1924);
nand U3885 (N_3885,In_2439,In_1946);
and U3886 (N_3886,In_39,In_1603);
xor U3887 (N_3887,In_465,In_2351);
and U3888 (N_3888,In_1499,In_1168);
nor U3889 (N_3889,In_1900,In_798);
or U3890 (N_3890,In_1798,In_862);
nor U3891 (N_3891,In_203,In_1163);
nor U3892 (N_3892,In_1793,In_1887);
xor U3893 (N_3893,In_2361,In_1910);
and U3894 (N_3894,In_261,In_1897);
or U3895 (N_3895,In_1044,In_771);
xnor U3896 (N_3896,In_1193,In_896);
or U3897 (N_3897,In_2119,In_1243);
xor U3898 (N_3898,In_616,In_724);
and U3899 (N_3899,In_1591,In_2022);
xor U3900 (N_3900,In_2275,In_1708);
xor U3901 (N_3901,In_1861,In_2473);
nand U3902 (N_3902,In_2447,In_486);
or U3903 (N_3903,In_1538,In_92);
nor U3904 (N_3904,In_2450,In_1215);
xnor U3905 (N_3905,In_1018,In_2138);
nand U3906 (N_3906,In_79,In_2310);
nand U3907 (N_3907,In_393,In_308);
nand U3908 (N_3908,In_1642,In_1462);
xnor U3909 (N_3909,In_2023,In_2298);
or U3910 (N_3910,In_1988,In_1161);
nor U3911 (N_3911,In_662,In_325);
xor U3912 (N_3912,In_2037,In_39);
nand U3913 (N_3913,In_115,In_451);
xnor U3914 (N_3914,In_2045,In_1364);
and U3915 (N_3915,In_1036,In_794);
or U3916 (N_3916,In_926,In_1573);
nand U3917 (N_3917,In_753,In_1348);
nand U3918 (N_3918,In_1164,In_1035);
and U3919 (N_3919,In_2357,In_882);
or U3920 (N_3920,In_1474,In_2045);
nor U3921 (N_3921,In_1404,In_1180);
xor U3922 (N_3922,In_2184,In_554);
xor U3923 (N_3923,In_1357,In_2375);
or U3924 (N_3924,In_2277,In_677);
or U3925 (N_3925,In_206,In_808);
and U3926 (N_3926,In_2479,In_2197);
nor U3927 (N_3927,In_2309,In_843);
and U3928 (N_3928,In_1059,In_53);
and U3929 (N_3929,In_1451,In_1703);
and U3930 (N_3930,In_1208,In_377);
xor U3931 (N_3931,In_372,In_916);
or U3932 (N_3932,In_1747,In_1280);
and U3933 (N_3933,In_1716,In_742);
xor U3934 (N_3934,In_421,In_788);
nor U3935 (N_3935,In_1265,In_118);
nand U3936 (N_3936,In_479,In_2202);
and U3937 (N_3937,In_1279,In_262);
nand U3938 (N_3938,In_1498,In_2009);
and U3939 (N_3939,In_1075,In_1906);
nor U3940 (N_3940,In_898,In_1022);
nor U3941 (N_3941,In_1128,In_1271);
nand U3942 (N_3942,In_1228,In_1137);
and U3943 (N_3943,In_841,In_1810);
nand U3944 (N_3944,In_2442,In_1821);
nand U3945 (N_3945,In_689,In_342);
xnor U3946 (N_3946,In_194,In_85);
nand U3947 (N_3947,In_978,In_34);
or U3948 (N_3948,In_2247,In_1484);
xor U3949 (N_3949,In_1809,In_2297);
or U3950 (N_3950,In_707,In_2025);
or U3951 (N_3951,In_138,In_1516);
nor U3952 (N_3952,In_2310,In_168);
or U3953 (N_3953,In_294,In_904);
and U3954 (N_3954,In_2359,In_1776);
or U3955 (N_3955,In_2447,In_1038);
and U3956 (N_3956,In_534,In_1496);
xnor U3957 (N_3957,In_2209,In_861);
nor U3958 (N_3958,In_241,In_1346);
or U3959 (N_3959,In_1705,In_1173);
and U3960 (N_3960,In_2457,In_1287);
xor U3961 (N_3961,In_2311,In_1555);
and U3962 (N_3962,In_1080,In_1565);
xor U3963 (N_3963,In_1911,In_1063);
nand U3964 (N_3964,In_2374,In_1335);
xor U3965 (N_3965,In_762,In_347);
and U3966 (N_3966,In_575,In_617);
and U3967 (N_3967,In_516,In_2311);
xor U3968 (N_3968,In_1431,In_1250);
xor U3969 (N_3969,In_458,In_1277);
and U3970 (N_3970,In_2392,In_1585);
and U3971 (N_3971,In_987,In_205);
nor U3972 (N_3972,In_413,In_1633);
nor U3973 (N_3973,In_1385,In_792);
or U3974 (N_3974,In_2138,In_1931);
nand U3975 (N_3975,In_2146,In_1391);
nand U3976 (N_3976,In_2252,In_794);
nor U3977 (N_3977,In_1498,In_1331);
nor U3978 (N_3978,In_1718,In_1349);
or U3979 (N_3979,In_470,In_531);
nand U3980 (N_3980,In_1976,In_1673);
nand U3981 (N_3981,In_598,In_329);
xnor U3982 (N_3982,In_585,In_1213);
xor U3983 (N_3983,In_988,In_1108);
and U3984 (N_3984,In_255,In_620);
and U3985 (N_3985,In_1497,In_1743);
nor U3986 (N_3986,In_1207,In_1958);
nand U3987 (N_3987,In_1555,In_629);
or U3988 (N_3988,In_18,In_629);
and U3989 (N_3989,In_817,In_743);
nor U3990 (N_3990,In_498,In_1138);
xor U3991 (N_3991,In_715,In_819);
or U3992 (N_3992,In_329,In_1749);
xnor U3993 (N_3993,In_573,In_269);
or U3994 (N_3994,In_1329,In_1331);
or U3995 (N_3995,In_1079,In_1802);
and U3996 (N_3996,In_705,In_1560);
nor U3997 (N_3997,In_1522,In_1680);
nor U3998 (N_3998,In_1656,In_2448);
xnor U3999 (N_3999,In_1789,In_494);
and U4000 (N_4000,In_1108,In_1582);
or U4001 (N_4001,In_2065,In_1509);
and U4002 (N_4002,In_793,In_2118);
and U4003 (N_4003,In_1228,In_1998);
or U4004 (N_4004,In_86,In_749);
nor U4005 (N_4005,In_163,In_1877);
or U4006 (N_4006,In_1724,In_1517);
and U4007 (N_4007,In_1096,In_383);
and U4008 (N_4008,In_2094,In_1921);
and U4009 (N_4009,In_784,In_1165);
or U4010 (N_4010,In_1486,In_738);
and U4011 (N_4011,In_2365,In_236);
nand U4012 (N_4012,In_1043,In_1065);
and U4013 (N_4013,In_1046,In_422);
or U4014 (N_4014,In_1609,In_657);
and U4015 (N_4015,In_857,In_1296);
nor U4016 (N_4016,In_752,In_630);
nand U4017 (N_4017,In_1596,In_1459);
xnor U4018 (N_4018,In_300,In_1293);
or U4019 (N_4019,In_374,In_676);
or U4020 (N_4020,In_1951,In_1623);
nand U4021 (N_4021,In_803,In_1760);
xnor U4022 (N_4022,In_899,In_1446);
nand U4023 (N_4023,In_1868,In_967);
nor U4024 (N_4024,In_126,In_1983);
xnor U4025 (N_4025,In_2079,In_2455);
xor U4026 (N_4026,In_459,In_898);
and U4027 (N_4027,In_2420,In_304);
or U4028 (N_4028,In_1261,In_1665);
or U4029 (N_4029,In_1383,In_1241);
nand U4030 (N_4030,In_1980,In_388);
nand U4031 (N_4031,In_1073,In_1394);
nor U4032 (N_4032,In_255,In_1539);
nor U4033 (N_4033,In_392,In_1645);
or U4034 (N_4034,In_1149,In_613);
or U4035 (N_4035,In_2413,In_1156);
nand U4036 (N_4036,In_73,In_2162);
or U4037 (N_4037,In_2234,In_1231);
and U4038 (N_4038,In_2069,In_966);
or U4039 (N_4039,In_1686,In_458);
or U4040 (N_4040,In_207,In_1412);
and U4041 (N_4041,In_176,In_924);
nand U4042 (N_4042,In_1114,In_2166);
xnor U4043 (N_4043,In_635,In_680);
xor U4044 (N_4044,In_1523,In_270);
or U4045 (N_4045,In_1231,In_1342);
xnor U4046 (N_4046,In_1703,In_610);
and U4047 (N_4047,In_1441,In_2470);
xor U4048 (N_4048,In_846,In_1331);
or U4049 (N_4049,In_939,In_1492);
nor U4050 (N_4050,In_1797,In_944);
nand U4051 (N_4051,In_33,In_872);
nand U4052 (N_4052,In_587,In_757);
and U4053 (N_4053,In_389,In_2454);
or U4054 (N_4054,In_1244,In_2290);
or U4055 (N_4055,In_1798,In_1482);
xnor U4056 (N_4056,In_745,In_2447);
xnor U4057 (N_4057,In_406,In_2357);
and U4058 (N_4058,In_107,In_2242);
and U4059 (N_4059,In_1745,In_937);
nor U4060 (N_4060,In_98,In_45);
nor U4061 (N_4061,In_161,In_2340);
and U4062 (N_4062,In_1884,In_1067);
or U4063 (N_4063,In_621,In_137);
or U4064 (N_4064,In_2331,In_90);
nor U4065 (N_4065,In_247,In_1360);
or U4066 (N_4066,In_579,In_312);
xnor U4067 (N_4067,In_307,In_1846);
and U4068 (N_4068,In_805,In_2465);
and U4069 (N_4069,In_1296,In_1963);
xnor U4070 (N_4070,In_1139,In_900);
xnor U4071 (N_4071,In_523,In_1981);
xor U4072 (N_4072,In_2105,In_928);
nand U4073 (N_4073,In_1696,In_1309);
nor U4074 (N_4074,In_41,In_805);
xnor U4075 (N_4075,In_631,In_1582);
nand U4076 (N_4076,In_2182,In_983);
and U4077 (N_4077,In_1233,In_2425);
xnor U4078 (N_4078,In_2254,In_1249);
nor U4079 (N_4079,In_1951,In_1256);
nor U4080 (N_4080,In_2059,In_2456);
xor U4081 (N_4081,In_2084,In_1111);
and U4082 (N_4082,In_254,In_59);
and U4083 (N_4083,In_332,In_1932);
nand U4084 (N_4084,In_1256,In_65);
or U4085 (N_4085,In_405,In_150);
and U4086 (N_4086,In_427,In_1259);
and U4087 (N_4087,In_358,In_746);
nand U4088 (N_4088,In_1354,In_1929);
xor U4089 (N_4089,In_366,In_757);
nor U4090 (N_4090,In_1700,In_457);
nand U4091 (N_4091,In_136,In_798);
nor U4092 (N_4092,In_1082,In_1925);
nand U4093 (N_4093,In_2207,In_1953);
xnor U4094 (N_4094,In_866,In_1611);
or U4095 (N_4095,In_2262,In_1321);
and U4096 (N_4096,In_432,In_124);
and U4097 (N_4097,In_1422,In_470);
nor U4098 (N_4098,In_680,In_2268);
xnor U4099 (N_4099,In_3,In_271);
and U4100 (N_4100,In_730,In_969);
nand U4101 (N_4101,In_1986,In_1608);
nor U4102 (N_4102,In_588,In_364);
nand U4103 (N_4103,In_1030,In_1959);
xor U4104 (N_4104,In_604,In_2118);
nor U4105 (N_4105,In_1676,In_1634);
and U4106 (N_4106,In_1983,In_1082);
or U4107 (N_4107,In_1756,In_1761);
and U4108 (N_4108,In_2389,In_254);
xnor U4109 (N_4109,In_1092,In_2358);
and U4110 (N_4110,In_2303,In_1590);
and U4111 (N_4111,In_1398,In_253);
nor U4112 (N_4112,In_789,In_1445);
or U4113 (N_4113,In_1300,In_1261);
and U4114 (N_4114,In_949,In_2366);
and U4115 (N_4115,In_1079,In_1949);
and U4116 (N_4116,In_433,In_1114);
and U4117 (N_4117,In_1627,In_1967);
and U4118 (N_4118,In_1258,In_388);
nand U4119 (N_4119,In_1204,In_390);
or U4120 (N_4120,In_1107,In_803);
nand U4121 (N_4121,In_80,In_300);
or U4122 (N_4122,In_1844,In_1489);
nor U4123 (N_4123,In_994,In_2481);
xnor U4124 (N_4124,In_1317,In_2327);
nand U4125 (N_4125,In_1707,In_1551);
nand U4126 (N_4126,In_80,In_1969);
or U4127 (N_4127,In_802,In_1483);
nor U4128 (N_4128,In_1711,In_2255);
nand U4129 (N_4129,In_880,In_2441);
and U4130 (N_4130,In_345,In_187);
or U4131 (N_4131,In_2217,In_55);
and U4132 (N_4132,In_1147,In_1325);
and U4133 (N_4133,In_439,In_2474);
nor U4134 (N_4134,In_2371,In_931);
nand U4135 (N_4135,In_365,In_1224);
nand U4136 (N_4136,In_1792,In_2149);
and U4137 (N_4137,In_729,In_2329);
nand U4138 (N_4138,In_1800,In_1964);
and U4139 (N_4139,In_439,In_1000);
and U4140 (N_4140,In_1508,In_853);
nor U4141 (N_4141,In_975,In_2417);
nor U4142 (N_4142,In_427,In_144);
nor U4143 (N_4143,In_907,In_711);
xor U4144 (N_4144,In_402,In_2108);
xor U4145 (N_4145,In_1081,In_981);
and U4146 (N_4146,In_247,In_1181);
nor U4147 (N_4147,In_1789,In_975);
and U4148 (N_4148,In_1915,In_1624);
and U4149 (N_4149,In_953,In_157);
nor U4150 (N_4150,In_1136,In_1740);
nor U4151 (N_4151,In_516,In_432);
or U4152 (N_4152,In_1730,In_900);
xnor U4153 (N_4153,In_1471,In_1511);
and U4154 (N_4154,In_1946,In_1796);
and U4155 (N_4155,In_1466,In_726);
nand U4156 (N_4156,In_2091,In_1103);
and U4157 (N_4157,In_1366,In_2162);
and U4158 (N_4158,In_1797,In_1920);
xnor U4159 (N_4159,In_1185,In_1200);
nor U4160 (N_4160,In_1515,In_1525);
nand U4161 (N_4161,In_969,In_2464);
and U4162 (N_4162,In_2408,In_1664);
or U4163 (N_4163,In_1159,In_495);
xnor U4164 (N_4164,In_1822,In_2471);
or U4165 (N_4165,In_2463,In_329);
and U4166 (N_4166,In_2098,In_624);
or U4167 (N_4167,In_1647,In_177);
and U4168 (N_4168,In_2046,In_72);
nor U4169 (N_4169,In_465,In_748);
or U4170 (N_4170,In_635,In_1302);
nand U4171 (N_4171,In_648,In_1058);
nor U4172 (N_4172,In_1578,In_1246);
and U4173 (N_4173,In_780,In_1719);
nand U4174 (N_4174,In_1121,In_1955);
xnor U4175 (N_4175,In_902,In_308);
or U4176 (N_4176,In_1518,In_1189);
xor U4177 (N_4177,In_1277,In_281);
nor U4178 (N_4178,In_1608,In_1266);
nand U4179 (N_4179,In_2341,In_642);
nor U4180 (N_4180,In_974,In_345);
nand U4181 (N_4181,In_2098,In_2341);
nand U4182 (N_4182,In_2002,In_431);
xor U4183 (N_4183,In_315,In_1874);
nand U4184 (N_4184,In_811,In_1825);
nor U4185 (N_4185,In_450,In_97);
nor U4186 (N_4186,In_2483,In_656);
and U4187 (N_4187,In_246,In_851);
nand U4188 (N_4188,In_1660,In_398);
xor U4189 (N_4189,In_957,In_1268);
and U4190 (N_4190,In_1556,In_1115);
nor U4191 (N_4191,In_1687,In_1294);
xor U4192 (N_4192,In_1746,In_2375);
nor U4193 (N_4193,In_554,In_1107);
nor U4194 (N_4194,In_74,In_1865);
or U4195 (N_4195,In_2266,In_2201);
nor U4196 (N_4196,In_806,In_2367);
nor U4197 (N_4197,In_1345,In_1672);
nor U4198 (N_4198,In_183,In_1337);
nor U4199 (N_4199,In_1229,In_1561);
and U4200 (N_4200,In_2370,In_2480);
and U4201 (N_4201,In_652,In_1625);
xor U4202 (N_4202,In_965,In_692);
xor U4203 (N_4203,In_1047,In_76);
nand U4204 (N_4204,In_2372,In_2478);
nand U4205 (N_4205,In_1994,In_111);
nand U4206 (N_4206,In_613,In_53);
nor U4207 (N_4207,In_2022,In_1935);
and U4208 (N_4208,In_1502,In_2341);
xor U4209 (N_4209,In_2010,In_2367);
and U4210 (N_4210,In_370,In_378);
xnor U4211 (N_4211,In_1456,In_1580);
nor U4212 (N_4212,In_1283,In_363);
xor U4213 (N_4213,In_1676,In_161);
xor U4214 (N_4214,In_865,In_137);
nand U4215 (N_4215,In_1854,In_1069);
or U4216 (N_4216,In_1141,In_181);
nand U4217 (N_4217,In_1808,In_1897);
nor U4218 (N_4218,In_2419,In_902);
nor U4219 (N_4219,In_1605,In_495);
nor U4220 (N_4220,In_1966,In_1128);
xor U4221 (N_4221,In_77,In_1379);
or U4222 (N_4222,In_1919,In_1778);
xor U4223 (N_4223,In_524,In_2396);
and U4224 (N_4224,In_1976,In_91);
nand U4225 (N_4225,In_2109,In_248);
or U4226 (N_4226,In_139,In_2461);
or U4227 (N_4227,In_2325,In_411);
nor U4228 (N_4228,In_1406,In_317);
xor U4229 (N_4229,In_430,In_420);
nor U4230 (N_4230,In_1086,In_979);
nand U4231 (N_4231,In_1037,In_15);
nor U4232 (N_4232,In_1650,In_526);
and U4233 (N_4233,In_1287,In_796);
nor U4234 (N_4234,In_836,In_2200);
and U4235 (N_4235,In_848,In_1575);
nor U4236 (N_4236,In_430,In_248);
and U4237 (N_4237,In_2483,In_2108);
or U4238 (N_4238,In_1536,In_714);
nand U4239 (N_4239,In_221,In_1591);
and U4240 (N_4240,In_547,In_2092);
and U4241 (N_4241,In_912,In_1008);
nor U4242 (N_4242,In_599,In_1936);
xor U4243 (N_4243,In_2377,In_146);
and U4244 (N_4244,In_2273,In_2470);
nor U4245 (N_4245,In_497,In_1510);
nand U4246 (N_4246,In_2218,In_256);
and U4247 (N_4247,In_864,In_367);
xnor U4248 (N_4248,In_342,In_321);
nand U4249 (N_4249,In_673,In_1676);
nand U4250 (N_4250,In_365,In_560);
and U4251 (N_4251,In_418,In_286);
or U4252 (N_4252,In_1826,In_2243);
or U4253 (N_4253,In_1730,In_2386);
nor U4254 (N_4254,In_2145,In_1003);
nor U4255 (N_4255,In_1714,In_1260);
nor U4256 (N_4256,In_608,In_791);
nor U4257 (N_4257,In_2021,In_1168);
nor U4258 (N_4258,In_449,In_677);
and U4259 (N_4259,In_890,In_274);
nor U4260 (N_4260,In_2445,In_1990);
nor U4261 (N_4261,In_875,In_1604);
or U4262 (N_4262,In_159,In_1987);
nand U4263 (N_4263,In_749,In_1328);
or U4264 (N_4264,In_1913,In_1990);
and U4265 (N_4265,In_2140,In_98);
xor U4266 (N_4266,In_455,In_974);
or U4267 (N_4267,In_1338,In_1982);
xnor U4268 (N_4268,In_202,In_1878);
or U4269 (N_4269,In_703,In_370);
xor U4270 (N_4270,In_2072,In_2355);
nor U4271 (N_4271,In_1898,In_228);
or U4272 (N_4272,In_2230,In_895);
xor U4273 (N_4273,In_1900,In_2109);
nand U4274 (N_4274,In_2150,In_1755);
or U4275 (N_4275,In_2045,In_386);
or U4276 (N_4276,In_1958,In_1084);
nand U4277 (N_4277,In_623,In_1801);
or U4278 (N_4278,In_1237,In_714);
or U4279 (N_4279,In_818,In_2370);
nor U4280 (N_4280,In_2221,In_2383);
or U4281 (N_4281,In_2208,In_786);
and U4282 (N_4282,In_1170,In_1838);
xnor U4283 (N_4283,In_679,In_495);
xor U4284 (N_4284,In_2485,In_1109);
nand U4285 (N_4285,In_2350,In_571);
xnor U4286 (N_4286,In_202,In_2262);
and U4287 (N_4287,In_1521,In_1265);
nor U4288 (N_4288,In_1224,In_2339);
or U4289 (N_4289,In_151,In_17);
nand U4290 (N_4290,In_1065,In_1538);
xnor U4291 (N_4291,In_767,In_1304);
xnor U4292 (N_4292,In_1221,In_508);
or U4293 (N_4293,In_1557,In_1834);
or U4294 (N_4294,In_1599,In_846);
or U4295 (N_4295,In_1133,In_74);
and U4296 (N_4296,In_371,In_535);
nor U4297 (N_4297,In_1544,In_976);
and U4298 (N_4298,In_1924,In_1212);
nand U4299 (N_4299,In_219,In_1577);
xnor U4300 (N_4300,In_2167,In_332);
and U4301 (N_4301,In_2430,In_456);
and U4302 (N_4302,In_1701,In_630);
nor U4303 (N_4303,In_2070,In_2482);
and U4304 (N_4304,In_309,In_2240);
nand U4305 (N_4305,In_2475,In_1658);
nand U4306 (N_4306,In_2295,In_812);
nand U4307 (N_4307,In_1100,In_843);
nor U4308 (N_4308,In_589,In_593);
and U4309 (N_4309,In_877,In_507);
nor U4310 (N_4310,In_131,In_693);
xnor U4311 (N_4311,In_296,In_2261);
or U4312 (N_4312,In_906,In_1792);
xnor U4313 (N_4313,In_1828,In_2014);
nor U4314 (N_4314,In_2360,In_2165);
nor U4315 (N_4315,In_1371,In_540);
nand U4316 (N_4316,In_1239,In_1066);
nand U4317 (N_4317,In_1994,In_2143);
nand U4318 (N_4318,In_963,In_431);
and U4319 (N_4319,In_2425,In_1733);
nand U4320 (N_4320,In_723,In_2079);
or U4321 (N_4321,In_1200,In_219);
nand U4322 (N_4322,In_633,In_995);
or U4323 (N_4323,In_1601,In_1839);
or U4324 (N_4324,In_2130,In_569);
and U4325 (N_4325,In_567,In_1684);
or U4326 (N_4326,In_164,In_1399);
xor U4327 (N_4327,In_1066,In_1646);
and U4328 (N_4328,In_1012,In_202);
and U4329 (N_4329,In_83,In_1480);
or U4330 (N_4330,In_1497,In_1371);
nand U4331 (N_4331,In_1903,In_514);
and U4332 (N_4332,In_1354,In_565);
and U4333 (N_4333,In_798,In_125);
or U4334 (N_4334,In_545,In_1970);
nor U4335 (N_4335,In_1214,In_1264);
nand U4336 (N_4336,In_1645,In_1194);
or U4337 (N_4337,In_1966,In_146);
nand U4338 (N_4338,In_2224,In_2252);
or U4339 (N_4339,In_2231,In_1323);
and U4340 (N_4340,In_1804,In_1505);
and U4341 (N_4341,In_1716,In_2047);
xor U4342 (N_4342,In_7,In_1474);
nand U4343 (N_4343,In_14,In_538);
and U4344 (N_4344,In_1208,In_1038);
xnor U4345 (N_4345,In_1096,In_635);
xnor U4346 (N_4346,In_806,In_1606);
nand U4347 (N_4347,In_1130,In_736);
nand U4348 (N_4348,In_1536,In_538);
nor U4349 (N_4349,In_1805,In_1015);
nand U4350 (N_4350,In_1211,In_791);
or U4351 (N_4351,In_1218,In_59);
xor U4352 (N_4352,In_1081,In_1493);
and U4353 (N_4353,In_1598,In_2246);
xor U4354 (N_4354,In_1320,In_1216);
or U4355 (N_4355,In_1933,In_2440);
xor U4356 (N_4356,In_1960,In_1012);
xor U4357 (N_4357,In_1769,In_2159);
nand U4358 (N_4358,In_1715,In_989);
or U4359 (N_4359,In_1556,In_1274);
and U4360 (N_4360,In_866,In_264);
xnor U4361 (N_4361,In_760,In_2396);
nor U4362 (N_4362,In_895,In_1669);
nor U4363 (N_4363,In_1993,In_705);
xor U4364 (N_4364,In_642,In_200);
nand U4365 (N_4365,In_2157,In_1467);
nor U4366 (N_4366,In_1259,In_1127);
or U4367 (N_4367,In_1735,In_904);
xor U4368 (N_4368,In_1977,In_465);
or U4369 (N_4369,In_1231,In_198);
nand U4370 (N_4370,In_2489,In_1334);
nand U4371 (N_4371,In_1724,In_486);
nand U4372 (N_4372,In_1550,In_122);
and U4373 (N_4373,In_1313,In_1375);
or U4374 (N_4374,In_263,In_1666);
and U4375 (N_4375,In_1813,In_408);
xnor U4376 (N_4376,In_2357,In_991);
nor U4377 (N_4377,In_1885,In_2223);
or U4378 (N_4378,In_2213,In_1179);
nor U4379 (N_4379,In_1898,In_2423);
nor U4380 (N_4380,In_329,In_1683);
nand U4381 (N_4381,In_741,In_356);
xnor U4382 (N_4382,In_918,In_1207);
xnor U4383 (N_4383,In_2295,In_295);
nand U4384 (N_4384,In_1549,In_541);
xor U4385 (N_4385,In_142,In_55);
xor U4386 (N_4386,In_949,In_1249);
and U4387 (N_4387,In_516,In_1462);
or U4388 (N_4388,In_1552,In_2043);
xnor U4389 (N_4389,In_616,In_227);
or U4390 (N_4390,In_2280,In_1248);
nor U4391 (N_4391,In_930,In_1761);
and U4392 (N_4392,In_1103,In_1382);
or U4393 (N_4393,In_689,In_2194);
nor U4394 (N_4394,In_74,In_2481);
nand U4395 (N_4395,In_2031,In_2446);
or U4396 (N_4396,In_7,In_713);
or U4397 (N_4397,In_819,In_1958);
xnor U4398 (N_4398,In_1070,In_2139);
xor U4399 (N_4399,In_138,In_1020);
nor U4400 (N_4400,In_472,In_2232);
xnor U4401 (N_4401,In_1437,In_2221);
nand U4402 (N_4402,In_1203,In_2102);
nand U4403 (N_4403,In_2246,In_462);
nor U4404 (N_4404,In_2290,In_1293);
nand U4405 (N_4405,In_431,In_2477);
nand U4406 (N_4406,In_1583,In_1217);
or U4407 (N_4407,In_704,In_762);
or U4408 (N_4408,In_2213,In_2400);
nand U4409 (N_4409,In_2199,In_1962);
nand U4410 (N_4410,In_2124,In_2441);
nand U4411 (N_4411,In_1224,In_519);
nand U4412 (N_4412,In_2332,In_2028);
and U4413 (N_4413,In_1683,In_1789);
and U4414 (N_4414,In_503,In_1708);
or U4415 (N_4415,In_2189,In_1039);
or U4416 (N_4416,In_518,In_596);
xnor U4417 (N_4417,In_2445,In_709);
nand U4418 (N_4418,In_1437,In_753);
or U4419 (N_4419,In_58,In_90);
xor U4420 (N_4420,In_257,In_2440);
or U4421 (N_4421,In_801,In_1452);
nor U4422 (N_4422,In_589,In_479);
nor U4423 (N_4423,In_607,In_413);
nand U4424 (N_4424,In_1386,In_1110);
xor U4425 (N_4425,In_1175,In_1817);
nor U4426 (N_4426,In_724,In_556);
and U4427 (N_4427,In_1949,In_1010);
nor U4428 (N_4428,In_2444,In_1629);
nor U4429 (N_4429,In_1946,In_1750);
and U4430 (N_4430,In_2417,In_717);
nor U4431 (N_4431,In_136,In_2162);
or U4432 (N_4432,In_374,In_1384);
nand U4433 (N_4433,In_1325,In_2316);
nor U4434 (N_4434,In_800,In_382);
or U4435 (N_4435,In_1998,In_2334);
or U4436 (N_4436,In_1798,In_2351);
nand U4437 (N_4437,In_1739,In_1569);
and U4438 (N_4438,In_303,In_591);
nand U4439 (N_4439,In_9,In_2044);
nand U4440 (N_4440,In_441,In_1358);
xnor U4441 (N_4441,In_2161,In_2127);
nor U4442 (N_4442,In_230,In_481);
and U4443 (N_4443,In_1329,In_1164);
or U4444 (N_4444,In_2085,In_355);
or U4445 (N_4445,In_2284,In_1989);
nor U4446 (N_4446,In_1622,In_1208);
nor U4447 (N_4447,In_785,In_1372);
nand U4448 (N_4448,In_893,In_2402);
xor U4449 (N_4449,In_1657,In_1962);
nor U4450 (N_4450,In_1028,In_228);
nand U4451 (N_4451,In_1629,In_52);
nor U4452 (N_4452,In_2256,In_773);
or U4453 (N_4453,In_234,In_1882);
or U4454 (N_4454,In_401,In_336);
nor U4455 (N_4455,In_1576,In_1464);
and U4456 (N_4456,In_121,In_885);
nor U4457 (N_4457,In_2179,In_190);
and U4458 (N_4458,In_96,In_2330);
nor U4459 (N_4459,In_1433,In_1813);
or U4460 (N_4460,In_327,In_598);
nand U4461 (N_4461,In_1258,In_1529);
nand U4462 (N_4462,In_1603,In_1551);
nand U4463 (N_4463,In_199,In_2112);
nand U4464 (N_4464,In_631,In_244);
xnor U4465 (N_4465,In_288,In_2351);
xnor U4466 (N_4466,In_1758,In_397);
xor U4467 (N_4467,In_730,In_1913);
nand U4468 (N_4468,In_648,In_1080);
and U4469 (N_4469,In_2257,In_1601);
and U4470 (N_4470,In_1631,In_1296);
xnor U4471 (N_4471,In_47,In_934);
or U4472 (N_4472,In_2233,In_1409);
and U4473 (N_4473,In_1877,In_554);
nand U4474 (N_4474,In_2054,In_2414);
nand U4475 (N_4475,In_1103,In_1013);
nor U4476 (N_4476,In_1573,In_2112);
nand U4477 (N_4477,In_883,In_2316);
nand U4478 (N_4478,In_2445,In_278);
xnor U4479 (N_4479,In_1931,In_508);
nand U4480 (N_4480,In_1188,In_2244);
xnor U4481 (N_4481,In_2029,In_2282);
nor U4482 (N_4482,In_385,In_1706);
and U4483 (N_4483,In_1521,In_547);
nand U4484 (N_4484,In_2282,In_394);
xor U4485 (N_4485,In_593,In_2130);
xnor U4486 (N_4486,In_673,In_300);
and U4487 (N_4487,In_2416,In_397);
and U4488 (N_4488,In_55,In_819);
nor U4489 (N_4489,In_1989,In_1606);
and U4490 (N_4490,In_120,In_2271);
nand U4491 (N_4491,In_315,In_2274);
or U4492 (N_4492,In_370,In_897);
xor U4493 (N_4493,In_17,In_1609);
and U4494 (N_4494,In_820,In_312);
or U4495 (N_4495,In_359,In_2399);
nor U4496 (N_4496,In_1878,In_926);
xor U4497 (N_4497,In_610,In_1193);
nor U4498 (N_4498,In_1053,In_446);
nand U4499 (N_4499,In_288,In_1067);
xor U4500 (N_4500,In_937,In_1435);
or U4501 (N_4501,In_77,In_2297);
nor U4502 (N_4502,In_697,In_546);
or U4503 (N_4503,In_2458,In_1358);
and U4504 (N_4504,In_646,In_1512);
nand U4505 (N_4505,In_2258,In_2380);
nand U4506 (N_4506,In_1394,In_668);
nand U4507 (N_4507,In_560,In_2230);
or U4508 (N_4508,In_2075,In_1139);
and U4509 (N_4509,In_1981,In_468);
and U4510 (N_4510,In_1362,In_2317);
xor U4511 (N_4511,In_1574,In_466);
or U4512 (N_4512,In_853,In_2247);
nand U4513 (N_4513,In_18,In_171);
and U4514 (N_4514,In_2449,In_1423);
nand U4515 (N_4515,In_1877,In_1182);
or U4516 (N_4516,In_1724,In_2270);
nor U4517 (N_4517,In_20,In_1070);
nor U4518 (N_4518,In_69,In_736);
nor U4519 (N_4519,In_59,In_1859);
nand U4520 (N_4520,In_1717,In_2236);
and U4521 (N_4521,In_811,In_1029);
nand U4522 (N_4522,In_498,In_567);
or U4523 (N_4523,In_208,In_1639);
or U4524 (N_4524,In_393,In_1577);
xnor U4525 (N_4525,In_67,In_2017);
or U4526 (N_4526,In_2437,In_2128);
or U4527 (N_4527,In_633,In_1718);
or U4528 (N_4528,In_2263,In_1020);
nor U4529 (N_4529,In_1881,In_1844);
or U4530 (N_4530,In_1031,In_1479);
nand U4531 (N_4531,In_1200,In_1148);
xnor U4532 (N_4532,In_96,In_2396);
or U4533 (N_4533,In_221,In_545);
or U4534 (N_4534,In_813,In_1887);
and U4535 (N_4535,In_1332,In_1924);
nand U4536 (N_4536,In_1582,In_643);
or U4537 (N_4537,In_2468,In_723);
nor U4538 (N_4538,In_2204,In_2068);
xor U4539 (N_4539,In_1692,In_2324);
or U4540 (N_4540,In_511,In_883);
nor U4541 (N_4541,In_1613,In_189);
and U4542 (N_4542,In_602,In_2224);
nand U4543 (N_4543,In_818,In_1266);
xnor U4544 (N_4544,In_1448,In_805);
nor U4545 (N_4545,In_300,In_1920);
xor U4546 (N_4546,In_1653,In_254);
nor U4547 (N_4547,In_1973,In_1026);
and U4548 (N_4548,In_1782,In_799);
or U4549 (N_4549,In_1648,In_1436);
nor U4550 (N_4550,In_219,In_1103);
nand U4551 (N_4551,In_1935,In_2327);
or U4552 (N_4552,In_1106,In_1608);
and U4553 (N_4553,In_1545,In_1312);
nor U4554 (N_4554,In_1073,In_1065);
or U4555 (N_4555,In_1835,In_1867);
xor U4556 (N_4556,In_1068,In_1275);
and U4557 (N_4557,In_1397,In_948);
or U4558 (N_4558,In_234,In_2340);
nor U4559 (N_4559,In_25,In_706);
or U4560 (N_4560,In_75,In_555);
xor U4561 (N_4561,In_2069,In_935);
nand U4562 (N_4562,In_1067,In_495);
and U4563 (N_4563,In_2486,In_1652);
or U4564 (N_4564,In_89,In_1059);
or U4565 (N_4565,In_2293,In_1501);
or U4566 (N_4566,In_1739,In_46);
nor U4567 (N_4567,In_612,In_522);
xnor U4568 (N_4568,In_1608,In_2321);
or U4569 (N_4569,In_1888,In_916);
xnor U4570 (N_4570,In_36,In_1087);
nor U4571 (N_4571,In_1304,In_1771);
nor U4572 (N_4572,In_1261,In_94);
nor U4573 (N_4573,In_1827,In_617);
or U4574 (N_4574,In_671,In_352);
and U4575 (N_4575,In_570,In_616);
nand U4576 (N_4576,In_1431,In_963);
or U4577 (N_4577,In_1970,In_962);
or U4578 (N_4578,In_910,In_1564);
xnor U4579 (N_4579,In_1216,In_647);
xnor U4580 (N_4580,In_1484,In_63);
nand U4581 (N_4581,In_1365,In_1841);
or U4582 (N_4582,In_2497,In_231);
nor U4583 (N_4583,In_225,In_1976);
and U4584 (N_4584,In_545,In_994);
xor U4585 (N_4585,In_1679,In_1714);
nor U4586 (N_4586,In_867,In_2404);
nor U4587 (N_4587,In_795,In_1248);
xor U4588 (N_4588,In_2360,In_510);
xnor U4589 (N_4589,In_333,In_605);
xor U4590 (N_4590,In_1624,In_902);
or U4591 (N_4591,In_2028,In_4);
nor U4592 (N_4592,In_651,In_928);
nor U4593 (N_4593,In_471,In_1448);
and U4594 (N_4594,In_888,In_235);
and U4595 (N_4595,In_1341,In_796);
or U4596 (N_4596,In_835,In_769);
nand U4597 (N_4597,In_91,In_963);
xor U4598 (N_4598,In_2109,In_1532);
or U4599 (N_4599,In_367,In_93);
nor U4600 (N_4600,In_1400,In_1837);
or U4601 (N_4601,In_623,In_196);
nand U4602 (N_4602,In_1631,In_2114);
xnor U4603 (N_4603,In_1987,In_847);
xor U4604 (N_4604,In_2276,In_1455);
nand U4605 (N_4605,In_1397,In_790);
xnor U4606 (N_4606,In_1514,In_620);
nand U4607 (N_4607,In_19,In_1775);
and U4608 (N_4608,In_1953,In_937);
nor U4609 (N_4609,In_1639,In_283);
nand U4610 (N_4610,In_1489,In_908);
nand U4611 (N_4611,In_1013,In_1248);
or U4612 (N_4612,In_1548,In_1230);
nand U4613 (N_4613,In_518,In_387);
nand U4614 (N_4614,In_1068,In_621);
and U4615 (N_4615,In_238,In_511);
nor U4616 (N_4616,In_1397,In_1743);
xor U4617 (N_4617,In_1360,In_1615);
nor U4618 (N_4618,In_2124,In_1797);
nand U4619 (N_4619,In_836,In_1481);
xnor U4620 (N_4620,In_206,In_707);
xor U4621 (N_4621,In_202,In_1672);
or U4622 (N_4622,In_1430,In_1087);
or U4623 (N_4623,In_358,In_980);
and U4624 (N_4624,In_1420,In_2392);
or U4625 (N_4625,In_165,In_145);
xnor U4626 (N_4626,In_2446,In_313);
or U4627 (N_4627,In_258,In_1047);
or U4628 (N_4628,In_1417,In_2006);
or U4629 (N_4629,In_2280,In_1566);
nand U4630 (N_4630,In_946,In_2231);
nand U4631 (N_4631,In_22,In_1760);
nand U4632 (N_4632,In_10,In_147);
nor U4633 (N_4633,In_2151,In_913);
and U4634 (N_4634,In_1245,In_2453);
xor U4635 (N_4635,In_1591,In_1504);
nand U4636 (N_4636,In_1621,In_1500);
and U4637 (N_4637,In_603,In_389);
nand U4638 (N_4638,In_2291,In_1586);
or U4639 (N_4639,In_1528,In_1962);
or U4640 (N_4640,In_1028,In_2341);
xnor U4641 (N_4641,In_1042,In_1641);
or U4642 (N_4642,In_388,In_2431);
xnor U4643 (N_4643,In_1809,In_1613);
and U4644 (N_4644,In_2295,In_191);
or U4645 (N_4645,In_715,In_1311);
and U4646 (N_4646,In_2218,In_2073);
or U4647 (N_4647,In_2415,In_1322);
nor U4648 (N_4648,In_1644,In_2293);
and U4649 (N_4649,In_734,In_329);
nand U4650 (N_4650,In_1791,In_1325);
or U4651 (N_4651,In_2037,In_1656);
and U4652 (N_4652,In_793,In_2241);
xor U4653 (N_4653,In_1414,In_162);
nor U4654 (N_4654,In_40,In_2415);
nor U4655 (N_4655,In_2467,In_552);
and U4656 (N_4656,In_1558,In_135);
and U4657 (N_4657,In_1645,In_1323);
or U4658 (N_4658,In_747,In_2024);
nor U4659 (N_4659,In_2287,In_1062);
and U4660 (N_4660,In_1550,In_1998);
xor U4661 (N_4661,In_263,In_718);
and U4662 (N_4662,In_355,In_254);
nor U4663 (N_4663,In_1359,In_750);
nor U4664 (N_4664,In_458,In_544);
or U4665 (N_4665,In_973,In_2372);
nor U4666 (N_4666,In_2499,In_679);
xnor U4667 (N_4667,In_2076,In_2389);
or U4668 (N_4668,In_945,In_326);
xor U4669 (N_4669,In_53,In_756);
xnor U4670 (N_4670,In_634,In_2379);
or U4671 (N_4671,In_1254,In_1015);
and U4672 (N_4672,In_355,In_224);
or U4673 (N_4673,In_1327,In_697);
nor U4674 (N_4674,In_681,In_1844);
or U4675 (N_4675,In_1648,In_1803);
nor U4676 (N_4676,In_2069,In_2400);
nor U4677 (N_4677,In_604,In_1875);
or U4678 (N_4678,In_1169,In_1342);
nor U4679 (N_4679,In_434,In_2197);
nand U4680 (N_4680,In_221,In_807);
nand U4681 (N_4681,In_2447,In_666);
nor U4682 (N_4682,In_585,In_322);
or U4683 (N_4683,In_2148,In_2496);
nand U4684 (N_4684,In_2349,In_2010);
nand U4685 (N_4685,In_807,In_634);
or U4686 (N_4686,In_774,In_1463);
nand U4687 (N_4687,In_2008,In_421);
or U4688 (N_4688,In_2423,In_1674);
or U4689 (N_4689,In_1653,In_2028);
nor U4690 (N_4690,In_2069,In_326);
nor U4691 (N_4691,In_1336,In_1225);
xor U4692 (N_4692,In_1637,In_416);
or U4693 (N_4693,In_751,In_839);
xnor U4694 (N_4694,In_1368,In_1542);
nand U4695 (N_4695,In_2018,In_697);
and U4696 (N_4696,In_818,In_1426);
nand U4697 (N_4697,In_844,In_1333);
and U4698 (N_4698,In_1840,In_1388);
or U4699 (N_4699,In_540,In_2427);
or U4700 (N_4700,In_1749,In_589);
and U4701 (N_4701,In_149,In_403);
nor U4702 (N_4702,In_1638,In_2448);
xor U4703 (N_4703,In_789,In_1460);
and U4704 (N_4704,In_1731,In_1295);
and U4705 (N_4705,In_722,In_1235);
or U4706 (N_4706,In_1529,In_2456);
xnor U4707 (N_4707,In_231,In_1671);
or U4708 (N_4708,In_80,In_2224);
nor U4709 (N_4709,In_2263,In_2366);
xnor U4710 (N_4710,In_2345,In_256);
xnor U4711 (N_4711,In_652,In_680);
xor U4712 (N_4712,In_1399,In_1682);
or U4713 (N_4713,In_106,In_1587);
nor U4714 (N_4714,In_972,In_515);
nand U4715 (N_4715,In_1855,In_933);
and U4716 (N_4716,In_499,In_1639);
nand U4717 (N_4717,In_1666,In_1183);
xor U4718 (N_4718,In_2008,In_1130);
or U4719 (N_4719,In_1202,In_2134);
nor U4720 (N_4720,In_472,In_1012);
nor U4721 (N_4721,In_1968,In_1663);
nand U4722 (N_4722,In_966,In_23);
nand U4723 (N_4723,In_1783,In_1092);
nand U4724 (N_4724,In_848,In_1245);
nand U4725 (N_4725,In_456,In_853);
nand U4726 (N_4726,In_2019,In_1928);
or U4727 (N_4727,In_728,In_167);
nor U4728 (N_4728,In_2141,In_1468);
or U4729 (N_4729,In_1412,In_706);
xnor U4730 (N_4730,In_511,In_2292);
and U4731 (N_4731,In_1571,In_984);
nor U4732 (N_4732,In_2112,In_1204);
nor U4733 (N_4733,In_2472,In_943);
nor U4734 (N_4734,In_946,In_677);
or U4735 (N_4735,In_2034,In_730);
nor U4736 (N_4736,In_473,In_221);
xor U4737 (N_4737,In_1843,In_1924);
nor U4738 (N_4738,In_1026,In_2349);
and U4739 (N_4739,In_250,In_2005);
nand U4740 (N_4740,In_1685,In_996);
nand U4741 (N_4741,In_1811,In_11);
or U4742 (N_4742,In_645,In_765);
nor U4743 (N_4743,In_1920,In_843);
and U4744 (N_4744,In_552,In_172);
and U4745 (N_4745,In_1070,In_2066);
nor U4746 (N_4746,In_1476,In_390);
nand U4747 (N_4747,In_1715,In_166);
nor U4748 (N_4748,In_1274,In_1292);
nand U4749 (N_4749,In_212,In_1821);
nor U4750 (N_4750,In_1797,In_2478);
and U4751 (N_4751,In_516,In_1492);
nor U4752 (N_4752,In_2485,In_1622);
and U4753 (N_4753,In_1762,In_147);
and U4754 (N_4754,In_1854,In_1965);
xnor U4755 (N_4755,In_1755,In_1951);
nor U4756 (N_4756,In_2163,In_1087);
xnor U4757 (N_4757,In_2003,In_1199);
xor U4758 (N_4758,In_1554,In_279);
and U4759 (N_4759,In_1247,In_126);
nand U4760 (N_4760,In_2426,In_1013);
nor U4761 (N_4761,In_1824,In_2422);
or U4762 (N_4762,In_1742,In_9);
or U4763 (N_4763,In_985,In_2401);
xnor U4764 (N_4764,In_1896,In_2101);
or U4765 (N_4765,In_1130,In_1156);
xor U4766 (N_4766,In_528,In_1457);
and U4767 (N_4767,In_142,In_387);
nor U4768 (N_4768,In_623,In_2416);
nand U4769 (N_4769,In_2232,In_1080);
and U4770 (N_4770,In_1507,In_2042);
nor U4771 (N_4771,In_975,In_1076);
xor U4772 (N_4772,In_426,In_2478);
nand U4773 (N_4773,In_461,In_609);
or U4774 (N_4774,In_746,In_2017);
nor U4775 (N_4775,In_606,In_562);
nor U4776 (N_4776,In_2464,In_1636);
or U4777 (N_4777,In_466,In_1781);
nor U4778 (N_4778,In_956,In_1643);
xnor U4779 (N_4779,In_1949,In_2156);
nor U4780 (N_4780,In_1923,In_497);
nand U4781 (N_4781,In_982,In_2253);
xnor U4782 (N_4782,In_2433,In_322);
or U4783 (N_4783,In_1834,In_1065);
and U4784 (N_4784,In_176,In_2121);
nor U4785 (N_4785,In_63,In_2127);
and U4786 (N_4786,In_1109,In_1541);
nand U4787 (N_4787,In_440,In_363);
nor U4788 (N_4788,In_757,In_1281);
or U4789 (N_4789,In_2042,In_828);
or U4790 (N_4790,In_415,In_2059);
or U4791 (N_4791,In_2498,In_1046);
nor U4792 (N_4792,In_446,In_1414);
xor U4793 (N_4793,In_2125,In_18);
nor U4794 (N_4794,In_508,In_1133);
and U4795 (N_4795,In_1637,In_708);
nor U4796 (N_4796,In_1123,In_269);
or U4797 (N_4797,In_1521,In_528);
nand U4798 (N_4798,In_1368,In_1723);
xnor U4799 (N_4799,In_1855,In_1211);
and U4800 (N_4800,In_1034,In_1409);
xnor U4801 (N_4801,In_1236,In_2390);
or U4802 (N_4802,In_2495,In_2180);
and U4803 (N_4803,In_2066,In_2127);
nor U4804 (N_4804,In_1679,In_2331);
nand U4805 (N_4805,In_1660,In_16);
xnor U4806 (N_4806,In_2463,In_2409);
nand U4807 (N_4807,In_477,In_2392);
xor U4808 (N_4808,In_2133,In_1228);
or U4809 (N_4809,In_1293,In_291);
xnor U4810 (N_4810,In_579,In_1907);
or U4811 (N_4811,In_1815,In_1980);
nor U4812 (N_4812,In_1551,In_26);
xor U4813 (N_4813,In_865,In_1158);
and U4814 (N_4814,In_2431,In_1097);
nor U4815 (N_4815,In_1086,In_829);
or U4816 (N_4816,In_489,In_225);
or U4817 (N_4817,In_2039,In_1457);
nand U4818 (N_4818,In_2282,In_943);
and U4819 (N_4819,In_2302,In_1507);
nand U4820 (N_4820,In_1409,In_2030);
xor U4821 (N_4821,In_2085,In_935);
nand U4822 (N_4822,In_1513,In_837);
nand U4823 (N_4823,In_464,In_460);
nor U4824 (N_4824,In_1773,In_1194);
or U4825 (N_4825,In_2452,In_1750);
nor U4826 (N_4826,In_476,In_2022);
nand U4827 (N_4827,In_1075,In_2052);
and U4828 (N_4828,In_228,In_754);
or U4829 (N_4829,In_1248,In_515);
xnor U4830 (N_4830,In_1132,In_226);
and U4831 (N_4831,In_843,In_396);
or U4832 (N_4832,In_1160,In_686);
nand U4833 (N_4833,In_1414,In_473);
xnor U4834 (N_4834,In_1217,In_339);
or U4835 (N_4835,In_2269,In_85);
nand U4836 (N_4836,In_2201,In_1578);
and U4837 (N_4837,In_586,In_908);
and U4838 (N_4838,In_2243,In_469);
or U4839 (N_4839,In_1798,In_1334);
and U4840 (N_4840,In_660,In_403);
and U4841 (N_4841,In_816,In_1291);
nor U4842 (N_4842,In_1260,In_217);
nand U4843 (N_4843,In_2136,In_1398);
xor U4844 (N_4844,In_766,In_1672);
and U4845 (N_4845,In_2470,In_85);
and U4846 (N_4846,In_2099,In_312);
xor U4847 (N_4847,In_9,In_1237);
xnor U4848 (N_4848,In_1410,In_2245);
xnor U4849 (N_4849,In_2341,In_999);
and U4850 (N_4850,In_1139,In_2397);
nor U4851 (N_4851,In_278,In_1262);
nor U4852 (N_4852,In_1929,In_2229);
nand U4853 (N_4853,In_574,In_1296);
xor U4854 (N_4854,In_1598,In_61);
and U4855 (N_4855,In_1265,In_1489);
nand U4856 (N_4856,In_1699,In_139);
xnor U4857 (N_4857,In_2086,In_1880);
nor U4858 (N_4858,In_234,In_1796);
and U4859 (N_4859,In_216,In_647);
nor U4860 (N_4860,In_2492,In_617);
nand U4861 (N_4861,In_1163,In_1389);
and U4862 (N_4862,In_373,In_1845);
nor U4863 (N_4863,In_1652,In_109);
or U4864 (N_4864,In_1022,In_980);
and U4865 (N_4865,In_1284,In_1121);
xnor U4866 (N_4866,In_2413,In_171);
nand U4867 (N_4867,In_234,In_1087);
nand U4868 (N_4868,In_859,In_1237);
or U4869 (N_4869,In_372,In_1084);
or U4870 (N_4870,In_848,In_696);
and U4871 (N_4871,In_1316,In_1837);
nand U4872 (N_4872,In_1280,In_698);
xnor U4873 (N_4873,In_829,In_865);
and U4874 (N_4874,In_284,In_2083);
xor U4875 (N_4875,In_1620,In_1585);
nor U4876 (N_4876,In_668,In_1894);
xor U4877 (N_4877,In_1981,In_2345);
nor U4878 (N_4878,In_1093,In_204);
nor U4879 (N_4879,In_1890,In_1036);
nor U4880 (N_4880,In_1528,In_301);
and U4881 (N_4881,In_468,In_1441);
or U4882 (N_4882,In_548,In_2010);
or U4883 (N_4883,In_916,In_433);
nor U4884 (N_4884,In_108,In_498);
and U4885 (N_4885,In_3,In_350);
and U4886 (N_4886,In_2108,In_977);
nor U4887 (N_4887,In_775,In_2240);
nor U4888 (N_4888,In_1896,In_2032);
and U4889 (N_4889,In_1377,In_1674);
nand U4890 (N_4890,In_1624,In_1058);
nand U4891 (N_4891,In_2186,In_271);
nor U4892 (N_4892,In_38,In_566);
nor U4893 (N_4893,In_1090,In_2225);
xor U4894 (N_4894,In_1805,In_191);
nor U4895 (N_4895,In_1953,In_1146);
nand U4896 (N_4896,In_865,In_639);
and U4897 (N_4897,In_282,In_2175);
nand U4898 (N_4898,In_2054,In_156);
and U4899 (N_4899,In_534,In_1328);
nor U4900 (N_4900,In_2426,In_490);
nand U4901 (N_4901,In_687,In_1118);
or U4902 (N_4902,In_2180,In_1239);
nor U4903 (N_4903,In_459,In_1884);
xnor U4904 (N_4904,In_2391,In_1047);
xnor U4905 (N_4905,In_2316,In_1225);
xor U4906 (N_4906,In_1008,In_2113);
nand U4907 (N_4907,In_593,In_201);
or U4908 (N_4908,In_808,In_2012);
nor U4909 (N_4909,In_2482,In_2371);
xor U4910 (N_4910,In_884,In_1904);
xnor U4911 (N_4911,In_1783,In_404);
or U4912 (N_4912,In_1989,In_232);
nor U4913 (N_4913,In_445,In_531);
xnor U4914 (N_4914,In_1515,In_1252);
and U4915 (N_4915,In_452,In_2253);
or U4916 (N_4916,In_1679,In_391);
or U4917 (N_4917,In_2013,In_2027);
xor U4918 (N_4918,In_2057,In_1324);
xnor U4919 (N_4919,In_1962,In_1472);
xnor U4920 (N_4920,In_1443,In_1576);
nor U4921 (N_4921,In_1195,In_665);
xnor U4922 (N_4922,In_896,In_1530);
nand U4923 (N_4923,In_2087,In_603);
and U4924 (N_4924,In_1491,In_1575);
or U4925 (N_4925,In_2044,In_1850);
and U4926 (N_4926,In_265,In_2423);
and U4927 (N_4927,In_1055,In_1635);
nand U4928 (N_4928,In_679,In_1943);
nor U4929 (N_4929,In_565,In_269);
and U4930 (N_4930,In_709,In_1108);
and U4931 (N_4931,In_2144,In_1603);
xor U4932 (N_4932,In_1974,In_2426);
and U4933 (N_4933,In_927,In_1499);
nand U4934 (N_4934,In_2133,In_2181);
or U4935 (N_4935,In_1695,In_1482);
xor U4936 (N_4936,In_975,In_1087);
nand U4937 (N_4937,In_2313,In_1226);
nor U4938 (N_4938,In_522,In_1822);
nor U4939 (N_4939,In_531,In_2107);
or U4940 (N_4940,In_2031,In_1621);
nand U4941 (N_4941,In_422,In_113);
nand U4942 (N_4942,In_48,In_1793);
xnor U4943 (N_4943,In_2127,In_2386);
and U4944 (N_4944,In_1878,In_211);
and U4945 (N_4945,In_52,In_332);
nand U4946 (N_4946,In_1975,In_586);
or U4947 (N_4947,In_1866,In_1074);
nor U4948 (N_4948,In_394,In_1058);
or U4949 (N_4949,In_1542,In_1070);
xnor U4950 (N_4950,In_1613,In_1047);
or U4951 (N_4951,In_2490,In_2294);
and U4952 (N_4952,In_2111,In_334);
or U4953 (N_4953,In_1481,In_655);
or U4954 (N_4954,In_546,In_1384);
xnor U4955 (N_4955,In_2330,In_771);
or U4956 (N_4956,In_150,In_2396);
xnor U4957 (N_4957,In_1864,In_2258);
nand U4958 (N_4958,In_1608,In_1341);
nand U4959 (N_4959,In_1424,In_1463);
and U4960 (N_4960,In_2201,In_1495);
nand U4961 (N_4961,In_2455,In_375);
xor U4962 (N_4962,In_2137,In_1022);
or U4963 (N_4963,In_775,In_338);
xor U4964 (N_4964,In_191,In_700);
xor U4965 (N_4965,In_661,In_752);
or U4966 (N_4966,In_827,In_29);
nand U4967 (N_4967,In_1837,In_1414);
or U4968 (N_4968,In_1558,In_2447);
and U4969 (N_4969,In_232,In_1730);
and U4970 (N_4970,In_2086,In_2342);
nor U4971 (N_4971,In_1299,In_1346);
xor U4972 (N_4972,In_1321,In_2047);
or U4973 (N_4973,In_108,In_2382);
xnor U4974 (N_4974,In_2249,In_852);
xnor U4975 (N_4975,In_1052,In_127);
or U4976 (N_4976,In_1134,In_542);
nand U4977 (N_4977,In_2333,In_159);
or U4978 (N_4978,In_1199,In_200);
nor U4979 (N_4979,In_340,In_767);
nand U4980 (N_4980,In_106,In_728);
xor U4981 (N_4981,In_2091,In_1728);
or U4982 (N_4982,In_91,In_1647);
and U4983 (N_4983,In_1125,In_547);
nand U4984 (N_4984,In_1139,In_596);
and U4985 (N_4985,In_2466,In_1814);
nand U4986 (N_4986,In_779,In_2167);
or U4987 (N_4987,In_2291,In_951);
xnor U4988 (N_4988,In_142,In_125);
nor U4989 (N_4989,In_1031,In_736);
and U4990 (N_4990,In_1994,In_1129);
nand U4991 (N_4991,In_1994,In_584);
nor U4992 (N_4992,In_2438,In_1917);
or U4993 (N_4993,In_1469,In_518);
nor U4994 (N_4994,In_167,In_994);
or U4995 (N_4995,In_1448,In_162);
nand U4996 (N_4996,In_889,In_2097);
xnor U4997 (N_4997,In_848,In_2464);
and U4998 (N_4998,In_2392,In_1063);
nor U4999 (N_4999,In_2043,In_103);
and U5000 (N_5000,N_2798,N_2547);
or U5001 (N_5001,N_1102,N_3324);
nand U5002 (N_5002,N_4896,N_1644);
xor U5003 (N_5003,N_923,N_477);
nand U5004 (N_5004,N_3915,N_1976);
nand U5005 (N_5005,N_2054,N_3707);
nor U5006 (N_5006,N_2626,N_2042);
or U5007 (N_5007,N_1145,N_4664);
nor U5008 (N_5008,N_371,N_1186);
or U5009 (N_5009,N_2279,N_154);
nor U5010 (N_5010,N_3431,N_1387);
xor U5011 (N_5011,N_3042,N_3019);
xor U5012 (N_5012,N_2311,N_145);
or U5013 (N_5013,N_2212,N_1446);
xor U5014 (N_5014,N_2616,N_626);
xnor U5015 (N_5015,N_3885,N_243);
and U5016 (N_5016,N_1935,N_1943);
nand U5017 (N_5017,N_1837,N_3457);
nand U5018 (N_5018,N_2312,N_2278);
xnor U5019 (N_5019,N_1472,N_3239);
xnor U5020 (N_5020,N_4613,N_771);
or U5021 (N_5021,N_1505,N_1423);
and U5022 (N_5022,N_1802,N_2562);
and U5023 (N_5023,N_619,N_1192);
or U5024 (N_5024,N_2618,N_3739);
nor U5025 (N_5025,N_4863,N_3180);
or U5026 (N_5026,N_4378,N_354);
nand U5027 (N_5027,N_3361,N_1888);
and U5028 (N_5028,N_4551,N_2836);
xor U5029 (N_5029,N_4190,N_3528);
nand U5030 (N_5030,N_2275,N_121);
or U5031 (N_5031,N_1316,N_2296);
or U5032 (N_5032,N_2088,N_3421);
nor U5033 (N_5033,N_1738,N_4418);
xor U5034 (N_5034,N_1353,N_4466);
and U5035 (N_5035,N_1609,N_2660);
nor U5036 (N_5036,N_2153,N_1494);
xnor U5037 (N_5037,N_3166,N_2635);
nand U5038 (N_5038,N_898,N_2335);
and U5039 (N_5039,N_1389,N_763);
and U5040 (N_5040,N_2773,N_4230);
nor U5041 (N_5041,N_1425,N_4710);
xnor U5042 (N_5042,N_179,N_3723);
and U5043 (N_5043,N_1143,N_1638);
xnor U5044 (N_5044,N_4020,N_4216);
or U5045 (N_5045,N_2307,N_991);
xor U5046 (N_5046,N_3246,N_556);
nor U5047 (N_5047,N_410,N_3720);
nand U5048 (N_5048,N_1700,N_377);
nor U5049 (N_5049,N_1601,N_3852);
or U5050 (N_5050,N_1891,N_3592);
xnor U5051 (N_5051,N_3458,N_1307);
and U5052 (N_5052,N_4552,N_1750);
xor U5053 (N_5053,N_2848,N_4958);
and U5054 (N_5054,N_3798,N_2041);
xnor U5055 (N_5055,N_3197,N_4559);
xnor U5056 (N_5056,N_1180,N_1722);
xnor U5057 (N_5057,N_1386,N_2707);
xnor U5058 (N_5058,N_1590,N_56);
xor U5059 (N_5059,N_3022,N_4725);
xor U5060 (N_5060,N_3749,N_3972);
nand U5061 (N_5061,N_645,N_170);
nand U5062 (N_5062,N_1944,N_2829);
xnor U5063 (N_5063,N_3814,N_3511);
nor U5064 (N_5064,N_3102,N_1206);
xor U5065 (N_5065,N_2959,N_4001);
nand U5066 (N_5066,N_1304,N_3564);
nor U5067 (N_5067,N_2583,N_3759);
or U5068 (N_5068,N_2516,N_2491);
xnor U5069 (N_5069,N_217,N_3202);
xnor U5070 (N_5070,N_840,N_242);
nor U5071 (N_5071,N_1685,N_4821);
nor U5072 (N_5072,N_1203,N_4882);
nand U5073 (N_5073,N_2542,N_3524);
xor U5074 (N_5074,N_4037,N_2853);
and U5075 (N_5075,N_1281,N_4206);
and U5076 (N_5076,N_4900,N_4726);
xor U5077 (N_5077,N_4212,N_2699);
nand U5078 (N_5078,N_3030,N_3868);
nand U5079 (N_5079,N_1319,N_764);
or U5080 (N_5080,N_4269,N_2692);
nand U5081 (N_5081,N_2104,N_1642);
nand U5082 (N_5082,N_2418,N_990);
or U5083 (N_5083,N_3628,N_1936);
and U5084 (N_5084,N_1634,N_825);
and U5085 (N_5085,N_1189,N_4445);
and U5086 (N_5086,N_1939,N_1262);
xnor U5087 (N_5087,N_1381,N_3178);
or U5088 (N_5088,N_4605,N_1463);
nor U5089 (N_5089,N_1451,N_3263);
nand U5090 (N_5090,N_1178,N_3125);
and U5091 (N_5091,N_3168,N_3669);
and U5092 (N_5092,N_306,N_401);
or U5093 (N_5093,N_1371,N_3136);
xnor U5094 (N_5094,N_2741,N_3403);
nand U5095 (N_5095,N_2937,N_4695);
or U5096 (N_5096,N_3615,N_2291);
nand U5097 (N_5097,N_3398,N_882);
nand U5098 (N_5098,N_1777,N_3394);
or U5099 (N_5099,N_2754,N_3786);
nor U5100 (N_5100,N_393,N_3179);
xnor U5101 (N_5101,N_3252,N_4012);
nand U5102 (N_5102,N_1465,N_2305);
nand U5103 (N_5103,N_2302,N_3445);
or U5104 (N_5104,N_3145,N_111);
nor U5105 (N_5105,N_4729,N_3186);
nand U5106 (N_5106,N_2118,N_1483);
nor U5107 (N_5107,N_1558,N_286);
xnor U5108 (N_5108,N_2914,N_2405);
nand U5109 (N_5109,N_4154,N_2316);
xnor U5110 (N_5110,N_4063,N_1064);
and U5111 (N_5111,N_1683,N_3591);
xor U5112 (N_5112,N_3718,N_4781);
and U5113 (N_5113,N_283,N_997);
and U5114 (N_5114,N_107,N_666);
nand U5115 (N_5115,N_3436,N_4129);
nand U5116 (N_5116,N_3839,N_129);
xor U5117 (N_5117,N_2513,N_2258);
or U5118 (N_5118,N_774,N_1833);
nand U5119 (N_5119,N_4356,N_106);
nand U5120 (N_5120,N_916,N_1690);
nor U5121 (N_5121,N_806,N_4243);
nor U5122 (N_5122,N_2889,N_3687);
and U5123 (N_5123,N_2095,N_1670);
nor U5124 (N_5124,N_159,N_2230);
nand U5125 (N_5125,N_1736,N_3031);
xor U5126 (N_5126,N_1537,N_4225);
and U5127 (N_5127,N_1500,N_1689);
xnor U5128 (N_5128,N_1331,N_4921);
nor U5129 (N_5129,N_365,N_2374);
or U5130 (N_5130,N_4032,N_4213);
nor U5131 (N_5131,N_1117,N_4130);
nand U5132 (N_5132,N_2991,N_1204);
xor U5133 (N_5133,N_4351,N_93);
and U5134 (N_5134,N_4066,N_4280);
nor U5135 (N_5135,N_531,N_3934);
nand U5136 (N_5136,N_4752,N_1202);
and U5137 (N_5137,N_2930,N_47);
nor U5138 (N_5138,N_4348,N_3649);
or U5139 (N_5139,N_262,N_2522);
nor U5140 (N_5140,N_3945,N_60);
and U5141 (N_5141,N_3510,N_2928);
nor U5142 (N_5142,N_1395,N_3905);
xnor U5143 (N_5143,N_3552,N_3167);
xor U5144 (N_5144,N_4463,N_4555);
or U5145 (N_5145,N_358,N_4302);
or U5146 (N_5146,N_3083,N_1497);
or U5147 (N_5147,N_4678,N_3531);
xor U5148 (N_5148,N_4282,N_1677);
xnor U5149 (N_5149,N_832,N_2744);
nand U5150 (N_5150,N_2675,N_2185);
nor U5151 (N_5151,N_736,N_3008);
nor U5152 (N_5152,N_2384,N_2841);
or U5153 (N_5153,N_4353,N_1025);
or U5154 (N_5154,N_1867,N_4202);
or U5155 (N_5155,N_1630,N_2619);
nand U5156 (N_5156,N_3610,N_1985);
and U5157 (N_5157,N_4777,N_2375);
xor U5158 (N_5158,N_4274,N_32);
or U5159 (N_5159,N_4713,N_1013);
nand U5160 (N_5160,N_3288,N_2685);
nor U5161 (N_5161,N_4341,N_431);
or U5162 (N_5162,N_610,N_1421);
xor U5163 (N_5163,N_658,N_3100);
nand U5164 (N_5164,N_4343,N_1829);
and U5165 (N_5165,N_1751,N_3032);
nand U5166 (N_5166,N_344,N_3910);
nor U5167 (N_5167,N_3353,N_3514);
nand U5168 (N_5168,N_415,N_314);
and U5169 (N_5169,N_2080,N_2998);
or U5170 (N_5170,N_178,N_1665);
or U5171 (N_5171,N_457,N_4279);
nor U5172 (N_5172,N_211,N_1139);
nor U5173 (N_5173,N_1323,N_357);
xor U5174 (N_5174,N_3000,N_3602);
xnor U5175 (N_5175,N_3208,N_3677);
xor U5176 (N_5176,N_230,N_407);
nand U5177 (N_5177,N_691,N_3236);
nand U5178 (N_5178,N_1627,N_1266);
xor U5179 (N_5179,N_2443,N_2689);
xnor U5180 (N_5180,N_1995,N_3352);
nor U5181 (N_5181,N_335,N_4727);
nor U5182 (N_5182,N_4270,N_4352);
and U5183 (N_5183,N_1199,N_4359);
or U5184 (N_5184,N_2023,N_3900);
xor U5185 (N_5185,N_1699,N_2622);
or U5186 (N_5186,N_3396,N_887);
or U5187 (N_5187,N_1545,N_674);
or U5188 (N_5188,N_257,N_1084);
nand U5189 (N_5189,N_77,N_1187);
or U5190 (N_5190,N_4671,N_594);
nor U5191 (N_5191,N_1855,N_3123);
xnor U5192 (N_5192,N_3325,N_3800);
nor U5193 (N_5193,N_2144,N_4857);
nor U5194 (N_5194,N_746,N_3689);
and U5195 (N_5195,N_1058,N_4705);
nor U5196 (N_5196,N_2434,N_1903);
nand U5197 (N_5197,N_4536,N_897);
xnor U5198 (N_5198,N_1093,N_9);
nand U5199 (N_5199,N_2832,N_2243);
xor U5200 (N_5200,N_1578,N_2543);
nor U5201 (N_5201,N_4080,N_1223);
or U5202 (N_5202,N_4928,N_4634);
nor U5203 (N_5203,N_3805,N_3829);
xnor U5204 (N_5204,N_4150,N_347);
and U5205 (N_5205,N_4662,N_4055);
and U5206 (N_5206,N_4048,N_2891);
and U5207 (N_5207,N_4415,N_4148);
nor U5208 (N_5208,N_812,N_3973);
and U5209 (N_5209,N_792,N_533);
or U5210 (N_5210,N_1278,N_3542);
and U5211 (N_5211,N_2136,N_2590);
and U5212 (N_5212,N_837,N_3115);
or U5213 (N_5213,N_1980,N_4217);
nand U5214 (N_5214,N_3066,N_418);
and U5215 (N_5215,N_1173,N_1863);
nor U5216 (N_5216,N_3381,N_3301);
nand U5217 (N_5217,N_947,N_2470);
nand U5218 (N_5218,N_4715,N_2645);
nor U5219 (N_5219,N_1660,N_2130);
or U5220 (N_5220,N_3705,N_863);
and U5221 (N_5221,N_4375,N_68);
and U5222 (N_5222,N_3266,N_1585);
and U5223 (N_5223,N_2141,N_3340);
or U5224 (N_5224,N_3496,N_2428);
xnor U5225 (N_5225,N_4438,N_4930);
nor U5226 (N_5226,N_3118,N_2849);
or U5227 (N_5227,N_1506,N_1466);
nor U5228 (N_5228,N_2568,N_4677);
nand U5229 (N_5229,N_1429,N_23);
or U5230 (N_5230,N_3721,N_3223);
xor U5231 (N_5231,N_2628,N_1551);
and U5232 (N_5232,N_1334,N_4510);
or U5233 (N_5233,N_4170,N_4983);
or U5234 (N_5234,N_2931,N_4108);
xnor U5235 (N_5235,N_970,N_993);
nor U5236 (N_5236,N_4594,N_1357);
xnor U5237 (N_5237,N_844,N_2961);
nor U5238 (N_5238,N_4446,N_2110);
and U5239 (N_5239,N_2170,N_1568);
and U5240 (N_5240,N_3029,N_4842);
xnor U5241 (N_5241,N_3439,N_4006);
xor U5242 (N_5242,N_215,N_1368);
xor U5243 (N_5243,N_482,N_4482);
and U5244 (N_5244,N_38,N_139);
xnor U5245 (N_5245,N_3751,N_3161);
nand U5246 (N_5246,N_805,N_2733);
and U5247 (N_5247,N_2775,N_1258);
xor U5248 (N_5248,N_566,N_1635);
xor U5249 (N_5249,N_2875,N_113);
nor U5250 (N_5250,N_1890,N_218);
nor U5251 (N_5251,N_384,N_4694);
and U5252 (N_5252,N_267,N_2532);
nand U5253 (N_5253,N_4593,N_3771);
nand U5254 (N_5254,N_1277,N_2032);
nor U5255 (N_5255,N_2360,N_2072);
xor U5256 (N_5256,N_4542,N_3138);
or U5257 (N_5257,N_828,N_3219);
and U5258 (N_5258,N_278,N_304);
xnor U5259 (N_5259,N_4519,N_3764);
nor U5260 (N_5260,N_3788,N_2455);
xor U5261 (N_5261,N_3311,N_3386);
xnor U5262 (N_5262,N_2046,N_315);
nand U5263 (N_5263,N_3221,N_3681);
nor U5264 (N_5264,N_4755,N_4679);
nor U5265 (N_5265,N_3757,N_938);
and U5266 (N_5266,N_4751,N_299);
nand U5267 (N_5267,N_2168,N_2276);
xor U5268 (N_5268,N_3304,N_1898);
xor U5269 (N_5269,N_3545,N_1375);
or U5270 (N_5270,N_1248,N_2815);
or U5271 (N_5271,N_3489,N_2833);
xor U5272 (N_5272,N_3670,N_2538);
nand U5273 (N_5273,N_744,N_3449);
nand U5274 (N_5274,N_4589,N_506);
xnor U5275 (N_5275,N_657,N_821);
and U5276 (N_5276,N_3404,N_2077);
nand U5277 (N_5277,N_3758,N_2843);
nor U5278 (N_5278,N_3565,N_3388);
and U5279 (N_5279,N_768,N_3152);
nand U5280 (N_5280,N_653,N_3026);
and U5281 (N_5281,N_3354,N_4905);
nand U5282 (N_5282,N_4918,N_1435);
and U5283 (N_5283,N_2245,N_4647);
or U5284 (N_5284,N_1827,N_4383);
or U5285 (N_5285,N_2482,N_1132);
nor U5286 (N_5286,N_3994,N_1716);
or U5287 (N_5287,N_185,N_2440);
nor U5288 (N_5288,N_2872,N_2386);
and U5289 (N_5289,N_1794,N_2356);
xnor U5290 (N_5290,N_2999,N_4616);
nand U5291 (N_5291,N_4068,N_553);
nand U5292 (N_5292,N_1150,N_3142);
or U5293 (N_5293,N_1507,N_3430);
nand U5294 (N_5294,N_4711,N_988);
and U5295 (N_5295,N_1174,N_3117);
xor U5296 (N_5296,N_1687,N_4826);
nand U5297 (N_5297,N_2942,N_497);
nor U5298 (N_5298,N_4574,N_1648);
or U5299 (N_5299,N_2385,N_224);
nand U5300 (N_5300,N_1619,N_3081);
xor U5301 (N_5301,N_1999,N_1061);
xnor U5302 (N_5302,N_3466,N_3819);
or U5303 (N_5303,N_3065,N_4408);
or U5304 (N_5304,N_4157,N_4088);
or U5305 (N_5305,N_849,N_3497);
xor U5306 (N_5306,N_875,N_3589);
nand U5307 (N_5307,N_690,N_3544);
nor U5308 (N_5308,N_4163,N_2329);
or U5309 (N_5309,N_4633,N_4911);
or U5310 (N_5310,N_3087,N_3237);
xnor U5311 (N_5311,N_1671,N_2755);
or U5312 (N_5312,N_555,N_601);
xnor U5313 (N_5313,N_3981,N_751);
xor U5314 (N_5314,N_3355,N_900);
nor U5315 (N_5315,N_2390,N_1808);
and U5316 (N_5316,N_1300,N_4123);
or U5317 (N_5317,N_4475,N_1523);
nand U5318 (N_5318,N_2975,N_148);
or U5319 (N_5319,N_1346,N_730);
nand U5320 (N_5320,N_2238,N_2973);
xnor U5321 (N_5321,N_4447,N_1873);
nand U5322 (N_5322,N_438,N_539);
nand U5323 (N_5323,N_3982,N_3068);
xor U5324 (N_5324,N_1439,N_4291);
and U5325 (N_5325,N_2309,N_4102);
xor U5326 (N_5326,N_2352,N_3257);
nand U5327 (N_5327,N_3777,N_2953);
and U5328 (N_5328,N_964,N_759);
nor U5329 (N_5329,N_4388,N_2525);
and U5330 (N_5330,N_2293,N_2608);
nand U5331 (N_5331,N_3663,N_2284);
or U5332 (N_5332,N_4702,N_274);
or U5333 (N_5333,N_1287,N_2079);
and U5334 (N_5334,N_4578,N_2936);
or U5335 (N_5335,N_785,N_3987);
nand U5336 (N_5336,N_3728,N_4231);
nor U5337 (N_5337,N_2581,N_4172);
nor U5338 (N_5338,N_2207,N_4053);
nand U5339 (N_5339,N_4128,N_2987);
or U5340 (N_5340,N_1596,N_4806);
nand U5341 (N_5341,N_4237,N_4606);
nand U5342 (N_5342,N_4234,N_1884);
and U5343 (N_5343,N_2036,N_4512);
and U5344 (N_5344,N_4743,N_1442);
nor U5345 (N_5345,N_3321,N_1851);
and U5346 (N_5346,N_295,N_1979);
nand U5347 (N_5347,N_2621,N_2711);
and U5348 (N_5348,N_979,N_4041);
nor U5349 (N_5349,N_2317,N_628);
nor U5350 (N_5350,N_4034,N_726);
and U5351 (N_5351,N_1495,N_2177);
nand U5352 (N_5352,N_1654,N_925);
nor U5353 (N_5353,N_3411,N_3743);
xor U5354 (N_5354,N_3172,N_4615);
and U5355 (N_5355,N_3604,N_340);
nand U5356 (N_5356,N_2518,N_307);
xor U5357 (N_5357,N_1901,N_3998);
and U5358 (N_5358,N_4016,N_2250);
nor U5359 (N_5359,N_99,N_864);
nor U5360 (N_5360,N_3909,N_4923);
xnor U5361 (N_5361,N_436,N_4372);
or U5362 (N_5362,N_190,N_2705);
and U5363 (N_5363,N_4203,N_4778);
and U5364 (N_5364,N_878,N_4908);
and U5365 (N_5365,N_752,N_1631);
and U5366 (N_5366,N_2857,N_2617);
nand U5367 (N_5367,N_1170,N_2641);
xnor U5368 (N_5368,N_237,N_4669);
nand U5369 (N_5369,N_3253,N_1790);
xnor U5370 (N_5370,N_3966,N_1260);
nor U5371 (N_5371,N_4953,N_2379);
and U5372 (N_5372,N_1356,N_1945);
nor U5373 (N_5373,N_2129,N_4252);
or U5374 (N_5374,N_2272,N_419);
nand U5375 (N_5375,N_2084,N_885);
nor U5376 (N_5376,N_3175,N_2520);
nor U5377 (N_5377,N_3995,N_3903);
and U5378 (N_5378,N_2392,N_1676);
nor U5379 (N_5379,N_4955,N_817);
or U5380 (N_5380,N_3182,N_81);
or U5381 (N_5381,N_2827,N_3048);
or U5382 (N_5382,N_2703,N_4061);
nor U5383 (N_5383,N_2753,N_3279);
nor U5384 (N_5384,N_2407,N_2657);
and U5385 (N_5385,N_3184,N_1309);
and U5386 (N_5386,N_4854,N_3317);
xnor U5387 (N_5387,N_4984,N_3918);
nor U5388 (N_5388,N_2447,N_289);
xor U5389 (N_5389,N_2219,N_3134);
and U5390 (N_5390,N_1768,N_2866);
nand U5391 (N_5391,N_3997,N_667);
or U5392 (N_5392,N_3285,N_1679);
xor U5393 (N_5393,N_4367,N_4666);
and U5394 (N_5394,N_4745,N_723);
and U5395 (N_5395,N_44,N_2123);
and U5396 (N_5396,N_310,N_4501);
and U5397 (N_5397,N_4637,N_1526);
nand U5398 (N_5398,N_3896,N_4509);
nand U5399 (N_5399,N_2623,N_2607);
nand U5400 (N_5400,N_188,N_4506);
or U5401 (N_5401,N_3699,N_3477);
or U5402 (N_5402,N_2499,N_2612);
nor U5403 (N_5403,N_4145,N_387);
xor U5404 (N_5404,N_3907,N_319);
nand U5405 (N_5405,N_984,N_1961);
nor U5406 (N_5406,N_1172,N_3472);
and U5407 (N_5407,N_2188,N_1055);
xnor U5408 (N_5408,N_3673,N_2728);
nand U5409 (N_5409,N_4884,N_3332);
or U5410 (N_5410,N_3756,N_1691);
and U5411 (N_5411,N_941,N_2341);
nand U5412 (N_5412,N_3974,N_1735);
nand U5413 (N_5413,N_982,N_4558);
and U5414 (N_5414,N_2464,N_1608);
nor U5415 (N_5415,N_2361,N_4158);
and U5416 (N_5416,N_1107,N_3011);
and U5417 (N_5417,N_3790,N_4043);
xor U5418 (N_5418,N_4720,N_239);
or U5419 (N_5419,N_3731,N_2887);
xnor U5420 (N_5420,N_3703,N_4364);
xnor U5421 (N_5421,N_487,N_4763);
nand U5422 (N_5422,N_2138,N_1940);
nand U5423 (N_5423,N_4808,N_784);
nand U5424 (N_5424,N_1407,N_4480);
or U5425 (N_5425,N_3349,N_1664);
and U5426 (N_5426,N_1938,N_2636);
xor U5427 (N_5427,N_1951,N_2571);
or U5428 (N_5428,N_4277,N_3928);
and U5429 (N_5429,N_2403,N_1096);
nand U5430 (N_5430,N_2481,N_1746);
and U5431 (N_5431,N_4389,N_1325);
xnor U5432 (N_5432,N_3712,N_921);
xnor U5433 (N_5433,N_2727,N_3760);
and U5434 (N_5434,N_1487,N_3665);
xnor U5435 (N_5435,N_1835,N_3432);
and U5436 (N_5436,N_1820,N_3948);
and U5437 (N_5437,N_2839,N_2181);
nand U5438 (N_5438,N_4174,N_4297);
xor U5439 (N_5439,N_2759,N_3519);
nor U5440 (N_5440,N_798,N_558);
xor U5441 (N_5441,N_3444,N_4377);
and U5442 (N_5442,N_2164,N_4073);
xor U5443 (N_5443,N_2395,N_1544);
xnor U5444 (N_5444,N_3601,N_4404);
xnor U5445 (N_5445,N_3890,N_3516);
or U5446 (N_5446,N_490,N_2974);
xnor U5447 (N_5447,N_21,N_485);
or U5448 (N_5448,N_1989,N_3877);
nor U5449 (N_5449,N_890,N_177);
xnor U5450 (N_5450,N_4619,N_4342);
or U5451 (N_5451,N_3916,N_29);
xnor U5452 (N_5452,N_4442,N_1052);
nor U5453 (N_5453,N_1434,N_4060);
xor U5454 (N_5454,N_836,N_1807);
or U5455 (N_5455,N_3043,N_4008);
nand U5456 (N_5456,N_3277,N_18);
xnor U5457 (N_5457,N_3787,N_2368);
nand U5458 (N_5458,N_4503,N_2512);
nor U5459 (N_5459,N_4897,N_4820);
and U5460 (N_5460,N_3268,N_1987);
nand U5461 (N_5461,N_3680,N_1522);
or U5462 (N_5462,N_108,N_2476);
or U5463 (N_5463,N_2005,N_3135);
xnor U5464 (N_5464,N_579,N_3379);
and U5465 (N_5465,N_670,N_2318);
and U5466 (N_5466,N_4429,N_1632);
xor U5467 (N_5467,N_3284,N_2659);
or U5468 (N_5468,N_2150,N_727);
or U5469 (N_5469,N_933,N_587);
or U5470 (N_5470,N_2061,N_2203);
nand U5471 (N_5471,N_1021,N_1729);
nand U5472 (N_5472,N_412,N_1211);
nor U5473 (N_5473,N_3679,N_4740);
xor U5474 (N_5474,N_4137,N_61);
xor U5475 (N_5475,N_408,N_1714);
nand U5476 (N_5476,N_2682,N_998);
and U5477 (N_5477,N_4511,N_4644);
nand U5478 (N_5478,N_1858,N_3232);
nand U5479 (N_5479,N_4192,N_3474);
and U5480 (N_5480,N_4126,N_2429);
and U5481 (N_5481,N_2591,N_4222);
and U5482 (N_5482,N_3770,N_1663);
xor U5483 (N_5483,N_1707,N_201);
nor U5484 (N_5484,N_623,N_4);
xor U5485 (N_5485,N_2415,N_4653);
nor U5486 (N_5486,N_1245,N_2022);
and U5487 (N_5487,N_3715,N_3181);
xor U5488 (N_5488,N_4609,N_2267);
nor U5489 (N_5489,N_3391,N_624);
or U5490 (N_5490,N_3855,N_1535);
nor U5491 (N_5491,N_4071,N_2157);
and U5492 (N_5492,N_4464,N_3200);
nor U5493 (N_5493,N_1928,N_4424);
or U5494 (N_5494,N_1074,N_1036);
xnor U5495 (N_5495,N_3275,N_816);
and U5496 (N_5496,N_4693,N_3062);
nor U5497 (N_5497,N_4879,N_2894);
nand U5498 (N_5498,N_4996,N_1039);
nor U5499 (N_5499,N_609,N_165);
nor U5500 (N_5500,N_1050,N_3120);
nand U5501 (N_5501,N_4046,N_67);
or U5502 (N_5502,N_84,N_3189);
and U5503 (N_5503,N_3682,N_327);
nand U5504 (N_5504,N_4608,N_1549);
and U5505 (N_5505,N_4259,N_2769);
xnor U5506 (N_5506,N_2015,N_4887);
and U5507 (N_5507,N_3023,N_4058);
nand U5508 (N_5508,N_2890,N_4161);
and U5509 (N_5509,N_4621,N_1196);
and U5510 (N_5510,N_492,N_336);
nand U5511 (N_5511,N_3639,N_3272);
or U5512 (N_5512,N_1006,N_4214);
or U5513 (N_5513,N_473,N_4290);
nand U5514 (N_5514,N_4931,N_4125);
and U5515 (N_5515,N_4455,N_434);
or U5516 (N_5516,N_2584,N_4205);
nor U5517 (N_5517,N_2346,N_1184);
xnor U5518 (N_5518,N_1000,N_4638);
nand U5519 (N_5519,N_4439,N_1040);
or U5520 (N_5520,N_22,N_4146);
and U5521 (N_5521,N_4612,N_3141);
or U5522 (N_5522,N_2073,N_895);
and U5523 (N_5523,N_1254,N_1821);
or U5524 (N_5524,N_2932,N_1090);
nor U5525 (N_5525,N_2465,N_4306);
xnor U5526 (N_5526,N_1744,N_720);
xor U5527 (N_5527,N_2760,N_413);
and U5528 (N_5528,N_4532,N_2630);
and U5529 (N_5529,N_2472,N_1268);
xor U5530 (N_5530,N_903,N_1498);
xor U5531 (N_5531,N_3571,N_101);
and U5532 (N_5532,N_1992,N_2174);
or U5533 (N_5533,N_3647,N_647);
and U5534 (N_5534,N_824,N_1809);
nor U5535 (N_5535,N_2693,N_2548);
xnor U5536 (N_5536,N_4982,N_1476);
and U5537 (N_5537,N_3148,N_879);
or U5538 (N_5538,N_3664,N_69);
and U5539 (N_5539,N_3440,N_3803);
nand U5540 (N_5540,N_4494,N_1237);
nand U5541 (N_5541,N_4479,N_3952);
nor U5542 (N_5542,N_4964,N_4948);
nor U5543 (N_5543,N_2126,N_4891);
and U5544 (N_5544,N_4758,N_3520);
nand U5545 (N_5545,N_1471,N_3280);
nand U5546 (N_5546,N_4260,N_1902);
and U5547 (N_5547,N_4913,N_2251);
xor U5548 (N_5548,N_2466,N_4696);
and U5549 (N_5549,N_2109,N_3625);
and U5550 (N_5550,N_298,N_2691);
nor U5551 (N_5551,N_738,N_1966);
nand U5552 (N_5552,N_1490,N_2572);
nand U5553 (N_5553,N_3072,N_3769);
and U5554 (N_5554,N_4014,N_912);
or U5555 (N_5555,N_3463,N_3911);
or U5556 (N_5556,N_2195,N_1123);
xnor U5557 (N_5557,N_332,N_1003);
nor U5558 (N_5558,N_4888,N_386);
nand U5559 (N_5559,N_4833,N_1034);
nand U5560 (N_5560,N_2217,N_756);
or U5561 (N_5561,N_1286,N_2970);
xnor U5562 (N_5562,N_2024,N_2190);
or U5563 (N_5563,N_4187,N_4036);
nand U5564 (N_5564,N_2864,N_3986);
nand U5565 (N_5565,N_4197,N_2915);
nand U5566 (N_5566,N_46,N_134);
and U5567 (N_5567,N_3162,N_2260);
nand U5568 (N_5568,N_2821,N_175);
or U5569 (N_5569,N_2546,N_4314);
and U5570 (N_5570,N_3261,N_544);
xor U5571 (N_5571,N_1711,N_1070);
or U5572 (N_5572,N_2738,N_2156);
nor U5573 (N_5573,N_1011,N_3385);
nor U5574 (N_5574,N_3082,N_4898);
nor U5575 (N_5575,N_4379,N_3674);
nand U5576 (N_5576,N_312,N_4529);
xor U5577 (N_5577,N_3061,N_193);
nand U5578 (N_5578,N_2381,N_2826);
xor U5579 (N_5579,N_1641,N_4468);
or U5580 (N_5580,N_2098,N_3825);
or U5581 (N_5581,N_4135,N_1885);
and U5582 (N_5582,N_2901,N_4837);
nor U5583 (N_5583,N_1154,N_1475);
xnor U5584 (N_5584,N_648,N_3719);
nor U5585 (N_5585,N_1511,N_695);
or U5586 (N_5586,N_395,N_2947);
and U5587 (N_5587,N_1610,N_4937);
or U5588 (N_5588,N_1591,N_144);
nor U5589 (N_5589,N_2698,N_2828);
nand U5590 (N_5590,N_4856,N_227);
or U5591 (N_5591,N_2069,N_3126);
nand U5592 (N_5592,N_949,N_2541);
nor U5593 (N_5593,N_2752,N_4050);
or U5594 (N_5594,N_4874,N_2117);
or U5595 (N_5595,N_3983,N_2913);
xor U5596 (N_5596,N_537,N_2202);
nor U5597 (N_5597,N_699,N_630);
nand U5598 (N_5598,N_4793,N_381);
xnor U5599 (N_5599,N_914,N_348);
and U5600 (N_5600,N_2160,N_2327);
nand U5601 (N_5601,N_430,N_1845);
nor U5602 (N_5602,N_2421,N_4030);
and U5603 (N_5603,N_2644,N_2736);
or U5604 (N_5604,N_3265,N_3468);
nor U5605 (N_5605,N_3633,N_1789);
nor U5606 (N_5606,N_402,N_507);
or U5607 (N_5607,N_173,N_1219);
or U5608 (N_5608,N_3395,N_935);
xor U5609 (N_5609,N_3638,N_2265);
and U5610 (N_5610,N_905,N_4827);
nor U5611 (N_5611,N_260,N_3849);
and U5612 (N_5612,N_4832,N_1493);
and U5613 (N_5613,N_4401,N_1194);
or U5614 (N_5614,N_3400,N_526);
xnor U5615 (N_5615,N_603,N_1388);
and U5616 (N_5616,N_3848,N_1524);
xnor U5617 (N_5617,N_4570,N_1942);
nand U5618 (N_5618,N_2445,N_3745);
nand U5619 (N_5619,N_3206,N_2480);
or U5620 (N_5620,N_3741,N_4200);
or U5621 (N_5621,N_503,N_491);
xnor U5622 (N_5622,N_1761,N_2940);
or U5623 (N_5623,N_280,N_4659);
nand U5624 (N_5624,N_4717,N_2977);
xnor U5625 (N_5625,N_4318,N_363);
xnor U5626 (N_5626,N_4209,N_3906);
nand U5627 (N_5627,N_3921,N_317);
and U5628 (N_5628,N_677,N_4005);
xnor U5629 (N_5629,N_4119,N_223);
or U5630 (N_5630,N_292,N_486);
nor U5631 (N_5631,N_4360,N_3558);
nand U5632 (N_5632,N_2663,N_4394);
xor U5633 (N_5633,N_3697,N_3807);
nand U5634 (N_5634,N_1452,N_2816);
and U5635 (N_5635,N_4077,N_4947);
or U5636 (N_5636,N_3384,N_3414);
nand U5637 (N_5637,N_452,N_2354);
and U5638 (N_5638,N_1704,N_4105);
nor U5639 (N_5639,N_17,N_1149);
nor U5640 (N_5640,N_1133,N_573);
and U5641 (N_5641,N_2763,N_2345);
nand U5642 (N_5642,N_4477,N_569);
nor U5643 (N_5643,N_367,N_3867);
nand U5644 (N_5644,N_2241,N_4554);
nand U5645 (N_5645,N_3962,N_4792);
and U5646 (N_5646,N_2175,N_4591);
nand U5647 (N_5647,N_3704,N_311);
nand U5648 (N_5648,N_686,N_813);
xnor U5649 (N_5649,N_1567,N_3348);
and U5650 (N_5650,N_323,N_356);
nand U5651 (N_5651,N_1385,N_4870);
and U5652 (N_5652,N_2114,N_4668);
xor U5653 (N_5653,N_4675,N_1467);
and U5654 (N_5654,N_1302,N_2344);
nand U5655 (N_5655,N_2349,N_3583);
or U5656 (N_5656,N_2782,N_4628);
nand U5657 (N_5657,N_2493,N_765);
xnor U5658 (N_5658,N_4334,N_4788);
and U5659 (N_5659,N_2633,N_4449);
nor U5660 (N_5660,N_819,N_3794);
and U5661 (N_5661,N_883,N_4822);
or U5662 (N_5662,N_3776,N_2063);
nor U5663 (N_5663,N_2722,N_3851);
nand U5664 (N_5664,N_4266,N_4284);
nor U5665 (N_5665,N_449,N_4708);
nor U5666 (N_5666,N_2536,N_2325);
nor U5667 (N_5667,N_4021,N_1811);
and U5668 (N_5668,N_1692,N_1105);
nor U5669 (N_5669,N_662,N_796);
or U5670 (N_5670,N_3747,N_3336);
or U5671 (N_5671,N_2173,N_2904);
nor U5672 (N_5672,N_814,N_2783);
xnor U5673 (N_5673,N_2059,N_4308);
nor U5674 (N_5674,N_166,N_1126);
or U5675 (N_5675,N_3199,N_1456);
or U5676 (N_5676,N_3410,N_4261);
nor U5677 (N_5677,N_2868,N_3557);
nor U5678 (N_5678,N_2824,N_169);
nand U5679 (N_5679,N_3260,N_3858);
and U5680 (N_5680,N_1019,N_271);
nor U5681 (N_5681,N_927,N_1810);
and U5682 (N_5682,N_3286,N_1763);
or U5683 (N_5683,N_4825,N_2225);
xor U5684 (N_5684,N_2952,N_1116);
xnor U5685 (N_5685,N_1419,N_1740);
xor U5686 (N_5686,N_1239,N_4070);
nor U5687 (N_5687,N_3131,N_1032);
xor U5688 (N_5688,N_4117,N_256);
nor U5689 (N_5689,N_2863,N_3211);
nor U5690 (N_5690,N_3887,N_1779);
xnor U5691 (N_5691,N_3201,N_598);
and U5692 (N_5692,N_3041,N_2021);
xor U5693 (N_5693,N_4766,N_1818);
nor U5694 (N_5694,N_4583,N_1303);
and U5695 (N_5695,N_4299,N_3536);
xnor U5696 (N_5696,N_4002,N_3282);
xnor U5697 (N_5697,N_1986,N_1250);
and U5698 (N_5698,N_4436,N_2730);
nor U5699 (N_5699,N_1795,N_4434);
nand U5700 (N_5700,N_92,N_301);
or U5701 (N_5701,N_2003,N_4681);
xor U5702 (N_5702,N_1892,N_3174);
or U5703 (N_5703,N_1043,N_4771);
and U5704 (N_5704,N_1168,N_2561);
nor U5705 (N_5705,N_461,N_3441);
or U5706 (N_5706,N_1361,N_2900);
nor U5707 (N_5707,N_3873,N_2310);
nand U5708 (N_5708,N_2478,N_4267);
and U5709 (N_5709,N_4999,N_3685);
nor U5710 (N_5710,N_2811,N_454);
xor U5711 (N_5711,N_3320,N_4687);
xnor U5712 (N_5712,N_4876,N_4538);
or U5713 (N_5713,N_2083,N_1166);
nor U5714 (N_5714,N_2357,N_1509);
nor U5715 (N_5715,N_3862,N_1846);
or U5716 (N_5716,N_3630,N_1153);
or U5717 (N_5717,N_3193,N_2876);
nor U5718 (N_5718,N_2473,N_1098);
xnor U5719 (N_5719,N_423,N_2001);
nor U5720 (N_5720,N_1376,N_3842);
nand U5721 (N_5721,N_4527,N_1825);
xnor U5722 (N_5722,N_987,N_1366);
or U5723 (N_5723,N_4845,N_3515);
or U5724 (N_5724,N_2554,N_1925);
and U5725 (N_5725,N_313,N_2762);
or U5726 (N_5726,N_416,N_2206);
and U5727 (N_5727,N_4818,N_383);
and U5728 (N_5728,N_1314,N_4772);
or U5729 (N_5729,N_2732,N_128);
xor U5730 (N_5730,N_3053,N_4657);
and U5731 (N_5731,N_1629,N_4207);
nor U5732 (N_5732,N_1169,N_1198);
nand U5733 (N_5733,N_1780,N_2809);
nand U5734 (N_5734,N_4847,N_2939);
nor U5735 (N_5735,N_3701,N_1176);
nor U5736 (N_5736,N_2962,N_4300);
and U5737 (N_5737,N_2264,N_4617);
nand U5738 (N_5738,N_3503,N_85);
or U5739 (N_5739,N_2640,N_1349);
and U5740 (N_5740,N_4361,N_4052);
nand U5741 (N_5741,N_2045,N_2819);
or U5742 (N_5742,N_2847,N_2056);
and U5743 (N_5743,N_793,N_3795);
xnor U5744 (N_5744,N_995,N_368);
and U5745 (N_5745,N_4571,N_3020);
and U5746 (N_5746,N_3572,N_1539);
or U5747 (N_5747,N_2948,N_1501);
and U5748 (N_5748,N_2982,N_4786);
or U5749 (N_5749,N_1351,N_1622);
nand U5750 (N_5750,N_2820,N_4627);
nor U5751 (N_5751,N_426,N_596);
or U5752 (N_5752,N_2789,N_3686);
nand U5753 (N_5753,N_4191,N_1322);
and U5754 (N_5754,N_959,N_515);
nand U5755 (N_5755,N_710,N_2433);
nand U5756 (N_5756,N_2492,N_4018);
or U5757 (N_5757,N_4487,N_3356);
or U5758 (N_5758,N_4895,N_3483);
nand U5759 (N_5759,N_2261,N_1606);
and U5760 (N_5760,N_251,N_236);
or U5761 (N_5761,N_4387,N_1159);
and U5762 (N_5762,N_1125,N_2283);
nand U5763 (N_5763,N_4839,N_458);
and U5764 (N_5764,N_4962,N_2090);
and U5765 (N_5765,N_1384,N_489);
nand U5766 (N_5766,N_1227,N_4180);
nor U5767 (N_5767,N_2570,N_25);
xor U5768 (N_5768,N_3996,N_2132);
or U5769 (N_5769,N_2993,N_3217);
nor U5770 (N_5770,N_4915,N_3314);
or U5771 (N_5771,N_4390,N_854);
and U5772 (N_5772,N_3375,N_3094);
nor U5773 (N_5773,N_2417,N_876);
and U5774 (N_5774,N_3024,N_513);
or U5775 (N_5775,N_4855,N_398);
and U5776 (N_5776,N_1165,N_975);
xnor U5777 (N_5777,N_4848,N_3331);
xor U5778 (N_5778,N_1294,N_1621);
nand U5779 (N_5779,N_3753,N_3054);
and U5780 (N_5780,N_2688,N_2879);
and U5781 (N_5781,N_359,N_1955);
nor U5782 (N_5782,N_4760,N_1124);
nor U5783 (N_5783,N_1066,N_3696);
and U5784 (N_5784,N_530,N_4169);
nand U5785 (N_5785,N_153,N_4366);
or U5786 (N_5786,N_3850,N_4090);
and U5787 (N_5787,N_3844,N_1212);
nand U5788 (N_5788,N_3821,N_3621);
nand U5789 (N_5789,N_4892,N_4471);
nand U5790 (N_5790,N_4398,N_3936);
nand U5791 (N_5791,N_973,N_1478);
nor U5792 (N_5792,N_2449,N_856);
xnor U5793 (N_5793,N_4699,N_1950);
or U5794 (N_5794,N_2595,N_4556);
or U5795 (N_5795,N_1355,N_631);
nor U5796 (N_5796,N_3836,N_1296);
nor U5797 (N_5797,N_2049,N_1119);
nor U5798 (N_5798,N_2859,N_3044);
nand U5799 (N_5799,N_15,N_1826);
and U5800 (N_5800,N_1848,N_1653);
or U5801 (N_5801,N_1510,N_1702);
or U5802 (N_5802,N_1042,N_2563);
xnor U5803 (N_5803,N_3541,N_3357);
nand U5804 (N_5804,N_1907,N_3713);
nand U5805 (N_5805,N_2496,N_2574);
nor U5806 (N_5806,N_3423,N_3377);
xnor U5807 (N_5807,N_206,N_3706);
and U5808 (N_5808,N_3941,N_155);
or U5809 (N_5809,N_2831,N_2718);
nand U5810 (N_5810,N_4196,N_1092);
nand U5811 (N_5811,N_2615,N_583);
or U5812 (N_5812,N_1378,N_716);
xnor U5813 (N_5813,N_1803,N_502);
nand U5814 (N_5814,N_3343,N_4176);
nand U5815 (N_5815,N_4860,N_599);
nor U5816 (N_5816,N_7,N_2351);
and U5817 (N_5817,N_2115,N_1785);
and U5818 (N_5818,N_4120,N_4661);
xnor U5819 (N_5819,N_1458,N_82);
and U5820 (N_5820,N_3233,N_3269);
and U5821 (N_5821,N_614,N_1282);
and U5822 (N_5822,N_2587,N_2226);
nand U5823 (N_5823,N_2147,N_4103);
nand U5824 (N_5824,N_1911,N_992);
nand U5825 (N_5825,N_1253,N_577);
or U5826 (N_5826,N_1428,N_2119);
nor U5827 (N_5827,N_3015,N_3487);
nor U5828 (N_5828,N_559,N_2979);
xor U5829 (N_5829,N_1252,N_4219);
nand U5830 (N_5830,N_1529,N_73);
or U5831 (N_5831,N_901,N_1409);
xnor U5832 (N_5832,N_24,N_3659);
and U5833 (N_5833,N_4272,N_635);
nor U5834 (N_5834,N_1367,N_4584);
nand U5835 (N_5835,N_66,N_1949);
xor U5836 (N_5836,N_1703,N_4013);
xor U5837 (N_5837,N_53,N_4087);
nand U5838 (N_5838,N_4650,N_4354);
nand U5839 (N_5839,N_1272,N_209);
nor U5840 (N_5840,N_552,N_1542);
and U5841 (N_5841,N_2923,N_839);
xor U5842 (N_5842,N_3700,N_918);
nor U5843 (N_5843,N_1489,N_4563);
nand U5844 (N_5844,N_373,N_3780);
and U5845 (N_5845,N_678,N_4444);
and U5846 (N_5846,N_4460,N_220);
nor U5847 (N_5847,N_2372,N_1135);
nand U5848 (N_5848,N_360,N_4152);
or U5849 (N_5849,N_130,N_1360);
xnor U5850 (N_5850,N_3976,N_3055);
nand U5851 (N_5851,N_3397,N_4309);
nor U5852 (N_5852,N_2501,N_1063);
nor U5853 (N_5853,N_4744,N_4968);
and U5854 (N_5854,N_2751,N_4904);
xnor U5855 (N_5855,N_288,N_2348);
and U5856 (N_5856,N_613,N_2441);
and U5857 (N_5857,N_4907,N_4315);
xnor U5858 (N_5858,N_1091,N_2614);
nor U5859 (N_5859,N_1264,N_3315);
nor U5860 (N_5860,N_3149,N_2460);
xnor U5861 (N_5861,N_888,N_1834);
nor U5862 (N_5862,N_1543,N_2837);
nor U5863 (N_5863,N_802,N_1033);
xor U5864 (N_5864,N_2187,N_4293);
xor U5865 (N_5865,N_4288,N_1636);
nand U5866 (N_5866,N_1962,N_2400);
or U5867 (N_5867,N_3539,N_1222);
and U5868 (N_5868,N_2624,N_1142);
or U5869 (N_5869,N_2228,N_4110);
and U5870 (N_5870,N_2106,N_4337);
xnor U5871 (N_5871,N_4718,N_4133);
nand U5872 (N_5872,N_1083,N_1548);
xor U5873 (N_5873,N_2720,N_2427);
nor U5874 (N_5874,N_4802,N_3727);
xnor U5875 (N_5875,N_767,N_2180);
xnor U5876 (N_5876,N_4906,N_361);
nand U5877 (N_5877,N_889,N_4654);
nand U5878 (N_5878,N_1138,N_3147);
xor U5879 (N_5879,N_2702,N_521);
nand U5880 (N_5880,N_536,N_2244);
nor U5881 (N_5881,N_1004,N_1733);
nor U5882 (N_5882,N_913,N_1841);
and U5883 (N_5883,N_3158,N_1918);
and U5884 (N_5884,N_440,N_4701);
and U5885 (N_5885,N_3616,N_20);
or U5886 (N_5886,N_1937,N_4952);
and U5887 (N_5887,N_3553,N_4890);
and U5888 (N_5888,N_3881,N_2081);
nor U5889 (N_5889,N_78,N_3939);
nor U5890 (N_5890,N_2116,N_2047);
or U5891 (N_5891,N_4499,N_1673);
and U5892 (N_5892,N_4655,N_4515);
and U5893 (N_5893,N_534,N_572);
and U5894 (N_5894,N_2764,N_4164);
or U5895 (N_5895,N_2885,N_3957);
nor U5896 (N_5896,N_4156,N_4859);
nand U5897 (N_5897,N_740,N_3450);
and U5898 (N_5898,N_2695,N_4167);
or U5899 (N_5899,N_591,N_70);
nand U5900 (N_5900,N_2189,N_3799);
xor U5901 (N_5901,N_3817,N_4142);
and U5902 (N_5902,N_789,N_4248);
and U5903 (N_5903,N_4189,N_3195);
and U5904 (N_5904,N_2287,N_2580);
and U5905 (N_5905,N_119,N_2599);
nand U5906 (N_5906,N_2342,N_2093);
and U5907 (N_5907,N_1875,N_2535);
and U5908 (N_5908,N_2239,N_542);
nand U5909 (N_5909,N_541,N_1257);
xnor U5910 (N_5910,N_2179,N_4097);
xor U5911 (N_5911,N_1321,N_1872);
nor U5912 (N_5912,N_3034,N_2896);
nor U5913 (N_5913,N_2785,N_4670);
and U5914 (N_5914,N_2709,N_2011);
or U5915 (N_5915,N_2176,N_320);
nand U5916 (N_5916,N_2780,N_2877);
nand U5917 (N_5917,N_4096,N_4263);
and U5918 (N_5918,N_589,N_2343);
or U5919 (N_5919,N_511,N_4652);
or U5920 (N_5920,N_2371,N_2221);
nand U5921 (N_5921,N_2601,N_4069);
nand U5922 (N_5922,N_4835,N_1285);
nand U5923 (N_5923,N_2503,N_2398);
nand U5924 (N_5924,N_3107,N_2280);
and U5925 (N_5925,N_140,N_3802);
nand U5926 (N_5926,N_3833,N_266);
and U5927 (N_5927,N_2012,N_3811);
and U5928 (N_5928,N_3303,N_818);
and U5929 (N_5929,N_3932,N_3922);
or U5930 (N_5930,N_868,N_4493);
nor U5931 (N_5931,N_3590,N_575);
xor U5932 (N_5932,N_939,N_4812);
and U5933 (N_5933,N_1,N_4346);
xnor U5934 (N_5934,N_3109,N_4155);
xnor U5935 (N_5935,N_4550,N_4265);
nor U5936 (N_5936,N_4592,N_4531);
or U5937 (N_5937,N_2076,N_3360);
or U5938 (N_5938,N_1362,N_2424);
or U5939 (N_5939,N_1562,N_3294);
or U5940 (N_5940,N_4371,N_39);
or U5941 (N_5941,N_4545,N_525);
or U5942 (N_5942,N_3634,N_946);
or U5943 (N_5943,N_1406,N_4179);
nor U5944 (N_5944,N_4933,N_1840);
nand U5945 (N_5945,N_2240,N_1695);
or U5946 (N_5946,N_3018,N_4684);
nand U5947 (N_5947,N_3600,N_1148);
or U5948 (N_5948,N_4345,N_1686);
or U5949 (N_5949,N_4543,N_893);
nor U5950 (N_5950,N_2662,N_1927);
xnor U5951 (N_5951,N_3342,N_2297);
nor U5952 (N_5952,N_232,N_3872);
xor U5953 (N_5953,N_1906,N_2687);
nand U5954 (N_5954,N_3380,N_1326);
or U5955 (N_5955,N_1647,N_1144);
nor U5956 (N_5956,N_1065,N_1730);
xor U5957 (N_5957,N_1231,N_3532);
xnor U5958 (N_5958,N_91,N_1433);
or U5959 (N_5959,N_1503,N_3392);
xnor U5960 (N_5960,N_1662,N_3215);
nand U5961 (N_5961,N_3021,N_2631);
or U5962 (N_5962,N_1109,N_557);
or U5963 (N_5963,N_1312,N_1584);
nor U5964 (N_5964,N_683,N_1828);
and U5965 (N_5965,N_334,N_2197);
nand U5966 (N_5966,N_2971,N_2406);
xnor U5967 (N_5967,N_4347,N_2674);
nand U5968 (N_5968,N_1878,N_4741);
or U5969 (N_5969,N_4500,N_3036);
xor U5970 (N_5970,N_4816,N_2273);
and U5971 (N_5971,N_127,N_414);
or U5972 (N_5972,N_4940,N_4513);
or U5973 (N_5973,N_221,N_4254);
nor U5974 (N_5974,N_162,N_2205);
xnor U5975 (N_5975,N_4047,N_1128);
nor U5976 (N_5976,N_4782,N_4803);
xnor U5977 (N_5977,N_4223,N_652);
nand U5978 (N_5978,N_3169,N_3132);
or U5979 (N_5979,N_1024,N_4596);
nand U5980 (N_5980,N_2167,N_1570);
nor U5981 (N_5981,N_4151,N_1812);
or U5982 (N_5982,N_1352,N_2845);
nand U5983 (N_5983,N_1905,N_3264);
and U5984 (N_5984,N_3578,N_1215);
nor U5985 (N_5985,N_4431,N_1358);
nand U5986 (N_5986,N_3287,N_1765);
and U5987 (N_5987,N_960,N_3775);
nor U5988 (N_5988,N_4296,N_4929);
xnor U5989 (N_5989,N_1909,N_245);
or U5990 (N_5990,N_3598,N_2967);
nor U5991 (N_5991,N_597,N_3879);
or U5992 (N_5992,N_4294,N_116);
xor U5993 (N_5993,N_3097,N_4547);
xnor U5994 (N_5994,N_1682,N_3341);
xnor U5995 (N_5995,N_4159,N_3014);
or U5996 (N_5996,N_406,N_4124);
xor U5997 (N_5997,N_3006,N_3116);
and U5998 (N_5998,N_3620,N_505);
and U5999 (N_5999,N_2786,N_3378);
nor U6000 (N_6000,N_2725,N_2714);
nand U6001 (N_6001,N_4430,N_2214);
xnor U6002 (N_6002,N_3946,N_2556);
nand U6003 (N_6003,N_202,N_1299);
and U6004 (N_6004,N_4369,N_4864);
nand U6005 (N_6005,N_2586,N_2968);
xor U6006 (N_6006,N_3114,N_1247);
nor U6007 (N_6007,N_2065,N_3190);
xor U6008 (N_6008,N_2322,N_773);
xor U6009 (N_6009,N_3292,N_681);
nor U6010 (N_6010,N_1881,N_3177);
xor U6011 (N_6011,N_3708,N_4283);
nor U6012 (N_6012,N_3585,N_3490);
nand U6013 (N_6013,N_126,N_1438);
or U6014 (N_6014,N_4188,N_1760);
xor U6015 (N_6015,N_4849,N_3975);
nor U6016 (N_6016,N_717,N_4785);
nor U6017 (N_6017,N_1798,N_1383);
and U6018 (N_6018,N_2534,N_2609);
nand U6019 (N_6019,N_2020,N_1364);
nand U6020 (N_6020,N_54,N_1053);
nand U6021 (N_6021,N_2377,N_1155);
nor U6022 (N_6022,N_1628,N_1680);
xnor U6023 (N_6023,N_4969,N_2880);
or U6024 (N_6024,N_3613,N_2313);
or U6025 (N_6025,N_4236,N_1400);
and U6026 (N_6026,N_3652,N_4843);
nor U6027 (N_6027,N_1459,N_3618);
or U6028 (N_6028,N_3859,N_2224);
nor U6029 (N_6029,N_2667,N_2366);
or U6030 (N_6030,N_4298,N_3838);
nand U6031 (N_6031,N_3205,N_3267);
nand U6032 (N_6032,N_2469,N_4814);
and U6033 (N_6033,N_1852,N_4285);
nor U6034 (N_6034,N_2694,N_2560);
nand U6035 (N_6035,N_3789,N_3912);
nand U6036 (N_6036,N_4228,N_831);
nand U6037 (N_6037,N_1566,N_4902);
nand U6038 (N_6038,N_2758,N_3347);
xor U6039 (N_6039,N_4396,N_4454);
xnor U6040 (N_6040,N_2860,N_3140);
nand U6041 (N_6041,N_3176,N_2025);
nand U6042 (N_6042,N_2912,N_2223);
or U6043 (N_6043,N_3506,N_2925);
nor U6044 (N_6044,N_2438,N_4405);
xnor U6045 (N_6045,N_3683,N_2781);
nand U6046 (N_6046,N_1508,N_2457);
and U6047 (N_6047,N_2281,N_3090);
nand U6048 (N_6048,N_3338,N_808);
or U6049 (N_6049,N_3128,N_803);
or U6050 (N_6050,N_1801,N_3980);
xor U6051 (N_6051,N_4040,N_137);
or U6052 (N_6052,N_634,N_4413);
nand U6053 (N_6053,N_3302,N_2564);
xor U6054 (N_6054,N_1581,N_3033);
xor U6055 (N_6055,N_909,N_1972);
nand U6056 (N_6056,N_983,N_3129);
nand U6057 (N_6057,N_3429,N_4985);
or U6058 (N_6058,N_2051,N_375);
xor U6059 (N_6059,N_1550,N_2596);
xor U6060 (N_6060,N_1921,N_3732);
nand U6061 (N_6061,N_4851,N_2350);
nand U6062 (N_6062,N_2431,N_769);
nand U6063 (N_6063,N_263,N_409);
nor U6064 (N_6064,N_151,N_3222);
nor U6065 (N_6065,N_3106,N_3908);
xor U6066 (N_6066,N_729,N_3722);
or U6067 (N_6067,N_189,N_4815);
nand U6068 (N_6068,N_3546,N_550);
or U6069 (N_6069,N_3954,N_2903);
or U6070 (N_6070,N_3078,N_1605);
nor U6071 (N_6071,N_1512,N_4787);
and U6072 (N_6072,N_3057,N_2101);
nor U6073 (N_6073,N_1216,N_1991);
nor U6074 (N_6074,N_4894,N_2743);
and U6075 (N_6075,N_2257,N_4004);
nor U6076 (N_6076,N_1073,N_3091);
nor U6077 (N_6077,N_1998,N_929);
or U6078 (N_6078,N_2634,N_1179);
or U6079 (N_6079,N_2569,N_3247);
or U6080 (N_6080,N_3276,N_3224);
xor U6081 (N_6081,N_922,N_1871);
and U6082 (N_6082,N_4799,N_543);
or U6083 (N_6083,N_3050,N_2474);
nand U6084 (N_6084,N_3698,N_4329);
nor U6085 (N_6085,N_2777,N_4754);
or U6086 (N_6086,N_3801,N_3990);
or U6087 (N_6087,N_3291,N_143);
or U6088 (N_6088,N_268,N_4764);
and U6089 (N_6089,N_3894,N_1577);
nor U6090 (N_6090,N_2514,N_2920);
nor U6091 (N_6091,N_860,N_1728);
xnor U6092 (N_6092,N_963,N_1849);
xnor U6093 (N_6093,N_4160,N_757);
nand U6094 (N_6094,N_3488,N_2739);
and U6095 (N_6095,N_4731,N_4522);
and U6096 (N_6096,N_464,N_1787);
nor U6097 (N_6097,N_3295,N_859);
or U6098 (N_6098,N_661,N_4566);
nand U6099 (N_6099,N_2166,N_2610);
nor U6100 (N_6100,N_753,N_1668);
nand U6101 (N_6101,N_1870,N_665);
and U6102 (N_6102,N_3530,N_3914);
and U6103 (N_6103,N_924,N_4355);
xor U6104 (N_6104,N_3290,N_331);
or U6105 (N_6105,N_2165,N_1756);
nand U6106 (N_6106,N_2078,N_3569);
xor U6107 (N_6107,N_493,N_627);
xnor U6108 (N_6108,N_1002,N_1249);
and U6109 (N_6109,N_1369,N_3576);
nor U6110 (N_6110,N_4412,N_3629);
nand U6111 (N_6111,N_3650,N_1045);
and U6112 (N_6112,N_3187,N_1565);
nor U6113 (N_6113,N_4224,N_1464);
xnor U6114 (N_6114,N_254,N_1924);
xnor U6115 (N_6115,N_2038,N_3089);
nand U6116 (N_6116,N_3782,N_640);
nand U6117 (N_6117,N_1726,N_2559);
xor U6118 (N_6118,N_2033,N_538);
xnor U6119 (N_6119,N_4604,N_439);
nand U6120 (N_6120,N_2990,N_830);
and U6121 (N_6121,N_3969,N_2684);
xor U6122 (N_6122,N_1617,N_1208);
or U6123 (N_6123,N_3104,N_4443);
and U6124 (N_6124,N_1623,N_2048);
nand U6125 (N_6125,N_1363,N_2383);
or U6126 (N_6126,N_2339,N_3538);
and U6127 (N_6127,N_4456,N_2331);
nor U6128 (N_6128,N_3560,N_1297);
nor U6129 (N_6129,N_3854,N_2740);
xor U6130 (N_6130,N_1146,N_3988);
and U6131 (N_6131,N_4875,N_1015);
nand U6132 (N_6132,N_3570,N_1965);
xor U6133 (N_6133,N_4648,N_2549);
or U6134 (N_6134,N_1424,N_1279);
or U6135 (N_6135,N_164,N_4572);
nand U6136 (N_6136,N_4910,N_1259);
nor U6137 (N_6137,N_3527,N_721);
xor U6138 (N_6138,N_1559,N_4791);
xnor U6139 (N_6139,N_2242,N_187);
nand U6140 (N_6140,N_1068,N_1311);
or U6141 (N_6141,N_3367,N_911);
nor U6142 (N_6142,N_1823,N_4278);
nand U6143 (N_6143,N_2508,N_3526);
and U6144 (N_6144,N_1041,N_1420);
xor U6145 (N_6145,N_906,N_3318);
or U6146 (N_6146,N_2716,N_390);
or U6147 (N_6147,N_2519,N_4029);
or U6148 (N_6148,N_4707,N_465);
or U6149 (N_6149,N_4730,N_1832);
nand U6150 (N_6150,N_225,N_1335);
xnor U6151 (N_6151,N_2874,N_4095);
or U6152 (N_6152,N_4031,N_3561);
nor U6153 (N_6153,N_2576,N_2461);
nand U6154 (N_6154,N_1440,N_3084);
nor U6155 (N_6155,N_1226,N_4689);
and U6156 (N_6156,N_755,N_2208);
nand U6157 (N_6157,N_1530,N_2545);
nand U6158 (N_6158,N_2137,N_3931);
and U6159 (N_6159,N_3039,N_374);
nand U6160 (N_6160,N_3717,N_4974);
and U6161 (N_6161,N_1100,N_3902);
or U6162 (N_6162,N_1269,N_115);
and U6163 (N_6163,N_761,N_3860);
nand U6164 (N_6164,N_689,N_3533);
and U6165 (N_6165,N_826,N_2807);
nand U6166 (N_6166,N_3407,N_4866);
xnor U6167 (N_6167,N_3130,N_181);
xor U6168 (N_6168,N_3895,N_3809);
and U6169 (N_6169,N_186,N_1588);
nor U6170 (N_6170,N_2198,N_31);
xor U6171 (N_6171,N_4138,N_2053);
or U6172 (N_6172,N_2103,N_355);
and U6173 (N_6173,N_3899,N_351);
nand U6174 (N_6174,N_2805,N_1720);
and U6175 (N_6175,N_1754,N_247);
nand U6176 (N_6176,N_3393,N_4023);
or U6177 (N_6177,N_633,N_58);
or U6178 (N_6178,N_1290,N_4195);
xor U6179 (N_6179,N_4313,N_229);
xnor U6180 (N_6180,N_2411,N_2285);
nor U6181 (N_6181,N_4414,N_2192);
nor U6182 (N_6182,N_96,N_43);
or U6183 (N_6183,N_52,N_2620);
nand U6184 (N_6184,N_2509,N_2462);
and U6185 (N_6185,N_1164,N_707);
nand U6186 (N_6186,N_4358,N_2911);
and U6187 (N_6187,N_920,N_1468);
nor U6188 (N_6188,N_972,N_1693);
and U6189 (N_6189,N_3146,N_2068);
or U6190 (N_6190,N_1427,N_1012);
or U6191 (N_6191,N_2918,N_3593);
nor U6192 (N_6192,N_866,N_2154);
or U6193 (N_6193,N_1380,N_4944);
and U6194 (N_6194,N_4813,N_1757);
and U6195 (N_6195,N_3358,N_1978);
xor U6196 (N_6196,N_3588,N_1137);
nand U6197 (N_6197,N_1436,N_1404);
and U6198 (N_6198,N_1327,N_4084);
nor U6199 (N_6199,N_4595,N_250);
nand U6200 (N_6200,N_4469,N_1684);
or U6201 (N_6201,N_2588,N_4765);
nand U6202 (N_6202,N_2336,N_770);
nor U6203 (N_6203,N_4432,N_3363);
and U6204 (N_6204,N_3978,N_786);
or U6205 (N_6205,N_518,N_3550);
and U6206 (N_6206,N_1225,N_110);
and U6207 (N_6207,N_3122,N_3103);
xnor U6208 (N_6208,N_2506,N_1791);
and U6209 (N_6209,N_3298,N_2817);
and U6210 (N_6210,N_1482,N_4045);
xnor U6211 (N_6211,N_4286,N_4185);
and U6212 (N_6212,N_654,N_2413);
nand U6213 (N_6213,N_3835,N_4722);
or U6214 (N_6214,N_2704,N_605);
nand U6215 (N_6215,N_743,N_3225);
or U6216 (N_6216,N_1869,N_4478);
nand U6217 (N_6217,N_1749,N_3864);
and U6218 (N_6218,N_2328,N_3063);
nand U6219 (N_6219,N_3313,N_705);
or U6220 (N_6220,N_4823,N_2027);
xnor U6221 (N_6221,N_1271,N_45);
xor U6222 (N_6222,N_207,N_950);
nand U6223 (N_6223,N_2102,N_1417);
xor U6224 (N_6224,N_200,N_198);
nand U6225 (N_6225,N_4924,N_4416);
and U6226 (N_6226,N_3399,N_2333);
nor U6227 (N_6227,N_1057,N_3766);
xor U6228 (N_6228,N_3234,N_3471);
nand U6229 (N_6229,N_3562,N_877);
nand U6230 (N_6230,N_86,N_2963);
xor U6231 (N_6231,N_4453,N_4757);
or U6232 (N_6232,N_2404,N_2039);
or U6233 (N_6233,N_943,N_2772);
or U6234 (N_6234,N_4458,N_3876);
nor U6235 (N_6235,N_1994,N_3012);
xnor U6236 (N_6236,N_664,N_957);
xnor U6237 (N_6237,N_444,N_63);
nand U6238 (N_6238,N_2477,N_3306);
nand U6239 (N_6239,N_3925,N_1432);
xor U6240 (N_6240,N_3750,N_520);
xnor U6241 (N_6241,N_150,N_483);
nand U6242 (N_6242,N_3351,N_4153);
nand U6243 (N_6243,N_2459,N_4523);
xnor U6244 (N_6244,N_1298,N_1624);
nand U6245 (N_6245,N_2653,N_3305);
and U6246 (N_6246,N_1240,N_655);
or U6247 (N_6247,N_3453,N_3748);
nand U6248 (N_6248,N_4007,N_4199);
and U6249 (N_6249,N_546,N_389);
or U6250 (N_6250,N_625,N_1183);
and U6251 (N_6251,N_1496,N_3003);
nand U6252 (N_6252,N_3017,N_1104);
or U6253 (N_6253,N_1657,N_1561);
nor U6254 (N_6254,N_4709,N_3964);
and U6255 (N_6255,N_3101,N_2355);
nand U6256 (N_6256,N_3826,N_4101);
nor U6257 (N_6257,N_3059,N_996);
or U6258 (N_6258,N_65,N_3672);
or U6259 (N_6259,N_2183,N_3543);
and U6260 (N_6260,N_604,N_4934);
nor U6261 (N_6261,N_2941,N_4742);
nor U6262 (N_6262,N_3307,N_1054);
or U6263 (N_6263,N_4186,N_3688);
nand U6264 (N_6264,N_1295,N_4310);
xor U6265 (N_6265,N_161,N_2908);
nand U6266 (N_6266,N_2489,N_74);
nand U6267 (N_6267,N_447,N_3726);
xor U6268 (N_6268,N_4440,N_3958);
xnor U6269 (N_6269,N_781,N_2256);
and U6270 (N_6270,N_1650,N_2426);
nor U6271 (N_6271,N_362,N_3606);
and U6272 (N_6272,N_174,N_3979);
and U6273 (N_6273,N_1592,N_3923);
xnor U6274 (N_6274,N_4165,N_2304);
nand U6275 (N_6275,N_2808,N_697);
nand U6276 (N_6276,N_3963,N_3242);
xor U6277 (N_6277,N_4534,N_4733);
or U6278 (N_6278,N_4525,N_3611);
xnor U6279 (N_6279,N_3535,N_1007);
nor U6280 (N_6280,N_3919,N_2058);
nand U6281 (N_6281,N_688,N_2184);
nor U6282 (N_6282,N_3500,N_1838);
or U6283 (N_6283,N_3970,N_1639);
or U6284 (N_6284,N_4530,N_231);
or U6285 (N_6285,N_3345,N_1318);
or U6286 (N_6286,N_4392,N_2498);
nor U6287 (N_6287,N_399,N_2746);
and U6288 (N_6288,N_324,N_3938);
or U6289 (N_6289,N_944,N_2706);
nor U6290 (N_6290,N_1228,N_1868);
and U6291 (N_6291,N_1712,N_122);
and U6292 (N_6292,N_1047,N_872);
or U6293 (N_6293,N_253,N_1339);
xnor U6294 (N_6294,N_3493,N_2253);
and U6295 (N_6295,N_4610,N_2007);
or U6296 (N_6296,N_3250,N_2681);
xor U6297 (N_6297,N_1973,N_1957);
and U6298 (N_6298,N_4391,N_11);
and U6299 (N_6299,N_4524,N_1044);
nor U6300 (N_6300,N_886,N_3666);
and U6301 (N_6301,N_1113,N_884);
and U6302 (N_6302,N_4957,N_1843);
and U6303 (N_6303,N_1932,N_2089);
or U6304 (N_6304,N_961,N_1461);
nand U6305 (N_6305,N_3929,N_4422);
and U6306 (N_6306,N_3296,N_1480);
xor U6307 (N_6307,N_1416,N_2254);
nor U6308 (N_6308,N_2237,N_4301);
nand U6309 (N_6309,N_3761,N_4692);
nor U6310 (N_6310,N_2439,N_2337);
xor U6311 (N_6311,N_2637,N_62);
nand U6312 (N_6312,N_1520,N_1370);
nor U6313 (N_6313,N_2249,N_4943);
nand U6314 (N_6314,N_1964,N_2878);
and U6315 (N_6315,N_1453,N_4998);
or U6316 (N_6316,N_650,N_142);
xor U6317 (N_6317,N_1860,N_1889);
and U6318 (N_6318,N_2897,N_2678);
nand U6319 (N_6319,N_346,N_3326);
nor U6320 (N_6320,N_1514,N_269);
xor U6321 (N_6321,N_1217,N_1175);
nor U6322 (N_6322,N_2274,N_2269);
and U6323 (N_6323,N_4611,N_3556);
and U6324 (N_6324,N_4840,N_2235);
nand U6325 (N_6325,N_1426,N_870);
or U6326 (N_6326,N_3469,N_1402);
or U6327 (N_6327,N_2840,N_2745);
nand U6328 (N_6328,N_4927,N_2127);
xor U6329 (N_6329,N_4465,N_4131);
xor U6330 (N_6330,N_2533,N_2870);
nand U6331 (N_6331,N_4516,N_4579);
nor U6332 (N_6332,N_2950,N_1706);
nand U6333 (N_6333,N_4320,N_480);
and U6334 (N_6334,N_3605,N_2389);
nand U6335 (N_6335,N_275,N_4990);
nor U6336 (N_6336,N_971,N_4817);
and U6337 (N_6337,N_2558,N_1850);
or U6338 (N_6338,N_745,N_3212);
xnor U6339 (N_6339,N_853,N_519);
nor U6340 (N_6340,N_3935,N_4922);
nor U6341 (N_6341,N_1681,N_660);
and U6342 (N_6342,N_3509,N_1340);
or U6343 (N_6343,N_1721,N_3563);
nor U6344 (N_6344,N_4451,N_501);
xor U6345 (N_6345,N_4093,N_2578);
or U6346 (N_6346,N_2067,N_1724);
nor U6347 (N_6347,N_27,N_4333);
or U6348 (N_6348,N_4409,N_3330);
nor U6349 (N_6349,N_962,N_2997);
nor U6350 (N_6350,N_3567,N_1112);
nand U6351 (N_6351,N_2976,N_1784);
nand U6352 (N_6352,N_4753,N_4783);
nand U6353 (N_6353,N_2883,N_4452);
or U6354 (N_6354,N_322,N_508);
nand U6355 (N_6355,N_3785,N_2822);
and U6356 (N_6356,N_2134,N_3121);
nand U6357 (N_6357,N_2050,N_235);
or U6358 (N_6358,N_4035,N_3641);
nand U6359 (N_6359,N_1333,N_3333);
nor U6360 (N_6360,N_1088,N_4909);
xor U6361 (N_6361,N_6,N_1655);
and U6362 (N_6362,N_3991,N_3213);
xnor U6363 (N_6363,N_4247,N_4100);
and U6364 (N_6364,N_1190,N_4553);
nor U6365 (N_6365,N_2670,N_1880);
or U6366 (N_6366,N_3889,N_1737);
nor U6367 (N_6367,N_4642,N_124);
and U6368 (N_6368,N_3243,N_4311);
nand U6369 (N_6369,N_4178,N_146);
xnor U6370 (N_6370,N_711,N_3076);
or U6371 (N_6371,N_3216,N_4533);
nand U6372 (N_6372,N_1020,N_475);
nor U6373 (N_6373,N_2218,N_1926);
and U6374 (N_6374,N_378,N_4569);
and U6375 (N_6375,N_3883,N_1916);
xor U6376 (N_6376,N_980,N_34);
xnor U6377 (N_6377,N_1755,N_3426);
xnor U6378 (N_6378,N_4025,N_2408);
nand U6379 (N_6379,N_1781,N_1001);
and U6380 (N_6380,N_3577,N_2029);
xnor U6381 (N_6381,N_3051,N_672);
and U6382 (N_6382,N_429,N_4242);
and U6383 (N_6383,N_4877,N_1292);
and U6384 (N_6384,N_2550,N_2995);
nand U6385 (N_6385,N_1320,N_467);
and U6386 (N_6386,N_1600,N_4989);
nand U6387 (N_6387,N_191,N_341);
nand U6388 (N_6388,N_2483,N_1181);
nor U6389 (N_6389,N_4873,N_3622);
nor U6390 (N_6390,N_1462,N_176);
nor U6391 (N_6391,N_2721,N_1027);
or U6392 (N_6392,N_517,N_3955);
nand U6393 (N_6393,N_64,N_2668);
nand U6394 (N_6394,N_3624,N_4719);
and U6395 (N_6395,N_3462,N_1365);
and U6396 (N_6396,N_3402,N_2353);
nor U6397 (N_6397,N_196,N_2113);
nor U6398 (N_6398,N_4240,N_2082);
and U6399 (N_6399,N_3278,N_1492);
or U6400 (N_6400,N_2437,N_2686);
nor U6401 (N_6401,N_1958,N_4861);
nand U6402 (N_6402,N_3837,N_1397);
and U6403 (N_6403,N_788,N_1016);
xor U6404 (N_6404,N_713,N_2747);
and U6405 (N_6405,N_3119,N_2016);
or U6406 (N_6406,N_1111,N_4656);
and U6407 (N_6407,N_2679,N_2803);
nand U6408 (N_6408,N_2954,N_1415);
nor U6409 (N_6409,N_1218,N_2402);
nor U6410 (N_6410,N_3831,N_4106);
xor U6411 (N_6411,N_2401,N_4967);
or U6412 (N_6412,N_3480,N_3417);
xor U6413 (N_6413,N_3791,N_1586);
nor U6414 (N_6414,N_2655,N_4330);
xor U6415 (N_6415,N_676,N_2737);
nand U6416 (N_6416,N_168,N_1831);
nor U6417 (N_6417,N_3203,N_4581);
and U6418 (N_6418,N_1752,N_4486);
nand U6419 (N_6419,N_2927,N_2540);
xnor U6420 (N_6420,N_2515,N_448);
and U6421 (N_6421,N_1576,N_3442);
or U6422 (N_6422,N_694,N_3999);
or U6423 (N_6423,N_2994,N_3428);
nand U6424 (N_6424,N_4427,N_2642);
and U6425 (N_6425,N_1470,N_255);
nor U6426 (N_6426,N_4565,N_1418);
and U6427 (N_6427,N_4732,N_592);
xnor U6428 (N_6428,N_2286,N_4582);
nor U6429 (N_6429,N_2524,N_4872);
nor U6430 (N_6430,N_1727,N_3334);
nand U6431 (N_6431,N_4198,N_3478);
xor U6432 (N_6432,N_2488,N_4977);
xor U6433 (N_6433,N_1643,N_4380);
xnor U6434 (N_6434,N_1997,N_4437);
nor U6435 (N_6435,N_3729,N_182);
nor U6436 (N_6436,N_4235,N_3387);
nor U6437 (N_6437,N_4227,N_965);
nand U6438 (N_6438,N_4978,N_704);
xor U6439 (N_6439,N_1023,N_89);
nand U6440 (N_6440,N_2467,N_421);
xor U6441 (N_6441,N_2592,N_72);
and U6442 (N_6442,N_1167,N_3812);
xor U6443 (N_6443,N_3793,N_241);
or U6444 (N_6444,N_1553,N_2397);
and U6445 (N_6445,N_3013,N_3626);
xor U6446 (N_6446,N_4241,N_3438);
and U6447 (N_6447,N_1207,N_4663);
nand U6448 (N_6448,N_1230,N_2186);
nor U6449 (N_6449,N_4368,N_4092);
or U6450 (N_6450,N_210,N_1574);
or U6451 (N_6451,N_1569,N_3832);
nor U6452 (N_6452,N_1430,N_2142);
and U6453 (N_6453,N_3856,N_1556);
nor U6454 (N_6454,N_3337,N_750);
or U6455 (N_6455,N_471,N_1813);
nor U6456 (N_6456,N_97,N_2893);
or U6457 (N_6457,N_120,N_1734);
xnor U6458 (N_6458,N_3191,N_2922);
nor U6459 (N_6459,N_4796,N_3940);
nand U6460 (N_6460,N_4402,N_3738);
and U6461 (N_6461,N_2112,N_1824);
xor U6462 (N_6462,N_3235,N_3820);
nor U6463 (N_6463,N_2986,N_4601);
or U6464 (N_6464,N_737,N_1910);
or U6465 (N_6465,N_2972,N_3678);
xor U6466 (N_6466,N_3644,N_2497);
xor U6467 (N_6467,N_3144,N_1626);
xnor U6468 (N_6468,N_2965,N_156);
xnor U6469 (N_6469,N_1934,N_2066);
nor U6470 (N_6470,N_2907,N_2155);
xor U6471 (N_6471,N_3435,N_2122);
nor U6472 (N_6472,N_2213,N_3052);
nor U6473 (N_6473,N_1947,N_3067);
nand U6474 (N_6474,N_4950,N_2494);
or U6475 (N_6475,N_4672,N_2529);
and U6476 (N_6476,N_2776,N_4936);
or U6477 (N_6477,N_3920,N_3259);
nand U6478 (N_6478,N_4210,N_2299);
or U6479 (N_6479,N_4972,N_4183);
nand U6480 (N_6480,N_3580,N_629);
nand U6481 (N_6481,N_442,N_468);
or U6482 (N_6482,N_2448,N_264);
and U6483 (N_6483,N_1587,N_4954);
nand U6484 (N_6484,N_3460,N_57);
or U6485 (N_6485,N_656,N_1745);
or U6486 (N_6486,N_715,N_3433);
nand U6487 (N_6487,N_1914,N_611);
nand U6488 (N_6488,N_2442,N_857);
and U6489 (N_6489,N_195,N_4370);
and U6490 (N_6490,N_4850,N_2135);
nand U6491 (N_6491,N_1563,N_3930);
nor U6492 (N_6492,N_3143,N_4340);
nand U6493 (N_6493,N_4598,N_1546);
nand U6494 (N_6494,N_2823,N_1718);
or U6495 (N_6495,N_4738,N_3744);
and U6496 (N_6496,N_4328,N_1147);
nor U6497 (N_6497,N_4316,N_30);
nor U6498 (N_6498,N_4912,N_1306);
nor U6499 (N_6499,N_4607,N_35);
nor U6500 (N_6500,N_3523,N_4144);
nor U6501 (N_6501,N_2490,N_1329);
nand U6502 (N_6502,N_3319,N_1345);
nor U6503 (N_6503,N_1193,N_4118);
nor U6504 (N_6504,N_1672,N_2665);
nor U6505 (N_6505,N_1081,N_867);
nand U6506 (N_6506,N_4549,N_4838);
nor U6507 (N_6507,N_1233,N_3382);
nor U6508 (N_6508,N_3494,N_3951);
nand U6509 (N_6509,N_4881,N_3074);
nor U6510 (N_6510,N_3891,N_4483);
nor U6511 (N_6511,N_4064,N_4181);
nand U6512 (N_6512,N_2742,N_2340);
or U6513 (N_6513,N_3599,N_1095);
nor U6514 (N_6514,N_1886,N_98);
or U6515 (N_6515,N_4520,N_1819);
and U6516 (N_6516,N_1996,N_643);
and U6517 (N_6517,N_2603,N_2854);
and U6518 (N_6518,N_285,N_3073);
xnor U6519 (N_6519,N_1026,N_758);
xnor U6520 (N_6520,N_2062,N_2938);
nand U6521 (N_6521,N_584,N_608);
or U6522 (N_6522,N_265,N_4767);
xor U6523 (N_6523,N_2671,N_3815);
nand U6524 (N_6524,N_948,N_2909);
xor U6525 (N_6525,N_616,N_2396);
and U6526 (N_6526,N_1134,N_2233);
or U6527 (N_6527,N_3781,N_2731);
nand U6528 (N_6528,N_4094,N_183);
or U6529 (N_6529,N_2646,N_4631);
and U6530 (N_6530,N_1210,N_1883);
nor U6531 (N_6531,N_420,N_1080);
nand U6532 (N_6532,N_1573,N_208);
nor U6533 (N_6533,N_2330,N_339);
nand U6534 (N_6534,N_858,N_2750);
and U6535 (N_6535,N_3204,N_999);
xnor U6536 (N_6536,N_692,N_772);
nor U6537 (N_6537,N_4641,N_4682);
or U6538 (N_6538,N_4423,N_4557);
nand U6539 (N_6539,N_510,N_2917);
or U6540 (N_6540,N_4665,N_2321);
nor U6541 (N_6541,N_2700,N_4099);
nand U6542 (N_6542,N_3157,N_582);
and U6543 (N_6543,N_2259,N_1555);
or U6544 (N_6544,N_1114,N_369);
xor U6545 (N_6545,N_1450,N_1077);
and U6546 (N_6546,N_3086,N_3245);
or U6547 (N_6547,N_2450,N_4287);
nand U6548 (N_6548,N_3210,N_2294);
or U6549 (N_6549,N_4253,N_3316);
nand U6550 (N_6550,N_4804,N_80);
nor U6551 (N_6551,N_3446,N_2487);
or U6552 (N_6552,N_4268,N_1688);
nor U6553 (N_6553,N_3454,N_1862);
and U6554 (N_6554,N_3362,N_4258);
nand U6555 (N_6555,N_3637,N_3427);
nand U6556 (N_6556,N_1141,N_4997);
nand U6557 (N_6557,N_3507,N_2861);
or U6558 (N_6558,N_899,N_4335);
and U6559 (N_6559,N_3586,N_3853);
or U6560 (N_6560,N_567,N_4649);
nor U6561 (N_6561,N_4697,N_4973);
nor U6562 (N_6562,N_4448,N_4878);
xnor U6563 (N_6563,N_4065,N_308);
or U6564 (N_6564,N_171,N_801);
nand U6565 (N_6565,N_2582,N_1059);
and U6566 (N_6566,N_2199,N_3607);
xor U6567 (N_6567,N_2055,N_4009);
nand U6568 (N_6568,N_2710,N_615);
nand U6569 (N_6569,N_4762,N_3961);
xor U6570 (N_6570,N_1280,N_4488);
and U6571 (N_6571,N_865,N_2399);
and U6572 (N_6572,N_3273,N_2300);
nor U6573 (N_6573,N_2654,N_1552);
xnor U6574 (N_6574,N_2182,N_484);
nor U6575 (N_6575,N_4056,N_3099);
or U6576 (N_6576,N_3575,N_790);
xnor U6577 (N_6577,N_4540,N_3840);
xor U6578 (N_6578,N_3724,N_3735);
or U6579 (N_6579,N_4173,N_1723);
nand U6580 (N_6580,N_366,N_4039);
or U6581 (N_6581,N_2031,N_104);
or U6582 (N_6582,N_1602,N_1403);
or U6583 (N_6583,N_2537,N_4470);
nand U6584 (N_6584,N_1338,N_1598);
nand U6585 (N_6585,N_328,N_1981);
nand U6586 (N_6586,N_3498,N_4585);
and U6587 (N_6587,N_2,N_352);
nor U6588 (N_6588,N_4749,N_2713);
nand U6589 (N_6589,N_3299,N_325);
xnor U6590 (N_6590,N_2347,N_3774);
nand U6591 (N_6591,N_3335,N_1970);
xor U6592 (N_6592,N_3448,N_1391);
nor U6593 (N_6593,N_1645,N_1513);
nor U6594 (N_6594,N_3004,N_2121);
and U6595 (N_6595,N_4769,N_3917);
xor U6596 (N_6596,N_2756,N_1354);
and U6597 (N_6597,N_4635,N_1637);
or U6598 (N_6598,N_2980,N_1122);
or U6599 (N_6599,N_2812,N_2794);
nand U6600 (N_6600,N_894,N_1694);
nand U6601 (N_6601,N_26,N_551);
xor U6602 (N_6602,N_3984,N_4504);
or U6603 (N_6603,N_2850,N_2652);
or U6604 (N_6604,N_1941,N_1162);
nand U6605 (N_6605,N_4397,N_3733);
nand U6606 (N_6606,N_1866,N_3495);
nor U6607 (N_6607,N_2696,N_646);
nor U6608 (N_6608,N_2766,N_1171);
nor U6609 (N_6609,N_3229,N_1454);
and U6610 (N_6610,N_4175,N_316);
nand U6611 (N_6611,N_2530,N_279);
xnor U6612 (N_6612,N_1086,N_2232);
or U6613 (N_6613,N_4132,N_2430);
nand U6614 (N_6614,N_2451,N_1238);
or U6615 (N_6615,N_4576,N_851);
and U6616 (N_6616,N_4033,N_4865);
nor U6617 (N_6617,N_2510,N_1896);
nor U6618 (N_6618,N_4215,N_2565);
xor U6619 (N_6619,N_3088,N_3619);
nand U6620 (N_6620,N_3804,N_2070);
nand U6621 (N_6621,N_3370,N_3691);
nand U6622 (N_6622,N_1182,N_4385);
nor U6623 (N_6623,N_966,N_3525);
or U6624 (N_6624,N_861,N_2151);
nor U6625 (N_6625,N_4903,N_3740);
and U6626 (N_6626,N_1983,N_3596);
and U6627 (N_6627,N_580,N_212);
or U6628 (N_6628,N_871,N_2597);
nand U6629 (N_6629,N_1589,N_3671);
and U6630 (N_6630,N_3093,N_3668);
nand U6631 (N_6631,N_3009,N_167);
and U6632 (N_6632,N_3772,N_741);
nand U6633 (N_6633,N_1516,N_4051);
nand U6634 (N_6634,N_4880,N_955);
nor U6635 (N_6635,N_2916,N_2996);
nor U6636 (N_6636,N_568,N_1110);
xor U6637 (N_6637,N_3371,N_2004);
and U6638 (N_6638,N_2507,N_4640);
xor U6639 (N_6639,N_3409,N_2935);
xnor U6640 (N_6640,N_4951,N_4420);
nor U6641 (N_6641,N_3165,N_4182);
and U6642 (N_6642,N_240,N_4304);
nor U6643 (N_6643,N_2458,N_1324);
nor U6644 (N_6644,N_669,N_919);
nand U6645 (N_6645,N_2598,N_1620);
nand U6646 (N_6646,N_3049,N_4204);
nor U6647 (N_6647,N_1788,N_2162);
nand U6648 (N_6648,N_1405,N_1197);
xnor U6649 (N_6649,N_3522,N_1477);
nand U6650 (N_6650,N_3254,N_4062);
nand U6651 (N_6651,N_4229,N_937);
and U6652 (N_6652,N_827,N_1267);
or U6653 (N_6653,N_4925,N_2432);
xor U6654 (N_6654,N_976,N_1705);
and U6655 (N_6655,N_4901,N_2475);
nor U6656 (N_6656,N_75,N_1920);
nand U6657 (N_6657,N_4780,N_1273);
nand U6658 (N_6658,N_4168,N_2531);
and U6659 (N_6659,N_514,N_3164);
and U6660 (N_6660,N_2882,N_3648);
or U6661 (N_6661,N_3274,N_2419);
and U6662 (N_6662,N_739,N_4484);
and U6663 (N_6663,N_725,N_2629);
or U6664 (N_6664,N_1082,N_3188);
or U6665 (N_6665,N_4588,N_4774);
nor U6666 (N_6666,N_3095,N_2800);
and U6667 (N_6667,N_4489,N_1649);
nand U6668 (N_6668,N_560,N_4704);
nor U6669 (N_6669,N_2034,N_2002);
xor U6670 (N_6670,N_3594,N_4122);
and U6671 (N_6671,N_3447,N_4400);
xnor U6672 (N_6672,N_2813,N_3762);
and U6673 (N_6673,N_4885,N_10);
or U6674 (N_6674,N_2210,N_4518);
xor U6675 (N_6675,N_4945,N_244);
or U6676 (N_6676,N_3667,N_4639);
or U6677 (N_6677,N_2774,N_563);
nand U6678 (N_6678,N_1804,N_2255);
and U6679 (N_6679,N_2844,N_3806);
and U6680 (N_6680,N_118,N_1669);
nor U6681 (N_6681,N_570,N_4028);
nand U6682 (N_6682,N_233,N_3573);
nor U6683 (N_6683,N_2715,N_3893);
or U6684 (N_6684,N_3475,N_3420);
nor U6685 (N_6685,N_3452,N_1519);
nand U6686 (N_6686,N_4244,N_3185);
and U6687 (N_6687,N_4706,N_4970);
or U6688 (N_6688,N_4026,N_4321);
xor U6689 (N_6689,N_4292,N_4580);
xnor U6690 (N_6690,N_1151,N_881);
and U6691 (N_6691,N_3482,N_2362);
and U6692 (N_6692,N_2194,N_422);
xnor U6693 (N_6693,N_989,N_719);
nand U6694 (N_6694,N_892,N_3822);
or U6695 (N_6695,N_4775,N_2527);
or U6696 (N_6696,N_2886,N_2052);
nor U6697 (N_6697,N_4564,N_4568);
nand U6698 (N_6698,N_1373,N_2028);
nand U6699 (N_6699,N_3657,N_4603);
xnor U6700 (N_6700,N_2215,N_249);
nand U6701 (N_6701,N_4425,N_3547);
or U6702 (N_6702,N_3977,N_4995);
or U6703 (N_6703,N_4597,N_3322);
and U6704 (N_6704,N_2734,N_1830);
and U6705 (N_6705,N_1557,N_4828);
xor U6706 (N_6706,N_4485,N_4177);
and U6707 (N_6707,N_2289,N_36);
nor U6708 (N_6708,N_1035,N_3300);
and U6709 (N_6709,N_807,N_4147);
or U6710 (N_6710,N_800,N_1915);
and U6711 (N_6711,N_396,N_117);
nand U6712 (N_6712,N_238,N_548);
and U6713 (N_6713,N_874,N_4981);
nor U6714 (N_6714,N_1715,N_3608);
nor U6715 (N_6715,N_4393,N_3096);
and U6716 (N_6716,N_940,N_1696);
or U6717 (N_6717,N_112,N_379);
and U6718 (N_6718,N_4462,N_494);
nand U6719 (N_6719,N_4098,N_4917);
nor U6720 (N_6720,N_3763,N_2270);
xnor U6721 (N_6721,N_1887,N_2526);
nor U6722 (N_6722,N_3654,N_3002);
and U6723 (N_6723,N_2765,N_3467);
nor U6724 (N_6724,N_2013,N_4403);
or U6725 (N_6725,N_4993,N_488);
or U6726 (N_6726,N_4942,N_4673);
and U6727 (N_6727,N_1484,N_3038);
nor U6728 (N_6728,N_3632,N_1658);
xor U6729 (N_6729,N_2960,N_273);
nor U6730 (N_6730,N_1611,N_3255);
and U6731 (N_6731,N_1414,N_1948);
nor U6732 (N_6732,N_1313,N_3827);
and U6733 (N_6733,N_562,N_4038);
or U6734 (N_6734,N_535,N_4010);
xor U6735 (N_6735,N_1069,N_593);
nand U6736 (N_6736,N_2757,N_1444);
and U6737 (N_6737,N_4127,N_4676);
xnor U6738 (N_6738,N_2669,N_4193);
nor U6739 (N_6739,N_4807,N_1275);
or U6740 (N_6740,N_3077,N_4797);
xnor U6741 (N_6741,N_4841,N_4226);
xnor U6742 (N_6742,N_2949,N_2555);
xor U6743 (N_6743,N_4636,N_994);
xnor U6744 (N_6744,N_2842,N_2989);
nand U6745 (N_6745,N_1129,N_2131);
xor U6746 (N_6746,N_3283,N_3173);
nand U6747 (N_6747,N_2724,N_3504);
and U6748 (N_6748,N_3071,N_606);
xor U6749 (N_6749,N_3692,N_1800);
and U6750 (N_6750,N_4920,N_203);
and U6751 (N_6751,N_4162,N_397);
nor U6752 (N_6752,N_3486,N_2367);
or U6753 (N_6753,N_1956,N_3112);
or U6754 (N_6754,N_637,N_2884);
nor U6755 (N_6755,N_685,N_463);
nand U6756 (N_6756,N_3834,N_1079);
xor U6757 (N_6757,N_4166,N_290);
nand U6758 (N_6758,N_2308,N_4467);
xor U6759 (N_6759,N_1060,N_3537);
nor U6760 (N_6760,N_3828,N_3584);
xnor U6761 (N_6761,N_4691,N_1799);
and U6762 (N_6762,N_545,N_2898);
nand U6763 (N_6763,N_4233,N_1968);
or U6764 (N_6764,N_4406,N_3170);
nor U6765 (N_6765,N_3959,N_303);
or U6766 (N_6766,N_4441,N_4971);
or U6767 (N_6767,N_2566,N_3434);
nand U6768 (N_6768,N_3559,N_3702);
nand U6769 (N_6769,N_3897,N_1101);
xor U6770 (N_6770,N_2338,N_2394);
or U6771 (N_6771,N_432,N_4295);
nor U6772 (N_6772,N_1076,N_4712);
nand U6773 (N_6773,N_3079,N_3778);
xnor U6774 (N_6774,N_2320,N_4734);
nor U6775 (N_6775,N_2365,N_3238);
nand U6776 (N_6776,N_3736,N_2108);
xor U6777 (N_6777,N_2649,N_476);
or U6778 (N_6778,N_3690,N_4083);
and U6779 (N_6779,N_3194,N_636);
nand U6780 (N_6780,N_3989,N_1121);
and U6781 (N_6781,N_3646,N_3160);
nand U6782 (N_6782,N_309,N_2158);
or U6783 (N_6783,N_3555,N_1037);
or U6784 (N_6784,N_4134,N_684);
nand U6785 (N_6785,N_1538,N_466);
or U6786 (N_6786,N_2680,N_3390);
xnor U6787 (N_6787,N_1748,N_277);
and U6788 (N_6788,N_869,N_3451);
xor U6789 (N_6789,N_4079,N_930);
xnor U6790 (N_6790,N_1625,N_4091);
nand U6791 (N_6791,N_1713,N_3830);
nand U6792 (N_6792,N_820,N_1457);
nor U6793 (N_6793,N_3933,N_3512);
xor U6794 (N_6794,N_838,N_3485);
or U6795 (N_6795,N_3374,N_3422);
and U6796 (N_6796,N_783,N_1046);
nand U6797 (N_6797,N_1666,N_2958);
and U6798 (N_6798,N_4852,N_4357);
or U6799 (N_6799,N_3693,N_540);
nand U6800 (N_6800,N_4326,N_1839);
xor U6801 (N_6801,N_4121,N_3716);
nand U6802 (N_6802,N_3226,N_4115);
xor U6803 (N_6803,N_1214,N_197);
xnor U6804 (N_6804,N_671,N_3270);
nand U6805 (N_6805,N_1856,N_2085);
or U6806 (N_6806,N_4790,N_3056);
and U6807 (N_6807,N_2594,N_2664);
nor U6808 (N_6808,N_986,N_3505);
and U6809 (N_6809,N_4054,N_2295);
or U6810 (N_6810,N_766,N_2363);
and U6811 (N_6811,N_3645,N_4748);
nor U6812 (N_6812,N_945,N_105);
nor U6813 (N_6813,N_2858,N_4331);
nand U6814 (N_6814,N_4113,N_852);
xor U6815 (N_6815,N_1315,N_478);
nand U6816 (N_6816,N_4805,N_3309);
nor U6817 (N_6817,N_1317,N_3695);
nand U6818 (N_6818,N_2964,N_907);
nand U6819 (N_6819,N_1038,N_403);
nand U6820 (N_6820,N_133,N_3105);
nand U6821 (N_6821,N_2677,N_2229);
xnor U6822 (N_6822,N_829,N_94);
or U6823 (N_6823,N_516,N_282);
and U6824 (N_6824,N_1431,N_1861);
and U6825 (N_6825,N_103,N_1030);
and U6826 (N_6826,N_2387,N_2589);
xor U6827 (N_6827,N_3413,N_3344);
and U6828 (N_6828,N_2712,N_2201);
xnor U6829 (N_6829,N_2236,N_4632);
xnor U6830 (N_6830,N_370,N_1652);
or U6831 (N_6831,N_2306,N_2479);
nand U6832 (N_6832,N_3046,N_2735);
or U6833 (N_6833,N_1773,N_3517);
or U6834 (N_6834,N_2298,N_969);
nand U6835 (N_6835,N_1815,N_2231);
nor U6836 (N_6836,N_3742,N_4059);
xor U6837 (N_6837,N_1241,N_700);
xnor U6838 (N_6838,N_3151,N_3937);
nand U6839 (N_6839,N_4976,N_3016);
xnor U6840 (N_6840,N_349,N_1731);
or U6841 (N_6841,N_850,N_3405);
nor U6842 (N_6842,N_394,N_981);
or U6843 (N_6843,N_1954,N_1103);
xor U6844 (N_6844,N_3947,N_1759);
xor U6845 (N_6845,N_3035,N_2463);
xnor U6846 (N_6846,N_968,N_2086);
xnor U6847 (N_6847,N_834,N_3548);
or U6848 (N_6848,N_1717,N_833);
nand U6849 (N_6849,N_847,N_794);
and U6850 (N_6850,N_4800,N_3231);
nand U6851 (N_6851,N_2074,N_1195);
xnor U6852 (N_6852,N_2600,N_1797);
nand U6853 (N_6853,N_3513,N_1982);
xnor U6854 (N_6854,N_1963,N_3470);
and U6855 (N_6855,N_1504,N_391);
xnor U6856 (N_6856,N_2373,N_219);
and U6857 (N_6857,N_3220,N_1372);
xnor U6858 (N_6858,N_1975,N_1067);
or U6859 (N_6859,N_296,N_3133);
or U6860 (N_6860,N_3070,N_4535);
nand U6861 (N_6861,N_1486,N_4075);
nand U6862 (N_6862,N_4899,N_428);
nor U6863 (N_6863,N_4809,N_2107);
or U6864 (N_6864,N_3111,N_1256);
nand U6865 (N_6865,N_1445,N_450);
nand U6866 (N_6866,N_1390,N_1633);
and U6867 (N_6867,N_135,N_2933);
or U6868 (N_6868,N_1130,N_4220);
nor U6869 (N_6869,N_3443,N_910);
xor U6870 (N_6870,N_3623,N_3658);
nand U6871 (N_6871,N_2370,N_2981);
nand U6872 (N_6872,N_3069,N_4473);
xnor U6873 (N_6873,N_1185,N_3656);
xor U6874 (N_6874,N_4773,N_1274);
and U6875 (N_6875,N_2919,N_1347);
or U6876 (N_6876,N_1969,N_1518);
xor U6877 (N_6877,N_79,N_967);
nand U6878 (N_6878,N_2951,N_4363);
xnor U6879 (N_6879,N_3455,N_3960);
or U6880 (N_6880,N_4831,N_1244);
nand U6881 (N_6881,N_2412,N_509);
xor U6882 (N_6882,N_300,N_2729);
and U6883 (N_6883,N_3993,N_3110);
nand U6884 (N_6884,N_2577,N_4700);
and U6885 (N_6885,N_3127,N_3579);
nand U6886 (N_6886,N_2749,N_4410);
or U6887 (N_6887,N_1118,N_4939);
xnor U6888 (N_6888,N_4966,N_2625);
nand U6889 (N_6889,N_1008,N_731);
and U6890 (N_6890,N_1502,N_3603);
or U6891 (N_6891,N_1778,N_2446);
or U6892 (N_6892,N_3534,N_318);
or U6893 (N_6893,N_523,N_2708);
nor U6894 (N_6894,N_4327,N_4003);
xnor U6895 (N_6895,N_2266,N_1330);
xor U6896 (N_6896,N_2030,N_4811);
nor U6897 (N_6897,N_2303,N_302);
nor U6898 (N_6898,N_4844,N_4577);
nand U6899 (N_6899,N_1922,N_673);
and U6900 (N_6900,N_4435,N_4362);
or U6901 (N_6901,N_618,N_4384);
xnor U6902 (N_6902,N_2425,N_754);
nand U6903 (N_6903,N_3359,N_1140);
and U6904 (N_6904,N_2485,N_2282);
or U6905 (N_6905,N_4257,N_880);
nand U6906 (N_6906,N_2778,N_3159);
nor U6907 (N_6907,N_762,N_2639);
nor U6908 (N_6908,N_2364,N_4756);
and U6909 (N_6909,N_1157,N_2075);
and U6910 (N_6910,N_2802,N_1900);
nand U6911 (N_6911,N_1284,N_1191);
or U6912 (N_6912,N_1597,N_1615);
and U6913 (N_6913,N_2673,N_1698);
or U6914 (N_6914,N_2382,N_3612);
nor U6915 (N_6915,N_524,N_4963);
xor U6916 (N_6916,N_4587,N_1382);
nand U6917 (N_6917,N_1893,N_4492);
and U6918 (N_6918,N_3155,N_1308);
or U6919 (N_6919,N_2902,N_3297);
and U6920 (N_6920,N_1594,N_855);
nor U6921 (N_6921,N_4685,N_1766);
nor U6922 (N_6922,N_1923,N_985);
nor U6923 (N_6923,N_680,N_343);
nor U6924 (N_6924,N_1742,N_372);
or U6925 (N_6925,N_2528,N_936);
nand U6926 (N_6926,N_2539,N_252);
xor U6927 (N_6927,N_4317,N_2838);
nor U6928 (N_6928,N_3025,N_4528);
or U6929 (N_6929,N_1697,N_3752);
or U6930 (N_6930,N_3456,N_3725);
and U6931 (N_6931,N_3784,N_1398);
nand U6932 (N_6932,N_293,N_3874);
nor U6933 (N_6933,N_1771,N_4561);
xor U6934 (N_6934,N_2606,N_3901);
xor U6935 (N_6935,N_3227,N_953);
nand U6936 (N_6936,N_2511,N_59);
or U6937 (N_6937,N_481,N_90);
xor U6938 (N_6938,N_621,N_1874);
nand U6939 (N_6939,N_1359,N_791);
or U6940 (N_6940,N_3346,N_4698);
xnor U6941 (N_6941,N_2992,N_3956);
nor U6942 (N_6942,N_4739,N_3529);
nor U6943 (N_6943,N_4459,N_1224);
or U6944 (N_6944,N_3308,N_3465);
nor U6945 (N_6945,N_1474,N_4218);
xnor U6946 (N_6946,N_4645,N_2788);
nand U6947 (N_6947,N_2204,N_472);
nand U6948 (N_6948,N_578,N_2799);
xor U6949 (N_6949,N_4171,N_2292);
nor U6950 (N_6950,N_845,N_2627);
nand U6951 (N_6951,N_3481,N_4688);
or U6952 (N_6952,N_321,N_952);
and U6953 (N_6953,N_2124,N_1485);
or U6954 (N_6954,N_2910,N_1094);
nor U6955 (N_6955,N_1967,N_2111);
nor U6956 (N_6956,N_3383,N_2768);
nor U6957 (N_6957,N_4599,N_3366);
xor U6958 (N_6958,N_4779,N_1022);
nor U6959 (N_6959,N_2209,N_3241);
nand U6960 (N_6960,N_2271,N_3878);
nand U6961 (N_6961,N_4965,N_2314);
xor U6962 (N_6962,N_1595,N_4411);
xnor U6963 (N_6963,N_95,N_2376);
nand U6964 (N_6964,N_1236,N_3289);
or U6965 (N_6965,N_3005,N_3461);
or U6966 (N_6966,N_4759,N_4262);
nor U6967 (N_6967,N_1408,N_1741);
nor U6968 (N_6968,N_3783,N_40);
and U6969 (N_6969,N_3950,N_3595);
or U6970 (N_6970,N_2835,N_1953);
and U6971 (N_6971,N_4381,N_3328);
xor U6972 (N_6972,N_1393,N_3218);
nand U6973 (N_6973,N_902,N_433);
and U6974 (N_6974,N_797,N_4776);
and U6975 (N_6975,N_600,N_2983);
nand U6976 (N_6976,N_404,N_4724);
nor U6977 (N_6977,N_284,N_2444);
nand U6978 (N_6978,N_4324,N_2779);
or U6979 (N_6979,N_1782,N_1392);
nand U6980 (N_6980,N_2611,N_364);
xnor U6981 (N_6981,N_848,N_2985);
nand U6982 (N_6982,N_4076,N_2690);
xor U6983 (N_6983,N_2099,N_4987);
and U6984 (N_6984,N_1929,N_1847);
nor U6985 (N_6985,N_4683,N_2454);
xnor U6986 (N_6986,N_576,N_842);
xnor U6987 (N_6987,N_4149,N_3064);
or U6988 (N_6988,N_2146,N_682);
xor U6989 (N_6989,N_4586,N_2651);
and U6990 (N_6990,N_19,N_1767);
nand U6991 (N_6991,N_4232,N_1108);
and U6992 (N_6992,N_3425,N_2087);
nor U6993 (N_6993,N_2723,N_272);
and U6994 (N_6994,N_350,N_1674);
or U6995 (N_6995,N_1413,N_4853);
nor U6996 (N_6996,N_2966,N_2830);
nand U6997 (N_6997,N_1048,N_742);
nand U6998 (N_6998,N_276,N_4208);
or U6999 (N_6999,N_1422,N_529);
nand U7000 (N_7000,N_2378,N_2262);
nor U7001 (N_7001,N_4714,N_500);
xor U7002 (N_7002,N_3971,N_4980);
xnor U7003 (N_7003,N_908,N_1310);
nor U7004 (N_7004,N_956,N_2873);
xnor U7005 (N_7005,N_4548,N_4184);
nor U7006 (N_7006,N_1805,N_1242);
or U7007 (N_7007,N_2956,N_4941);
and U7008 (N_7008,N_4011,N_747);
nand U7009 (N_7009,N_2672,N_733);
nor U7010 (N_7010,N_1200,N_2846);
or U7011 (N_7011,N_2697,N_3714);
xor U7012 (N_7012,N_3737,N_2216);
or U7013 (N_7013,N_496,N_4750);
and U7014 (N_7014,N_2579,N_4433);
nand U7015 (N_7015,N_3568,N_3293);
nor U7016 (N_7016,N_4721,N_4626);
nand U7017 (N_7017,N_1908,N_1769);
nor U7018 (N_7018,N_4000,N_2178);
xor U7019 (N_7019,N_136,N_3631);
nor U7020 (N_7020,N_456,N_3209);
or U7021 (N_7021,N_3499,N_659);
nand U7022 (N_7022,N_1719,N_958);
nand U7023 (N_7023,N_4049,N_424);
and U7024 (N_7024,N_2040,N_405);
and U7025 (N_7025,N_2019,N_194);
xnor U7026 (N_7026,N_4686,N_4271);
and U7027 (N_7027,N_3060,N_3473);
nor U7028 (N_7028,N_2771,N_2761);
nor U7029 (N_7029,N_1816,N_3871);
xor U7030 (N_7030,N_4836,N_843);
nand U7031 (N_7031,N_1532,N_778);
or U7032 (N_7032,N_3985,N_1859);
xor U7033 (N_7033,N_1974,N_1904);
or U7034 (N_7034,N_4946,N_3150);
or U7035 (N_7035,N_2748,N_1455);
nor U7036 (N_7036,N_4824,N_586);
xor U7037 (N_7037,N_4421,N_4325);
xnor U7038 (N_7038,N_4728,N_795);
and U7039 (N_7039,N_1952,N_3711);
xnor U7040 (N_7040,N_3389,N_1822);
or U7041 (N_7041,N_1201,N_3240);
nor U7042 (N_7042,N_1018,N_2008);
and U7043 (N_7043,N_3554,N_2551);
xnor U7044 (N_7044,N_2453,N_172);
xor U7045 (N_7045,N_4276,N_4660);
xnor U7046 (N_7046,N_2200,N_2388);
and U7047 (N_7047,N_564,N_3968);
nor U7048 (N_7048,N_2717,N_2806);
and U7049 (N_7049,N_4868,N_1793);
or U7050 (N_7050,N_2105,N_787);
and U7051 (N_7051,N_4560,N_3424);
xor U7052 (N_7052,N_4419,N_1120);
or U7053 (N_7053,N_2334,N_270);
nand U7054 (N_7054,N_896,N_199);
xor U7055 (N_7055,N_2043,N_2009);
nand U7056 (N_7056,N_2926,N_4376);
xnor U7057 (N_7057,N_3137,N_3765);
and U7058 (N_7058,N_522,N_474);
and U7059 (N_7059,N_2862,N_3437);
nor U7060 (N_7060,N_4502,N_125);
nor U7061 (N_7061,N_33,N_158);
or U7062 (N_7062,N_3880,N_4139);
xor U7063 (N_7063,N_1243,N_1469);
and U7064 (N_7064,N_392,N_3479);
or U7065 (N_7065,N_2573,N_4926);
xnor U7066 (N_7066,N_617,N_4338);
nor U7067 (N_7067,N_2818,N_1536);
or U7068 (N_7068,N_1960,N_4893);
xnor U7069 (N_7069,N_2523,N_1772);
or U7070 (N_7070,N_1071,N_2881);
nand U7071 (N_7071,N_565,N_417);
nand U7072 (N_7072,N_1276,N_4476);
xor U7073 (N_7073,N_3271,N_3312);
or U7074 (N_7074,N_3230,N_1533);
nand U7075 (N_7075,N_2359,N_4956);
nor U7076 (N_7076,N_4201,N_3808);
nand U7077 (N_7077,N_3007,N_4716);
and U7078 (N_7078,N_4938,N_4798);
nand U7079 (N_7079,N_2410,N_862);
nor U7080 (N_7080,N_3627,N_4305);
or U7081 (N_7081,N_4975,N_574);
and U7082 (N_7082,N_261,N_216);
and U7083 (N_7083,N_4747,N_2944);
or U7084 (N_7084,N_2632,N_3080);
and U7085 (N_7085,N_3635,N_799);
xor U7086 (N_7086,N_607,N_4810);
or U7087 (N_7087,N_3540,N_3248);
nor U7088 (N_7088,N_2504,N_2468);
nand U7089 (N_7089,N_4085,N_2120);
xor U7090 (N_7090,N_3549,N_668);
or U7091 (N_7091,N_3813,N_4869);
and U7092 (N_7092,N_152,N_3792);
nand U7093 (N_7093,N_775,N_4490);
nand U7094 (N_7094,N_2957,N_1531);
nor U7095 (N_7095,N_3228,N_917);
or U7096 (N_7096,N_1616,N_2795);
nand U7097 (N_7097,N_2014,N_1865);
nor U7098 (N_7098,N_41,N_2921);
nor U7099 (N_7099,N_0,N_2852);
nand U7100 (N_7100,N_4457,N_8);
and U7101 (N_7101,N_4507,N_1659);
nor U7102 (N_7102,N_1087,N_3884);
nor U7103 (N_7103,N_1527,N_3281);
and U7104 (N_7104,N_1876,N_1062);
nor U7105 (N_7105,N_3258,N_4886);
or U7106 (N_7106,N_2159,N_2784);
nand U7107 (N_7107,N_3949,N_732);
nand U7108 (N_7108,N_4322,N_1342);
xnor U7109 (N_7109,N_4498,N_3369);
xnor U7110 (N_7110,N_3256,N_1332);
nor U7111 (N_7111,N_2290,N_3108);
nor U7112 (N_7112,N_4395,N_1933);
xor U7113 (N_7113,N_4770,N_4986);
nor U7114 (N_7114,N_3927,N_2148);
and U7115 (N_7115,N_1675,N_4992);
or U7116 (N_7116,N_2945,N_3244);
or U7117 (N_7117,N_1739,N_693);
nor U7118 (N_7118,N_1521,N_2145);
or U7119 (N_7119,N_451,N_1554);
nand U7120 (N_7120,N_329,N_205);
or U7121 (N_7121,N_934,N_2683);
or U7122 (N_7122,N_4323,N_1560);
nor U7123 (N_7123,N_1161,N_622);
and U7124 (N_7124,N_4690,N_1770);
xnor U7125 (N_7125,N_2471,N_291);
and U7126 (N_7126,N_4273,N_4082);
and U7127 (N_7127,N_3944,N_2978);
or U7128 (N_7128,N_2553,N_2502);
nand U7129 (N_7129,N_1078,N_1337);
or U7130 (N_7130,N_2369,N_28);
nor U7131 (N_7131,N_4382,N_4022);
nor U7132 (N_7132,N_4374,N_1481);
and U7133 (N_7133,N_712,N_4736);
and U7134 (N_7134,N_4784,N_1651);
and U7135 (N_7135,N_4194,N_3675);
nand U7136 (N_7136,N_4251,N_4281);
nor U7137 (N_7137,N_2435,N_4883);
xnor U7138 (N_7138,N_1776,N_2211);
nand U7139 (N_7139,N_4674,N_3754);
xor U7140 (N_7140,N_1261,N_760);
nand U7141 (N_7141,N_1017,N_4703);
nor U7142 (N_7142,N_1152,N_1580);
nor U7143 (N_7143,N_4350,N_2161);
or U7144 (N_7144,N_1350,N_297);
or U7145 (N_7145,N_385,N_1575);
nor U7146 (N_7146,N_1009,N_3124);
nor U7147 (N_7147,N_931,N_3843);
nor U7148 (N_7148,N_4919,N_532);
nor U7149 (N_7149,N_228,N_3368);
nand U7150 (N_7150,N_3416,N_1774);
nand U7151 (N_7151,N_1618,N_2044);
and U7152 (N_7152,N_2094,N_3);
nor U7153 (N_7153,N_3710,N_512);
nand U7154 (N_7154,N_2825,N_3329);
nand U7155 (N_7155,N_2793,N_3651);
nor U7156 (N_7156,N_3865,N_4461);
xnor U7157 (N_7157,N_638,N_1990);
nand U7158 (N_7158,N_4600,N_157);
xnor U7159 (N_7159,N_3617,N_1221);
nand U7160 (N_7160,N_4526,N_709);
nor U7161 (N_7161,N_1399,N_2315);
nor U7162 (N_7162,N_2895,N_2010);
xor U7163 (N_7163,N_1579,N_459);
xnor U7164 (N_7164,N_4651,N_3171);
xnor U7165 (N_7165,N_55,N_3196);
and U7166 (N_7166,N_706,N_4537);
and U7167 (N_7167,N_338,N_4834);
nand U7168 (N_7168,N_581,N_435);
or U7169 (N_7169,N_1604,N_702);
nor U7170 (N_7170,N_3823,N_4116);
or U7171 (N_7171,N_83,N_1213);
nand U7172 (N_7172,N_1817,N_3953);
xor U7173 (N_7173,N_3841,N_1255);
and U7174 (N_7174,N_1491,N_149);
and U7175 (N_7175,N_4255,N_3924);
or U7176 (N_7176,N_3508,N_644);
nand U7177 (N_7177,N_3047,N_37);
nand U7178 (N_7178,N_1528,N_718);
xnor U7179 (N_7179,N_1234,N_4630);
nor U7180 (N_7180,N_3967,N_3640);
nor U7181 (N_7181,N_1336,N_1783);
nor U7182 (N_7182,N_2719,N_71);
and U7183 (N_7183,N_1895,N_2247);
nand U7184 (N_7184,N_4015,N_1097);
and U7185 (N_7185,N_2277,N_3824);
xnor U7186 (N_7186,N_3310,N_427);
xnor U7187 (N_7187,N_2658,N_4339);
xnor U7188 (N_7188,N_3521,N_1917);
nand U7189 (N_7189,N_3816,N_4319);
nor U7190 (N_7190,N_4889,N_810);
xnor U7191 (N_7191,N_651,N_1541);
nor U7192 (N_7192,N_2650,N_4994);
or U7193 (N_7193,N_3709,N_4312);
nand U7194 (N_7194,N_1473,N_1678);
nand U7195 (N_7195,N_809,N_2393);
xnor U7196 (N_7196,N_2726,N_1899);
and U7197 (N_7197,N_1246,N_1056);
xnor U7198 (N_7198,N_2605,N_4590);
nor U7199 (N_7199,N_333,N_213);
or U7200 (N_7200,N_258,N_1443);
or U7201 (N_7201,N_4143,N_3262);
nand U7202 (N_7202,N_1984,N_1479);
nor U7203 (N_7203,N_2416,N_2552);
xor U7204 (N_7204,N_1607,N_1377);
nand U7205 (N_7205,N_3847,N_3746);
and U7206 (N_7206,N_1499,N_281);
nand U7207 (N_7207,N_4081,N_163);
xnor U7208 (N_7208,N_3581,N_2924);
xor U7209 (N_7209,N_734,N_978);
nand U7210 (N_7210,N_4768,N_1156);
nand U7211 (N_7211,N_4959,N_1857);
xnor U7212 (N_7212,N_1572,N_3926);
and U7213 (N_7213,N_3582,N_1571);
nand U7214 (N_7214,N_376,N_3662);
or U7215 (N_7215,N_504,N_248);
and U7216 (N_7216,N_1930,N_4829);
nor U7217 (N_7217,N_1764,N_1796);
or U7218 (N_7218,N_2648,N_1646);
nand U7219 (N_7219,N_1614,N_1305);
nor U7220 (N_7220,N_3518,N_1051);
xor U7221 (N_7221,N_4623,N_1897);
nand U7222 (N_7222,N_2324,N_141);
nand U7223 (N_7223,N_3730,N_2263);
nand U7224 (N_7224,N_2505,N_4303);
nor U7225 (N_7225,N_776,N_4497);
or U7226 (N_7226,N_400,N_411);
nand U7227 (N_7227,N_2661,N_4428);
xnor U7228 (N_7228,N_823,N_3156);
nand U7229 (N_7229,N_954,N_3214);
nand U7230 (N_7230,N_1163,N_3965);
nand U7231 (N_7231,N_4867,N_2234);
xor U7232 (N_7232,N_3412,N_3846);
xnor U7233 (N_7233,N_123,N_822);
xnor U7234 (N_7234,N_2452,N_4140);
and U7235 (N_7235,N_3372,N_1401);
nand U7236 (N_7236,N_2602,N_2097);
and U7237 (N_7237,N_815,N_2196);
or U7238 (N_7238,N_1072,N_1177);
or U7239 (N_7239,N_2856,N_846);
nand U7240 (N_7240,N_3207,N_1854);
nor U7241 (N_7241,N_3092,N_2414);
xor U7242 (N_7242,N_2000,N_2984);
or U7243 (N_7243,N_3027,N_4646);
and U7244 (N_7244,N_4789,N_3614);
and U7245 (N_7245,N_4332,N_1341);
nand U7246 (N_7246,N_1488,N_3870);
nor U7247 (N_7247,N_2332,N_1288);
or U7248 (N_7248,N_3845,N_2676);
and U7249 (N_7249,N_1394,N_4112);
and U7250 (N_7250,N_2125,N_1411);
and U7251 (N_7251,N_1603,N_3863);
or U7252 (N_7252,N_446,N_3251);
and U7253 (N_7253,N_4667,N_460);
xor U7254 (N_7254,N_3198,N_4211);
xor U7255 (N_7255,N_287,N_2100);
nor U7256 (N_7256,N_3734,N_1806);
xnor U7257 (N_7257,N_3768,N_1160);
nor U7258 (N_7258,N_632,N_1209);
nor U7259 (N_7259,N_1842,N_1410);
or U7260 (N_7260,N_1447,N_1708);
nor U7261 (N_7261,N_4399,N_3365);
xor U7262 (N_7262,N_2017,N_4916);
nand U7263 (N_7263,N_1613,N_3408);
and U7264 (N_7264,N_3491,N_811);
nand U7265 (N_7265,N_4407,N_4336);
nand U7266 (N_7266,N_3779,N_1913);
and U7267 (N_7267,N_4794,N_2892);
or U7268 (N_7268,N_138,N_2128);
and U7269 (N_7269,N_3661,N_3684);
xor U7270 (N_7270,N_337,N_259);
xnor U7271 (N_7271,N_3415,N_904);
nand U7272 (N_7272,N_192,N_2071);
nor U7273 (N_7273,N_4567,N_779);
nor U7274 (N_7274,N_147,N_2420);
or U7275 (N_7275,N_2666,N_2969);
nor U7276 (N_7276,N_4067,N_4539);
nand U7277 (N_7277,N_184,N_4622);
and U7278 (N_7278,N_932,N_441);
or U7279 (N_7279,N_1701,N_2319);
xor U7280 (N_7280,N_1988,N_696);
nand U7281 (N_7281,N_479,N_2169);
xor U7282 (N_7282,N_2585,N_2899);
nor U7283 (N_7283,N_3755,N_1540);
or U7284 (N_7284,N_1775,N_1993);
xor U7285 (N_7285,N_4508,N_4914);
and U7286 (N_7286,N_3797,N_1853);
and U7287 (N_7287,N_1534,N_4658);
or U7288 (N_7288,N_1115,N_4349);
nor U7289 (N_7289,N_2171,N_3373);
nand U7290 (N_7290,N_777,N_234);
nand U7291 (N_7291,N_1301,N_437);
xnor U7292 (N_7292,N_3943,N_462);
and U7293 (N_7293,N_2787,N_2358);
and U7294 (N_7294,N_2801,N_3327);
or U7295 (N_7295,N_1449,N_3642);
nand U7296 (N_7296,N_2220,N_639);
xor U7297 (N_7297,N_3484,N_2422);
or U7298 (N_7298,N_3888,N_4250);
and U7299 (N_7299,N_3587,N_1263);
nand U7300 (N_7300,N_1593,N_2252);
and U7301 (N_7301,N_4141,N_4344);
nor U7302 (N_7302,N_4111,N_722);
nor U7303 (N_7303,N_2867,N_1235);
and U7304 (N_7304,N_4044,N_443);
or U7305 (N_7305,N_109,N_1251);
xor U7306 (N_7306,N_4256,N_2037);
xnor U7307 (N_7307,N_3459,N_4949);
nor U7308 (N_7308,N_1814,N_841);
and U7309 (N_7309,N_1188,N_4932);
nand U7310 (N_7310,N_3192,N_4472);
or U7311 (N_7311,N_4249,N_2888);
nand U7312 (N_7312,N_2701,N_873);
and U7313 (N_7313,N_12,N_4935);
and U7314 (N_7314,N_3085,N_4373);
xnor U7315 (N_7315,N_4801,N_305);
or U7316 (N_7316,N_226,N_3492);
and U7317 (N_7317,N_714,N_3001);
or U7318 (N_7318,N_891,N_1732);
and U7319 (N_7319,N_380,N_1583);
and U7320 (N_7320,N_1049,N_2149);
nor U7321 (N_7321,N_620,N_701);
nand U7322 (N_7322,N_342,N_3886);
nand U7323 (N_7323,N_2484,N_2767);
and U7324 (N_7324,N_804,N_782);
xnor U7325 (N_7325,N_4238,N_4275);
xnor U7326 (N_7326,N_2851,N_1089);
or U7327 (N_7327,N_1136,N_1412);
xnor U7328 (N_7328,N_4795,N_2380);
and U7329 (N_7329,N_2436,N_4221);
xor U7330 (N_7330,N_679,N_4495);
nor U7331 (N_7331,N_2613,N_1289);
xor U7332 (N_7332,N_527,N_2006);
nand U7333 (N_7333,N_1099,N_3818);
nand U7334 (N_7334,N_4505,N_2557);
and U7335 (N_7335,N_2323,N_2139);
xor U7336 (N_7336,N_1564,N_1912);
or U7337 (N_7337,N_2495,N_1205);
or U7338 (N_7338,N_1640,N_3636);
or U7339 (N_7339,N_3875,N_2456);
nand U7340 (N_7340,N_455,N_1836);
nand U7341 (N_7341,N_2409,N_2906);
xor U7342 (N_7342,N_87,N_698);
nand U7343 (N_7343,N_3694,N_4961);
nor U7344 (N_7344,N_1127,N_3913);
and U7345 (N_7345,N_2500,N_445);
or U7346 (N_7346,N_728,N_4074);
nand U7347 (N_7347,N_2593,N_4624);
nand U7348 (N_7348,N_2988,N_1029);
nor U7349 (N_7349,N_13,N_2191);
nor U7350 (N_7350,N_3992,N_4573);
xnor U7351 (N_7351,N_4136,N_2955);
nand U7352 (N_7352,N_2326,N_735);
and U7353 (N_7353,N_4107,N_51);
or U7354 (N_7354,N_3058,N_1844);
nand U7355 (N_7355,N_951,N_3350);
nand U7356 (N_7356,N_1515,N_1441);
xor U7357 (N_7357,N_1220,N_641);
or U7358 (N_7358,N_3037,N_3810);
and U7359 (N_7359,N_1010,N_588);
nand U7360 (N_7360,N_4819,N_3339);
nor U7361 (N_7361,N_1283,N_1786);
and U7362 (N_7362,N_4625,N_835);
nand U7363 (N_7363,N_4562,N_4017);
nand U7364 (N_7364,N_4491,N_222);
or U7365 (N_7365,N_4680,N_1931);
xnor U7366 (N_7366,N_4846,N_4365);
nor U7367 (N_7367,N_3098,N_4114);
nand U7368 (N_7368,N_114,N_2792);
nand U7369 (N_7369,N_3406,N_3419);
nand U7370 (N_7370,N_1525,N_2517);
nor U7371 (N_7371,N_4735,N_4618);
nand U7372 (N_7372,N_547,N_595);
or U7373 (N_7373,N_3660,N_1348);
xor U7374 (N_7374,N_160,N_2797);
nor U7375 (N_7375,N_1882,N_2946);
xnor U7376 (N_7376,N_4862,N_3676);
and U7377 (N_7377,N_3857,N_4104);
xnor U7378 (N_7378,N_2905,N_4450);
xnor U7379 (N_7379,N_4245,N_246);
xnor U7380 (N_7380,N_2770,N_3154);
or U7381 (N_7381,N_2222,N_2423);
nor U7382 (N_7382,N_1758,N_2172);
nor U7383 (N_7383,N_2391,N_3010);
nor U7384 (N_7384,N_2643,N_703);
and U7385 (N_7385,N_4057,N_470);
or U7386 (N_7386,N_3942,N_2521);
nand U7387 (N_7387,N_345,N_2064);
and U7388 (N_7388,N_1667,N_1599);
and U7389 (N_7389,N_3401,N_2647);
nand U7390 (N_7390,N_498,N_1131);
or U7391 (N_7391,N_2057,N_4723);
xor U7392 (N_7392,N_3597,N_294);
nand U7393 (N_7393,N_1075,N_4089);
nor U7394 (N_7394,N_4830,N_3364);
xnor U7395 (N_7395,N_649,N_49);
nor U7396 (N_7396,N_4289,N_3249);
xnor U7397 (N_7397,N_3643,N_2486);
or U7398 (N_7398,N_4988,N_3904);
and U7399 (N_7399,N_2638,N_2943);
or U7400 (N_7400,N_76,N_2026);
or U7401 (N_7401,N_585,N_2871);
xor U7402 (N_7402,N_1396,N_3869);
and U7403 (N_7403,N_642,N_3028);
and U7404 (N_7404,N_1946,N_388);
or U7405 (N_7405,N_3183,N_1747);
xor U7406 (N_7406,N_3153,N_3551);
nor U7407 (N_7407,N_2855,N_3139);
xor U7408 (N_7408,N_1864,N_48);
and U7409 (N_7409,N_2791,N_214);
xnor U7410 (N_7410,N_1005,N_1547);
xnor U7411 (N_7411,N_1106,N_3040);
nand U7412 (N_7412,N_1919,N_1710);
nand U7413 (N_7413,N_4042,N_1328);
xor U7414 (N_7414,N_4991,N_2814);
nand U7415 (N_7415,N_1232,N_4481);
nand U7416 (N_7416,N_2193,N_1612);
nor U7417 (N_7417,N_663,N_3892);
and U7418 (N_7418,N_180,N_590);
and U7419 (N_7419,N_4960,N_1265);
and U7420 (N_7420,N_2140,N_4072);
nand U7421 (N_7421,N_2143,N_4979);
xor U7422 (N_7422,N_3767,N_5);
and U7423 (N_7423,N_1344,N_326);
nand U7424 (N_7424,N_554,N_3323);
xnor U7425 (N_7425,N_2929,N_353);
nor U7426 (N_7426,N_3773,N_4546);
nor U7427 (N_7427,N_4474,N_4239);
nand U7428 (N_7428,N_2934,N_204);
or U7429 (N_7429,N_1031,N_4514);
nor U7430 (N_7430,N_42,N_2018);
nand U7431 (N_7431,N_2656,N_3655);
and U7432 (N_7432,N_4496,N_4761);
or U7433 (N_7433,N_102,N_602);
nor U7434 (N_7434,N_1877,N_1291);
xnor U7435 (N_7435,N_16,N_1374);
or U7436 (N_7436,N_3861,N_4521);
nand U7437 (N_7437,N_4746,N_3866);
or U7438 (N_7438,N_3075,N_2790);
nand U7439 (N_7439,N_132,N_2133);
xnor U7440 (N_7440,N_2796,N_571);
nor U7441 (N_7441,N_1379,N_3882);
or U7442 (N_7442,N_977,N_780);
nand U7443 (N_7443,N_4517,N_4246);
xor U7444 (N_7444,N_3502,N_2268);
or U7445 (N_7445,N_330,N_1959);
or U7446 (N_7446,N_2567,N_2091);
nand U7447 (N_7447,N_2152,N_675);
xnor U7448 (N_7448,N_3574,N_4307);
nor U7449 (N_7449,N_1028,N_1229);
or U7450 (N_7450,N_382,N_1743);
nand U7451 (N_7451,N_3898,N_2246);
or U7452 (N_7452,N_1460,N_88);
nor U7453 (N_7453,N_748,N_612);
xor U7454 (N_7454,N_131,N_2060);
and U7455 (N_7455,N_749,N_528);
nor U7456 (N_7456,N_499,N_1437);
and U7457 (N_7457,N_2810,N_1971);
nand U7458 (N_7458,N_3796,N_915);
or U7459 (N_7459,N_2865,N_549);
or U7460 (N_7460,N_2544,N_4426);
and U7461 (N_7461,N_926,N_1879);
nand U7462 (N_7462,N_4643,N_50);
nand U7463 (N_7463,N_4417,N_3501);
nor U7464 (N_7464,N_3113,N_4575);
nor U7465 (N_7465,N_3045,N_4386);
and U7466 (N_7466,N_4871,N_3418);
nand U7467 (N_7467,N_2834,N_1725);
xnor U7468 (N_7468,N_2575,N_495);
and U7469 (N_7469,N_425,N_1158);
nor U7470 (N_7470,N_1656,N_4737);
and U7471 (N_7471,N_1894,N_1792);
or U7472 (N_7472,N_4541,N_2869);
or U7473 (N_7473,N_1582,N_561);
xor U7474 (N_7474,N_3566,N_4078);
and U7475 (N_7475,N_3476,N_2804);
nand U7476 (N_7476,N_4019,N_469);
nand U7477 (N_7477,N_1014,N_4109);
and U7478 (N_7478,N_3653,N_4024);
or U7479 (N_7479,N_4264,N_2288);
or U7480 (N_7480,N_4544,N_4629);
and U7481 (N_7481,N_1448,N_3376);
nor U7482 (N_7482,N_4614,N_942);
nor U7483 (N_7483,N_3609,N_4620);
nor U7484 (N_7484,N_974,N_2035);
and U7485 (N_7485,N_2604,N_1293);
xor U7486 (N_7486,N_2163,N_100);
or U7487 (N_7487,N_3464,N_724);
xnor U7488 (N_7488,N_2301,N_687);
nand U7489 (N_7489,N_1343,N_1661);
nand U7490 (N_7490,N_2248,N_1753);
or U7491 (N_7491,N_2227,N_2092);
and U7492 (N_7492,N_4602,N_1085);
or U7493 (N_7493,N_2096,N_1977);
and U7494 (N_7494,N_1762,N_1709);
xor U7495 (N_7495,N_1517,N_708);
nor U7496 (N_7496,N_3163,N_453);
nor U7497 (N_7497,N_928,N_1270);
xor U7498 (N_7498,N_4027,N_4086);
xnor U7499 (N_7499,N_14,N_4858);
and U7500 (N_7500,N_3491,N_211);
xnor U7501 (N_7501,N_613,N_3005);
xnor U7502 (N_7502,N_1498,N_3030);
and U7503 (N_7503,N_3949,N_3578);
nor U7504 (N_7504,N_3026,N_3607);
and U7505 (N_7505,N_1161,N_4891);
nand U7506 (N_7506,N_1460,N_2047);
nand U7507 (N_7507,N_4299,N_1387);
nor U7508 (N_7508,N_3194,N_2627);
nor U7509 (N_7509,N_718,N_3862);
nand U7510 (N_7510,N_528,N_4414);
or U7511 (N_7511,N_4929,N_1589);
or U7512 (N_7512,N_2306,N_3320);
or U7513 (N_7513,N_3702,N_3150);
nand U7514 (N_7514,N_3516,N_463);
or U7515 (N_7515,N_586,N_1730);
and U7516 (N_7516,N_264,N_4064);
nor U7517 (N_7517,N_1412,N_2067);
nor U7518 (N_7518,N_2107,N_186);
nor U7519 (N_7519,N_5,N_4184);
xor U7520 (N_7520,N_2896,N_1030);
or U7521 (N_7521,N_3717,N_1242);
nand U7522 (N_7522,N_3520,N_3563);
nor U7523 (N_7523,N_3377,N_3508);
nand U7524 (N_7524,N_19,N_4505);
nor U7525 (N_7525,N_2930,N_4962);
and U7526 (N_7526,N_713,N_3783);
or U7527 (N_7527,N_3424,N_1112);
nor U7528 (N_7528,N_3819,N_3195);
xnor U7529 (N_7529,N_4529,N_1683);
nor U7530 (N_7530,N_327,N_4791);
or U7531 (N_7531,N_3420,N_2234);
or U7532 (N_7532,N_1396,N_3166);
and U7533 (N_7533,N_2410,N_2060);
nand U7534 (N_7534,N_1463,N_3753);
nor U7535 (N_7535,N_1211,N_3930);
xnor U7536 (N_7536,N_2013,N_1065);
nand U7537 (N_7537,N_2736,N_2860);
nor U7538 (N_7538,N_1368,N_2057);
xnor U7539 (N_7539,N_31,N_2108);
nand U7540 (N_7540,N_663,N_2990);
nand U7541 (N_7541,N_807,N_2646);
nor U7542 (N_7542,N_1429,N_340);
nand U7543 (N_7543,N_4024,N_1278);
xnor U7544 (N_7544,N_1777,N_4349);
or U7545 (N_7545,N_3473,N_264);
or U7546 (N_7546,N_72,N_70);
or U7547 (N_7547,N_4738,N_1123);
or U7548 (N_7548,N_3951,N_112);
or U7549 (N_7549,N_3780,N_4402);
nor U7550 (N_7550,N_3843,N_995);
nor U7551 (N_7551,N_571,N_1327);
and U7552 (N_7552,N_2217,N_4143);
and U7553 (N_7553,N_4284,N_4743);
nand U7554 (N_7554,N_3429,N_530);
and U7555 (N_7555,N_3810,N_2750);
xor U7556 (N_7556,N_2494,N_1109);
xor U7557 (N_7557,N_124,N_3559);
nor U7558 (N_7558,N_3615,N_1262);
and U7559 (N_7559,N_2143,N_1057);
and U7560 (N_7560,N_4145,N_2049);
nand U7561 (N_7561,N_4678,N_3635);
xnor U7562 (N_7562,N_2994,N_2665);
or U7563 (N_7563,N_1308,N_3116);
nand U7564 (N_7564,N_599,N_71);
nor U7565 (N_7565,N_2887,N_3519);
or U7566 (N_7566,N_1323,N_4939);
and U7567 (N_7567,N_2186,N_1316);
nor U7568 (N_7568,N_4946,N_1773);
and U7569 (N_7569,N_2128,N_4519);
nor U7570 (N_7570,N_1332,N_4998);
and U7571 (N_7571,N_2414,N_2247);
nor U7572 (N_7572,N_1747,N_4356);
or U7573 (N_7573,N_4001,N_4511);
or U7574 (N_7574,N_2463,N_3493);
and U7575 (N_7575,N_3895,N_2016);
and U7576 (N_7576,N_3731,N_3612);
and U7577 (N_7577,N_2949,N_1368);
nor U7578 (N_7578,N_1936,N_531);
xnor U7579 (N_7579,N_1642,N_1885);
xnor U7580 (N_7580,N_2287,N_509);
or U7581 (N_7581,N_2707,N_1507);
xnor U7582 (N_7582,N_1864,N_766);
nand U7583 (N_7583,N_159,N_3538);
and U7584 (N_7584,N_2562,N_1923);
nand U7585 (N_7585,N_4793,N_553);
and U7586 (N_7586,N_1635,N_1627);
nand U7587 (N_7587,N_4218,N_522);
or U7588 (N_7588,N_3257,N_1193);
and U7589 (N_7589,N_4750,N_1621);
nor U7590 (N_7590,N_3952,N_775);
nor U7591 (N_7591,N_3238,N_4537);
nand U7592 (N_7592,N_607,N_4292);
and U7593 (N_7593,N_923,N_1489);
xnor U7594 (N_7594,N_892,N_1536);
nand U7595 (N_7595,N_3223,N_2856);
and U7596 (N_7596,N_336,N_261);
and U7597 (N_7597,N_713,N_1132);
xnor U7598 (N_7598,N_2920,N_4101);
and U7599 (N_7599,N_1344,N_2104);
nor U7600 (N_7600,N_3124,N_4880);
xnor U7601 (N_7601,N_4980,N_4789);
nor U7602 (N_7602,N_2774,N_15);
and U7603 (N_7603,N_2886,N_3985);
nor U7604 (N_7604,N_2018,N_4245);
nand U7605 (N_7605,N_1878,N_1741);
and U7606 (N_7606,N_4095,N_4007);
and U7607 (N_7607,N_3930,N_1229);
nor U7608 (N_7608,N_853,N_206);
and U7609 (N_7609,N_1375,N_3786);
xnor U7610 (N_7610,N_1969,N_1350);
xor U7611 (N_7611,N_2396,N_2006);
or U7612 (N_7612,N_5,N_2294);
or U7613 (N_7613,N_4036,N_4708);
xnor U7614 (N_7614,N_75,N_3914);
and U7615 (N_7615,N_1904,N_4333);
xnor U7616 (N_7616,N_4631,N_2299);
nand U7617 (N_7617,N_3517,N_2567);
or U7618 (N_7618,N_3281,N_3322);
xor U7619 (N_7619,N_893,N_1697);
and U7620 (N_7620,N_3019,N_2840);
xor U7621 (N_7621,N_116,N_4960);
nand U7622 (N_7622,N_3336,N_1318);
and U7623 (N_7623,N_868,N_1935);
nand U7624 (N_7624,N_4573,N_2078);
and U7625 (N_7625,N_383,N_576);
xnor U7626 (N_7626,N_4433,N_981);
and U7627 (N_7627,N_3508,N_4524);
nand U7628 (N_7628,N_4739,N_3035);
nand U7629 (N_7629,N_587,N_3095);
and U7630 (N_7630,N_1945,N_1510);
and U7631 (N_7631,N_125,N_938);
nor U7632 (N_7632,N_1260,N_4169);
xnor U7633 (N_7633,N_1342,N_636);
nor U7634 (N_7634,N_1818,N_3320);
nor U7635 (N_7635,N_2247,N_757);
nand U7636 (N_7636,N_760,N_3236);
xor U7637 (N_7637,N_53,N_837);
nand U7638 (N_7638,N_3210,N_999);
nand U7639 (N_7639,N_2058,N_1234);
and U7640 (N_7640,N_3056,N_45);
nand U7641 (N_7641,N_3384,N_4518);
xnor U7642 (N_7642,N_4708,N_2103);
or U7643 (N_7643,N_3405,N_954);
nand U7644 (N_7644,N_4145,N_351);
and U7645 (N_7645,N_4252,N_2851);
and U7646 (N_7646,N_578,N_58);
nor U7647 (N_7647,N_1327,N_912);
nand U7648 (N_7648,N_638,N_2674);
nor U7649 (N_7649,N_4088,N_4016);
xor U7650 (N_7650,N_4937,N_1468);
and U7651 (N_7651,N_3389,N_2615);
nor U7652 (N_7652,N_1386,N_2153);
nand U7653 (N_7653,N_1778,N_2365);
or U7654 (N_7654,N_752,N_3361);
nor U7655 (N_7655,N_1450,N_1653);
or U7656 (N_7656,N_2759,N_187);
and U7657 (N_7657,N_3206,N_1987);
nand U7658 (N_7658,N_4701,N_3880);
or U7659 (N_7659,N_3390,N_1390);
and U7660 (N_7660,N_236,N_1258);
and U7661 (N_7661,N_2287,N_2038);
or U7662 (N_7662,N_1542,N_1360);
xnor U7663 (N_7663,N_4376,N_1759);
and U7664 (N_7664,N_421,N_3950);
or U7665 (N_7665,N_2015,N_4778);
nor U7666 (N_7666,N_2271,N_2343);
xnor U7667 (N_7667,N_3924,N_1010);
and U7668 (N_7668,N_649,N_2850);
or U7669 (N_7669,N_3951,N_721);
and U7670 (N_7670,N_3369,N_4524);
or U7671 (N_7671,N_1283,N_3470);
and U7672 (N_7672,N_3018,N_2623);
or U7673 (N_7673,N_1272,N_543);
xor U7674 (N_7674,N_2469,N_1770);
xor U7675 (N_7675,N_1389,N_1175);
and U7676 (N_7676,N_2721,N_2152);
nand U7677 (N_7677,N_159,N_4457);
or U7678 (N_7678,N_3192,N_1494);
and U7679 (N_7679,N_4944,N_2283);
nand U7680 (N_7680,N_1657,N_2422);
and U7681 (N_7681,N_3428,N_1348);
xor U7682 (N_7682,N_4987,N_52);
and U7683 (N_7683,N_2679,N_1849);
nand U7684 (N_7684,N_3831,N_2043);
nor U7685 (N_7685,N_3865,N_3730);
or U7686 (N_7686,N_2625,N_2044);
and U7687 (N_7687,N_1547,N_971);
nand U7688 (N_7688,N_4904,N_21);
and U7689 (N_7689,N_3389,N_947);
nor U7690 (N_7690,N_4918,N_3251);
or U7691 (N_7691,N_1110,N_4776);
nor U7692 (N_7692,N_4548,N_262);
nor U7693 (N_7693,N_2640,N_4379);
and U7694 (N_7694,N_2018,N_3012);
nand U7695 (N_7695,N_3452,N_2867);
nand U7696 (N_7696,N_3799,N_4032);
nor U7697 (N_7697,N_4704,N_591);
nor U7698 (N_7698,N_493,N_2615);
xor U7699 (N_7699,N_1808,N_782);
nor U7700 (N_7700,N_1394,N_141);
nand U7701 (N_7701,N_700,N_628);
nand U7702 (N_7702,N_879,N_4188);
nor U7703 (N_7703,N_2728,N_147);
nor U7704 (N_7704,N_1070,N_4322);
nor U7705 (N_7705,N_3831,N_4471);
xnor U7706 (N_7706,N_2060,N_4714);
or U7707 (N_7707,N_3549,N_4250);
nand U7708 (N_7708,N_1007,N_4250);
xor U7709 (N_7709,N_2460,N_3925);
xnor U7710 (N_7710,N_956,N_4335);
nor U7711 (N_7711,N_3555,N_516);
xnor U7712 (N_7712,N_3360,N_3270);
nor U7713 (N_7713,N_32,N_4830);
nand U7714 (N_7714,N_751,N_1913);
nor U7715 (N_7715,N_2435,N_3469);
or U7716 (N_7716,N_4276,N_3343);
or U7717 (N_7717,N_3512,N_4734);
nand U7718 (N_7718,N_4149,N_2598);
and U7719 (N_7719,N_1028,N_3135);
and U7720 (N_7720,N_1159,N_2277);
nor U7721 (N_7721,N_2757,N_4328);
and U7722 (N_7722,N_3234,N_4348);
nand U7723 (N_7723,N_4179,N_863);
nor U7724 (N_7724,N_1270,N_837);
nand U7725 (N_7725,N_1012,N_2453);
and U7726 (N_7726,N_4833,N_3125);
xor U7727 (N_7727,N_4940,N_947);
nand U7728 (N_7728,N_2030,N_3924);
nor U7729 (N_7729,N_4408,N_3932);
and U7730 (N_7730,N_2495,N_682);
or U7731 (N_7731,N_820,N_1827);
or U7732 (N_7732,N_1421,N_3951);
xnor U7733 (N_7733,N_2680,N_4226);
xor U7734 (N_7734,N_2040,N_1058);
nand U7735 (N_7735,N_4043,N_4335);
and U7736 (N_7736,N_1584,N_2495);
nand U7737 (N_7737,N_4151,N_663);
or U7738 (N_7738,N_4941,N_301);
nand U7739 (N_7739,N_4315,N_1437);
or U7740 (N_7740,N_1296,N_3358);
and U7741 (N_7741,N_4694,N_2578);
and U7742 (N_7742,N_3010,N_196);
nor U7743 (N_7743,N_1461,N_154);
and U7744 (N_7744,N_37,N_4524);
nor U7745 (N_7745,N_3635,N_2579);
nand U7746 (N_7746,N_1859,N_80);
nor U7747 (N_7747,N_4218,N_1877);
and U7748 (N_7748,N_4146,N_3982);
and U7749 (N_7749,N_1144,N_21);
and U7750 (N_7750,N_1682,N_3860);
or U7751 (N_7751,N_555,N_771);
or U7752 (N_7752,N_2733,N_674);
or U7753 (N_7753,N_465,N_4174);
nor U7754 (N_7754,N_949,N_1551);
xnor U7755 (N_7755,N_2387,N_4693);
and U7756 (N_7756,N_3866,N_163);
nor U7757 (N_7757,N_2667,N_1275);
nand U7758 (N_7758,N_1814,N_3784);
nor U7759 (N_7759,N_3260,N_1877);
nor U7760 (N_7760,N_177,N_3406);
xnor U7761 (N_7761,N_3621,N_3345);
or U7762 (N_7762,N_2449,N_2737);
and U7763 (N_7763,N_4303,N_1946);
xor U7764 (N_7764,N_106,N_3630);
or U7765 (N_7765,N_189,N_1347);
and U7766 (N_7766,N_2942,N_3220);
nand U7767 (N_7767,N_3674,N_4595);
nand U7768 (N_7768,N_4469,N_4002);
nor U7769 (N_7769,N_4445,N_2384);
xnor U7770 (N_7770,N_3817,N_915);
and U7771 (N_7771,N_2100,N_2563);
xor U7772 (N_7772,N_2774,N_399);
nand U7773 (N_7773,N_1886,N_2295);
nor U7774 (N_7774,N_339,N_3139);
nor U7775 (N_7775,N_2283,N_2586);
and U7776 (N_7776,N_3534,N_3017);
and U7777 (N_7777,N_2445,N_2622);
nand U7778 (N_7778,N_3440,N_4807);
nand U7779 (N_7779,N_4807,N_599);
nor U7780 (N_7780,N_644,N_4010);
and U7781 (N_7781,N_3043,N_4762);
nand U7782 (N_7782,N_3425,N_1336);
xnor U7783 (N_7783,N_3920,N_998);
xnor U7784 (N_7784,N_3251,N_4715);
nand U7785 (N_7785,N_2720,N_4149);
nand U7786 (N_7786,N_692,N_4432);
xor U7787 (N_7787,N_1319,N_2563);
xnor U7788 (N_7788,N_661,N_1071);
or U7789 (N_7789,N_3295,N_301);
nand U7790 (N_7790,N_2811,N_3864);
nand U7791 (N_7791,N_4968,N_214);
or U7792 (N_7792,N_3803,N_3475);
nand U7793 (N_7793,N_4183,N_4662);
and U7794 (N_7794,N_1686,N_1315);
nor U7795 (N_7795,N_30,N_3496);
or U7796 (N_7796,N_2945,N_504);
nand U7797 (N_7797,N_3778,N_1555);
nor U7798 (N_7798,N_4223,N_2577);
or U7799 (N_7799,N_1703,N_3943);
and U7800 (N_7800,N_3794,N_2605);
xnor U7801 (N_7801,N_2819,N_3151);
xor U7802 (N_7802,N_165,N_2716);
nor U7803 (N_7803,N_554,N_2700);
nor U7804 (N_7804,N_2078,N_1280);
nand U7805 (N_7805,N_4122,N_3537);
and U7806 (N_7806,N_884,N_1909);
and U7807 (N_7807,N_1004,N_2984);
nand U7808 (N_7808,N_421,N_821);
nor U7809 (N_7809,N_383,N_63);
or U7810 (N_7810,N_3826,N_4618);
or U7811 (N_7811,N_1495,N_871);
and U7812 (N_7812,N_4485,N_1103);
or U7813 (N_7813,N_4253,N_4492);
or U7814 (N_7814,N_685,N_2725);
and U7815 (N_7815,N_4187,N_2508);
nor U7816 (N_7816,N_3407,N_3559);
nand U7817 (N_7817,N_1092,N_2419);
xnor U7818 (N_7818,N_4063,N_66);
nand U7819 (N_7819,N_510,N_97);
or U7820 (N_7820,N_3424,N_3821);
or U7821 (N_7821,N_4143,N_583);
nor U7822 (N_7822,N_670,N_1189);
nor U7823 (N_7823,N_3482,N_1227);
or U7824 (N_7824,N_3321,N_588);
nor U7825 (N_7825,N_4891,N_3450);
or U7826 (N_7826,N_4114,N_757);
xor U7827 (N_7827,N_2821,N_1015);
or U7828 (N_7828,N_2538,N_3634);
or U7829 (N_7829,N_1792,N_1316);
or U7830 (N_7830,N_2869,N_995);
nor U7831 (N_7831,N_2314,N_223);
or U7832 (N_7832,N_3251,N_792);
xnor U7833 (N_7833,N_142,N_4972);
or U7834 (N_7834,N_3317,N_15);
nand U7835 (N_7835,N_863,N_4843);
and U7836 (N_7836,N_1576,N_1942);
nor U7837 (N_7837,N_648,N_1406);
or U7838 (N_7838,N_575,N_3218);
nand U7839 (N_7839,N_2850,N_4127);
and U7840 (N_7840,N_4571,N_835);
or U7841 (N_7841,N_3538,N_1348);
or U7842 (N_7842,N_4081,N_4492);
nand U7843 (N_7843,N_51,N_3022);
xor U7844 (N_7844,N_4601,N_3848);
nand U7845 (N_7845,N_2659,N_279);
or U7846 (N_7846,N_1142,N_3303);
nor U7847 (N_7847,N_3028,N_1645);
nor U7848 (N_7848,N_4460,N_3320);
xnor U7849 (N_7849,N_1853,N_3533);
nor U7850 (N_7850,N_1087,N_671);
and U7851 (N_7851,N_3899,N_4674);
nor U7852 (N_7852,N_1869,N_2118);
and U7853 (N_7853,N_4431,N_4980);
nand U7854 (N_7854,N_1351,N_702);
and U7855 (N_7855,N_3889,N_4556);
or U7856 (N_7856,N_95,N_2128);
or U7857 (N_7857,N_1033,N_1890);
xnor U7858 (N_7858,N_774,N_3209);
xor U7859 (N_7859,N_4468,N_4597);
nor U7860 (N_7860,N_254,N_1431);
nand U7861 (N_7861,N_1167,N_1234);
xor U7862 (N_7862,N_3412,N_3744);
nand U7863 (N_7863,N_3872,N_4241);
and U7864 (N_7864,N_3250,N_4318);
and U7865 (N_7865,N_1344,N_2260);
or U7866 (N_7866,N_3680,N_3606);
nand U7867 (N_7867,N_4549,N_91);
or U7868 (N_7868,N_479,N_2322);
nand U7869 (N_7869,N_60,N_4407);
or U7870 (N_7870,N_654,N_2306);
or U7871 (N_7871,N_3367,N_4641);
or U7872 (N_7872,N_2132,N_3265);
and U7873 (N_7873,N_2204,N_4478);
nor U7874 (N_7874,N_1731,N_323);
nand U7875 (N_7875,N_1901,N_3623);
nor U7876 (N_7876,N_3524,N_698);
and U7877 (N_7877,N_4580,N_314);
nor U7878 (N_7878,N_2510,N_4450);
nor U7879 (N_7879,N_3010,N_2838);
nand U7880 (N_7880,N_1078,N_3579);
xor U7881 (N_7881,N_3043,N_1770);
or U7882 (N_7882,N_2692,N_3901);
nor U7883 (N_7883,N_2703,N_2457);
and U7884 (N_7884,N_2415,N_3338);
or U7885 (N_7885,N_1019,N_2389);
nor U7886 (N_7886,N_388,N_2338);
xnor U7887 (N_7887,N_1347,N_3875);
and U7888 (N_7888,N_1124,N_534);
and U7889 (N_7889,N_558,N_4734);
and U7890 (N_7890,N_3873,N_3351);
nand U7891 (N_7891,N_4909,N_2904);
and U7892 (N_7892,N_1688,N_1697);
and U7893 (N_7893,N_2343,N_1362);
nor U7894 (N_7894,N_547,N_468);
xor U7895 (N_7895,N_187,N_3039);
xor U7896 (N_7896,N_1075,N_2412);
nand U7897 (N_7897,N_3260,N_4757);
or U7898 (N_7898,N_1237,N_1947);
or U7899 (N_7899,N_4775,N_2454);
xor U7900 (N_7900,N_677,N_2908);
nor U7901 (N_7901,N_2514,N_1346);
or U7902 (N_7902,N_2003,N_1504);
nand U7903 (N_7903,N_2199,N_1476);
xor U7904 (N_7904,N_3377,N_1296);
and U7905 (N_7905,N_4298,N_462);
or U7906 (N_7906,N_4943,N_952);
and U7907 (N_7907,N_238,N_159);
xnor U7908 (N_7908,N_3318,N_3776);
nor U7909 (N_7909,N_4146,N_2279);
and U7910 (N_7910,N_3514,N_2998);
xnor U7911 (N_7911,N_2458,N_1936);
xnor U7912 (N_7912,N_1503,N_2138);
xnor U7913 (N_7913,N_1449,N_1893);
or U7914 (N_7914,N_3024,N_1682);
nor U7915 (N_7915,N_4481,N_1848);
and U7916 (N_7916,N_4562,N_1148);
nand U7917 (N_7917,N_4694,N_1585);
nand U7918 (N_7918,N_4967,N_3700);
and U7919 (N_7919,N_1310,N_3097);
nor U7920 (N_7920,N_3807,N_3912);
xnor U7921 (N_7921,N_540,N_2382);
or U7922 (N_7922,N_196,N_3383);
nor U7923 (N_7923,N_3750,N_2234);
nor U7924 (N_7924,N_3001,N_4286);
or U7925 (N_7925,N_1142,N_2736);
or U7926 (N_7926,N_3877,N_779);
xnor U7927 (N_7927,N_4996,N_3705);
nand U7928 (N_7928,N_4077,N_3387);
nor U7929 (N_7929,N_481,N_4388);
nand U7930 (N_7930,N_3853,N_3541);
and U7931 (N_7931,N_1272,N_4142);
and U7932 (N_7932,N_447,N_3116);
xnor U7933 (N_7933,N_1709,N_2114);
xnor U7934 (N_7934,N_3322,N_3812);
nor U7935 (N_7935,N_3365,N_3803);
and U7936 (N_7936,N_1282,N_3731);
or U7937 (N_7937,N_2229,N_435);
nand U7938 (N_7938,N_4298,N_1510);
or U7939 (N_7939,N_3601,N_4959);
nor U7940 (N_7940,N_4987,N_4634);
nor U7941 (N_7941,N_3570,N_3835);
nand U7942 (N_7942,N_3148,N_2907);
or U7943 (N_7943,N_352,N_4209);
or U7944 (N_7944,N_1398,N_3383);
or U7945 (N_7945,N_2508,N_3172);
and U7946 (N_7946,N_757,N_3208);
and U7947 (N_7947,N_4433,N_2088);
and U7948 (N_7948,N_1616,N_994);
nand U7949 (N_7949,N_1527,N_4471);
nand U7950 (N_7950,N_3327,N_711);
or U7951 (N_7951,N_84,N_2406);
and U7952 (N_7952,N_908,N_1529);
nand U7953 (N_7953,N_2999,N_1568);
or U7954 (N_7954,N_854,N_3243);
and U7955 (N_7955,N_2500,N_1838);
xor U7956 (N_7956,N_1410,N_4876);
xnor U7957 (N_7957,N_694,N_2396);
and U7958 (N_7958,N_265,N_4055);
xor U7959 (N_7959,N_2440,N_3951);
nor U7960 (N_7960,N_3153,N_1564);
and U7961 (N_7961,N_1198,N_141);
xnor U7962 (N_7962,N_4184,N_1904);
or U7963 (N_7963,N_157,N_1936);
xor U7964 (N_7964,N_155,N_4261);
nor U7965 (N_7965,N_1283,N_2188);
nand U7966 (N_7966,N_1795,N_1849);
nand U7967 (N_7967,N_4128,N_1908);
nand U7968 (N_7968,N_4723,N_1699);
xor U7969 (N_7969,N_2205,N_1204);
and U7970 (N_7970,N_786,N_4174);
xnor U7971 (N_7971,N_4395,N_4647);
nand U7972 (N_7972,N_3905,N_1113);
nand U7973 (N_7973,N_438,N_3902);
and U7974 (N_7974,N_2889,N_950);
or U7975 (N_7975,N_2703,N_4281);
xnor U7976 (N_7976,N_4718,N_4722);
nand U7977 (N_7977,N_2097,N_4942);
or U7978 (N_7978,N_4388,N_1718);
nor U7979 (N_7979,N_4621,N_970);
nand U7980 (N_7980,N_4447,N_3422);
nor U7981 (N_7981,N_3658,N_1772);
nand U7982 (N_7982,N_3648,N_1613);
or U7983 (N_7983,N_572,N_3105);
nor U7984 (N_7984,N_658,N_4327);
nand U7985 (N_7985,N_1015,N_4664);
nand U7986 (N_7986,N_4153,N_1922);
nor U7987 (N_7987,N_4418,N_3330);
or U7988 (N_7988,N_3930,N_4821);
xnor U7989 (N_7989,N_1507,N_4688);
nand U7990 (N_7990,N_1415,N_952);
and U7991 (N_7991,N_1990,N_3647);
nor U7992 (N_7992,N_1683,N_2105);
nor U7993 (N_7993,N_4499,N_438);
or U7994 (N_7994,N_154,N_4576);
nand U7995 (N_7995,N_2713,N_146);
nor U7996 (N_7996,N_2350,N_2906);
xor U7997 (N_7997,N_1586,N_1911);
or U7998 (N_7998,N_66,N_141);
xor U7999 (N_7999,N_3827,N_3325);
nor U8000 (N_8000,N_18,N_2813);
nand U8001 (N_8001,N_2714,N_3137);
xnor U8002 (N_8002,N_4545,N_988);
nand U8003 (N_8003,N_2538,N_2074);
nor U8004 (N_8004,N_4239,N_1259);
xor U8005 (N_8005,N_3324,N_4019);
xnor U8006 (N_8006,N_605,N_2017);
nand U8007 (N_8007,N_1176,N_1619);
nand U8008 (N_8008,N_1940,N_3955);
or U8009 (N_8009,N_960,N_3873);
or U8010 (N_8010,N_3598,N_4825);
and U8011 (N_8011,N_240,N_4249);
and U8012 (N_8012,N_641,N_4412);
nand U8013 (N_8013,N_4478,N_3657);
or U8014 (N_8014,N_4734,N_4992);
xor U8015 (N_8015,N_4388,N_4510);
xnor U8016 (N_8016,N_1381,N_2959);
nor U8017 (N_8017,N_3170,N_512);
and U8018 (N_8018,N_2949,N_402);
or U8019 (N_8019,N_312,N_4783);
xor U8020 (N_8020,N_2288,N_1310);
xnor U8021 (N_8021,N_4565,N_4259);
nor U8022 (N_8022,N_221,N_72);
nand U8023 (N_8023,N_918,N_4597);
and U8024 (N_8024,N_4499,N_4960);
or U8025 (N_8025,N_3277,N_3209);
or U8026 (N_8026,N_698,N_1490);
or U8027 (N_8027,N_4358,N_124);
and U8028 (N_8028,N_1197,N_2937);
or U8029 (N_8029,N_4628,N_4953);
and U8030 (N_8030,N_3460,N_1552);
nand U8031 (N_8031,N_1380,N_544);
nor U8032 (N_8032,N_493,N_4202);
and U8033 (N_8033,N_96,N_954);
xor U8034 (N_8034,N_2413,N_2837);
and U8035 (N_8035,N_4904,N_571);
or U8036 (N_8036,N_703,N_2068);
or U8037 (N_8037,N_603,N_1834);
and U8038 (N_8038,N_1531,N_344);
and U8039 (N_8039,N_3503,N_190);
or U8040 (N_8040,N_1786,N_185);
nand U8041 (N_8041,N_2935,N_775);
or U8042 (N_8042,N_2468,N_3942);
nor U8043 (N_8043,N_2936,N_1273);
and U8044 (N_8044,N_1915,N_691);
xnor U8045 (N_8045,N_1007,N_999);
xor U8046 (N_8046,N_1720,N_2665);
xor U8047 (N_8047,N_1654,N_1619);
and U8048 (N_8048,N_4288,N_4333);
and U8049 (N_8049,N_4492,N_2204);
and U8050 (N_8050,N_1313,N_3250);
and U8051 (N_8051,N_327,N_4419);
xor U8052 (N_8052,N_918,N_2620);
nor U8053 (N_8053,N_179,N_3855);
nand U8054 (N_8054,N_1411,N_1630);
and U8055 (N_8055,N_425,N_3357);
and U8056 (N_8056,N_817,N_3450);
or U8057 (N_8057,N_4352,N_3745);
xnor U8058 (N_8058,N_2709,N_2963);
or U8059 (N_8059,N_3292,N_1739);
or U8060 (N_8060,N_3449,N_1639);
xnor U8061 (N_8061,N_1029,N_2841);
xor U8062 (N_8062,N_2057,N_732);
nand U8063 (N_8063,N_4828,N_2527);
or U8064 (N_8064,N_3909,N_4527);
nor U8065 (N_8065,N_4010,N_500);
nor U8066 (N_8066,N_2944,N_930);
nor U8067 (N_8067,N_1538,N_3666);
xor U8068 (N_8068,N_717,N_698);
or U8069 (N_8069,N_2814,N_1279);
nor U8070 (N_8070,N_3493,N_4330);
nand U8071 (N_8071,N_4050,N_1893);
nand U8072 (N_8072,N_1744,N_2783);
or U8073 (N_8073,N_2459,N_531);
nand U8074 (N_8074,N_4990,N_4326);
and U8075 (N_8075,N_51,N_87);
and U8076 (N_8076,N_2601,N_96);
or U8077 (N_8077,N_4294,N_3576);
xor U8078 (N_8078,N_247,N_1435);
and U8079 (N_8079,N_346,N_4838);
xor U8080 (N_8080,N_1496,N_4740);
and U8081 (N_8081,N_3789,N_1591);
nand U8082 (N_8082,N_2517,N_3702);
or U8083 (N_8083,N_1330,N_305);
and U8084 (N_8084,N_4130,N_2773);
nand U8085 (N_8085,N_4691,N_820);
and U8086 (N_8086,N_539,N_889);
and U8087 (N_8087,N_2151,N_3276);
nand U8088 (N_8088,N_1829,N_4458);
and U8089 (N_8089,N_3760,N_338);
nand U8090 (N_8090,N_2223,N_3987);
nor U8091 (N_8091,N_3335,N_3249);
and U8092 (N_8092,N_1058,N_4296);
xnor U8093 (N_8093,N_2440,N_1156);
xnor U8094 (N_8094,N_1883,N_2030);
or U8095 (N_8095,N_2610,N_502);
xor U8096 (N_8096,N_4077,N_3822);
or U8097 (N_8097,N_3759,N_2130);
and U8098 (N_8098,N_2399,N_3261);
nand U8099 (N_8099,N_2687,N_288);
nand U8100 (N_8100,N_3096,N_78);
and U8101 (N_8101,N_3711,N_2866);
and U8102 (N_8102,N_114,N_4758);
nand U8103 (N_8103,N_3554,N_502);
and U8104 (N_8104,N_1278,N_4652);
or U8105 (N_8105,N_2723,N_3092);
and U8106 (N_8106,N_4080,N_263);
nand U8107 (N_8107,N_623,N_219);
nor U8108 (N_8108,N_3746,N_1584);
and U8109 (N_8109,N_169,N_2207);
or U8110 (N_8110,N_1649,N_3217);
nor U8111 (N_8111,N_4093,N_4783);
nor U8112 (N_8112,N_4851,N_4937);
or U8113 (N_8113,N_1353,N_1640);
and U8114 (N_8114,N_4862,N_3479);
or U8115 (N_8115,N_2479,N_4976);
or U8116 (N_8116,N_4560,N_4641);
or U8117 (N_8117,N_2031,N_4741);
nand U8118 (N_8118,N_29,N_3563);
nand U8119 (N_8119,N_1984,N_330);
nand U8120 (N_8120,N_3056,N_2384);
or U8121 (N_8121,N_1545,N_498);
xor U8122 (N_8122,N_4134,N_168);
and U8123 (N_8123,N_3057,N_4375);
or U8124 (N_8124,N_3932,N_2147);
nor U8125 (N_8125,N_4566,N_4650);
xnor U8126 (N_8126,N_4717,N_2472);
xnor U8127 (N_8127,N_188,N_2326);
and U8128 (N_8128,N_3882,N_1704);
and U8129 (N_8129,N_3376,N_313);
and U8130 (N_8130,N_2244,N_1113);
xor U8131 (N_8131,N_1408,N_1266);
xnor U8132 (N_8132,N_2609,N_1006);
nor U8133 (N_8133,N_1134,N_720);
or U8134 (N_8134,N_3722,N_4606);
nand U8135 (N_8135,N_1817,N_3348);
nor U8136 (N_8136,N_1162,N_4337);
xnor U8137 (N_8137,N_3677,N_2620);
xor U8138 (N_8138,N_1335,N_2638);
and U8139 (N_8139,N_3007,N_2131);
and U8140 (N_8140,N_3360,N_4231);
nor U8141 (N_8141,N_3265,N_4513);
nand U8142 (N_8142,N_4632,N_1673);
or U8143 (N_8143,N_3060,N_1406);
nor U8144 (N_8144,N_4171,N_1173);
xnor U8145 (N_8145,N_929,N_206);
or U8146 (N_8146,N_2885,N_1114);
and U8147 (N_8147,N_3560,N_2638);
and U8148 (N_8148,N_3984,N_142);
and U8149 (N_8149,N_1773,N_3772);
and U8150 (N_8150,N_977,N_3951);
and U8151 (N_8151,N_3414,N_163);
and U8152 (N_8152,N_4240,N_742);
nand U8153 (N_8153,N_4151,N_2834);
or U8154 (N_8154,N_1801,N_3786);
xnor U8155 (N_8155,N_4622,N_4511);
nor U8156 (N_8156,N_4089,N_3881);
and U8157 (N_8157,N_4155,N_4484);
and U8158 (N_8158,N_1588,N_3123);
nand U8159 (N_8159,N_4456,N_789);
or U8160 (N_8160,N_1688,N_2103);
nand U8161 (N_8161,N_3912,N_4393);
nand U8162 (N_8162,N_3030,N_2447);
nand U8163 (N_8163,N_4798,N_2088);
and U8164 (N_8164,N_2538,N_2089);
xor U8165 (N_8165,N_365,N_4029);
xnor U8166 (N_8166,N_1765,N_3497);
nor U8167 (N_8167,N_1814,N_2531);
nor U8168 (N_8168,N_3336,N_3180);
or U8169 (N_8169,N_2011,N_3178);
nor U8170 (N_8170,N_3945,N_731);
and U8171 (N_8171,N_1767,N_3995);
nor U8172 (N_8172,N_1826,N_1581);
xor U8173 (N_8173,N_3808,N_3982);
and U8174 (N_8174,N_2338,N_1356);
nor U8175 (N_8175,N_1574,N_2446);
or U8176 (N_8176,N_4688,N_551);
and U8177 (N_8177,N_3281,N_2265);
xor U8178 (N_8178,N_4854,N_4452);
nand U8179 (N_8179,N_4388,N_3535);
or U8180 (N_8180,N_3713,N_3430);
and U8181 (N_8181,N_4258,N_2035);
nor U8182 (N_8182,N_1091,N_3327);
and U8183 (N_8183,N_355,N_2465);
xnor U8184 (N_8184,N_804,N_244);
nand U8185 (N_8185,N_375,N_2477);
nand U8186 (N_8186,N_1760,N_528);
and U8187 (N_8187,N_1268,N_4087);
and U8188 (N_8188,N_2672,N_4564);
nor U8189 (N_8189,N_4609,N_3049);
and U8190 (N_8190,N_4061,N_3231);
or U8191 (N_8191,N_2267,N_3942);
nor U8192 (N_8192,N_4572,N_3845);
nand U8193 (N_8193,N_3174,N_4333);
xnor U8194 (N_8194,N_3431,N_3274);
or U8195 (N_8195,N_4480,N_3751);
or U8196 (N_8196,N_3082,N_4221);
and U8197 (N_8197,N_4667,N_3253);
nand U8198 (N_8198,N_2428,N_4826);
and U8199 (N_8199,N_4130,N_1344);
nand U8200 (N_8200,N_948,N_3819);
xor U8201 (N_8201,N_680,N_4027);
xor U8202 (N_8202,N_414,N_4728);
nand U8203 (N_8203,N_811,N_4393);
and U8204 (N_8204,N_4333,N_222);
nor U8205 (N_8205,N_1150,N_793);
xnor U8206 (N_8206,N_1032,N_1769);
nor U8207 (N_8207,N_1074,N_4652);
or U8208 (N_8208,N_1277,N_3869);
and U8209 (N_8209,N_3369,N_1751);
nand U8210 (N_8210,N_635,N_1401);
xnor U8211 (N_8211,N_544,N_2737);
or U8212 (N_8212,N_2361,N_1333);
nand U8213 (N_8213,N_2860,N_253);
nand U8214 (N_8214,N_2934,N_2787);
and U8215 (N_8215,N_1353,N_2535);
nor U8216 (N_8216,N_2405,N_3217);
xnor U8217 (N_8217,N_4320,N_4136);
or U8218 (N_8218,N_4536,N_244);
and U8219 (N_8219,N_1071,N_4759);
or U8220 (N_8220,N_680,N_486);
nor U8221 (N_8221,N_639,N_3354);
or U8222 (N_8222,N_1751,N_626);
or U8223 (N_8223,N_1591,N_3975);
nor U8224 (N_8224,N_4068,N_3332);
or U8225 (N_8225,N_1131,N_246);
or U8226 (N_8226,N_2858,N_557);
or U8227 (N_8227,N_4111,N_4811);
and U8228 (N_8228,N_2568,N_3697);
xor U8229 (N_8229,N_3686,N_4427);
nand U8230 (N_8230,N_1668,N_4188);
or U8231 (N_8231,N_983,N_4039);
or U8232 (N_8232,N_1448,N_1485);
nand U8233 (N_8233,N_2727,N_1538);
or U8234 (N_8234,N_232,N_4592);
nand U8235 (N_8235,N_3927,N_4315);
nand U8236 (N_8236,N_4841,N_1459);
nand U8237 (N_8237,N_1040,N_4310);
nor U8238 (N_8238,N_3530,N_1920);
xnor U8239 (N_8239,N_1693,N_4948);
xor U8240 (N_8240,N_4818,N_739);
nand U8241 (N_8241,N_1441,N_3816);
xnor U8242 (N_8242,N_1601,N_353);
xnor U8243 (N_8243,N_1994,N_1210);
xnor U8244 (N_8244,N_595,N_1823);
nor U8245 (N_8245,N_4812,N_1473);
or U8246 (N_8246,N_1244,N_1666);
and U8247 (N_8247,N_2708,N_2726);
nand U8248 (N_8248,N_2198,N_61);
nand U8249 (N_8249,N_4228,N_2255);
or U8250 (N_8250,N_748,N_4856);
nand U8251 (N_8251,N_805,N_3213);
xor U8252 (N_8252,N_3221,N_516);
nand U8253 (N_8253,N_4427,N_14);
nand U8254 (N_8254,N_2215,N_4857);
xnor U8255 (N_8255,N_4373,N_3721);
nand U8256 (N_8256,N_4059,N_142);
xor U8257 (N_8257,N_4369,N_2217);
xnor U8258 (N_8258,N_975,N_3621);
nor U8259 (N_8259,N_3410,N_4319);
or U8260 (N_8260,N_3624,N_3988);
or U8261 (N_8261,N_3535,N_3099);
nand U8262 (N_8262,N_3633,N_2831);
and U8263 (N_8263,N_3391,N_4708);
or U8264 (N_8264,N_181,N_1146);
nand U8265 (N_8265,N_2111,N_4514);
nand U8266 (N_8266,N_4683,N_4228);
nor U8267 (N_8267,N_381,N_3939);
or U8268 (N_8268,N_999,N_684);
nand U8269 (N_8269,N_4991,N_3024);
and U8270 (N_8270,N_1512,N_1370);
nor U8271 (N_8271,N_2400,N_1547);
or U8272 (N_8272,N_3909,N_2256);
and U8273 (N_8273,N_3539,N_1538);
xor U8274 (N_8274,N_2569,N_2109);
nor U8275 (N_8275,N_2607,N_823);
nand U8276 (N_8276,N_3445,N_4933);
xor U8277 (N_8277,N_574,N_2066);
and U8278 (N_8278,N_1311,N_4826);
and U8279 (N_8279,N_2271,N_2425);
nor U8280 (N_8280,N_283,N_2782);
nand U8281 (N_8281,N_4463,N_4744);
xnor U8282 (N_8282,N_4454,N_2223);
and U8283 (N_8283,N_4466,N_1322);
xnor U8284 (N_8284,N_357,N_1072);
or U8285 (N_8285,N_3557,N_1550);
nand U8286 (N_8286,N_113,N_1363);
xnor U8287 (N_8287,N_3271,N_204);
nor U8288 (N_8288,N_3312,N_3780);
xnor U8289 (N_8289,N_4845,N_2961);
xnor U8290 (N_8290,N_1396,N_478);
or U8291 (N_8291,N_2941,N_2994);
xnor U8292 (N_8292,N_1201,N_325);
xor U8293 (N_8293,N_4550,N_2540);
or U8294 (N_8294,N_2551,N_2861);
nor U8295 (N_8295,N_3344,N_769);
and U8296 (N_8296,N_666,N_2007);
xnor U8297 (N_8297,N_4709,N_518);
or U8298 (N_8298,N_2862,N_4540);
xor U8299 (N_8299,N_4305,N_1531);
and U8300 (N_8300,N_2013,N_4841);
nand U8301 (N_8301,N_1224,N_243);
xnor U8302 (N_8302,N_1868,N_3028);
or U8303 (N_8303,N_4298,N_975);
nand U8304 (N_8304,N_1972,N_1311);
nand U8305 (N_8305,N_864,N_1111);
and U8306 (N_8306,N_616,N_3600);
and U8307 (N_8307,N_4688,N_1727);
nor U8308 (N_8308,N_969,N_3164);
nor U8309 (N_8309,N_3530,N_1357);
or U8310 (N_8310,N_3650,N_984);
xnor U8311 (N_8311,N_2183,N_972);
or U8312 (N_8312,N_4324,N_3367);
xnor U8313 (N_8313,N_3795,N_4471);
or U8314 (N_8314,N_4160,N_1492);
or U8315 (N_8315,N_4646,N_1312);
nand U8316 (N_8316,N_3162,N_962);
and U8317 (N_8317,N_4570,N_586);
nor U8318 (N_8318,N_1736,N_2867);
or U8319 (N_8319,N_400,N_3045);
nor U8320 (N_8320,N_3912,N_3367);
nor U8321 (N_8321,N_3680,N_3205);
or U8322 (N_8322,N_2423,N_4711);
nor U8323 (N_8323,N_3170,N_392);
nand U8324 (N_8324,N_3433,N_3250);
nand U8325 (N_8325,N_609,N_105);
or U8326 (N_8326,N_2844,N_2165);
or U8327 (N_8327,N_2182,N_2820);
and U8328 (N_8328,N_3053,N_2391);
nand U8329 (N_8329,N_4588,N_3604);
or U8330 (N_8330,N_4441,N_723);
nand U8331 (N_8331,N_53,N_511);
and U8332 (N_8332,N_9,N_4632);
xor U8333 (N_8333,N_4174,N_1046);
nand U8334 (N_8334,N_1873,N_4576);
xnor U8335 (N_8335,N_3880,N_4087);
and U8336 (N_8336,N_807,N_4717);
nand U8337 (N_8337,N_134,N_4639);
or U8338 (N_8338,N_1501,N_920);
nor U8339 (N_8339,N_4917,N_950);
nand U8340 (N_8340,N_2555,N_1289);
and U8341 (N_8341,N_4755,N_1323);
or U8342 (N_8342,N_76,N_67);
and U8343 (N_8343,N_2959,N_3004);
xnor U8344 (N_8344,N_178,N_780);
nor U8345 (N_8345,N_2848,N_3359);
xor U8346 (N_8346,N_4261,N_3001);
xor U8347 (N_8347,N_3483,N_739);
xnor U8348 (N_8348,N_4102,N_2190);
nand U8349 (N_8349,N_4684,N_2505);
nand U8350 (N_8350,N_1838,N_1774);
or U8351 (N_8351,N_4781,N_4971);
xor U8352 (N_8352,N_822,N_1753);
nand U8353 (N_8353,N_879,N_638);
nand U8354 (N_8354,N_1405,N_83);
nor U8355 (N_8355,N_3642,N_1781);
nand U8356 (N_8356,N_1572,N_4657);
and U8357 (N_8357,N_286,N_4442);
nand U8358 (N_8358,N_344,N_3144);
or U8359 (N_8359,N_3531,N_2997);
and U8360 (N_8360,N_1513,N_3915);
nand U8361 (N_8361,N_2796,N_4086);
nand U8362 (N_8362,N_677,N_2744);
and U8363 (N_8363,N_2032,N_2);
xnor U8364 (N_8364,N_4816,N_1743);
xor U8365 (N_8365,N_4710,N_4715);
xor U8366 (N_8366,N_326,N_4376);
or U8367 (N_8367,N_509,N_2507);
or U8368 (N_8368,N_2504,N_1531);
nand U8369 (N_8369,N_4301,N_1181);
nor U8370 (N_8370,N_4591,N_569);
and U8371 (N_8371,N_1524,N_937);
or U8372 (N_8372,N_2875,N_3254);
or U8373 (N_8373,N_4401,N_872);
xor U8374 (N_8374,N_3345,N_3786);
or U8375 (N_8375,N_3484,N_2722);
nand U8376 (N_8376,N_4889,N_2126);
nor U8377 (N_8377,N_3771,N_3606);
nor U8378 (N_8378,N_2425,N_2435);
or U8379 (N_8379,N_1167,N_3634);
nand U8380 (N_8380,N_334,N_1582);
and U8381 (N_8381,N_1365,N_4881);
nor U8382 (N_8382,N_2962,N_2154);
xor U8383 (N_8383,N_3303,N_458);
nor U8384 (N_8384,N_711,N_3036);
xor U8385 (N_8385,N_3874,N_3245);
and U8386 (N_8386,N_4432,N_4410);
nand U8387 (N_8387,N_3733,N_3365);
nor U8388 (N_8388,N_3335,N_851);
xor U8389 (N_8389,N_3438,N_4357);
nor U8390 (N_8390,N_890,N_1475);
or U8391 (N_8391,N_315,N_4551);
xor U8392 (N_8392,N_4734,N_3612);
and U8393 (N_8393,N_1301,N_1204);
nand U8394 (N_8394,N_4851,N_1348);
nor U8395 (N_8395,N_3158,N_2094);
or U8396 (N_8396,N_2434,N_1664);
or U8397 (N_8397,N_4189,N_4237);
nand U8398 (N_8398,N_3521,N_21);
nand U8399 (N_8399,N_1175,N_4155);
and U8400 (N_8400,N_3053,N_1546);
nor U8401 (N_8401,N_4138,N_3086);
or U8402 (N_8402,N_260,N_4550);
nor U8403 (N_8403,N_1316,N_3050);
nand U8404 (N_8404,N_4615,N_962);
nand U8405 (N_8405,N_4621,N_3134);
or U8406 (N_8406,N_4051,N_5);
nor U8407 (N_8407,N_3369,N_4196);
or U8408 (N_8408,N_4532,N_2077);
and U8409 (N_8409,N_3194,N_4098);
and U8410 (N_8410,N_1082,N_911);
or U8411 (N_8411,N_4388,N_1630);
or U8412 (N_8412,N_4896,N_2738);
nor U8413 (N_8413,N_626,N_2346);
nor U8414 (N_8414,N_322,N_722);
nand U8415 (N_8415,N_4245,N_3703);
nand U8416 (N_8416,N_4111,N_4173);
nand U8417 (N_8417,N_4348,N_2380);
nor U8418 (N_8418,N_4741,N_3595);
and U8419 (N_8419,N_2911,N_3176);
or U8420 (N_8420,N_3149,N_4741);
xnor U8421 (N_8421,N_1711,N_971);
xor U8422 (N_8422,N_1657,N_4921);
or U8423 (N_8423,N_2082,N_305);
and U8424 (N_8424,N_3415,N_1621);
or U8425 (N_8425,N_500,N_2603);
nand U8426 (N_8426,N_2276,N_2018);
or U8427 (N_8427,N_1746,N_3645);
nand U8428 (N_8428,N_4557,N_3821);
xnor U8429 (N_8429,N_4420,N_2294);
nor U8430 (N_8430,N_387,N_4543);
nor U8431 (N_8431,N_4531,N_1373);
xor U8432 (N_8432,N_4581,N_3815);
xnor U8433 (N_8433,N_4324,N_3453);
xnor U8434 (N_8434,N_4959,N_1392);
or U8435 (N_8435,N_817,N_3683);
or U8436 (N_8436,N_2007,N_2522);
and U8437 (N_8437,N_110,N_238);
nand U8438 (N_8438,N_4161,N_1699);
nor U8439 (N_8439,N_4093,N_4000);
or U8440 (N_8440,N_2696,N_4230);
nor U8441 (N_8441,N_3062,N_872);
xnor U8442 (N_8442,N_4953,N_1590);
xor U8443 (N_8443,N_1322,N_1757);
nand U8444 (N_8444,N_4212,N_2735);
nand U8445 (N_8445,N_3049,N_1219);
and U8446 (N_8446,N_1336,N_3778);
nor U8447 (N_8447,N_1941,N_1515);
nand U8448 (N_8448,N_3519,N_501);
xor U8449 (N_8449,N_1852,N_10);
nand U8450 (N_8450,N_2357,N_289);
xor U8451 (N_8451,N_4672,N_3225);
nor U8452 (N_8452,N_2880,N_3762);
or U8453 (N_8453,N_3414,N_3035);
and U8454 (N_8454,N_1651,N_666);
nand U8455 (N_8455,N_4798,N_4229);
xnor U8456 (N_8456,N_943,N_2793);
or U8457 (N_8457,N_565,N_84);
xnor U8458 (N_8458,N_4160,N_2254);
and U8459 (N_8459,N_1030,N_186);
or U8460 (N_8460,N_3508,N_2823);
or U8461 (N_8461,N_3373,N_3751);
and U8462 (N_8462,N_427,N_4864);
nor U8463 (N_8463,N_4803,N_1335);
or U8464 (N_8464,N_4068,N_3324);
and U8465 (N_8465,N_4758,N_1827);
and U8466 (N_8466,N_2870,N_10);
and U8467 (N_8467,N_2422,N_80);
or U8468 (N_8468,N_2864,N_4567);
nor U8469 (N_8469,N_3416,N_2581);
and U8470 (N_8470,N_817,N_2128);
nor U8471 (N_8471,N_313,N_4468);
or U8472 (N_8472,N_350,N_900);
and U8473 (N_8473,N_4737,N_1649);
or U8474 (N_8474,N_3558,N_2165);
xnor U8475 (N_8475,N_4707,N_2993);
nor U8476 (N_8476,N_2942,N_4929);
and U8477 (N_8477,N_4048,N_2126);
xor U8478 (N_8478,N_2885,N_2872);
and U8479 (N_8479,N_1306,N_3947);
or U8480 (N_8480,N_1348,N_4228);
and U8481 (N_8481,N_2543,N_239);
and U8482 (N_8482,N_4409,N_603);
and U8483 (N_8483,N_199,N_4061);
xnor U8484 (N_8484,N_438,N_2236);
xnor U8485 (N_8485,N_3892,N_1538);
xnor U8486 (N_8486,N_464,N_1775);
and U8487 (N_8487,N_2387,N_79);
and U8488 (N_8488,N_77,N_4765);
xor U8489 (N_8489,N_2559,N_2659);
xor U8490 (N_8490,N_1464,N_1242);
or U8491 (N_8491,N_110,N_3300);
or U8492 (N_8492,N_3423,N_4755);
or U8493 (N_8493,N_4285,N_1910);
xor U8494 (N_8494,N_148,N_573);
nand U8495 (N_8495,N_45,N_4226);
xor U8496 (N_8496,N_2384,N_1772);
and U8497 (N_8497,N_2869,N_1387);
and U8498 (N_8498,N_1126,N_1782);
nand U8499 (N_8499,N_578,N_3708);
nand U8500 (N_8500,N_3732,N_3124);
xnor U8501 (N_8501,N_4894,N_1502);
and U8502 (N_8502,N_3426,N_1197);
nor U8503 (N_8503,N_3635,N_4917);
nand U8504 (N_8504,N_944,N_2296);
nor U8505 (N_8505,N_2927,N_3861);
xnor U8506 (N_8506,N_1204,N_4565);
nand U8507 (N_8507,N_4794,N_87);
xnor U8508 (N_8508,N_2056,N_4618);
nor U8509 (N_8509,N_37,N_2537);
or U8510 (N_8510,N_637,N_518);
nand U8511 (N_8511,N_3078,N_2);
xor U8512 (N_8512,N_4137,N_4244);
nor U8513 (N_8513,N_4025,N_4271);
and U8514 (N_8514,N_2856,N_2773);
nor U8515 (N_8515,N_1212,N_1262);
and U8516 (N_8516,N_2574,N_422);
xor U8517 (N_8517,N_2894,N_1809);
xnor U8518 (N_8518,N_726,N_3228);
and U8519 (N_8519,N_982,N_3163);
xor U8520 (N_8520,N_3867,N_4256);
nand U8521 (N_8521,N_471,N_2717);
nor U8522 (N_8522,N_3421,N_569);
nand U8523 (N_8523,N_3803,N_1818);
xor U8524 (N_8524,N_2827,N_4265);
nor U8525 (N_8525,N_1236,N_1540);
nor U8526 (N_8526,N_2091,N_3320);
or U8527 (N_8527,N_2344,N_564);
nand U8528 (N_8528,N_831,N_4613);
nor U8529 (N_8529,N_3670,N_1636);
nor U8530 (N_8530,N_2404,N_2773);
nand U8531 (N_8531,N_2054,N_821);
and U8532 (N_8532,N_800,N_297);
and U8533 (N_8533,N_2788,N_1008);
or U8534 (N_8534,N_3047,N_382);
or U8535 (N_8535,N_905,N_4683);
nand U8536 (N_8536,N_3914,N_4586);
nand U8537 (N_8537,N_2960,N_1888);
nor U8538 (N_8538,N_3397,N_4013);
nor U8539 (N_8539,N_4851,N_2307);
nor U8540 (N_8540,N_2997,N_614);
or U8541 (N_8541,N_1166,N_2479);
nor U8542 (N_8542,N_3228,N_840);
and U8543 (N_8543,N_3980,N_4711);
xor U8544 (N_8544,N_4722,N_2950);
xor U8545 (N_8545,N_1482,N_2633);
nand U8546 (N_8546,N_3344,N_1070);
xor U8547 (N_8547,N_2690,N_4417);
and U8548 (N_8548,N_4763,N_1689);
xnor U8549 (N_8549,N_4458,N_4828);
nor U8550 (N_8550,N_857,N_2918);
xnor U8551 (N_8551,N_2764,N_4020);
and U8552 (N_8552,N_1664,N_2681);
nand U8553 (N_8553,N_3934,N_2384);
and U8554 (N_8554,N_2226,N_1649);
nor U8555 (N_8555,N_4703,N_4965);
and U8556 (N_8556,N_3243,N_1766);
nand U8557 (N_8557,N_943,N_34);
and U8558 (N_8558,N_4422,N_608);
and U8559 (N_8559,N_1060,N_4797);
and U8560 (N_8560,N_867,N_2982);
and U8561 (N_8561,N_4161,N_4497);
or U8562 (N_8562,N_679,N_2894);
and U8563 (N_8563,N_438,N_3151);
nand U8564 (N_8564,N_2617,N_963);
nor U8565 (N_8565,N_2137,N_2389);
and U8566 (N_8566,N_1891,N_2306);
and U8567 (N_8567,N_4525,N_4245);
nor U8568 (N_8568,N_3966,N_2171);
nor U8569 (N_8569,N_4100,N_4494);
or U8570 (N_8570,N_2707,N_1024);
nor U8571 (N_8571,N_174,N_4809);
and U8572 (N_8572,N_540,N_313);
or U8573 (N_8573,N_3702,N_2023);
or U8574 (N_8574,N_4377,N_4302);
or U8575 (N_8575,N_905,N_2348);
nor U8576 (N_8576,N_3688,N_1564);
nand U8577 (N_8577,N_36,N_3873);
nor U8578 (N_8578,N_2190,N_2974);
nand U8579 (N_8579,N_754,N_3765);
nand U8580 (N_8580,N_1947,N_947);
nor U8581 (N_8581,N_2838,N_2537);
or U8582 (N_8582,N_2470,N_622);
nand U8583 (N_8583,N_294,N_1575);
and U8584 (N_8584,N_3938,N_2493);
or U8585 (N_8585,N_4109,N_4558);
and U8586 (N_8586,N_988,N_1707);
nor U8587 (N_8587,N_4800,N_1820);
xor U8588 (N_8588,N_2931,N_1170);
nand U8589 (N_8589,N_905,N_2249);
nand U8590 (N_8590,N_3018,N_442);
or U8591 (N_8591,N_4344,N_206);
nand U8592 (N_8592,N_282,N_1189);
xnor U8593 (N_8593,N_234,N_3871);
xnor U8594 (N_8594,N_1946,N_122);
nand U8595 (N_8595,N_3074,N_544);
and U8596 (N_8596,N_2237,N_3972);
nand U8597 (N_8597,N_3203,N_1131);
or U8598 (N_8598,N_3354,N_2046);
nor U8599 (N_8599,N_3088,N_239);
nand U8600 (N_8600,N_190,N_1715);
and U8601 (N_8601,N_1582,N_1354);
nor U8602 (N_8602,N_1589,N_607);
nand U8603 (N_8603,N_2059,N_3453);
or U8604 (N_8604,N_129,N_1032);
xnor U8605 (N_8605,N_945,N_3127);
or U8606 (N_8606,N_206,N_4996);
nor U8607 (N_8607,N_3194,N_2137);
nand U8608 (N_8608,N_3669,N_511);
and U8609 (N_8609,N_95,N_2937);
or U8610 (N_8610,N_900,N_981);
xor U8611 (N_8611,N_1282,N_4045);
xnor U8612 (N_8612,N_1705,N_1926);
nor U8613 (N_8613,N_3116,N_1995);
and U8614 (N_8614,N_640,N_3302);
and U8615 (N_8615,N_3294,N_1207);
xnor U8616 (N_8616,N_3886,N_2931);
xor U8617 (N_8617,N_3947,N_3291);
and U8618 (N_8618,N_2966,N_3475);
xor U8619 (N_8619,N_2542,N_4524);
xor U8620 (N_8620,N_1249,N_4845);
xnor U8621 (N_8621,N_3807,N_266);
or U8622 (N_8622,N_1751,N_1015);
and U8623 (N_8623,N_1408,N_2110);
nor U8624 (N_8624,N_254,N_2619);
or U8625 (N_8625,N_1032,N_3146);
nand U8626 (N_8626,N_2653,N_1783);
or U8627 (N_8627,N_3877,N_4100);
nand U8628 (N_8628,N_1282,N_4570);
nor U8629 (N_8629,N_2888,N_2666);
and U8630 (N_8630,N_3845,N_306);
nand U8631 (N_8631,N_2410,N_2514);
and U8632 (N_8632,N_1622,N_3625);
xnor U8633 (N_8633,N_3944,N_3633);
nor U8634 (N_8634,N_1627,N_1667);
or U8635 (N_8635,N_1096,N_1155);
nand U8636 (N_8636,N_3440,N_3902);
or U8637 (N_8637,N_1663,N_2741);
nand U8638 (N_8638,N_1176,N_2961);
nor U8639 (N_8639,N_487,N_2113);
xor U8640 (N_8640,N_3290,N_3063);
and U8641 (N_8641,N_2099,N_1248);
nor U8642 (N_8642,N_4757,N_2865);
xor U8643 (N_8643,N_2169,N_3997);
nand U8644 (N_8644,N_4799,N_3407);
nand U8645 (N_8645,N_3375,N_2105);
nor U8646 (N_8646,N_4321,N_1690);
nand U8647 (N_8647,N_3462,N_1380);
xnor U8648 (N_8648,N_1439,N_1205);
xnor U8649 (N_8649,N_2662,N_3355);
xnor U8650 (N_8650,N_2676,N_3059);
nand U8651 (N_8651,N_3358,N_1890);
xnor U8652 (N_8652,N_1368,N_2874);
and U8653 (N_8653,N_4687,N_205);
xor U8654 (N_8654,N_2571,N_548);
xor U8655 (N_8655,N_1764,N_4335);
and U8656 (N_8656,N_149,N_2013);
and U8657 (N_8657,N_1667,N_4247);
nand U8658 (N_8658,N_4401,N_2423);
xor U8659 (N_8659,N_4655,N_2647);
and U8660 (N_8660,N_3520,N_367);
xnor U8661 (N_8661,N_1660,N_3176);
nor U8662 (N_8662,N_4585,N_694);
and U8663 (N_8663,N_499,N_487);
nor U8664 (N_8664,N_3772,N_3327);
xnor U8665 (N_8665,N_1591,N_1499);
xor U8666 (N_8666,N_4939,N_3114);
xor U8667 (N_8667,N_2035,N_4746);
and U8668 (N_8668,N_1002,N_3548);
and U8669 (N_8669,N_262,N_1301);
nor U8670 (N_8670,N_1523,N_3411);
and U8671 (N_8671,N_627,N_3058);
nor U8672 (N_8672,N_709,N_408);
xnor U8673 (N_8673,N_1061,N_1587);
xor U8674 (N_8674,N_3784,N_632);
xnor U8675 (N_8675,N_1235,N_1400);
nor U8676 (N_8676,N_3482,N_1215);
xor U8677 (N_8677,N_3329,N_3506);
nor U8678 (N_8678,N_4773,N_1512);
xnor U8679 (N_8679,N_4882,N_663);
or U8680 (N_8680,N_4784,N_4344);
or U8681 (N_8681,N_791,N_4659);
nand U8682 (N_8682,N_152,N_3844);
or U8683 (N_8683,N_1419,N_2857);
or U8684 (N_8684,N_98,N_1956);
nand U8685 (N_8685,N_4162,N_910);
or U8686 (N_8686,N_3197,N_1914);
or U8687 (N_8687,N_4593,N_4334);
and U8688 (N_8688,N_2094,N_1575);
and U8689 (N_8689,N_3325,N_2069);
nand U8690 (N_8690,N_4487,N_1434);
nor U8691 (N_8691,N_4620,N_526);
and U8692 (N_8692,N_472,N_1568);
nand U8693 (N_8693,N_2189,N_3104);
nand U8694 (N_8694,N_2432,N_3165);
and U8695 (N_8695,N_4431,N_975);
nand U8696 (N_8696,N_4480,N_1003);
xnor U8697 (N_8697,N_1888,N_2583);
nand U8698 (N_8698,N_1707,N_4898);
nor U8699 (N_8699,N_311,N_4084);
or U8700 (N_8700,N_3962,N_3155);
nor U8701 (N_8701,N_2347,N_272);
xnor U8702 (N_8702,N_4405,N_4463);
xnor U8703 (N_8703,N_378,N_1079);
nand U8704 (N_8704,N_4246,N_177);
and U8705 (N_8705,N_4481,N_626);
nand U8706 (N_8706,N_4730,N_967);
nor U8707 (N_8707,N_4645,N_2801);
xor U8708 (N_8708,N_3501,N_2712);
nand U8709 (N_8709,N_4027,N_4569);
nand U8710 (N_8710,N_952,N_4103);
xor U8711 (N_8711,N_3704,N_2510);
nor U8712 (N_8712,N_2161,N_2350);
xnor U8713 (N_8713,N_3068,N_1292);
nor U8714 (N_8714,N_1109,N_3572);
xnor U8715 (N_8715,N_1245,N_249);
nor U8716 (N_8716,N_3239,N_3935);
xor U8717 (N_8717,N_2997,N_435);
or U8718 (N_8718,N_995,N_4723);
and U8719 (N_8719,N_2867,N_2813);
or U8720 (N_8720,N_3278,N_3081);
or U8721 (N_8721,N_144,N_2450);
xor U8722 (N_8722,N_3590,N_4008);
nand U8723 (N_8723,N_3420,N_2546);
and U8724 (N_8724,N_4509,N_1078);
and U8725 (N_8725,N_2587,N_4341);
xnor U8726 (N_8726,N_4886,N_2477);
or U8727 (N_8727,N_1857,N_2012);
xnor U8728 (N_8728,N_4616,N_3924);
nor U8729 (N_8729,N_2653,N_3956);
and U8730 (N_8730,N_1249,N_2861);
nor U8731 (N_8731,N_3966,N_2073);
nand U8732 (N_8732,N_2233,N_2853);
nor U8733 (N_8733,N_3578,N_3619);
or U8734 (N_8734,N_4878,N_4072);
nor U8735 (N_8735,N_4071,N_2672);
xnor U8736 (N_8736,N_329,N_2873);
nand U8737 (N_8737,N_4426,N_3009);
and U8738 (N_8738,N_2424,N_3352);
nor U8739 (N_8739,N_4328,N_1031);
and U8740 (N_8740,N_3726,N_313);
xor U8741 (N_8741,N_3955,N_842);
nand U8742 (N_8742,N_637,N_1199);
nor U8743 (N_8743,N_1327,N_2055);
or U8744 (N_8744,N_1489,N_2081);
nand U8745 (N_8745,N_910,N_4904);
or U8746 (N_8746,N_2592,N_2013);
xor U8747 (N_8747,N_2751,N_4084);
nor U8748 (N_8748,N_4018,N_4538);
nand U8749 (N_8749,N_3724,N_2994);
and U8750 (N_8750,N_2324,N_3996);
nand U8751 (N_8751,N_3738,N_1791);
nor U8752 (N_8752,N_1827,N_3162);
xnor U8753 (N_8753,N_510,N_2880);
or U8754 (N_8754,N_633,N_1432);
xnor U8755 (N_8755,N_3022,N_1423);
nor U8756 (N_8756,N_2768,N_3996);
nor U8757 (N_8757,N_4759,N_3136);
nand U8758 (N_8758,N_117,N_3148);
and U8759 (N_8759,N_2532,N_2339);
and U8760 (N_8760,N_768,N_3690);
nand U8761 (N_8761,N_4013,N_4111);
xor U8762 (N_8762,N_2764,N_1930);
and U8763 (N_8763,N_3814,N_324);
or U8764 (N_8764,N_3740,N_806);
nor U8765 (N_8765,N_2952,N_354);
nor U8766 (N_8766,N_3212,N_4831);
and U8767 (N_8767,N_3233,N_2774);
nor U8768 (N_8768,N_1961,N_4958);
nor U8769 (N_8769,N_2975,N_880);
nand U8770 (N_8770,N_614,N_3947);
nand U8771 (N_8771,N_2849,N_4390);
or U8772 (N_8772,N_3978,N_554);
and U8773 (N_8773,N_3489,N_4921);
nand U8774 (N_8774,N_635,N_1513);
nor U8775 (N_8775,N_868,N_1221);
nand U8776 (N_8776,N_1798,N_928);
nand U8777 (N_8777,N_666,N_4392);
nor U8778 (N_8778,N_2684,N_531);
nand U8779 (N_8779,N_2282,N_3895);
xor U8780 (N_8780,N_1007,N_4993);
nor U8781 (N_8781,N_1907,N_3103);
nand U8782 (N_8782,N_3830,N_3011);
or U8783 (N_8783,N_780,N_2801);
nand U8784 (N_8784,N_1653,N_4976);
nand U8785 (N_8785,N_3262,N_2086);
nand U8786 (N_8786,N_4814,N_4214);
and U8787 (N_8787,N_3981,N_2915);
xor U8788 (N_8788,N_1406,N_2746);
nor U8789 (N_8789,N_412,N_2653);
or U8790 (N_8790,N_4581,N_1468);
and U8791 (N_8791,N_4495,N_39);
or U8792 (N_8792,N_2573,N_4760);
nand U8793 (N_8793,N_2757,N_1646);
or U8794 (N_8794,N_666,N_3433);
nand U8795 (N_8795,N_1176,N_1415);
nand U8796 (N_8796,N_4790,N_3462);
xnor U8797 (N_8797,N_851,N_1961);
nor U8798 (N_8798,N_3152,N_2776);
and U8799 (N_8799,N_4379,N_4452);
nor U8800 (N_8800,N_4336,N_1876);
nor U8801 (N_8801,N_2471,N_1545);
or U8802 (N_8802,N_3613,N_4410);
or U8803 (N_8803,N_4815,N_4149);
and U8804 (N_8804,N_1379,N_4192);
xnor U8805 (N_8805,N_3513,N_3436);
and U8806 (N_8806,N_660,N_119);
xnor U8807 (N_8807,N_1753,N_3009);
nor U8808 (N_8808,N_1493,N_100);
nor U8809 (N_8809,N_471,N_176);
nor U8810 (N_8810,N_1966,N_3185);
xor U8811 (N_8811,N_1949,N_4133);
nor U8812 (N_8812,N_2496,N_1669);
and U8813 (N_8813,N_4121,N_3881);
xor U8814 (N_8814,N_8,N_1111);
nand U8815 (N_8815,N_3238,N_4903);
nand U8816 (N_8816,N_904,N_227);
or U8817 (N_8817,N_2551,N_980);
xnor U8818 (N_8818,N_2030,N_4526);
nand U8819 (N_8819,N_1684,N_3492);
nor U8820 (N_8820,N_3293,N_4898);
and U8821 (N_8821,N_4106,N_1417);
xor U8822 (N_8822,N_3576,N_4242);
nor U8823 (N_8823,N_3124,N_714);
or U8824 (N_8824,N_3165,N_4636);
nand U8825 (N_8825,N_1716,N_179);
nor U8826 (N_8826,N_231,N_3558);
nor U8827 (N_8827,N_4411,N_2864);
or U8828 (N_8828,N_1028,N_4495);
and U8829 (N_8829,N_4741,N_2254);
or U8830 (N_8830,N_1581,N_115);
nor U8831 (N_8831,N_3117,N_4990);
and U8832 (N_8832,N_1315,N_803);
or U8833 (N_8833,N_3140,N_4552);
xor U8834 (N_8834,N_1049,N_1324);
xor U8835 (N_8835,N_4574,N_3148);
xor U8836 (N_8836,N_546,N_1580);
or U8837 (N_8837,N_4184,N_1419);
nor U8838 (N_8838,N_3971,N_832);
or U8839 (N_8839,N_598,N_4089);
or U8840 (N_8840,N_4398,N_2110);
and U8841 (N_8841,N_4755,N_4939);
or U8842 (N_8842,N_3016,N_3928);
nand U8843 (N_8843,N_867,N_2533);
nor U8844 (N_8844,N_224,N_3432);
or U8845 (N_8845,N_2070,N_2531);
nor U8846 (N_8846,N_3742,N_2667);
xnor U8847 (N_8847,N_4849,N_1007);
or U8848 (N_8848,N_4152,N_3895);
or U8849 (N_8849,N_4469,N_635);
or U8850 (N_8850,N_2223,N_3933);
xnor U8851 (N_8851,N_2018,N_1794);
xnor U8852 (N_8852,N_4103,N_1336);
nand U8853 (N_8853,N_1576,N_4985);
xnor U8854 (N_8854,N_2686,N_4957);
xor U8855 (N_8855,N_1083,N_1538);
xnor U8856 (N_8856,N_4819,N_4639);
and U8857 (N_8857,N_692,N_1345);
nand U8858 (N_8858,N_2699,N_355);
nand U8859 (N_8859,N_2021,N_4178);
xor U8860 (N_8860,N_1844,N_4108);
nand U8861 (N_8861,N_2218,N_1317);
nand U8862 (N_8862,N_2532,N_3381);
nor U8863 (N_8863,N_4647,N_450);
nor U8864 (N_8864,N_3336,N_3079);
xor U8865 (N_8865,N_503,N_3313);
xnor U8866 (N_8866,N_1064,N_206);
nor U8867 (N_8867,N_346,N_2076);
or U8868 (N_8868,N_4702,N_467);
nand U8869 (N_8869,N_4058,N_2175);
nand U8870 (N_8870,N_4276,N_924);
xnor U8871 (N_8871,N_3094,N_1405);
xnor U8872 (N_8872,N_1528,N_1629);
and U8873 (N_8873,N_870,N_4741);
xor U8874 (N_8874,N_1070,N_3506);
or U8875 (N_8875,N_3899,N_2624);
nand U8876 (N_8876,N_1415,N_1162);
nand U8877 (N_8877,N_1931,N_3649);
xor U8878 (N_8878,N_3203,N_4073);
nand U8879 (N_8879,N_834,N_2005);
or U8880 (N_8880,N_4943,N_1399);
nor U8881 (N_8881,N_1169,N_4781);
or U8882 (N_8882,N_2779,N_1058);
nand U8883 (N_8883,N_4442,N_1754);
or U8884 (N_8884,N_4776,N_953);
nor U8885 (N_8885,N_1291,N_4593);
nand U8886 (N_8886,N_2454,N_3638);
nand U8887 (N_8887,N_2806,N_3161);
and U8888 (N_8888,N_1576,N_3165);
and U8889 (N_8889,N_1834,N_4360);
and U8890 (N_8890,N_2231,N_1627);
or U8891 (N_8891,N_1311,N_4140);
xnor U8892 (N_8892,N_1337,N_4689);
and U8893 (N_8893,N_84,N_4875);
nor U8894 (N_8894,N_883,N_235);
nand U8895 (N_8895,N_1610,N_2914);
nand U8896 (N_8896,N_3027,N_4164);
nor U8897 (N_8897,N_4385,N_99);
and U8898 (N_8898,N_3122,N_3237);
nand U8899 (N_8899,N_108,N_390);
and U8900 (N_8900,N_3529,N_4935);
and U8901 (N_8901,N_942,N_4954);
xnor U8902 (N_8902,N_2795,N_4450);
xnor U8903 (N_8903,N_3968,N_378);
nand U8904 (N_8904,N_1560,N_4654);
and U8905 (N_8905,N_1580,N_3679);
or U8906 (N_8906,N_1515,N_2511);
or U8907 (N_8907,N_1707,N_701);
nand U8908 (N_8908,N_3809,N_3847);
xor U8909 (N_8909,N_3645,N_3306);
nor U8910 (N_8910,N_365,N_3531);
nand U8911 (N_8911,N_3794,N_558);
nand U8912 (N_8912,N_2643,N_4837);
xnor U8913 (N_8913,N_4551,N_2626);
and U8914 (N_8914,N_823,N_2868);
nand U8915 (N_8915,N_4140,N_3054);
or U8916 (N_8916,N_4007,N_4248);
nor U8917 (N_8917,N_4729,N_3663);
and U8918 (N_8918,N_3391,N_1663);
nor U8919 (N_8919,N_2309,N_353);
xor U8920 (N_8920,N_1849,N_3422);
or U8921 (N_8921,N_4976,N_3522);
xor U8922 (N_8922,N_746,N_3347);
and U8923 (N_8923,N_4626,N_2194);
nor U8924 (N_8924,N_1921,N_411);
nand U8925 (N_8925,N_153,N_3610);
xnor U8926 (N_8926,N_1810,N_2941);
or U8927 (N_8927,N_4500,N_2900);
or U8928 (N_8928,N_353,N_908);
nor U8929 (N_8929,N_614,N_1208);
nand U8930 (N_8930,N_2849,N_726);
xnor U8931 (N_8931,N_4267,N_3896);
xor U8932 (N_8932,N_1295,N_1418);
xor U8933 (N_8933,N_2037,N_4411);
and U8934 (N_8934,N_1545,N_2149);
and U8935 (N_8935,N_4921,N_4833);
nor U8936 (N_8936,N_1299,N_4456);
nor U8937 (N_8937,N_287,N_267);
or U8938 (N_8938,N_2265,N_2680);
or U8939 (N_8939,N_1555,N_2845);
nand U8940 (N_8940,N_338,N_4258);
or U8941 (N_8941,N_175,N_2258);
or U8942 (N_8942,N_2850,N_3101);
nor U8943 (N_8943,N_4946,N_4437);
and U8944 (N_8944,N_466,N_1116);
nand U8945 (N_8945,N_2629,N_1719);
nor U8946 (N_8946,N_2426,N_263);
or U8947 (N_8947,N_1026,N_1518);
xnor U8948 (N_8948,N_2573,N_4414);
nor U8949 (N_8949,N_3672,N_140);
xnor U8950 (N_8950,N_2882,N_4465);
nand U8951 (N_8951,N_1867,N_1516);
and U8952 (N_8952,N_289,N_3703);
and U8953 (N_8953,N_432,N_2133);
nand U8954 (N_8954,N_2510,N_430);
or U8955 (N_8955,N_4718,N_4549);
and U8956 (N_8956,N_3423,N_553);
nand U8957 (N_8957,N_408,N_767);
xor U8958 (N_8958,N_1670,N_4188);
and U8959 (N_8959,N_2267,N_4821);
xnor U8960 (N_8960,N_2536,N_641);
nor U8961 (N_8961,N_129,N_4861);
or U8962 (N_8962,N_810,N_2002);
nor U8963 (N_8963,N_3425,N_2938);
and U8964 (N_8964,N_2855,N_2283);
nand U8965 (N_8965,N_4770,N_4988);
nand U8966 (N_8966,N_360,N_1273);
nor U8967 (N_8967,N_494,N_4062);
and U8968 (N_8968,N_4934,N_1411);
and U8969 (N_8969,N_3645,N_299);
xnor U8970 (N_8970,N_2293,N_1639);
and U8971 (N_8971,N_3548,N_2354);
or U8972 (N_8972,N_117,N_3296);
or U8973 (N_8973,N_1865,N_2055);
and U8974 (N_8974,N_1503,N_884);
or U8975 (N_8975,N_3778,N_1313);
xor U8976 (N_8976,N_2581,N_630);
or U8977 (N_8977,N_4039,N_1558);
nor U8978 (N_8978,N_2858,N_2355);
xor U8979 (N_8979,N_3022,N_2340);
or U8980 (N_8980,N_3645,N_858);
nand U8981 (N_8981,N_1411,N_374);
or U8982 (N_8982,N_2283,N_484);
and U8983 (N_8983,N_4369,N_1457);
and U8984 (N_8984,N_4834,N_136);
nor U8985 (N_8985,N_296,N_2249);
or U8986 (N_8986,N_2548,N_3448);
xnor U8987 (N_8987,N_3509,N_2744);
xnor U8988 (N_8988,N_3948,N_3003);
xor U8989 (N_8989,N_2596,N_1455);
nor U8990 (N_8990,N_4838,N_2250);
nor U8991 (N_8991,N_3544,N_3997);
nand U8992 (N_8992,N_906,N_2379);
nor U8993 (N_8993,N_1823,N_3796);
nor U8994 (N_8994,N_4354,N_667);
xnor U8995 (N_8995,N_2970,N_1215);
and U8996 (N_8996,N_537,N_3751);
nor U8997 (N_8997,N_1131,N_2962);
nand U8998 (N_8998,N_1877,N_4869);
nand U8999 (N_8999,N_2330,N_1890);
nand U9000 (N_9000,N_579,N_1070);
or U9001 (N_9001,N_4741,N_1720);
nand U9002 (N_9002,N_4903,N_1407);
xnor U9003 (N_9003,N_901,N_2323);
and U9004 (N_9004,N_3756,N_35);
nand U9005 (N_9005,N_1921,N_3729);
nand U9006 (N_9006,N_858,N_3782);
nand U9007 (N_9007,N_3648,N_3998);
nand U9008 (N_9008,N_3454,N_1562);
and U9009 (N_9009,N_4305,N_3138);
and U9010 (N_9010,N_3848,N_2464);
nand U9011 (N_9011,N_1964,N_2501);
xnor U9012 (N_9012,N_4632,N_4346);
xor U9013 (N_9013,N_188,N_2088);
xnor U9014 (N_9014,N_3002,N_811);
nor U9015 (N_9015,N_2209,N_3344);
nor U9016 (N_9016,N_3390,N_3795);
nand U9017 (N_9017,N_355,N_4742);
xor U9018 (N_9018,N_3991,N_1191);
nor U9019 (N_9019,N_2604,N_515);
xor U9020 (N_9020,N_2030,N_1728);
and U9021 (N_9021,N_1003,N_4402);
and U9022 (N_9022,N_4175,N_2772);
or U9023 (N_9023,N_400,N_135);
xor U9024 (N_9024,N_3862,N_4272);
xnor U9025 (N_9025,N_2470,N_3164);
and U9026 (N_9026,N_4780,N_3892);
or U9027 (N_9027,N_2981,N_3321);
or U9028 (N_9028,N_358,N_1923);
xnor U9029 (N_9029,N_850,N_1681);
or U9030 (N_9030,N_701,N_1651);
and U9031 (N_9031,N_4998,N_4605);
nor U9032 (N_9032,N_1493,N_4958);
xor U9033 (N_9033,N_313,N_4293);
or U9034 (N_9034,N_778,N_2592);
or U9035 (N_9035,N_2279,N_4509);
and U9036 (N_9036,N_2064,N_1501);
and U9037 (N_9037,N_4640,N_1699);
xor U9038 (N_9038,N_2210,N_1121);
or U9039 (N_9039,N_1494,N_510);
or U9040 (N_9040,N_1047,N_993);
and U9041 (N_9041,N_1195,N_3503);
or U9042 (N_9042,N_2717,N_2768);
or U9043 (N_9043,N_1287,N_901);
nand U9044 (N_9044,N_812,N_2246);
and U9045 (N_9045,N_2282,N_4032);
xnor U9046 (N_9046,N_1606,N_3167);
nor U9047 (N_9047,N_1030,N_845);
nand U9048 (N_9048,N_4011,N_469);
xor U9049 (N_9049,N_4515,N_978);
and U9050 (N_9050,N_52,N_3855);
or U9051 (N_9051,N_2154,N_3688);
and U9052 (N_9052,N_264,N_1041);
nand U9053 (N_9053,N_3103,N_3525);
nor U9054 (N_9054,N_1592,N_710);
or U9055 (N_9055,N_4336,N_2230);
nor U9056 (N_9056,N_34,N_3785);
nand U9057 (N_9057,N_1606,N_4456);
nand U9058 (N_9058,N_1938,N_4229);
and U9059 (N_9059,N_3788,N_1514);
nand U9060 (N_9060,N_3117,N_2144);
and U9061 (N_9061,N_3576,N_2213);
nor U9062 (N_9062,N_2298,N_223);
or U9063 (N_9063,N_3348,N_2003);
xor U9064 (N_9064,N_3253,N_3937);
or U9065 (N_9065,N_3909,N_3033);
nand U9066 (N_9066,N_393,N_522);
nand U9067 (N_9067,N_4731,N_2160);
nor U9068 (N_9068,N_980,N_1902);
nand U9069 (N_9069,N_895,N_3575);
nand U9070 (N_9070,N_1470,N_2281);
or U9071 (N_9071,N_1950,N_2206);
nand U9072 (N_9072,N_4162,N_2551);
and U9073 (N_9073,N_2282,N_971);
xor U9074 (N_9074,N_3595,N_4790);
xor U9075 (N_9075,N_1421,N_1966);
xor U9076 (N_9076,N_2343,N_2652);
nand U9077 (N_9077,N_2302,N_1188);
xor U9078 (N_9078,N_593,N_4207);
and U9079 (N_9079,N_450,N_1222);
nor U9080 (N_9080,N_4063,N_2465);
xor U9081 (N_9081,N_1888,N_2619);
xor U9082 (N_9082,N_2986,N_1174);
xnor U9083 (N_9083,N_1956,N_1389);
nor U9084 (N_9084,N_3965,N_3403);
xor U9085 (N_9085,N_2988,N_2057);
or U9086 (N_9086,N_977,N_915);
nand U9087 (N_9087,N_3244,N_4145);
and U9088 (N_9088,N_3247,N_3324);
and U9089 (N_9089,N_2835,N_4254);
xnor U9090 (N_9090,N_2138,N_3792);
and U9091 (N_9091,N_2466,N_899);
and U9092 (N_9092,N_860,N_326);
and U9093 (N_9093,N_2668,N_4799);
or U9094 (N_9094,N_1949,N_4911);
nand U9095 (N_9095,N_369,N_4550);
xor U9096 (N_9096,N_3539,N_3117);
nor U9097 (N_9097,N_4298,N_1017);
xnor U9098 (N_9098,N_4639,N_3165);
nor U9099 (N_9099,N_729,N_1657);
xnor U9100 (N_9100,N_2184,N_2246);
nor U9101 (N_9101,N_1893,N_2949);
nor U9102 (N_9102,N_3094,N_4320);
nand U9103 (N_9103,N_1092,N_4767);
xnor U9104 (N_9104,N_495,N_4239);
nand U9105 (N_9105,N_983,N_965);
and U9106 (N_9106,N_1592,N_1845);
xor U9107 (N_9107,N_2137,N_1706);
nand U9108 (N_9108,N_3064,N_2230);
nor U9109 (N_9109,N_2256,N_2975);
or U9110 (N_9110,N_1555,N_1001);
nor U9111 (N_9111,N_3340,N_3575);
or U9112 (N_9112,N_4995,N_1875);
nand U9113 (N_9113,N_2929,N_1095);
nand U9114 (N_9114,N_3064,N_4484);
or U9115 (N_9115,N_612,N_2157);
nand U9116 (N_9116,N_4365,N_4704);
nand U9117 (N_9117,N_1859,N_970);
and U9118 (N_9118,N_2848,N_2668);
xnor U9119 (N_9119,N_2944,N_1410);
nor U9120 (N_9120,N_3012,N_1898);
xor U9121 (N_9121,N_3353,N_1340);
nor U9122 (N_9122,N_2764,N_4791);
xnor U9123 (N_9123,N_4160,N_837);
nand U9124 (N_9124,N_1048,N_2001);
or U9125 (N_9125,N_3948,N_1474);
nor U9126 (N_9126,N_3272,N_3380);
nand U9127 (N_9127,N_4838,N_2085);
nor U9128 (N_9128,N_2330,N_4325);
nand U9129 (N_9129,N_91,N_4895);
or U9130 (N_9130,N_2129,N_3827);
and U9131 (N_9131,N_2759,N_1688);
and U9132 (N_9132,N_3748,N_4558);
nand U9133 (N_9133,N_1805,N_3407);
xor U9134 (N_9134,N_1357,N_3117);
and U9135 (N_9135,N_2533,N_2996);
nor U9136 (N_9136,N_1085,N_4270);
or U9137 (N_9137,N_4389,N_1814);
nor U9138 (N_9138,N_2676,N_4358);
xnor U9139 (N_9139,N_1779,N_3394);
nand U9140 (N_9140,N_4922,N_2433);
xor U9141 (N_9141,N_3497,N_2742);
or U9142 (N_9142,N_2320,N_1690);
or U9143 (N_9143,N_1880,N_209);
nand U9144 (N_9144,N_3180,N_583);
nand U9145 (N_9145,N_13,N_4859);
or U9146 (N_9146,N_1251,N_3064);
xnor U9147 (N_9147,N_2853,N_1603);
nor U9148 (N_9148,N_1054,N_3526);
and U9149 (N_9149,N_2300,N_4692);
nor U9150 (N_9150,N_4984,N_4128);
xor U9151 (N_9151,N_2078,N_4510);
nand U9152 (N_9152,N_1896,N_4527);
or U9153 (N_9153,N_4415,N_4140);
and U9154 (N_9154,N_2680,N_3703);
nor U9155 (N_9155,N_3427,N_3304);
or U9156 (N_9156,N_1630,N_2228);
or U9157 (N_9157,N_62,N_3418);
nor U9158 (N_9158,N_4933,N_2349);
or U9159 (N_9159,N_2304,N_2425);
and U9160 (N_9160,N_4192,N_3397);
nor U9161 (N_9161,N_2482,N_1330);
nor U9162 (N_9162,N_1802,N_2785);
nand U9163 (N_9163,N_2159,N_2605);
xnor U9164 (N_9164,N_2315,N_480);
nand U9165 (N_9165,N_2989,N_3567);
or U9166 (N_9166,N_3959,N_1532);
nand U9167 (N_9167,N_117,N_4723);
nand U9168 (N_9168,N_4159,N_4286);
or U9169 (N_9169,N_4816,N_3026);
xnor U9170 (N_9170,N_3718,N_421);
nor U9171 (N_9171,N_344,N_2746);
or U9172 (N_9172,N_3080,N_107);
nor U9173 (N_9173,N_4669,N_3232);
nor U9174 (N_9174,N_4683,N_2397);
or U9175 (N_9175,N_3464,N_3960);
and U9176 (N_9176,N_1684,N_242);
and U9177 (N_9177,N_1151,N_781);
nand U9178 (N_9178,N_1857,N_796);
nand U9179 (N_9179,N_2912,N_1967);
and U9180 (N_9180,N_4605,N_3843);
or U9181 (N_9181,N_1893,N_850);
xor U9182 (N_9182,N_3591,N_4320);
nand U9183 (N_9183,N_2407,N_4581);
nand U9184 (N_9184,N_1390,N_979);
xnor U9185 (N_9185,N_4276,N_4336);
xnor U9186 (N_9186,N_4293,N_2004);
nor U9187 (N_9187,N_556,N_3029);
xnor U9188 (N_9188,N_2529,N_1897);
nand U9189 (N_9189,N_4538,N_62);
nand U9190 (N_9190,N_3183,N_4343);
or U9191 (N_9191,N_954,N_4657);
xnor U9192 (N_9192,N_887,N_3111);
and U9193 (N_9193,N_4221,N_3599);
or U9194 (N_9194,N_1093,N_2634);
nor U9195 (N_9195,N_2286,N_3156);
xor U9196 (N_9196,N_3789,N_3921);
nor U9197 (N_9197,N_4413,N_3760);
nand U9198 (N_9198,N_3012,N_4561);
xnor U9199 (N_9199,N_99,N_2569);
or U9200 (N_9200,N_4401,N_4384);
and U9201 (N_9201,N_2847,N_1405);
and U9202 (N_9202,N_3712,N_4086);
xor U9203 (N_9203,N_2088,N_102);
nor U9204 (N_9204,N_2574,N_3241);
or U9205 (N_9205,N_1349,N_4042);
nand U9206 (N_9206,N_1278,N_486);
or U9207 (N_9207,N_4464,N_172);
nor U9208 (N_9208,N_3532,N_3280);
and U9209 (N_9209,N_2787,N_2220);
and U9210 (N_9210,N_3348,N_2692);
or U9211 (N_9211,N_1374,N_227);
nor U9212 (N_9212,N_3656,N_4438);
nor U9213 (N_9213,N_4293,N_2324);
nor U9214 (N_9214,N_4118,N_4019);
nor U9215 (N_9215,N_4769,N_2395);
xnor U9216 (N_9216,N_3000,N_1850);
xnor U9217 (N_9217,N_3474,N_1096);
or U9218 (N_9218,N_930,N_1591);
nand U9219 (N_9219,N_3379,N_64);
and U9220 (N_9220,N_778,N_4105);
nand U9221 (N_9221,N_3070,N_2701);
and U9222 (N_9222,N_1324,N_2363);
nand U9223 (N_9223,N_3904,N_2589);
or U9224 (N_9224,N_1462,N_3813);
nor U9225 (N_9225,N_1329,N_562);
xor U9226 (N_9226,N_226,N_2472);
or U9227 (N_9227,N_2750,N_2895);
or U9228 (N_9228,N_577,N_2763);
and U9229 (N_9229,N_89,N_4448);
nor U9230 (N_9230,N_3954,N_1199);
nor U9231 (N_9231,N_56,N_555);
or U9232 (N_9232,N_688,N_544);
nand U9233 (N_9233,N_4311,N_4142);
or U9234 (N_9234,N_3240,N_96);
nand U9235 (N_9235,N_4639,N_1097);
nand U9236 (N_9236,N_4535,N_4005);
or U9237 (N_9237,N_974,N_2406);
nor U9238 (N_9238,N_2559,N_2339);
or U9239 (N_9239,N_2807,N_2503);
and U9240 (N_9240,N_4373,N_483);
xnor U9241 (N_9241,N_904,N_2426);
xor U9242 (N_9242,N_2473,N_2143);
nor U9243 (N_9243,N_3089,N_3362);
nand U9244 (N_9244,N_1908,N_4441);
or U9245 (N_9245,N_799,N_3872);
nor U9246 (N_9246,N_3235,N_645);
nor U9247 (N_9247,N_3713,N_4662);
xnor U9248 (N_9248,N_4781,N_2941);
and U9249 (N_9249,N_960,N_3860);
nand U9250 (N_9250,N_2459,N_2696);
nand U9251 (N_9251,N_1091,N_666);
or U9252 (N_9252,N_3531,N_3159);
nand U9253 (N_9253,N_3639,N_3830);
or U9254 (N_9254,N_2440,N_2079);
xor U9255 (N_9255,N_330,N_2355);
nand U9256 (N_9256,N_1498,N_2029);
nor U9257 (N_9257,N_4359,N_3240);
nand U9258 (N_9258,N_2302,N_4020);
and U9259 (N_9259,N_4484,N_1648);
and U9260 (N_9260,N_4315,N_2152);
nand U9261 (N_9261,N_3115,N_3943);
or U9262 (N_9262,N_144,N_4502);
nand U9263 (N_9263,N_2251,N_1476);
and U9264 (N_9264,N_3895,N_4405);
nand U9265 (N_9265,N_1131,N_1216);
or U9266 (N_9266,N_2072,N_4460);
xor U9267 (N_9267,N_4968,N_4786);
or U9268 (N_9268,N_3158,N_755);
or U9269 (N_9269,N_965,N_2786);
nor U9270 (N_9270,N_1748,N_4514);
xor U9271 (N_9271,N_1963,N_689);
or U9272 (N_9272,N_2299,N_2981);
and U9273 (N_9273,N_3678,N_161);
and U9274 (N_9274,N_2281,N_4565);
and U9275 (N_9275,N_2325,N_2776);
nand U9276 (N_9276,N_3729,N_3132);
nor U9277 (N_9277,N_4035,N_1685);
nand U9278 (N_9278,N_1394,N_4654);
nand U9279 (N_9279,N_1643,N_1193);
nor U9280 (N_9280,N_1818,N_4915);
nand U9281 (N_9281,N_4319,N_2947);
xor U9282 (N_9282,N_3872,N_226);
nand U9283 (N_9283,N_1571,N_2633);
xnor U9284 (N_9284,N_4251,N_2200);
nand U9285 (N_9285,N_1494,N_4487);
nor U9286 (N_9286,N_1729,N_622);
or U9287 (N_9287,N_3947,N_4888);
nand U9288 (N_9288,N_954,N_3249);
nand U9289 (N_9289,N_770,N_2590);
nand U9290 (N_9290,N_568,N_4682);
nor U9291 (N_9291,N_117,N_900);
nor U9292 (N_9292,N_1511,N_3863);
nand U9293 (N_9293,N_2021,N_4978);
nor U9294 (N_9294,N_2520,N_3134);
nand U9295 (N_9295,N_992,N_2222);
nor U9296 (N_9296,N_635,N_3800);
xor U9297 (N_9297,N_2278,N_3034);
and U9298 (N_9298,N_1293,N_4030);
nand U9299 (N_9299,N_4033,N_2374);
nor U9300 (N_9300,N_3763,N_3987);
nand U9301 (N_9301,N_927,N_1725);
and U9302 (N_9302,N_3820,N_4134);
nand U9303 (N_9303,N_3133,N_2880);
xor U9304 (N_9304,N_1940,N_2742);
or U9305 (N_9305,N_3243,N_533);
xor U9306 (N_9306,N_1998,N_1065);
and U9307 (N_9307,N_67,N_4112);
and U9308 (N_9308,N_2704,N_1151);
nand U9309 (N_9309,N_3332,N_4782);
and U9310 (N_9310,N_455,N_1523);
nand U9311 (N_9311,N_1933,N_3838);
or U9312 (N_9312,N_3537,N_4674);
nand U9313 (N_9313,N_2676,N_1793);
and U9314 (N_9314,N_4231,N_3144);
and U9315 (N_9315,N_1493,N_1030);
xnor U9316 (N_9316,N_4130,N_3100);
and U9317 (N_9317,N_4759,N_1132);
xor U9318 (N_9318,N_1078,N_3055);
nor U9319 (N_9319,N_3245,N_3452);
nand U9320 (N_9320,N_1235,N_1664);
and U9321 (N_9321,N_3040,N_4359);
nor U9322 (N_9322,N_4837,N_2776);
or U9323 (N_9323,N_4956,N_2579);
and U9324 (N_9324,N_3848,N_3306);
and U9325 (N_9325,N_4887,N_2802);
xnor U9326 (N_9326,N_4843,N_223);
nor U9327 (N_9327,N_3126,N_897);
nand U9328 (N_9328,N_3486,N_2852);
and U9329 (N_9329,N_3651,N_2132);
or U9330 (N_9330,N_2382,N_2735);
xor U9331 (N_9331,N_2930,N_285);
and U9332 (N_9332,N_4537,N_787);
or U9333 (N_9333,N_4513,N_1281);
nand U9334 (N_9334,N_2511,N_643);
nor U9335 (N_9335,N_799,N_519);
or U9336 (N_9336,N_3831,N_1376);
xnor U9337 (N_9337,N_4867,N_757);
and U9338 (N_9338,N_3344,N_3632);
nor U9339 (N_9339,N_3571,N_2997);
nand U9340 (N_9340,N_1961,N_3087);
xor U9341 (N_9341,N_4713,N_1442);
and U9342 (N_9342,N_1048,N_1714);
or U9343 (N_9343,N_2663,N_1924);
xor U9344 (N_9344,N_3107,N_4366);
nand U9345 (N_9345,N_3127,N_3158);
nor U9346 (N_9346,N_1558,N_1192);
xnor U9347 (N_9347,N_4622,N_697);
or U9348 (N_9348,N_1313,N_4453);
nor U9349 (N_9349,N_1790,N_3436);
and U9350 (N_9350,N_3071,N_3724);
nand U9351 (N_9351,N_4003,N_589);
or U9352 (N_9352,N_4973,N_1423);
and U9353 (N_9353,N_266,N_2657);
nand U9354 (N_9354,N_4758,N_1141);
xnor U9355 (N_9355,N_1367,N_2961);
or U9356 (N_9356,N_2286,N_4271);
or U9357 (N_9357,N_1342,N_4767);
nand U9358 (N_9358,N_3864,N_4606);
or U9359 (N_9359,N_4539,N_37);
nor U9360 (N_9360,N_3452,N_3605);
or U9361 (N_9361,N_1163,N_3799);
nor U9362 (N_9362,N_4509,N_1294);
nand U9363 (N_9363,N_1494,N_3604);
nor U9364 (N_9364,N_3878,N_2138);
nor U9365 (N_9365,N_2944,N_2921);
xnor U9366 (N_9366,N_2138,N_1360);
or U9367 (N_9367,N_3147,N_694);
xnor U9368 (N_9368,N_4686,N_3469);
nor U9369 (N_9369,N_4337,N_813);
nand U9370 (N_9370,N_3737,N_3142);
or U9371 (N_9371,N_662,N_4462);
nand U9372 (N_9372,N_3601,N_1156);
or U9373 (N_9373,N_1058,N_2732);
xnor U9374 (N_9374,N_2718,N_2411);
nor U9375 (N_9375,N_1001,N_4430);
xor U9376 (N_9376,N_3545,N_3460);
and U9377 (N_9377,N_4564,N_1513);
nor U9378 (N_9378,N_1501,N_973);
xnor U9379 (N_9379,N_3644,N_763);
xnor U9380 (N_9380,N_1990,N_2698);
or U9381 (N_9381,N_277,N_578);
and U9382 (N_9382,N_4229,N_3997);
nand U9383 (N_9383,N_2239,N_2730);
or U9384 (N_9384,N_282,N_3268);
nor U9385 (N_9385,N_1552,N_2820);
nor U9386 (N_9386,N_1730,N_4419);
nor U9387 (N_9387,N_4848,N_437);
or U9388 (N_9388,N_4094,N_2640);
or U9389 (N_9389,N_2288,N_4861);
nor U9390 (N_9390,N_703,N_2478);
or U9391 (N_9391,N_1315,N_1611);
or U9392 (N_9392,N_880,N_4125);
xnor U9393 (N_9393,N_594,N_1377);
nor U9394 (N_9394,N_4245,N_942);
or U9395 (N_9395,N_2920,N_1817);
xnor U9396 (N_9396,N_2808,N_566);
nand U9397 (N_9397,N_802,N_3078);
nand U9398 (N_9398,N_4408,N_100);
nor U9399 (N_9399,N_2809,N_257);
and U9400 (N_9400,N_2690,N_2232);
nand U9401 (N_9401,N_2444,N_2602);
nand U9402 (N_9402,N_4670,N_3605);
nand U9403 (N_9403,N_679,N_3871);
nor U9404 (N_9404,N_584,N_2966);
nand U9405 (N_9405,N_415,N_4648);
xnor U9406 (N_9406,N_769,N_4305);
nand U9407 (N_9407,N_4080,N_377);
xor U9408 (N_9408,N_1162,N_4313);
or U9409 (N_9409,N_944,N_4083);
nor U9410 (N_9410,N_3698,N_2142);
or U9411 (N_9411,N_2381,N_3509);
nand U9412 (N_9412,N_2881,N_3521);
and U9413 (N_9413,N_3858,N_2191);
xnor U9414 (N_9414,N_1148,N_2000);
or U9415 (N_9415,N_4958,N_4706);
nor U9416 (N_9416,N_2854,N_894);
nor U9417 (N_9417,N_4685,N_694);
or U9418 (N_9418,N_3618,N_2249);
or U9419 (N_9419,N_1934,N_2535);
and U9420 (N_9420,N_3530,N_1946);
and U9421 (N_9421,N_1934,N_3422);
or U9422 (N_9422,N_3546,N_4004);
and U9423 (N_9423,N_2593,N_2194);
and U9424 (N_9424,N_2840,N_680);
nor U9425 (N_9425,N_4066,N_3694);
nor U9426 (N_9426,N_1930,N_2805);
or U9427 (N_9427,N_4819,N_2757);
nand U9428 (N_9428,N_1338,N_296);
and U9429 (N_9429,N_1838,N_1884);
or U9430 (N_9430,N_4576,N_3310);
nand U9431 (N_9431,N_2009,N_4527);
nor U9432 (N_9432,N_1753,N_81);
nor U9433 (N_9433,N_2453,N_1436);
nor U9434 (N_9434,N_1043,N_2972);
nand U9435 (N_9435,N_4376,N_1064);
nor U9436 (N_9436,N_3612,N_582);
and U9437 (N_9437,N_2065,N_4607);
xor U9438 (N_9438,N_3407,N_3904);
nor U9439 (N_9439,N_4956,N_3799);
and U9440 (N_9440,N_193,N_1094);
and U9441 (N_9441,N_1982,N_4375);
and U9442 (N_9442,N_1096,N_2549);
or U9443 (N_9443,N_4758,N_215);
xor U9444 (N_9444,N_159,N_3415);
or U9445 (N_9445,N_3320,N_4851);
and U9446 (N_9446,N_2064,N_2909);
and U9447 (N_9447,N_3433,N_1255);
nand U9448 (N_9448,N_3725,N_4786);
nand U9449 (N_9449,N_849,N_4032);
nor U9450 (N_9450,N_4568,N_1234);
nor U9451 (N_9451,N_591,N_2659);
xor U9452 (N_9452,N_555,N_4196);
nand U9453 (N_9453,N_967,N_1171);
xnor U9454 (N_9454,N_2269,N_2675);
xnor U9455 (N_9455,N_755,N_3427);
nand U9456 (N_9456,N_4601,N_4012);
nor U9457 (N_9457,N_2819,N_544);
nand U9458 (N_9458,N_2801,N_2351);
nand U9459 (N_9459,N_2800,N_1036);
xor U9460 (N_9460,N_4566,N_4811);
nor U9461 (N_9461,N_1550,N_1241);
nand U9462 (N_9462,N_2911,N_3731);
nand U9463 (N_9463,N_851,N_1203);
and U9464 (N_9464,N_784,N_474);
xnor U9465 (N_9465,N_4884,N_3195);
xnor U9466 (N_9466,N_1999,N_4650);
nand U9467 (N_9467,N_338,N_121);
and U9468 (N_9468,N_2805,N_4695);
nand U9469 (N_9469,N_1986,N_3935);
and U9470 (N_9470,N_3713,N_2317);
xor U9471 (N_9471,N_4547,N_4536);
nor U9472 (N_9472,N_4501,N_4559);
nand U9473 (N_9473,N_3640,N_1745);
nand U9474 (N_9474,N_3531,N_1026);
xnor U9475 (N_9475,N_1352,N_127);
or U9476 (N_9476,N_3075,N_3025);
nand U9477 (N_9477,N_4524,N_4827);
nor U9478 (N_9478,N_3490,N_4940);
nor U9479 (N_9479,N_3581,N_4002);
xnor U9480 (N_9480,N_398,N_4182);
or U9481 (N_9481,N_2123,N_1715);
nor U9482 (N_9482,N_3465,N_740);
xnor U9483 (N_9483,N_1829,N_3104);
or U9484 (N_9484,N_3947,N_678);
nor U9485 (N_9485,N_2412,N_475);
and U9486 (N_9486,N_1085,N_1694);
nor U9487 (N_9487,N_4091,N_1079);
or U9488 (N_9488,N_609,N_3084);
or U9489 (N_9489,N_1629,N_3282);
and U9490 (N_9490,N_1123,N_2093);
nand U9491 (N_9491,N_4303,N_172);
and U9492 (N_9492,N_3228,N_3123);
or U9493 (N_9493,N_1713,N_3339);
or U9494 (N_9494,N_1528,N_116);
nor U9495 (N_9495,N_4931,N_903);
and U9496 (N_9496,N_3331,N_211);
xnor U9497 (N_9497,N_3674,N_4320);
xor U9498 (N_9498,N_1253,N_4685);
or U9499 (N_9499,N_1178,N_53);
nor U9500 (N_9500,N_3931,N_641);
nand U9501 (N_9501,N_4834,N_4052);
or U9502 (N_9502,N_2916,N_257);
nor U9503 (N_9503,N_1897,N_3234);
nand U9504 (N_9504,N_4685,N_45);
nor U9505 (N_9505,N_2958,N_2176);
xnor U9506 (N_9506,N_365,N_2545);
xor U9507 (N_9507,N_3281,N_597);
nor U9508 (N_9508,N_4046,N_2988);
and U9509 (N_9509,N_2496,N_4044);
xor U9510 (N_9510,N_2646,N_1832);
xnor U9511 (N_9511,N_3022,N_3100);
nor U9512 (N_9512,N_3158,N_583);
or U9513 (N_9513,N_1670,N_2475);
or U9514 (N_9514,N_4094,N_4126);
xor U9515 (N_9515,N_569,N_4673);
xor U9516 (N_9516,N_4870,N_1485);
nor U9517 (N_9517,N_350,N_4017);
nand U9518 (N_9518,N_782,N_1051);
xnor U9519 (N_9519,N_1123,N_1748);
nor U9520 (N_9520,N_385,N_4957);
nor U9521 (N_9521,N_4822,N_2317);
and U9522 (N_9522,N_2387,N_3690);
nand U9523 (N_9523,N_1706,N_1645);
or U9524 (N_9524,N_2445,N_3767);
xor U9525 (N_9525,N_1087,N_4734);
nand U9526 (N_9526,N_1434,N_4581);
nor U9527 (N_9527,N_76,N_574);
nor U9528 (N_9528,N_2954,N_2613);
and U9529 (N_9529,N_3586,N_4190);
and U9530 (N_9530,N_3108,N_3287);
xor U9531 (N_9531,N_2911,N_917);
nor U9532 (N_9532,N_336,N_2392);
nor U9533 (N_9533,N_229,N_480);
xor U9534 (N_9534,N_2889,N_2845);
or U9535 (N_9535,N_2291,N_1996);
nand U9536 (N_9536,N_1085,N_4896);
nand U9537 (N_9537,N_4637,N_864);
or U9538 (N_9538,N_659,N_2585);
nor U9539 (N_9539,N_3253,N_767);
or U9540 (N_9540,N_4255,N_4978);
xor U9541 (N_9541,N_3445,N_100);
and U9542 (N_9542,N_2343,N_18);
xnor U9543 (N_9543,N_559,N_4316);
xor U9544 (N_9544,N_3207,N_1459);
nor U9545 (N_9545,N_3649,N_3651);
nand U9546 (N_9546,N_3592,N_4431);
and U9547 (N_9547,N_2642,N_2653);
and U9548 (N_9548,N_3098,N_4322);
nand U9549 (N_9549,N_4884,N_2631);
nor U9550 (N_9550,N_4713,N_4505);
nand U9551 (N_9551,N_4361,N_3518);
xor U9552 (N_9552,N_4712,N_73);
or U9553 (N_9553,N_714,N_2837);
or U9554 (N_9554,N_1234,N_443);
nand U9555 (N_9555,N_3608,N_2139);
or U9556 (N_9556,N_3034,N_2418);
xnor U9557 (N_9557,N_2968,N_4437);
and U9558 (N_9558,N_3793,N_2319);
and U9559 (N_9559,N_3,N_2292);
and U9560 (N_9560,N_3583,N_3279);
nor U9561 (N_9561,N_1671,N_2686);
xor U9562 (N_9562,N_81,N_2185);
xor U9563 (N_9563,N_1502,N_524);
nor U9564 (N_9564,N_3820,N_1867);
xor U9565 (N_9565,N_1666,N_1054);
xor U9566 (N_9566,N_2934,N_4487);
or U9567 (N_9567,N_362,N_1785);
nand U9568 (N_9568,N_4600,N_267);
nand U9569 (N_9569,N_60,N_178);
nand U9570 (N_9570,N_4756,N_1375);
xor U9571 (N_9571,N_3518,N_2435);
nor U9572 (N_9572,N_4532,N_700);
or U9573 (N_9573,N_1185,N_223);
and U9574 (N_9574,N_3041,N_990);
nand U9575 (N_9575,N_4318,N_2074);
xnor U9576 (N_9576,N_1888,N_898);
xnor U9577 (N_9577,N_4287,N_1075);
xnor U9578 (N_9578,N_909,N_1785);
nand U9579 (N_9579,N_3998,N_4976);
nand U9580 (N_9580,N_4976,N_2702);
nand U9581 (N_9581,N_511,N_2346);
nor U9582 (N_9582,N_409,N_4608);
or U9583 (N_9583,N_4229,N_804);
or U9584 (N_9584,N_3125,N_2788);
xor U9585 (N_9585,N_2087,N_3356);
nor U9586 (N_9586,N_1656,N_3802);
nand U9587 (N_9587,N_4029,N_4417);
nand U9588 (N_9588,N_3478,N_800);
nand U9589 (N_9589,N_4744,N_3905);
or U9590 (N_9590,N_2886,N_3450);
nand U9591 (N_9591,N_2702,N_3733);
and U9592 (N_9592,N_289,N_4247);
nor U9593 (N_9593,N_353,N_1442);
and U9594 (N_9594,N_4595,N_1464);
xnor U9595 (N_9595,N_1153,N_3150);
xor U9596 (N_9596,N_3827,N_751);
xor U9597 (N_9597,N_372,N_521);
and U9598 (N_9598,N_348,N_494);
nand U9599 (N_9599,N_3905,N_4834);
nand U9600 (N_9600,N_3945,N_103);
xnor U9601 (N_9601,N_2980,N_538);
nand U9602 (N_9602,N_3211,N_3056);
or U9603 (N_9603,N_1088,N_4536);
xor U9604 (N_9604,N_4352,N_547);
nor U9605 (N_9605,N_4123,N_2291);
xor U9606 (N_9606,N_3223,N_566);
and U9607 (N_9607,N_3877,N_3747);
xor U9608 (N_9608,N_4646,N_1487);
nand U9609 (N_9609,N_1170,N_2530);
xnor U9610 (N_9610,N_4746,N_3708);
and U9611 (N_9611,N_3636,N_2542);
or U9612 (N_9612,N_2613,N_4241);
and U9613 (N_9613,N_776,N_1376);
and U9614 (N_9614,N_281,N_3788);
nor U9615 (N_9615,N_2642,N_2527);
nor U9616 (N_9616,N_731,N_2849);
nand U9617 (N_9617,N_1668,N_4904);
nand U9618 (N_9618,N_534,N_2429);
nand U9619 (N_9619,N_2548,N_1371);
xnor U9620 (N_9620,N_1588,N_2049);
and U9621 (N_9621,N_28,N_2598);
xor U9622 (N_9622,N_3989,N_576);
xnor U9623 (N_9623,N_2624,N_2405);
nand U9624 (N_9624,N_3278,N_783);
and U9625 (N_9625,N_1105,N_3418);
xnor U9626 (N_9626,N_1101,N_1488);
and U9627 (N_9627,N_4977,N_640);
xor U9628 (N_9628,N_4965,N_4482);
or U9629 (N_9629,N_3390,N_3009);
or U9630 (N_9630,N_3379,N_1462);
nor U9631 (N_9631,N_2623,N_2168);
nor U9632 (N_9632,N_2023,N_1879);
nor U9633 (N_9633,N_3650,N_4983);
and U9634 (N_9634,N_1466,N_1966);
nand U9635 (N_9635,N_2127,N_682);
and U9636 (N_9636,N_2409,N_1142);
nor U9637 (N_9637,N_3394,N_1290);
and U9638 (N_9638,N_1210,N_4662);
nand U9639 (N_9639,N_4491,N_3963);
nor U9640 (N_9640,N_3906,N_4980);
nor U9641 (N_9641,N_4640,N_4129);
and U9642 (N_9642,N_40,N_1040);
or U9643 (N_9643,N_4963,N_2070);
nand U9644 (N_9644,N_1120,N_3620);
nand U9645 (N_9645,N_4812,N_203);
or U9646 (N_9646,N_1673,N_851);
xnor U9647 (N_9647,N_2719,N_207);
or U9648 (N_9648,N_2400,N_4208);
xnor U9649 (N_9649,N_2233,N_4061);
nand U9650 (N_9650,N_1451,N_217);
and U9651 (N_9651,N_3108,N_4017);
and U9652 (N_9652,N_4407,N_280);
and U9653 (N_9653,N_1426,N_4618);
nor U9654 (N_9654,N_4897,N_2777);
nand U9655 (N_9655,N_1691,N_615);
nand U9656 (N_9656,N_1602,N_23);
nand U9657 (N_9657,N_1474,N_3207);
xor U9658 (N_9658,N_2028,N_1997);
or U9659 (N_9659,N_2546,N_4752);
xnor U9660 (N_9660,N_1500,N_3260);
or U9661 (N_9661,N_3801,N_3796);
nor U9662 (N_9662,N_4760,N_3569);
or U9663 (N_9663,N_1725,N_3689);
nand U9664 (N_9664,N_4319,N_2828);
and U9665 (N_9665,N_2663,N_4776);
xnor U9666 (N_9666,N_1654,N_877);
xor U9667 (N_9667,N_2266,N_598);
nor U9668 (N_9668,N_1906,N_2141);
xnor U9669 (N_9669,N_4387,N_4873);
xnor U9670 (N_9670,N_107,N_4963);
xnor U9671 (N_9671,N_3540,N_3282);
xnor U9672 (N_9672,N_4294,N_2361);
xnor U9673 (N_9673,N_4053,N_4337);
xnor U9674 (N_9674,N_4446,N_4943);
nand U9675 (N_9675,N_4665,N_4925);
xor U9676 (N_9676,N_3254,N_476);
xor U9677 (N_9677,N_3026,N_4512);
xor U9678 (N_9678,N_4709,N_4008);
nand U9679 (N_9679,N_4183,N_2355);
and U9680 (N_9680,N_4743,N_1550);
and U9681 (N_9681,N_3673,N_3492);
and U9682 (N_9682,N_3950,N_2854);
and U9683 (N_9683,N_735,N_1481);
nand U9684 (N_9684,N_2158,N_1827);
nand U9685 (N_9685,N_698,N_2784);
and U9686 (N_9686,N_1515,N_729);
nand U9687 (N_9687,N_4790,N_1121);
nor U9688 (N_9688,N_4035,N_3837);
and U9689 (N_9689,N_3487,N_630);
and U9690 (N_9690,N_2625,N_3501);
and U9691 (N_9691,N_2929,N_3822);
nor U9692 (N_9692,N_2776,N_4005);
and U9693 (N_9693,N_2733,N_1337);
xor U9694 (N_9694,N_3987,N_1783);
nand U9695 (N_9695,N_3857,N_2102);
or U9696 (N_9696,N_4893,N_3884);
or U9697 (N_9697,N_628,N_2426);
nand U9698 (N_9698,N_4620,N_2083);
xor U9699 (N_9699,N_3162,N_3830);
or U9700 (N_9700,N_2053,N_416);
or U9701 (N_9701,N_75,N_1257);
or U9702 (N_9702,N_4066,N_4020);
xnor U9703 (N_9703,N_1306,N_1841);
nand U9704 (N_9704,N_4919,N_585);
and U9705 (N_9705,N_3952,N_2538);
nand U9706 (N_9706,N_382,N_700);
or U9707 (N_9707,N_1505,N_770);
or U9708 (N_9708,N_4986,N_988);
nand U9709 (N_9709,N_4226,N_4640);
or U9710 (N_9710,N_1477,N_775);
xor U9711 (N_9711,N_2877,N_1809);
nand U9712 (N_9712,N_4539,N_332);
nand U9713 (N_9713,N_4881,N_2522);
nand U9714 (N_9714,N_3038,N_1000);
nor U9715 (N_9715,N_1159,N_3964);
nor U9716 (N_9716,N_3317,N_3931);
and U9717 (N_9717,N_3799,N_1574);
nor U9718 (N_9718,N_1339,N_4656);
xor U9719 (N_9719,N_666,N_4430);
or U9720 (N_9720,N_4004,N_416);
xnor U9721 (N_9721,N_2132,N_1658);
nand U9722 (N_9722,N_841,N_2176);
nor U9723 (N_9723,N_2550,N_1270);
nand U9724 (N_9724,N_689,N_1240);
xor U9725 (N_9725,N_4960,N_2687);
xor U9726 (N_9726,N_1658,N_2776);
nand U9727 (N_9727,N_708,N_3635);
xnor U9728 (N_9728,N_3497,N_2764);
nand U9729 (N_9729,N_4498,N_1582);
nand U9730 (N_9730,N_4664,N_4682);
nor U9731 (N_9731,N_1771,N_4917);
nor U9732 (N_9732,N_3393,N_1871);
nand U9733 (N_9733,N_1921,N_3235);
xor U9734 (N_9734,N_4067,N_4336);
nand U9735 (N_9735,N_4176,N_4600);
xnor U9736 (N_9736,N_4748,N_4694);
xnor U9737 (N_9737,N_4188,N_2569);
and U9738 (N_9738,N_4370,N_4849);
or U9739 (N_9739,N_618,N_1708);
and U9740 (N_9740,N_144,N_2423);
or U9741 (N_9741,N_1635,N_2503);
and U9742 (N_9742,N_811,N_631);
xnor U9743 (N_9743,N_4319,N_2326);
xnor U9744 (N_9744,N_519,N_3075);
nand U9745 (N_9745,N_4345,N_2956);
nand U9746 (N_9746,N_3027,N_4332);
xor U9747 (N_9747,N_4022,N_2846);
and U9748 (N_9748,N_1043,N_4966);
xor U9749 (N_9749,N_4616,N_3077);
nor U9750 (N_9750,N_4992,N_2103);
or U9751 (N_9751,N_4358,N_3755);
xnor U9752 (N_9752,N_3185,N_4721);
and U9753 (N_9753,N_4247,N_2719);
xor U9754 (N_9754,N_2036,N_909);
and U9755 (N_9755,N_916,N_3211);
and U9756 (N_9756,N_96,N_3619);
and U9757 (N_9757,N_4619,N_2450);
and U9758 (N_9758,N_4411,N_274);
nand U9759 (N_9759,N_3069,N_2900);
nor U9760 (N_9760,N_483,N_2015);
xnor U9761 (N_9761,N_4942,N_2203);
and U9762 (N_9762,N_597,N_3562);
nor U9763 (N_9763,N_3000,N_2718);
or U9764 (N_9764,N_4630,N_477);
and U9765 (N_9765,N_2805,N_4001);
nand U9766 (N_9766,N_3833,N_1579);
and U9767 (N_9767,N_4069,N_3968);
and U9768 (N_9768,N_1757,N_1806);
nand U9769 (N_9769,N_1201,N_225);
or U9770 (N_9770,N_2023,N_1441);
xnor U9771 (N_9771,N_2982,N_970);
nand U9772 (N_9772,N_3024,N_2095);
nor U9773 (N_9773,N_2049,N_1260);
or U9774 (N_9774,N_4339,N_832);
nor U9775 (N_9775,N_3297,N_4852);
or U9776 (N_9776,N_484,N_392);
and U9777 (N_9777,N_1757,N_3424);
and U9778 (N_9778,N_555,N_2024);
nand U9779 (N_9779,N_1669,N_2656);
nand U9780 (N_9780,N_1626,N_4895);
xnor U9781 (N_9781,N_513,N_3302);
nand U9782 (N_9782,N_4409,N_4256);
or U9783 (N_9783,N_2629,N_3201);
or U9784 (N_9784,N_1132,N_167);
nand U9785 (N_9785,N_974,N_1110);
or U9786 (N_9786,N_2247,N_4396);
xnor U9787 (N_9787,N_980,N_4953);
and U9788 (N_9788,N_1098,N_2720);
xnor U9789 (N_9789,N_4605,N_3461);
nand U9790 (N_9790,N_3194,N_1529);
nor U9791 (N_9791,N_4112,N_1998);
or U9792 (N_9792,N_1331,N_4996);
or U9793 (N_9793,N_1067,N_2728);
or U9794 (N_9794,N_1842,N_3073);
and U9795 (N_9795,N_292,N_816);
nor U9796 (N_9796,N_1601,N_978);
xor U9797 (N_9797,N_2189,N_732);
or U9798 (N_9798,N_2470,N_2625);
nand U9799 (N_9799,N_4568,N_1315);
xor U9800 (N_9800,N_1664,N_2972);
nor U9801 (N_9801,N_4874,N_2386);
nor U9802 (N_9802,N_4414,N_1210);
nor U9803 (N_9803,N_890,N_2661);
nor U9804 (N_9804,N_2312,N_1802);
and U9805 (N_9805,N_4390,N_1304);
nand U9806 (N_9806,N_3066,N_963);
or U9807 (N_9807,N_192,N_573);
xor U9808 (N_9808,N_23,N_4444);
nor U9809 (N_9809,N_1957,N_2236);
nand U9810 (N_9810,N_3018,N_4280);
nand U9811 (N_9811,N_1161,N_3191);
xnor U9812 (N_9812,N_2540,N_3999);
or U9813 (N_9813,N_3481,N_4494);
nand U9814 (N_9814,N_283,N_736);
nor U9815 (N_9815,N_3635,N_3617);
xnor U9816 (N_9816,N_1425,N_3237);
and U9817 (N_9817,N_3651,N_3589);
or U9818 (N_9818,N_4361,N_487);
xnor U9819 (N_9819,N_2931,N_505);
or U9820 (N_9820,N_4968,N_230);
or U9821 (N_9821,N_1226,N_1255);
and U9822 (N_9822,N_3952,N_1053);
xnor U9823 (N_9823,N_3564,N_2392);
nor U9824 (N_9824,N_1644,N_966);
and U9825 (N_9825,N_3497,N_826);
xor U9826 (N_9826,N_445,N_4737);
xnor U9827 (N_9827,N_1908,N_544);
nand U9828 (N_9828,N_3596,N_4641);
nor U9829 (N_9829,N_2890,N_4774);
xor U9830 (N_9830,N_3058,N_1787);
or U9831 (N_9831,N_4599,N_4846);
xnor U9832 (N_9832,N_2307,N_359);
xor U9833 (N_9833,N_4800,N_3186);
nor U9834 (N_9834,N_3856,N_3170);
or U9835 (N_9835,N_2327,N_4014);
and U9836 (N_9836,N_2858,N_1924);
nor U9837 (N_9837,N_1155,N_4063);
and U9838 (N_9838,N_4591,N_3226);
and U9839 (N_9839,N_76,N_388);
xor U9840 (N_9840,N_1318,N_791);
xnor U9841 (N_9841,N_3728,N_4047);
and U9842 (N_9842,N_2133,N_2609);
nand U9843 (N_9843,N_1113,N_759);
or U9844 (N_9844,N_4001,N_4454);
nand U9845 (N_9845,N_4583,N_1559);
or U9846 (N_9846,N_2365,N_4018);
and U9847 (N_9847,N_2402,N_2700);
xor U9848 (N_9848,N_1517,N_3116);
xnor U9849 (N_9849,N_4458,N_2833);
or U9850 (N_9850,N_3541,N_4418);
nor U9851 (N_9851,N_4691,N_4238);
or U9852 (N_9852,N_2908,N_4645);
nand U9853 (N_9853,N_3108,N_1984);
and U9854 (N_9854,N_4870,N_4949);
and U9855 (N_9855,N_2361,N_2176);
or U9856 (N_9856,N_3047,N_4478);
xor U9857 (N_9857,N_694,N_3509);
or U9858 (N_9858,N_3143,N_4498);
nand U9859 (N_9859,N_3746,N_973);
nor U9860 (N_9860,N_1432,N_2543);
and U9861 (N_9861,N_794,N_177);
xor U9862 (N_9862,N_78,N_4999);
nor U9863 (N_9863,N_4785,N_2759);
or U9864 (N_9864,N_2044,N_4950);
and U9865 (N_9865,N_1699,N_2253);
or U9866 (N_9866,N_299,N_1375);
or U9867 (N_9867,N_743,N_1111);
or U9868 (N_9868,N_2028,N_1014);
and U9869 (N_9869,N_1076,N_4234);
and U9870 (N_9870,N_213,N_1588);
or U9871 (N_9871,N_2417,N_4659);
nand U9872 (N_9872,N_1805,N_1567);
xnor U9873 (N_9873,N_4830,N_4639);
xor U9874 (N_9874,N_1609,N_1473);
xor U9875 (N_9875,N_1590,N_1107);
and U9876 (N_9876,N_4383,N_829);
nand U9877 (N_9877,N_841,N_4364);
nor U9878 (N_9878,N_1172,N_158);
xor U9879 (N_9879,N_3784,N_877);
nor U9880 (N_9880,N_3145,N_499);
nor U9881 (N_9881,N_2042,N_501);
xor U9882 (N_9882,N_1634,N_4247);
nor U9883 (N_9883,N_919,N_3279);
xor U9884 (N_9884,N_1953,N_3708);
xor U9885 (N_9885,N_1818,N_913);
xnor U9886 (N_9886,N_1936,N_1451);
nand U9887 (N_9887,N_1732,N_2443);
and U9888 (N_9888,N_3259,N_1993);
xnor U9889 (N_9889,N_4904,N_1114);
and U9890 (N_9890,N_3485,N_3535);
or U9891 (N_9891,N_3421,N_1194);
xnor U9892 (N_9892,N_2096,N_2039);
nand U9893 (N_9893,N_1490,N_1958);
xnor U9894 (N_9894,N_3722,N_4787);
or U9895 (N_9895,N_3136,N_658);
or U9896 (N_9896,N_4474,N_114);
xnor U9897 (N_9897,N_3660,N_954);
or U9898 (N_9898,N_1329,N_1568);
nand U9899 (N_9899,N_3209,N_809);
nand U9900 (N_9900,N_3438,N_75);
nor U9901 (N_9901,N_1641,N_2573);
nor U9902 (N_9902,N_2883,N_4590);
nand U9903 (N_9903,N_3954,N_4383);
nor U9904 (N_9904,N_4592,N_4982);
nor U9905 (N_9905,N_4879,N_4964);
and U9906 (N_9906,N_2310,N_821);
xnor U9907 (N_9907,N_2103,N_592);
or U9908 (N_9908,N_3784,N_1768);
and U9909 (N_9909,N_2001,N_3679);
or U9910 (N_9910,N_4075,N_114);
nand U9911 (N_9911,N_1606,N_646);
or U9912 (N_9912,N_1282,N_928);
xor U9913 (N_9913,N_12,N_720);
or U9914 (N_9914,N_290,N_891);
and U9915 (N_9915,N_2596,N_1210);
or U9916 (N_9916,N_1258,N_1998);
or U9917 (N_9917,N_1355,N_572);
xor U9918 (N_9918,N_889,N_3043);
nor U9919 (N_9919,N_3582,N_2695);
or U9920 (N_9920,N_2,N_1186);
xor U9921 (N_9921,N_4579,N_2095);
nand U9922 (N_9922,N_1026,N_4937);
xnor U9923 (N_9923,N_1251,N_3419);
and U9924 (N_9924,N_887,N_596);
nor U9925 (N_9925,N_4920,N_468);
or U9926 (N_9926,N_3470,N_611);
or U9927 (N_9927,N_4826,N_3239);
nor U9928 (N_9928,N_1560,N_4353);
or U9929 (N_9929,N_4229,N_2820);
xor U9930 (N_9930,N_4875,N_892);
nor U9931 (N_9931,N_3130,N_2869);
or U9932 (N_9932,N_3984,N_1886);
and U9933 (N_9933,N_2536,N_1296);
or U9934 (N_9934,N_786,N_3635);
and U9935 (N_9935,N_4425,N_3441);
or U9936 (N_9936,N_1690,N_4196);
nand U9937 (N_9937,N_4648,N_3747);
nor U9938 (N_9938,N_3840,N_3425);
xor U9939 (N_9939,N_3066,N_2574);
nand U9940 (N_9940,N_2848,N_169);
or U9941 (N_9941,N_4853,N_1522);
xor U9942 (N_9942,N_4211,N_844);
and U9943 (N_9943,N_3041,N_749);
nand U9944 (N_9944,N_1866,N_4191);
and U9945 (N_9945,N_2687,N_2820);
nor U9946 (N_9946,N_3952,N_993);
xor U9947 (N_9947,N_4506,N_4554);
nand U9948 (N_9948,N_3369,N_3918);
nand U9949 (N_9949,N_331,N_4622);
and U9950 (N_9950,N_4348,N_836);
nor U9951 (N_9951,N_686,N_2101);
or U9952 (N_9952,N_2065,N_2897);
xor U9953 (N_9953,N_3850,N_272);
nor U9954 (N_9954,N_2087,N_2224);
xnor U9955 (N_9955,N_4422,N_1812);
nor U9956 (N_9956,N_3816,N_3244);
xor U9957 (N_9957,N_3144,N_4491);
xor U9958 (N_9958,N_2895,N_2848);
xnor U9959 (N_9959,N_2100,N_1831);
nand U9960 (N_9960,N_4726,N_1999);
and U9961 (N_9961,N_4122,N_1980);
nand U9962 (N_9962,N_2605,N_602);
nand U9963 (N_9963,N_1451,N_70);
and U9964 (N_9964,N_4636,N_2823);
or U9965 (N_9965,N_2913,N_1535);
or U9966 (N_9966,N_3271,N_2301);
or U9967 (N_9967,N_3280,N_4724);
xnor U9968 (N_9968,N_770,N_1138);
nor U9969 (N_9969,N_18,N_62);
or U9970 (N_9970,N_4900,N_1580);
nand U9971 (N_9971,N_4717,N_748);
nand U9972 (N_9972,N_937,N_4516);
nand U9973 (N_9973,N_1564,N_2777);
xnor U9974 (N_9974,N_959,N_4428);
or U9975 (N_9975,N_978,N_2104);
and U9976 (N_9976,N_802,N_366);
nand U9977 (N_9977,N_3540,N_398);
xnor U9978 (N_9978,N_2830,N_3115);
nor U9979 (N_9979,N_1704,N_4393);
xnor U9980 (N_9980,N_4692,N_1474);
or U9981 (N_9981,N_655,N_3658);
xor U9982 (N_9982,N_1581,N_270);
nand U9983 (N_9983,N_158,N_1383);
nor U9984 (N_9984,N_3307,N_1276);
xnor U9985 (N_9985,N_3273,N_1768);
xnor U9986 (N_9986,N_2627,N_3628);
nand U9987 (N_9987,N_4797,N_3333);
and U9988 (N_9988,N_3613,N_1673);
xor U9989 (N_9989,N_760,N_3914);
nor U9990 (N_9990,N_4296,N_930);
xnor U9991 (N_9991,N_1719,N_2479);
or U9992 (N_9992,N_2052,N_3059);
xor U9993 (N_9993,N_677,N_3501);
xor U9994 (N_9994,N_702,N_2781);
xnor U9995 (N_9995,N_1910,N_3737);
or U9996 (N_9996,N_3755,N_1516);
nand U9997 (N_9997,N_4068,N_4642);
nand U9998 (N_9998,N_2213,N_4816);
xor U9999 (N_9999,N_3442,N_3867);
or U10000 (N_10000,N_6792,N_9206);
and U10001 (N_10001,N_9872,N_9921);
nand U10002 (N_10002,N_6421,N_8681);
xnor U10003 (N_10003,N_9256,N_8467);
and U10004 (N_10004,N_8171,N_7967);
nand U10005 (N_10005,N_5983,N_6270);
nand U10006 (N_10006,N_8134,N_6349);
nand U10007 (N_10007,N_6373,N_6916);
xor U10008 (N_10008,N_5741,N_7480);
or U10009 (N_10009,N_9927,N_5321);
and U10010 (N_10010,N_7655,N_6292);
or U10011 (N_10011,N_6629,N_5817);
nand U10012 (N_10012,N_8400,N_8052);
and U10013 (N_10013,N_6648,N_7428);
or U10014 (N_10014,N_6485,N_9634);
and U10015 (N_10015,N_5623,N_6508);
or U10016 (N_10016,N_7035,N_8252);
nand U10017 (N_10017,N_7081,N_7797);
nand U10018 (N_10018,N_6841,N_7041);
xor U10019 (N_10019,N_8254,N_9429);
or U10020 (N_10020,N_9825,N_6249);
xor U10021 (N_10021,N_6877,N_9625);
xnor U10022 (N_10022,N_5457,N_8465);
nor U10023 (N_10023,N_7146,N_8256);
or U10024 (N_10024,N_8345,N_5052);
nand U10025 (N_10025,N_7503,N_7373);
xor U10026 (N_10026,N_8539,N_8119);
or U10027 (N_10027,N_9434,N_9166);
or U10028 (N_10028,N_8383,N_5782);
nand U10029 (N_10029,N_9842,N_6973);
nor U10030 (N_10030,N_5501,N_6983);
xnor U10031 (N_10031,N_7025,N_5757);
and U10032 (N_10032,N_7910,N_6026);
xnor U10033 (N_10033,N_5354,N_5152);
or U10034 (N_10034,N_6119,N_5833);
nand U10035 (N_10035,N_7892,N_9865);
xnor U10036 (N_10036,N_6427,N_6492);
or U10037 (N_10037,N_9751,N_7579);
and U10038 (N_10038,N_7999,N_6780);
nand U10039 (N_10039,N_5430,N_8165);
or U10040 (N_10040,N_7852,N_7196);
nor U10041 (N_10041,N_9248,N_8379);
xor U10042 (N_10042,N_8904,N_5558);
and U10043 (N_10043,N_7119,N_5766);
nor U10044 (N_10044,N_6263,N_8663);
nand U10045 (N_10045,N_6674,N_8194);
and U10046 (N_10046,N_7569,N_6147);
or U10047 (N_10047,N_6075,N_6250);
nor U10048 (N_10048,N_8109,N_7430);
nand U10049 (N_10049,N_6472,N_7710);
or U10050 (N_10050,N_6616,N_6244);
xnor U10051 (N_10051,N_6891,N_8514);
xor U10052 (N_10052,N_5909,N_7681);
nand U10053 (N_10053,N_9241,N_5407);
nand U10054 (N_10054,N_6441,N_8577);
nand U10055 (N_10055,N_8455,N_5281);
xnor U10056 (N_10056,N_8750,N_9738);
nor U10057 (N_10057,N_5703,N_7664);
nand U10058 (N_10058,N_9397,N_5953);
and U10059 (N_10059,N_8812,N_9762);
nand U10060 (N_10060,N_5298,N_9257);
nand U10061 (N_10061,N_5557,N_8759);
nand U10062 (N_10062,N_9601,N_6676);
nand U10063 (N_10063,N_9294,N_8805);
or U10064 (N_10064,N_7175,N_6788);
nand U10065 (N_10065,N_8836,N_9792);
and U10066 (N_10066,N_8468,N_7193);
nor U10067 (N_10067,N_9887,N_5569);
nand U10068 (N_10068,N_6863,N_7406);
and U10069 (N_10069,N_8800,N_6582);
or U10070 (N_10070,N_8235,N_5022);
xnor U10071 (N_10071,N_9804,N_9377);
or U10072 (N_10072,N_9716,N_7236);
xor U10073 (N_10073,N_6672,N_7676);
and U10074 (N_10074,N_7606,N_7169);
nand U10075 (N_10075,N_7050,N_9300);
and U10076 (N_10076,N_5979,N_7089);
or U10077 (N_10077,N_7743,N_5872);
nor U10078 (N_10078,N_7624,N_6623);
nand U10079 (N_10079,N_8788,N_5305);
and U10080 (N_10080,N_5846,N_5273);
xnor U10081 (N_10081,N_6769,N_9516);
nor U10082 (N_10082,N_5366,N_7549);
nor U10083 (N_10083,N_6044,N_7673);
nand U10084 (N_10084,N_9866,N_8907);
xnor U10085 (N_10085,N_5311,N_6282);
nand U10086 (N_10086,N_9492,N_6241);
nor U10087 (N_10087,N_6897,N_6014);
or U10088 (N_10088,N_7899,N_8353);
nand U10089 (N_10089,N_8689,N_9345);
or U10090 (N_10090,N_5451,N_6318);
or U10091 (N_10091,N_5274,N_6275);
xor U10092 (N_10092,N_6573,N_8857);
or U10093 (N_10093,N_7591,N_7446);
xnor U10094 (N_10094,N_9899,N_8363);
xor U10095 (N_10095,N_6999,N_7161);
or U10096 (N_10096,N_7943,N_7507);
or U10097 (N_10097,N_5509,N_8080);
or U10098 (N_10098,N_8984,N_8493);
xor U10099 (N_10099,N_7329,N_5986);
nor U10100 (N_10100,N_8470,N_6193);
or U10101 (N_10101,N_7415,N_8967);
xor U10102 (N_10102,N_8160,N_7307);
nand U10103 (N_10103,N_8098,N_9066);
nor U10104 (N_10104,N_7590,N_5885);
or U10105 (N_10105,N_9994,N_8614);
and U10106 (N_10106,N_6050,N_7901);
or U10107 (N_10107,N_8613,N_8576);
nand U10108 (N_10108,N_9026,N_7885);
xor U10109 (N_10109,N_9616,N_8022);
nand U10110 (N_10110,N_5510,N_9262);
and U10111 (N_10111,N_9694,N_8694);
nor U10112 (N_10112,N_9822,N_7473);
and U10113 (N_10113,N_7074,N_8270);
and U10114 (N_10114,N_7038,N_8722);
nand U10115 (N_10115,N_8257,N_9309);
xor U10116 (N_10116,N_7408,N_5495);
and U10117 (N_10117,N_8763,N_6569);
xnor U10118 (N_10118,N_8996,N_6604);
xor U10119 (N_10119,N_7971,N_5016);
or U10120 (N_10120,N_7711,N_8617);
nor U10121 (N_10121,N_9853,N_5243);
xor U10122 (N_10122,N_6405,N_9708);
nand U10123 (N_10123,N_6021,N_7270);
or U10124 (N_10124,N_8999,N_5362);
and U10125 (N_10125,N_6418,N_5756);
nand U10126 (N_10126,N_6781,N_9096);
and U10127 (N_10127,N_9321,N_5376);
nor U10128 (N_10128,N_8975,N_5419);
nor U10129 (N_10129,N_5278,N_5206);
nand U10130 (N_10130,N_9043,N_6593);
and U10131 (N_10131,N_9232,N_7722);
or U10132 (N_10132,N_6203,N_8233);
xnor U10133 (N_10133,N_9020,N_5694);
xnor U10134 (N_10134,N_6984,N_8602);
xor U10135 (N_10135,N_6425,N_9289);
nand U10136 (N_10136,N_6536,N_7564);
nand U10137 (N_10137,N_9117,N_7115);
nand U10138 (N_10138,N_6366,N_6268);
or U10139 (N_10139,N_9846,N_8889);
nand U10140 (N_10140,N_8348,N_5739);
and U10141 (N_10141,N_7343,N_6439);
nor U10142 (N_10142,N_6804,N_5559);
or U10143 (N_10143,N_5011,N_6309);
and U10144 (N_10144,N_7738,N_6884);
nand U10145 (N_10145,N_5265,N_8987);
or U10146 (N_10146,N_8683,N_8097);
or U10147 (N_10147,N_9912,N_6710);
and U10148 (N_10148,N_6542,N_6936);
nor U10149 (N_10149,N_8971,N_7529);
or U10150 (N_10150,N_5004,N_8776);
or U10151 (N_10151,N_5093,N_6225);
xor U10152 (N_10152,N_7519,N_5748);
nand U10153 (N_10153,N_5353,N_9889);
or U10154 (N_10154,N_6528,N_6566);
or U10155 (N_10155,N_9324,N_8606);
or U10156 (N_10156,N_6533,N_9267);
and U10157 (N_10157,N_9868,N_6335);
xor U10158 (N_10158,N_5484,N_7036);
nor U10159 (N_10159,N_5654,N_5740);
nand U10160 (N_10160,N_6029,N_6783);
nor U10161 (N_10161,N_8169,N_6041);
or U10162 (N_10162,N_6188,N_8272);
xnor U10163 (N_10163,N_6819,N_7809);
xor U10164 (N_10164,N_7979,N_8205);
nand U10165 (N_10165,N_7874,N_7709);
nor U10166 (N_10166,N_8968,N_7166);
and U10167 (N_10167,N_6015,N_9226);
or U10168 (N_10168,N_7754,N_8553);
and U10169 (N_10169,N_6993,N_5742);
and U10170 (N_10170,N_9452,N_6455);
nor U10171 (N_10171,N_8226,N_8020);
nand U10172 (N_10172,N_5306,N_6267);
nand U10173 (N_10173,N_8179,N_6880);
or U10174 (N_10174,N_8089,N_9688);
nor U10175 (N_10175,N_9263,N_6946);
or U10176 (N_10176,N_5819,N_7099);
nand U10177 (N_10177,N_8802,N_8253);
nand U10178 (N_10178,N_6033,N_6661);
nand U10179 (N_10179,N_6698,N_9657);
nand U10180 (N_10180,N_5255,N_8624);
or U10181 (N_10181,N_9967,N_5075);
xor U10182 (N_10182,N_5294,N_9908);
nand U10183 (N_10183,N_9031,N_8669);
or U10184 (N_10184,N_8598,N_7812);
nand U10185 (N_10185,N_8564,N_5364);
xor U10186 (N_10186,N_9619,N_6729);
nand U10187 (N_10187,N_9075,N_7842);
or U10188 (N_10188,N_9834,N_9756);
nand U10189 (N_10189,N_9587,N_9763);
xor U10190 (N_10190,N_9340,N_8186);
and U10191 (N_10191,N_6401,N_8401);
and U10192 (N_10192,N_5677,N_9126);
xnor U10193 (N_10193,N_9288,N_7800);
or U10194 (N_10194,N_7188,N_5965);
nand U10195 (N_10195,N_7894,N_9080);
nand U10196 (N_10196,N_7692,N_9204);
xor U10197 (N_10197,N_6525,N_7474);
nor U10198 (N_10198,N_9201,N_9609);
xor U10199 (N_10199,N_5417,N_9656);
nor U10200 (N_10200,N_8610,N_9906);
xnor U10201 (N_10201,N_7652,N_9273);
nand U10202 (N_10202,N_8712,N_8691);
or U10203 (N_10203,N_7588,N_8976);
nand U10204 (N_10204,N_9455,N_9951);
and U10205 (N_10205,N_5606,N_6590);
nand U10206 (N_10206,N_9766,N_9060);
nand U10207 (N_10207,N_6693,N_7926);
nand U10208 (N_10208,N_9001,N_8828);
nand U10209 (N_10209,N_6010,N_6459);
xnor U10210 (N_10210,N_5539,N_9322);
or U10211 (N_10211,N_8740,N_7921);
nand U10212 (N_10212,N_6468,N_6925);
xnor U10213 (N_10213,N_9356,N_8833);
xor U10214 (N_10214,N_8023,N_8132);
or U10215 (N_10215,N_6555,N_9505);
xnor U10216 (N_10216,N_8359,N_5977);
and U10217 (N_10217,N_6078,N_6944);
nor U10218 (N_10218,N_5429,N_7765);
xnor U10219 (N_10219,N_9140,N_8068);
or U10220 (N_10220,N_8579,N_8879);
nor U10221 (N_10221,N_6645,N_5512);
nor U10222 (N_10222,N_5967,N_9513);
nand U10223 (N_10223,N_9675,N_6939);
xnor U10224 (N_10224,N_6449,N_5711);
nand U10225 (N_10225,N_9233,N_9493);
or U10226 (N_10226,N_5119,N_9975);
nor U10227 (N_10227,N_8101,N_7530);
nand U10228 (N_10228,N_5709,N_9683);
xor U10229 (N_10229,N_7327,N_7001);
or U10230 (N_10230,N_9895,N_5828);
nand U10231 (N_10231,N_8085,N_5780);
or U10232 (N_10232,N_6256,N_5589);
nand U10233 (N_10233,N_6248,N_7330);
nand U10234 (N_10234,N_7679,N_7631);
and U10235 (N_10235,N_7172,N_5603);
or U10236 (N_10236,N_5355,N_6887);
nand U10237 (N_10237,N_5823,N_5796);
or U10238 (N_10238,N_9213,N_5891);
nand U10239 (N_10239,N_9151,N_7278);
nand U10240 (N_10240,N_8912,N_5026);
or U10241 (N_10241,N_9401,N_8679);
nand U10242 (N_10242,N_5221,N_9574);
and U10243 (N_10243,N_9424,N_5018);
xnor U10244 (N_10244,N_6370,N_5050);
or U10245 (N_10245,N_7241,N_8141);
nand U10246 (N_10246,N_8005,N_5876);
or U10247 (N_10247,N_9642,N_8842);
and U10248 (N_10248,N_6357,N_9948);
nor U10249 (N_10249,N_7731,N_7142);
nand U10250 (N_10250,N_7831,N_5947);
nor U10251 (N_10251,N_6608,N_5277);
and U10252 (N_10252,N_9501,N_6251);
xnor U10253 (N_10253,N_6640,N_7888);
and U10254 (N_10254,N_8027,N_8185);
or U10255 (N_10255,N_5081,N_9245);
xor U10256 (N_10256,N_5544,N_9431);
nand U10257 (N_10257,N_7012,N_8018);
nand U10258 (N_10258,N_5655,N_6931);
and U10259 (N_10259,N_6673,N_6101);
nor U10260 (N_10260,N_7750,N_9076);
nor U10261 (N_10261,N_7532,N_7880);
and U10262 (N_10262,N_8178,N_8964);
nor U10263 (N_10263,N_7411,N_8238);
and U10264 (N_10264,N_7699,N_5793);
and U10265 (N_10265,N_5945,N_6156);
or U10266 (N_10266,N_5341,N_7575);
nor U10267 (N_10267,N_6721,N_7251);
nand U10268 (N_10268,N_6883,N_7363);
xor U10269 (N_10269,N_8757,N_9779);
nand U10270 (N_10270,N_6012,N_7200);
nand U10271 (N_10271,N_7127,N_6894);
nor U10272 (N_10272,N_6609,N_6926);
nor U10273 (N_10273,N_7006,N_6641);
xnor U10274 (N_10274,N_8674,N_8596);
nor U10275 (N_10275,N_5181,N_7249);
nand U10276 (N_10276,N_8590,N_9029);
xnor U10277 (N_10277,N_7381,N_6386);
xor U10278 (N_10278,N_7953,N_5297);
and U10279 (N_10279,N_5525,N_7392);
nand U10280 (N_10280,N_7977,N_5747);
nor U10281 (N_10281,N_6283,N_8523);
nand U10282 (N_10282,N_7825,N_8482);
or U10283 (N_10283,N_9510,N_6212);
nor U10284 (N_10284,N_5056,N_9099);
and U10285 (N_10285,N_8931,N_7433);
nor U10286 (N_10286,N_7997,N_5227);
nor U10287 (N_10287,N_9805,N_6583);
and U10288 (N_10288,N_9438,N_9674);
xnor U10289 (N_10289,N_5726,N_7833);
nand U10290 (N_10290,N_7956,N_8130);
nor U10291 (N_10291,N_6109,N_6820);
nor U10292 (N_10292,N_6712,N_5785);
and U10293 (N_10293,N_5573,N_7133);
or U10294 (N_10294,N_8137,N_8959);
nand U10295 (N_10295,N_7317,N_8569);
xor U10296 (N_10296,N_5130,N_6214);
and U10297 (N_10297,N_6007,N_5122);
and U10298 (N_10298,N_6351,N_7752);
nor U10299 (N_10299,N_7222,N_5129);
and U10300 (N_10300,N_6818,N_6023);
and U10301 (N_10301,N_6746,N_7031);
nand U10302 (N_10302,N_8618,N_8871);
and U10303 (N_10303,N_9087,N_6980);
xor U10304 (N_10304,N_8526,N_7778);
and U10305 (N_10305,N_9149,N_5566);
or U10306 (N_10306,N_9422,N_5849);
xnor U10307 (N_10307,N_8983,N_5204);
or U10308 (N_10308,N_5914,N_5394);
and U10309 (N_10309,N_7887,N_7088);
nor U10310 (N_10310,N_8373,N_8507);
xor U10311 (N_10311,N_8449,N_9067);
and U10312 (N_10312,N_8572,N_7286);
nand U10313 (N_10313,N_8738,N_7048);
and U10314 (N_10314,N_8813,N_8657);
nor U10315 (N_10315,N_7262,N_9451);
or U10316 (N_10316,N_6682,N_7379);
and U10317 (N_10317,N_5966,N_5155);
xor U10318 (N_10318,N_6378,N_9668);
xnor U10319 (N_10319,N_8649,N_7816);
nor U10320 (N_10320,N_6865,N_8295);
or U10321 (N_10321,N_7737,N_8121);
nor U10322 (N_10322,N_7653,N_6517);
nor U10323 (N_10323,N_7534,N_8397);
nor U10324 (N_10324,N_6165,N_6065);
xor U10325 (N_10325,N_6098,N_8860);
xor U10326 (N_10326,N_7266,N_9700);
nor U10327 (N_10327,N_6070,N_6141);
xnor U10328 (N_10328,N_8670,N_8037);
nand U10329 (N_10329,N_6148,N_6557);
xor U10330 (N_10330,N_8905,N_5031);
nand U10331 (N_10331,N_8412,N_5337);
xor U10332 (N_10332,N_7980,N_6679);
nor U10333 (N_10333,N_8673,N_8753);
or U10334 (N_10334,N_9650,N_7570);
nand U10335 (N_10335,N_7360,N_8744);
xnor U10336 (N_10336,N_5957,N_8297);
xnor U10337 (N_10337,N_8170,N_9896);
or U10338 (N_10338,N_8547,N_5459);
nor U10339 (N_10339,N_7390,N_8399);
and U10340 (N_10340,N_7380,N_5436);
nor U10341 (N_10341,N_8214,N_8269);
or U10342 (N_10342,N_5871,N_6361);
nand U10343 (N_10343,N_8422,N_7422);
nand U10344 (N_10344,N_6368,N_5729);
and U10345 (N_10345,N_5970,N_7045);
and U10346 (N_10346,N_5345,N_5550);
nand U10347 (N_10347,N_9542,N_6649);
xor U10348 (N_10348,N_5285,N_9890);
and U10349 (N_10349,N_7767,N_9531);
xnor U10350 (N_10350,N_8311,N_6008);
xnor U10351 (N_10351,N_7219,N_5955);
xnor U10352 (N_10352,N_7501,N_8275);
xor U10353 (N_10353,N_7730,N_8219);
or U10354 (N_10354,N_5621,N_5843);
and U10355 (N_10355,N_5188,N_6892);
xor U10356 (N_10356,N_8044,N_5611);
xnor U10357 (N_10357,N_9945,N_5236);
and U10358 (N_10358,N_6257,N_7720);
and U10359 (N_10359,N_6400,N_7341);
xor U10360 (N_10360,N_6900,N_6090);
and U10361 (N_10361,N_5618,N_8946);
xor U10362 (N_10362,N_7460,N_7596);
xor U10363 (N_10363,N_6358,N_7867);
nand U10364 (N_10364,N_9770,N_7167);
or U10365 (N_10365,N_8011,N_9507);
xnor U10366 (N_10366,N_6417,N_7156);
nand U10367 (N_10367,N_6363,N_7086);
nor U10368 (N_10368,N_5094,N_6458);
nand U10369 (N_10369,N_9722,N_6597);
and U10370 (N_10370,N_6110,N_9595);
nand U10371 (N_10371,N_8172,N_8259);
nor U10372 (N_10372,N_6724,N_6374);
and U10373 (N_10373,N_8700,N_8123);
or U10374 (N_10374,N_5176,N_9044);
xor U10375 (N_10375,N_9807,N_9318);
or U10376 (N_10376,N_9009,N_9843);
nand U10377 (N_10377,N_6667,N_9049);
nand U10378 (N_10378,N_8661,N_9836);
nand U10379 (N_10379,N_6186,N_9800);
xor U10380 (N_10380,N_5749,N_9054);
xor U10381 (N_10381,N_8333,N_9871);
nor U10382 (N_10382,N_8352,N_9386);
or U10383 (N_10383,N_5024,N_5395);
or U10384 (N_10384,N_5490,N_7578);
xor U10385 (N_10385,N_9030,N_9023);
xor U10386 (N_10386,N_7204,N_5912);
or U10387 (N_10387,N_7000,N_6732);
nor U10388 (N_10388,N_6848,N_9174);
xnor U10389 (N_10389,N_7108,N_6680);
nand U10390 (N_10390,N_6172,N_5824);
xnor U10391 (N_10391,N_8660,N_8183);
and U10392 (N_10392,N_9279,N_9025);
xnor U10393 (N_10393,N_8903,N_9956);
or U10394 (N_10394,N_6354,N_5505);
nand U10395 (N_10395,N_5172,N_6086);
and U10396 (N_10396,N_6396,N_8492);
nor U10397 (N_10397,N_5144,N_9113);
and U10398 (N_10398,N_5528,N_5857);
or U10399 (N_10399,N_9995,N_6838);
nor U10400 (N_10400,N_8858,N_7497);
or U10401 (N_10401,N_9922,N_5032);
xnor U10402 (N_10402,N_9439,N_8427);
and U10403 (N_10403,N_5140,N_5521);
nor U10404 (N_10404,N_7764,N_5882);
nand U10405 (N_10405,N_7684,N_8111);
nand U10406 (N_10406,N_9714,N_7668);
nor U10407 (N_10407,N_6379,N_9019);
nand U10408 (N_10408,N_8719,N_9709);
nor U10409 (N_10409,N_9400,N_5097);
and U10410 (N_10410,N_9447,N_5699);
xor U10411 (N_10411,N_7677,N_8586);
nand U10412 (N_10412,N_7511,N_7678);
nand U10413 (N_10413,N_7871,N_5995);
nand U10414 (N_10414,N_8303,N_8034);
nor U10415 (N_10415,N_7966,N_7808);
and U10416 (N_10416,N_7060,N_5474);
nand U10417 (N_10417,N_5806,N_8300);
or U10418 (N_10418,N_9687,N_5530);
nand U10419 (N_10419,N_7316,N_5279);
and U10420 (N_10420,N_7491,N_9543);
xnor U10421 (N_10421,N_8442,N_9523);
nor U10422 (N_10422,N_6384,N_5064);
nand U10423 (N_10423,N_9525,N_9357);
nand U10424 (N_10424,N_9209,N_6191);
or U10425 (N_10425,N_5452,N_8450);
or U10426 (N_10426,N_9022,N_6253);
or U10427 (N_10427,N_5496,N_7245);
and U10428 (N_10428,N_8599,N_5881);
and U10429 (N_10429,N_6678,N_7919);
and U10430 (N_10430,N_7359,N_6947);
or U10431 (N_10431,N_5534,N_8914);
xor U10432 (N_10432,N_6652,N_6963);
nand U10433 (N_10433,N_8619,N_6096);
and U10434 (N_10434,N_6153,N_6025);
nand U10435 (N_10435,N_9533,N_6580);
xnor U10436 (N_10436,N_6493,N_6540);
and U10437 (N_10437,N_8633,N_5039);
xnor U10438 (N_10438,N_9235,N_8073);
and U10439 (N_10439,N_7914,N_8524);
nor U10440 (N_10440,N_9468,N_8196);
and U10441 (N_10441,N_9027,N_9100);
nor U10442 (N_10442,N_7047,N_9246);
nor U10443 (N_10443,N_5943,N_5842);
xor U10444 (N_10444,N_9137,N_6761);
or U10445 (N_10445,N_7429,N_5162);
nand U10446 (N_10446,N_7822,N_5923);
or U10447 (N_10447,N_9568,N_7478);
nand U10448 (N_10448,N_8429,N_5272);
nor U10449 (N_10449,N_8851,N_9572);
or U10450 (N_10450,N_7296,N_7536);
and U10451 (N_10451,N_6945,N_8500);
and U10452 (N_10452,N_7464,N_8671);
xor U10453 (N_10453,N_8372,N_6893);
and U10454 (N_10454,N_5269,N_9767);
or U10455 (N_10455,N_5367,N_9600);
and U10456 (N_10456,N_9179,N_7597);
and U10457 (N_10457,N_8543,N_5900);
and U10458 (N_10458,N_7069,N_5313);
nor U10459 (N_10459,N_9071,N_9878);
xor U10460 (N_10460,N_8486,N_6511);
or U10461 (N_10461,N_6992,N_6395);
nor U10462 (N_10462,N_6719,N_7093);
xor U10463 (N_10463,N_6986,N_8846);
or U10464 (N_10464,N_9184,N_6072);
xor U10465 (N_10465,N_8197,N_6815);
or U10466 (N_10466,N_7659,N_9791);
or U10467 (N_10467,N_7016,N_7993);
nor U10468 (N_10468,N_6477,N_5982);
xnor U10469 (N_10469,N_8201,N_5439);
and U10470 (N_10470,N_7671,N_9503);
or U10471 (N_10471,N_9215,N_8881);
or U10472 (N_10472,N_9712,N_6650);
and U10473 (N_10473,N_9303,N_5184);
and U10474 (N_10474,N_6494,N_6469);
nand U10475 (N_10475,N_9223,N_6830);
and U10476 (N_10476,N_5720,N_8809);
nor U10477 (N_10477,N_6930,N_8331);
and U10478 (N_10478,N_5687,N_5751);
nor U10479 (N_10479,N_5722,N_9885);
and U10480 (N_10480,N_9391,N_8032);
nor U10481 (N_10481,N_7883,N_9632);
nor U10482 (N_10482,N_7636,N_5454);
nor U10483 (N_10483,N_8510,N_5858);
and U10484 (N_10484,N_8338,N_9854);
xor U10485 (N_10485,N_5217,N_9320);
nor U10486 (N_10486,N_6084,N_9942);
or U10487 (N_10487,N_9584,N_6482);
nand U10488 (N_10488,N_5259,N_6562);
or U10489 (N_10489,N_9740,N_6226);
or U10490 (N_10490,N_6474,N_5638);
and U10491 (N_10491,N_6372,N_6857);
xor U10492 (N_10492,N_6496,N_9146);
nand U10493 (N_10493,N_6530,N_8454);
xor U10494 (N_10494,N_8279,N_6596);
or U10495 (N_10495,N_6638,N_8768);
and U10496 (N_10496,N_9664,N_9477);
nand U10497 (N_10497,N_8292,N_9932);
and U10498 (N_10498,N_7402,N_8534);
xnor U10499 (N_10499,N_7994,N_7203);
nand U10500 (N_10500,N_6778,N_6032);
nor U10501 (N_10501,N_6798,N_7616);
nand U10502 (N_10502,N_8994,N_5820);
and U10503 (N_10503,N_5875,N_8783);
or U10504 (N_10504,N_9944,N_6013);
and U10505 (N_10505,N_7320,N_5365);
xnor U10506 (N_10506,N_7477,N_9486);
xnor U10507 (N_10507,N_9521,N_8578);
xor U10508 (N_10508,N_8806,N_8724);
or U10509 (N_10509,N_8824,N_8451);
xnor U10510 (N_10510,N_7639,N_8898);
xnor U10511 (N_10511,N_6951,N_5601);
and U10512 (N_10512,N_7313,N_8726);
or U10513 (N_10513,N_8035,N_9560);
and U10514 (N_10514,N_5946,N_6619);
nor U10515 (N_10515,N_7122,N_6406);
xor U10516 (N_10516,N_7173,N_9719);
nor U10517 (N_10517,N_8225,N_9189);
or U10518 (N_10518,N_6625,N_7044);
xnor U10519 (N_10519,N_5320,N_5017);
nor U10520 (N_10520,N_8497,N_7527);
xnor U10521 (N_10521,N_8736,N_6207);
xnor U10522 (N_10522,N_6959,N_7384);
and U10523 (N_10523,N_7632,N_7070);
xnor U10524 (N_10524,N_6409,N_6755);
nand U10525 (N_10525,N_7144,N_5033);
nor U10526 (N_10526,N_7331,N_7103);
nand U10527 (N_10527,N_7500,N_7846);
or U10528 (N_10528,N_5164,N_8487);
nand U10529 (N_10529,N_7062,N_9382);
nor U10530 (N_10530,N_8952,N_9435);
nor U10531 (N_10531,N_7817,N_6129);
nand U10532 (N_10532,N_8820,N_7011);
xor U10533 (N_10533,N_8202,N_9573);
nor U10534 (N_10534,N_8142,N_9925);
nand U10535 (N_10535,N_7234,N_9396);
or U10536 (N_10536,N_8106,N_7785);
or U10537 (N_10537,N_5698,N_7004);
xor U10538 (N_10538,N_8108,N_8264);
nor U10539 (N_10539,N_8153,N_9898);
xor U10540 (N_10540,N_5497,N_9405);
nor U10541 (N_10541,N_8296,N_7281);
or U10542 (N_10542,N_8735,N_7955);
or U10543 (N_10543,N_8139,N_8853);
or U10544 (N_10544,N_9884,N_7189);
nand U10545 (N_10545,N_5230,N_6303);
or U10546 (N_10546,N_9544,N_6310);
nor U10547 (N_10547,N_9250,N_5079);
and U10548 (N_10548,N_8629,N_6711);
nor U10549 (N_10549,N_6383,N_5494);
nand U10550 (N_10550,N_8852,N_7180);
xnor U10551 (N_10551,N_7283,N_9661);
nand U10552 (N_10552,N_5218,N_5812);
nand U10553 (N_10553,N_8926,N_9597);
nand U10554 (N_10554,N_9776,N_8955);
and U10555 (N_10555,N_6103,N_5627);
and U10556 (N_10556,N_9375,N_7264);
xor U10557 (N_10557,N_7982,N_7213);
and U10558 (N_10558,N_8878,N_9721);
nand U10559 (N_10559,N_7061,N_6338);
or U10560 (N_10560,N_8200,N_6803);
nand U10561 (N_10561,N_5469,N_9727);
nand U10562 (N_10562,N_9880,N_5964);
nand U10563 (N_10563,N_8894,N_8181);
and U10564 (N_10564,N_6797,N_8839);
and U10565 (N_10565,N_6890,N_8391);
and U10566 (N_10566,N_7969,N_9109);
and U10567 (N_10567,N_6954,N_8848);
and U10568 (N_10568,N_9745,N_8739);
and U10569 (N_10569,N_8872,N_6076);
nand U10570 (N_10570,N_5317,N_5169);
nor U10571 (N_10571,N_5483,N_6905);
nand U10572 (N_10572,N_5821,N_6331);
nor U10573 (N_10573,N_7055,N_6208);
nor U10574 (N_10574,N_5418,N_7423);
nor U10575 (N_10575,N_5049,N_9710);
xor U10576 (N_10576,N_8001,N_7453);
or U10577 (N_10577,N_9660,N_6066);
xor U10578 (N_10578,N_9496,N_7742);
or U10579 (N_10579,N_7257,N_6908);
xor U10580 (N_10580,N_5554,N_8815);
or U10581 (N_10581,N_6653,N_8046);
nand U10582 (N_10582,N_9796,N_8755);
xor U10583 (N_10583,N_7290,N_5128);
nand U10584 (N_10584,N_8120,N_6773);
or U10585 (N_10585,N_8773,N_5800);
or U10586 (N_10586,N_7927,N_9015);
or U10587 (N_10587,N_6671,N_6553);
or U10588 (N_10588,N_9655,N_9789);
and U10589 (N_10589,N_6223,N_9374);
xnor U10590 (N_10590,N_6683,N_8685);
or U10591 (N_10591,N_7116,N_6463);
or U10592 (N_10592,N_8410,N_9870);
nand U10593 (N_10593,N_7159,N_6972);
and U10594 (N_10594,N_7246,N_8807);
nor U10595 (N_10595,N_6432,N_7903);
nand U10596 (N_10596,N_7838,N_6105);
xor U10597 (N_10597,N_8855,N_8516);
or U10598 (N_10598,N_7418,N_9268);
nor U10599 (N_10599,N_9089,N_6476);
and U10600 (N_10600,N_9202,N_9440);
nor U10601 (N_10601,N_9784,N_8559);
nor U10602 (N_10602,N_8702,N_8446);
xor U10603 (N_10603,N_6160,N_7090);
nand U10604 (N_10604,N_6575,N_6860);
nor U10605 (N_10605,N_7521,N_5335);
and U10606 (N_10606,N_5944,N_6842);
nor U10607 (N_10607,N_8387,N_9436);
and U10608 (N_10608,N_6464,N_8389);
and U10609 (N_10609,N_8533,N_6631);
or U10610 (N_10610,N_5391,N_8826);
or U10611 (N_10611,N_5254,N_6564);
and U10612 (N_10612,N_6751,N_7149);
nand U10613 (N_10613,N_9933,N_9812);
and U10614 (N_10614,N_8949,N_6272);
or U10615 (N_10615,N_5545,N_6437);
nor U10616 (N_10616,N_5814,N_9658);
xnor U10617 (N_10617,N_8728,N_8033);
nand U10618 (N_10618,N_6549,N_7207);
xnor U10619 (N_10619,N_5574,N_5148);
nand U10620 (N_10620,N_8703,N_8887);
or U10621 (N_10621,N_5005,N_9630);
and U10622 (N_10622,N_5115,N_9644);
nand U10623 (N_10623,N_9869,N_7868);
nand U10624 (N_10624,N_8519,N_7902);
nor U10625 (N_10625,N_5063,N_9393);
nor U10626 (N_10626,N_8140,N_7010);
or U10627 (N_10627,N_6359,N_7125);
and U10628 (N_10628,N_6487,N_7904);
nor U10629 (N_10629,N_5223,N_6876);
and U10630 (N_10630,N_7915,N_7552);
nand U10631 (N_10631,N_5382,N_5658);
xor U10632 (N_10632,N_7802,N_6998);
nand U10633 (N_10633,N_5704,N_7123);
nor U10634 (N_10634,N_8609,N_5706);
nor U10635 (N_10635,N_9244,N_6019);
and U10636 (N_10636,N_5473,N_5383);
and U10637 (N_10637,N_6265,N_5175);
nor U10638 (N_10638,N_5767,N_6541);
nor U10639 (N_10639,N_8969,N_8438);
xnor U10640 (N_10640,N_8896,N_9408);
nand U10641 (N_10641,N_7261,N_8893);
or U10642 (N_10642,N_7908,N_5462);
xor U10643 (N_10643,N_9628,N_8597);
or U10644 (N_10644,N_6937,N_5695);
nor U10645 (N_10645,N_9349,N_5734);
xor U10646 (N_10646,N_6277,N_6182);
or U10647 (N_10647,N_5962,N_8616);
nand U10648 (N_10648,N_9051,N_6091);
nand U10649 (N_10649,N_7988,N_9774);
and U10650 (N_10650,N_6911,N_8845);
xor U10651 (N_10651,N_6849,N_9808);
and U10652 (N_10652,N_7944,N_5609);
and U10653 (N_10653,N_6981,N_5935);
nand U10654 (N_10654,N_9614,N_7912);
and U10655 (N_10655,N_7928,N_6434);
and U10656 (N_10656,N_5551,N_9504);
xor U10657 (N_10657,N_6605,N_6006);
or U10658 (N_10658,N_6247,N_5797);
nand U10659 (N_10659,N_6896,N_5404);
and U10660 (N_10660,N_8977,N_5515);
xnor U10661 (N_10661,N_8795,N_7924);
nor U10662 (N_10662,N_8951,N_7391);
nand U10663 (N_10663,N_5841,N_6127);
and U10664 (N_10664,N_9463,N_6591);
and U10665 (N_10665,N_9005,N_6659);
and U10666 (N_10666,N_7933,N_5894);
and U10667 (N_10667,N_8642,N_7248);
or U10668 (N_10668,N_7961,N_7925);
nand U10669 (N_10669,N_8627,N_8834);
and U10670 (N_10670,N_7340,N_8167);
nand U10671 (N_10671,N_6758,N_7629);
and U10672 (N_10672,N_8091,N_8594);
nor U10673 (N_10673,N_7790,N_6545);
and U10674 (N_10674,N_5338,N_8261);
nand U10675 (N_10675,N_9594,N_7670);
xnor U10676 (N_10676,N_5133,N_8000);
xor U10677 (N_10677,N_7255,N_8248);
xor U10678 (N_10678,N_5560,N_5020);
nor U10679 (N_10679,N_5025,N_7505);
or U10680 (N_10680,N_6962,N_9406);
and U10681 (N_10681,N_7152,N_7023);
and U10682 (N_10682,N_7389,N_9631);
nor U10683 (N_10683,N_9670,N_9689);
xor U10684 (N_10684,N_9859,N_7913);
nor U10685 (N_10685,N_8758,N_9425);
xnor U10686 (N_10686,N_7163,N_7513);
and U10687 (N_10687,N_5746,N_7020);
or U10688 (N_10688,N_6844,N_5831);
or U10689 (N_10689,N_9203,N_5087);
nor U10690 (N_10690,N_7968,N_7856);
or U10691 (N_10691,N_9222,N_8250);
nand U10692 (N_10692,N_9480,N_9141);
nor U10693 (N_10693,N_8948,N_9491);
nand U10694 (N_10694,N_8138,N_8069);
or U10695 (N_10695,N_8332,N_5542);
or U10696 (N_10696,N_9613,N_9915);
nand U10697 (N_10697,N_9562,N_7656);
nand U10698 (N_10698,N_8532,N_5477);
and U10699 (N_10699,N_5786,N_8835);
xnor U10700 (N_10700,N_8818,N_5633);
xor U10701 (N_10701,N_8560,N_5480);
or U10702 (N_10702,N_7907,N_5117);
xnor U10703 (N_10703,N_5697,N_8286);
nor U10704 (N_10704,N_8615,N_8762);
and U10705 (N_10705,N_6594,N_8072);
xor U10706 (N_10706,N_7857,N_9541);
xnor U10707 (N_10707,N_6462,N_9537);
nor U10708 (N_10708,N_5778,N_7806);
xnor U10709 (N_10709,N_5527,N_6713);
nor U10710 (N_10710,N_8803,N_9696);
and U10711 (N_10711,N_7046,N_6161);
or U10712 (N_10712,N_8045,N_9638);
nor U10713 (N_10713,N_8210,N_6823);
xor U10714 (N_10714,N_5082,N_8943);
nand U10715 (N_10715,N_8528,N_6391);
nand U10716 (N_10716,N_8304,N_8199);
nor U10717 (N_10717,N_6699,N_5333);
xor U10718 (N_10718,N_8411,N_6600);
nor U10719 (N_10719,N_6606,N_8229);
nand U10720 (N_10720,N_5151,N_9296);
nor U10721 (N_10721,N_5347,N_5877);
xnor U10722 (N_10722,N_6791,N_9620);
or U10723 (N_10723,N_6410,N_7168);
nor U10724 (N_10724,N_6304,N_7512);
nor U10725 (N_10725,N_7398,N_5810);
xor U10726 (N_10726,N_6122,N_8369);
and U10727 (N_10727,N_6957,N_8794);
or U10728 (N_10728,N_6055,N_6722);
nand U10729 (N_10729,N_5636,N_9058);
nor U10730 (N_10730,N_6325,N_5180);
or U10731 (N_10731,N_8058,N_5195);
and U10732 (N_10732,N_8690,N_5379);
nor U10733 (N_10733,N_9336,N_9021);
or U10734 (N_10734,N_7247,N_7268);
and U10735 (N_10735,N_7284,N_6737);
and U10736 (N_10736,N_6202,N_9182);
and U10737 (N_10737,N_8693,N_8066);
nor U10738 (N_10738,N_5038,N_7009);
nor U10739 (N_10739,N_7949,N_8094);
or U10740 (N_10740,N_7403,N_6213);
nor U10741 (N_10741,N_9221,N_6301);
or U10742 (N_10742,N_7356,N_7242);
nor U10743 (N_10743,N_5916,N_9618);
nor U10744 (N_10744,N_9342,N_5092);
nor U10745 (N_10745,N_9554,N_5951);
nand U10746 (N_10746,N_5596,N_9042);
or U10747 (N_10747,N_5318,N_6875);
xor U10748 (N_10748,N_9467,N_7881);
or U10749 (N_10749,N_8289,N_7344);
nor U10750 (N_10750,N_8155,N_9064);
and U10751 (N_10751,N_5994,N_5728);
xnor U10752 (N_10752,N_7057,N_9828);
and U10753 (N_10753,N_7784,N_6853);
nand U10754 (N_10754,N_9535,N_5235);
xnor U10755 (N_10755,N_6516,N_5755);
nand U10756 (N_10756,N_5617,N_5442);
and U10757 (N_10757,N_6336,N_6124);
xor U10758 (N_10758,N_7282,N_9540);
and U10759 (N_10759,N_6262,N_8112);
or U10760 (N_10760,N_9579,N_8688);
nand U10761 (N_10761,N_5103,N_9479);
or U10762 (N_10762,N_9198,N_7658);
xor U10763 (N_10763,N_7014,N_8158);
nand U10764 (N_10764,N_9610,N_7865);
nor U10765 (N_10765,N_8495,N_5753);
nand U10766 (N_10766,N_7660,N_5619);
xnor U10767 (N_10767,N_9164,N_5389);
xor U10768 (N_10768,N_9886,N_7083);
nand U10769 (N_10769,N_5867,N_5062);
xor U10770 (N_10770,N_7504,N_7984);
nand U10771 (N_10771,N_5641,N_8393);
nor U10772 (N_10772,N_8575,N_5193);
nand U10773 (N_10773,N_9316,N_7452);
or U10774 (N_10774,N_6423,N_6402);
and U10775 (N_10775,N_5194,N_6020);
and U10776 (N_10776,N_6062,N_8584);
and U10777 (N_10777,N_5763,N_8869);
or U10778 (N_10778,N_8849,N_9665);
or U10779 (N_10779,N_5624,N_5628);
nand U10780 (N_10780,N_8917,N_6489);
xor U10781 (N_10781,N_5201,N_6027);
or U10782 (N_10782,N_8231,N_7974);
nor U10783 (N_10783,N_9500,N_9955);
nor U10784 (N_10784,N_5972,N_9962);
nor U10785 (N_10785,N_8184,N_6157);
xnor U10786 (N_10786,N_7067,N_8376);
nor U10787 (N_10787,N_5363,N_5918);
nor U10788 (N_10788,N_6173,N_8965);
and U10789 (N_10789,N_7026,N_9363);
nor U10790 (N_10790,N_6748,N_7986);
xor U10791 (N_10791,N_6833,N_9063);
or U10792 (N_10792,N_5980,N_6967);
nor U10793 (N_10793,N_8654,N_9806);
or U10794 (N_10794,N_8322,N_9265);
or U10795 (N_10795,N_7727,N_7141);
and U10796 (N_10796,N_9916,N_9012);
nand U10797 (N_10797,N_6707,N_8318);
or U10798 (N_10798,N_8294,N_5445);
or U10799 (N_10799,N_9793,N_7814);
xor U10800 (N_10800,N_7326,N_8319);
nor U10801 (N_10801,N_8148,N_7263);
xor U10802 (N_10802,N_5934,N_8781);
or U10803 (N_10803,N_7224,N_8041);
nor U10804 (N_10804,N_9008,N_9464);
xnor U10805 (N_10805,N_5396,N_7465);
and U10806 (N_10806,N_8827,N_7531);
xor U10807 (N_10807,N_9964,N_5683);
nand U10808 (N_10808,N_8263,N_7039);
and U10809 (N_10809,N_7486,N_8924);
xnor U10810 (N_10810,N_6414,N_5159);
or U10811 (N_10811,N_8423,N_8634);
nand U10812 (N_10812,N_5985,N_7337);
xnor U10813 (N_10813,N_8116,N_9055);
xnor U10814 (N_10814,N_5225,N_6341);
nand U10815 (N_10815,N_5237,N_6736);
nand U10816 (N_10816,N_7365,N_7922);
xnor U10817 (N_10817,N_5901,N_7308);
or U10818 (N_10818,N_5897,N_9603);
nand U10819 (N_10819,N_5229,N_9083);
nor U10820 (N_10820,N_9903,N_7492);
nand U10821 (N_10821,N_9947,N_5286);
nor U10822 (N_10822,N_7717,N_6847);
xor U10823 (N_10823,N_6227,N_8891);
or U10824 (N_10824,N_6559,N_7891);
xnor U10825 (N_10825,N_9627,N_9135);
or U10826 (N_10826,N_5686,N_9739);
xor U10827 (N_10827,N_9857,N_7801);
xnor U10828 (N_10828,N_7107,N_5708);
nand U10829 (N_10829,N_5453,N_5399);
and U10830 (N_10830,N_5802,N_7092);
xnor U10831 (N_10831,N_9755,N_7544);
xnor U10832 (N_10832,N_7342,N_6834);
nor U10833 (N_10833,N_9741,N_8445);
xnor U10834 (N_10834,N_6690,N_6685);
or U10835 (N_10835,N_7823,N_9494);
xnor U10836 (N_10836,N_8288,N_7736);
nand U10837 (N_10837,N_8635,N_8293);
nor U10838 (N_10838,N_9867,N_6067);
nor U10839 (N_10839,N_7996,N_8542);
and U10840 (N_10840,N_8821,N_6403);
xnor U10841 (N_10841,N_5023,N_9466);
nor U10842 (N_10842,N_9018,N_5114);
xnor U10843 (N_10843,N_5779,N_6979);
nand U10844 (N_10844,N_8843,N_8431);
xnor U10845 (N_10845,N_9989,N_9979);
and U10846 (N_10846,N_8503,N_6376);
and U10847 (N_10847,N_9389,N_6158);
and U10848 (N_10848,N_5482,N_5427);
or U10849 (N_10849,N_6587,N_6603);
xor U10850 (N_10850,N_7332,N_6703);
nand U10851 (N_10851,N_5116,N_5292);
or U10852 (N_10852,N_6466,N_6330);
xnor U10853 (N_10853,N_8592,N_7299);
nor U10854 (N_10854,N_7854,N_9765);
or U10855 (N_10855,N_9509,N_7068);
xor U10856 (N_10856,N_7335,N_7483);
xnor U10857 (N_10857,N_6747,N_6958);
and U10858 (N_10858,N_7441,N_5701);
xor U10859 (N_10859,N_8234,N_9570);
or U10860 (N_10860,N_8822,N_6922);
nand U10861 (N_10861,N_9353,N_7058);
or U10862 (N_10862,N_5437,N_9413);
nand U10863 (N_10863,N_5887,N_7560);
xnor U10864 (N_10864,N_6206,N_5765);
or U10865 (N_10865,N_7454,N_8972);
nand U10866 (N_10866,N_6507,N_7378);
and U10867 (N_10867,N_9197,N_9596);
nand U10868 (N_10868,N_9682,N_6935);
nor U10869 (N_10869,N_6776,N_8008);
or U10870 (N_10870,N_7312,N_8093);
xor U10871 (N_10871,N_5607,N_6387);
and U10872 (N_10872,N_8817,N_7368);
and U10873 (N_10873,N_6639,N_6348);
xor U10874 (N_10874,N_5620,N_7484);
and U10875 (N_10875,N_6821,N_9259);
or U10876 (N_10876,N_7084,N_7420);
xnor U10877 (N_10877,N_5238,N_7424);
nand U10878 (N_10878,N_7540,N_8460);
xnor U10879 (N_10879,N_6904,N_7064);
nand U10880 (N_10880,N_8650,N_9971);
nand U10881 (N_10881,N_7981,N_5141);
and U10882 (N_10882,N_5984,N_9437);
and U10883 (N_10883,N_6497,N_7085);
and U10884 (N_10884,N_8723,N_9187);
xnor U10885 (N_10885,N_6851,N_9972);
xnor U10886 (N_10886,N_7030,N_9368);
xor U10887 (N_10887,N_7834,N_7462);
and U10888 (N_10888,N_9536,N_5302);
or U10889 (N_10889,N_9788,N_5070);
nand U10890 (N_10890,N_8527,N_5295);
nor U10891 (N_10891,N_5853,N_5003);
nor U10892 (N_10892,N_6305,N_9163);
nor U10893 (N_10893,N_7394,N_5602);
nor U10894 (N_10894,N_5375,N_6231);
xor U10895 (N_10895,N_8191,N_8471);
xnor U10896 (N_10896,N_5937,N_6293);
nand U10897 (N_10897,N_9621,N_7417);
nor U10898 (N_10898,N_7469,N_8779);
and U10899 (N_10899,N_7644,N_5673);
and U10900 (N_10900,N_7457,N_7129);
and U10901 (N_10901,N_6170,N_7795);
xnor U10902 (N_10902,N_8481,N_8135);
xnor U10903 (N_10903,N_5325,N_9144);
nor U10904 (N_10904,N_7598,N_6978);
xnor U10905 (N_10905,N_7882,N_9308);
nand U10906 (N_10906,N_7072,N_9155);
nor U10907 (N_10907,N_5089,N_5346);
or U10908 (N_10908,N_7932,N_8159);
xor U10909 (N_10909,N_7451,N_9409);
or U10910 (N_10910,N_5848,N_6539);
or U10911 (N_10911,N_7223,N_8936);
nor U10912 (N_10912,N_9592,N_6689);
nor U10913 (N_10913,N_5296,N_6708);
xor U10914 (N_10914,N_7447,N_9365);
xor U10915 (N_10915,N_8090,N_6011);
nor U10916 (N_10916,N_8938,N_6131);
and U10917 (N_10917,N_8646,N_5762);
or U10918 (N_10918,N_5645,N_9518);
xnor U10919 (N_10919,N_6632,N_5138);
and U10920 (N_10920,N_9526,N_7049);
xor U10921 (N_10921,N_7574,N_5570);
or U10922 (N_10922,N_7114,N_6779);
xnor U10923 (N_10923,N_7900,N_7063);
and U10924 (N_10924,N_8873,N_7976);
xor U10925 (N_10925,N_5595,N_5666);
or U10926 (N_10926,N_5905,N_5275);
and U10927 (N_10927,N_6334,N_9104);
nor U10928 (N_10928,N_7237,N_9116);
xor U10929 (N_10929,N_7111,N_8143);
nor U10930 (N_10930,N_6415,N_8215);
and U10931 (N_10931,N_9894,N_7151);
or U10932 (N_10932,N_7620,N_9487);
nor U10933 (N_10933,N_9195,N_9565);
xor U10934 (N_10934,N_9011,N_7916);
xor U10935 (N_10935,N_7950,N_7080);
nand U10936 (N_10936,N_7594,N_7279);
nor U10937 (N_10937,N_9462,N_8862);
nor U10938 (N_10938,N_5435,N_5349);
nand U10939 (N_10939,N_6491,N_5811);
nor U10940 (N_10940,N_7350,N_9551);
nand U10941 (N_10941,N_9210,N_5795);
nand U10942 (N_10942,N_9818,N_5370);
and U10943 (N_10943,N_9640,N_6168);
xnor U10944 (N_10944,N_8919,N_9419);
or U10945 (N_10945,N_5423,N_8443);
nor U10946 (N_10946,N_6345,N_9855);
xor U10947 (N_10947,N_9407,N_9553);
or U10948 (N_10948,N_7863,N_6687);
and U10949 (N_10949,N_5915,N_8273);
and U10950 (N_10950,N_7466,N_9815);
or U10951 (N_10951,N_5160,N_9841);
or U10952 (N_10952,N_6118,N_9230);
and U10953 (N_10953,N_7295,N_9775);
nor U10954 (N_10954,N_9965,N_9082);
or U10955 (N_10955,N_8435,N_7905);
nand U10956 (N_10956,N_8306,N_5649);
nor U10957 (N_10957,N_9092,N_5899);
nor U10958 (N_10958,N_9936,N_9037);
nand U10959 (N_10959,N_5440,N_8189);
xnor U10960 (N_10960,N_7397,N_9410);
xor U10961 (N_10961,N_8854,N_5731);
and U10962 (N_10962,N_5585,N_6933);
nand U10963 (N_10963,N_6167,N_6456);
or U10964 (N_10964,N_7476,N_5053);
or U10965 (N_10965,N_9685,N_9225);
nand U10966 (N_10966,N_8997,N_7539);
nor U10967 (N_10967,N_6752,N_9810);
and U10968 (N_10968,N_8039,N_9598);
nand U10969 (N_10969,N_5134,N_9833);
xnor U10970 (N_10970,N_5219,N_9347);
and U10971 (N_10971,N_6985,N_9794);
nand U10972 (N_10972,N_6176,N_7726);
or U10973 (N_10973,N_9901,N_7761);
or U10974 (N_10974,N_7254,N_8071);
and U10975 (N_10975,N_7077,N_9605);
xor U10976 (N_10976,N_9838,N_7162);
nor U10977 (N_10977,N_6145,N_6835);
and U10978 (N_10978,N_9415,N_6077);
or U10979 (N_10979,N_7855,N_8177);
and U10980 (N_10980,N_9986,N_8081);
nor U10981 (N_10981,N_8874,N_7669);
and U10982 (N_10982,N_9939,N_6100);
or U10983 (N_10983,N_8605,N_8620);
or U10984 (N_10984,N_9443,N_5426);
xnor U10985 (N_10985,N_7917,N_6934);
xnor U10986 (N_10986,N_5948,N_8886);
xor U10987 (N_10987,N_7647,N_7421);
or U10988 (N_10988,N_7321,N_7828);
nand U10989 (N_10989,N_6288,N_8499);
nor U10990 (N_10990,N_5386,N_8491);
nor U10991 (N_10991,N_6327,N_5234);
xnor U10992 (N_10992,N_5692,N_9319);
xor U10993 (N_10993,N_7110,N_8337);
and U10994 (N_10994,N_7733,N_5499);
nor U10995 (N_10995,N_6187,N_7935);
xnor U10996 (N_10996,N_8954,N_6717);
or U10997 (N_10997,N_8283,N_7027);
nor U10998 (N_10998,N_5715,N_8444);
or U10999 (N_10999,N_7829,N_6237);
and U11000 (N_11000,N_7375,N_5443);
nor U11001 (N_11001,N_8307,N_8677);
or U11002 (N_11002,N_8866,N_7297);
xnor U11003 (N_11003,N_8911,N_7554);
nor U11004 (N_11004,N_9599,N_7059);
nor U11005 (N_11005,N_9914,N_7695);
nand U11006 (N_11006,N_8720,N_6574);
and U11007 (N_11007,N_9626,N_6784);
nand U11008 (N_11008,N_5299,N_8741);
xnor U11009 (N_11009,N_8102,N_5205);
and U11010 (N_11010,N_7654,N_8466);
xor U11011 (N_11011,N_8974,N_9219);
or U11012 (N_11012,N_7939,N_6766);
nand U11013 (N_11013,N_9931,N_7137);
and U11014 (N_11014,N_9339,N_8124);
nand U11015 (N_11015,N_9152,N_5202);
nor U11016 (N_11016,N_9534,N_7164);
nor U11017 (N_11017,N_7745,N_7217);
xnor U11018 (N_11018,N_8727,N_9953);
xnor U11019 (N_11019,N_8204,N_7936);
nand U11020 (N_11020,N_7682,N_9652);
and U11021 (N_11021,N_6831,N_9907);
and U11022 (N_11022,N_7989,N_8419);
and U11023 (N_11023,N_7715,N_9061);
nand U11024 (N_11024,N_7220,N_7506);
or U11025 (N_11025,N_9178,N_8019);
nor U11026 (N_11026,N_5209,N_9282);
xnor U11027 (N_11027,N_8772,N_7314);
and U11028 (N_11028,N_5647,N_7769);
xor U11029 (N_11029,N_8114,N_9110);
xor U11030 (N_11030,N_8706,N_9470);
nor U11031 (N_11031,N_8464,N_8237);
nand U11032 (N_11032,N_7425,N_9969);
nor U11033 (N_11033,N_8582,N_9520);
nand U11034 (N_11034,N_6216,N_7087);
nand U11035 (N_11035,N_6886,N_5874);
and U11036 (N_11036,N_7877,N_6047);
or U11037 (N_11037,N_8796,N_7489);
and U11038 (N_11038,N_5065,N_6164);
nand U11039 (N_11039,N_7827,N_9361);
and U11040 (N_11040,N_5860,N_6061);
or U11041 (N_11041,N_5716,N_9449);
xnor U11042 (N_11042,N_6484,N_6620);
or U11043 (N_11043,N_8638,N_8062);
and U11044 (N_11044,N_5113,N_8010);
nand U11045 (N_11045,N_7260,N_6910);
nand U11046 (N_11046,N_7239,N_9254);
and U11047 (N_11047,N_7583,N_6928);
and U11048 (N_11048,N_7520,N_6867);
nor U11049 (N_11049,N_9237,N_7983);
xor U11050 (N_11050,N_5592,N_7572);
and U11051 (N_11051,N_6224,N_8365);
xnor U11052 (N_11052,N_8641,N_7543);
nor U11053 (N_11053,N_7309,N_5608);
and U11054 (N_11054,N_5048,N_9251);
or U11055 (N_11055,N_9264,N_6996);
xor U11056 (N_11056,N_6135,N_7713);
nand U11057 (N_11057,N_5233,N_6994);
nor U11058 (N_11058,N_5583,N_6813);
nand U11059 (N_11059,N_8003,N_9819);
nor U11060 (N_11060,N_7942,N_9980);
or U11061 (N_11061,N_7448,N_8374);
xor U11062 (N_11062,N_9811,N_9006);
or U11063 (N_11063,N_6184,N_8368);
nand U11064 (N_11064,N_9556,N_5425);
nand U11065 (N_11065,N_5283,N_9453);
and U11066 (N_11066,N_5156,N_8163);
xnor U11067 (N_11067,N_5118,N_8061);
xnor U11068 (N_11068,N_7171,N_6829);
nand U11069 (N_11069,N_9913,N_5975);
nor U11070 (N_11070,N_5840,N_6614);
and U11071 (N_11071,N_5126,N_5174);
nor U11072 (N_11072,N_6795,N_5835);
xnor U11073 (N_11073,N_5931,N_8051);
xnor U11074 (N_11074,N_8301,N_5319);
or U11075 (N_11075,N_6279,N_6929);
and U11076 (N_11076,N_9193,N_6907);
xnor U11077 (N_11077,N_7563,N_9293);
and U11078 (N_11078,N_6281,N_8801);
nor U11079 (N_11079,N_8459,N_8786);
or U11080 (N_11080,N_7227,N_9845);
xnor U11081 (N_11081,N_5546,N_6215);
and U11082 (N_11082,N_8474,N_6081);
and U11083 (N_11083,N_8511,N_8054);
and U11084 (N_11084,N_9729,N_7471);
or U11085 (N_11085,N_8207,N_6787);
nor U11086 (N_11086,N_8082,N_9337);
or U11087 (N_11087,N_8222,N_8298);
nand U11088 (N_11088,N_6287,N_7218);
nor U11089 (N_11089,N_6326,N_5458);
or U11090 (N_11090,N_5378,N_8217);
or U11091 (N_11091,N_8305,N_5342);
and U11092 (N_11092,N_9849,N_7043);
xnor U11093 (N_11093,N_6734,N_9239);
nor U11094 (N_11094,N_9519,N_8562);
nor U11095 (N_11095,N_8861,N_5197);
or U11096 (N_11096,N_5096,N_8944);
and U11097 (N_11097,N_5541,N_9093);
or U11098 (N_11098,N_8325,N_7930);
nor U11099 (N_11099,N_5166,N_7065);
and U11100 (N_11100,N_8692,N_7557);
nand U11101 (N_11101,N_7605,N_7698);
nor U11102 (N_11102,N_5859,N_9180);
nor U11103 (N_11103,N_7837,N_5198);
nor U11104 (N_11104,N_6444,N_8371);
and U11105 (N_11105,N_5942,N_6302);
and U11106 (N_11106,N_9985,N_6175);
nand U11107 (N_11107,N_8136,N_5723);
nand U11108 (N_11108,N_8505,N_6974);
or U11109 (N_11109,N_8731,N_8129);
nand U11110 (N_11110,N_6192,N_7215);
xnor U11111 (N_11111,N_6140,N_9999);
and U11112 (N_11112,N_6438,N_9783);
xor U11113 (N_11113,N_7526,N_8607);
nand U11114 (N_11114,N_9469,N_9813);
nor U11115 (N_11115,N_9840,N_6520);
nor U11116 (N_11116,N_8405,N_8730);
and U11117 (N_11117,N_8963,N_9988);
nand U11118 (N_11118,N_9711,N_5906);
xnor U11119 (N_11119,N_7667,N_5712);
or U11120 (N_11120,N_9960,N_6668);
xnor U11121 (N_11121,N_6042,N_9332);
and U11122 (N_11122,N_9879,N_6194);
xor U11123 (N_11123,N_5178,N_5315);
or U11124 (N_11124,N_8535,N_8567);
or U11125 (N_11125,N_8260,N_9132);
nand U11126 (N_11126,N_6038,N_7528);
and U11127 (N_11127,N_7770,N_7839);
or U11128 (N_11128,N_7138,N_5997);
and U11129 (N_11129,N_5069,N_6049);
xnor U11130 (N_11130,N_9743,N_5939);
and U11131 (N_11131,N_7285,N_7608);
nand U11132 (N_11132,N_5813,N_7721);
nor U11133 (N_11133,N_5304,N_7177);
or U11134 (N_11134,N_9414,N_5921);
nand U11135 (N_11135,N_7818,N_6504);
nor U11136 (N_11136,N_6285,N_7621);
nand U11137 (N_11137,N_8378,N_9105);
or U11138 (N_11138,N_7324,N_9646);
and U11139 (N_11139,N_8144,N_9888);
or U11140 (N_11140,N_5745,N_7291);
nor U11141 (N_11141,N_9143,N_8933);
xnor U11142 (N_11142,N_9718,N_6633);
nor U11143 (N_11143,N_9680,N_6328);
nor U11144 (N_11144,N_9170,N_9428);
nor U11145 (N_11145,N_8705,N_6450);
and U11146 (N_11146,N_9456,N_9576);
nand U11147 (N_11147,N_6162,N_8485);
nand U11148 (N_11148,N_6537,N_6342);
xnor U11149 (N_11149,N_9997,N_6741);
nand U11150 (N_11150,N_9669,N_9056);
and U11151 (N_11151,N_6684,N_6022);
nand U11152 (N_11152,N_6607,N_7269);
nand U11153 (N_11153,N_5700,N_5303);
xnor U11154 (N_11154,N_8104,N_5034);
and U11155 (N_11155,N_5888,N_6056);
xor U11156 (N_11156,N_6117,N_7370);
and U11157 (N_11157,N_8566,N_5777);
or U11158 (N_11158,N_6064,N_9938);
nand U11159 (N_11159,N_8007,N_7182);
nand U11160 (N_11160,N_7388,N_6498);
or U11161 (N_11161,N_8218,N_7288);
or U11162 (N_11162,N_7427,N_6572);
nand U11163 (N_11163,N_6700,N_9306);
nor U11164 (N_11164,N_7638,N_5646);
nor U11165 (N_11165,N_7523,N_8885);
or U11166 (N_11166,N_8816,N_5352);
or U11167 (N_11167,N_5466,N_7187);
or U11168 (N_11168,N_6388,N_6120);
xor U11169 (N_11169,N_9362,N_7346);
nand U11170 (N_11170,N_7622,N_9935);
nand U11171 (N_11171,N_6807,N_7853);
and U11172 (N_11172,N_5925,N_5657);
nand U11173 (N_11173,N_8956,N_9346);
and U11174 (N_11174,N_7252,N_5447);
and U11175 (N_11175,N_6024,N_6181);
or U11176 (N_11176,N_8985,N_5536);
nor U11177 (N_11177,N_7805,N_9730);
or U11178 (N_11178,N_5424,N_8390);
nor U11179 (N_11179,N_6503,N_5422);
nand U11180 (N_11180,N_6744,N_9747);
xor U11181 (N_11181,N_7964,N_5691);
nand U11182 (N_11182,N_5464,N_9016);
nand U11183 (N_11183,N_5973,N_5384);
and U11184 (N_11184,N_5752,N_7651);
nor U11185 (N_11185,N_6968,N_6666);
and U11186 (N_11186,N_7923,N_8243);
xnor U11187 (N_11187,N_5878,N_9378);
and U11188 (N_11188,N_8746,N_9112);
or U11189 (N_11189,N_9473,N_7134);
and U11190 (N_11190,N_5167,N_9748);
and U11191 (N_11191,N_6706,N_5903);
xor U11192 (N_11192,N_8187,N_8509);
and U11193 (N_11193,N_6490,N_9403);
nor U11194 (N_11194,N_7960,N_9583);
nor U11195 (N_11195,N_6940,N_6845);
and U11196 (N_11196,N_7845,N_8335);
nor U11197 (N_11197,N_5326,N_7276);
or U11198 (N_11198,N_6111,N_7176);
xnor U11199 (N_11199,N_7558,N_7096);
nor U11200 (N_11200,N_8265,N_7703);
nand U11201 (N_11201,N_7712,N_5405);
and U11202 (N_11202,N_8382,N_5717);
nor U11203 (N_11203,N_6870,N_7697);
and U11204 (N_11204,N_5434,N_9459);
nor U11205 (N_11205,N_6451,N_9946);
nand U11206 (N_11206,N_5974,N_6435);
and U11207 (N_11207,N_9313,N_6627);
nor U11208 (N_11208,N_9271,N_7821);
xor U11209 (N_11209,N_5750,N_7199);
or U11210 (N_11210,N_5251,N_8867);
nand U11211 (N_11211,N_5228,N_6218);
nand U11212 (N_11212,N_5879,N_9157);
nand U11213 (N_11213,N_9381,N_9961);
and U11214 (N_11214,N_8324,N_7851);
nor U11215 (N_11215,N_6577,N_7595);
xor U11216 (N_11216,N_7396,N_7216);
or U11217 (N_11217,N_7395,N_6046);
and U11218 (N_11218,N_8056,N_7319);
nand U11219 (N_11219,N_8585,N_9963);
xor U11220 (N_11220,N_7198,N_7858);
or U11221 (N_11221,N_9371,N_6806);
nand U11222 (N_11222,N_8156,N_5516);
or U11223 (N_11223,N_5725,N_7586);
or U11224 (N_11224,N_9527,N_8545);
and U11225 (N_11225,N_6130,N_7338);
nand U11226 (N_11226,N_6355,N_9512);
or U11227 (N_11227,N_7929,N_6888);
nand U11228 (N_11228,N_9476,N_6329);
or U11229 (N_11229,N_9617,N_6209);
nand U11230 (N_11230,N_5862,N_8356);
nand U11231 (N_11231,N_5519,N_9284);
nand U11232 (N_11232,N_9883,N_6960);
and U11233 (N_11233,N_5616,N_9973);
and U11234 (N_11234,N_6291,N_9676);
and U11235 (N_11235,N_6428,N_5579);
xor U11236 (N_11236,N_7566,N_8751);
and U11237 (N_11237,N_5444,N_6273);
nor U11238 (N_11238,N_5908,N_9162);
nor U11239 (N_11239,N_5415,N_8536);
nor U11240 (N_11240,N_6234,N_6483);
xor U11241 (N_11241,N_8734,N_7287);
or U11242 (N_11242,N_6997,N_8309);
or U11243 (N_11243,N_8344,N_8125);
or U11244 (N_11244,N_8518,N_8937);
nand U11245 (N_11245,N_8384,N_5578);
xnor U11246 (N_11246,N_7728,N_9681);
or U11247 (N_11247,N_9474,N_5572);
nor U11248 (N_11248,N_5058,N_9552);
or U11249 (N_11249,N_8447,N_7824);
xnor U11250 (N_11250,N_8711,N_6869);
xor U11251 (N_11251,N_6369,N_9827);
nand U11252 (N_11252,N_8767,N_9882);
nand U11253 (N_11253,N_8877,N_5773);
xnor U11254 (N_11254,N_9902,N_7082);
and U11255 (N_11255,N_7562,N_8213);
or U11256 (N_11256,N_8016,N_7191);
nor U11257 (N_11257,N_6767,N_9731);
nand U11258 (N_11258,N_5865,N_5968);
or U11259 (N_11259,N_9448,N_7788);
or U11260 (N_11260,N_9127,N_9138);
or U11261 (N_11261,N_8440,N_6488);
nor U11262 (N_11262,N_7627,N_6058);
nor U11263 (N_11263,N_7559,N_8381);
nor U11264 (N_11264,N_5330,N_7179);
or U11265 (N_11265,N_5226,N_7524);
nor U11266 (N_11266,N_8637,N_8921);
xnor U11267 (N_11267,N_5108,N_6881);
or U11268 (N_11268,N_9243,N_5127);
and U11269 (N_11269,N_9892,N_6501);
nand U11270 (N_11270,N_8648,N_7548);
xnor U11271 (N_11271,N_8059,N_8882);
and U11272 (N_11272,N_6017,N_7197);
nor U11273 (N_11273,N_5987,N_5580);
or U11274 (N_11274,N_9372,N_7318);
xor U11275 (N_11275,N_5804,N_7589);
nor U11276 (N_11276,N_8992,N_5632);
or U11277 (N_11277,N_6323,N_8847);
nor U11278 (N_11278,N_7952,N_6448);
and U11279 (N_11279,N_9258,N_7112);
and U11280 (N_11280,N_5960,N_8180);
or U11281 (N_11281,N_5460,N_8055);
nor U11282 (N_11282,N_5555,N_6526);
and U11283 (N_11283,N_5713,N_6656);
or U11284 (N_11284,N_7604,N_9593);
or U11285 (N_11285,N_5414,N_7768);
and U11286 (N_11286,N_8198,N_9421);
nor U11287 (N_11287,N_5242,N_6424);
xor U11288 (N_11288,N_8426,N_6198);
or U11289 (N_11289,N_8725,N_6663);
xor U11290 (N_11290,N_8255,N_9647);
nand U11291 (N_11291,N_5291,N_9072);
nor U11292 (N_11292,N_6045,N_7987);
or U11293 (N_11293,N_5832,N_8947);
or U11294 (N_11294,N_6952,N_8580);
nand U11295 (N_11295,N_5106,N_9508);
xnor U11296 (N_11296,N_5051,N_5969);
xor U11297 (N_11297,N_5936,N_5993);
nand U11298 (N_11298,N_6696,N_7170);
nor U11299 (N_11299,N_8096,N_6258);
nand U11300 (N_11300,N_6005,N_9653);
nand U11301 (N_11301,N_7759,N_5416);
xnor U11302 (N_11302,N_8026,N_5798);
or U11303 (N_11303,N_7861,N_6864);
and U11304 (N_11304,N_9968,N_6245);
nand U11305 (N_11305,N_7895,N_7160);
nor U11306 (N_11306,N_9773,N_6786);
or U11307 (N_11307,N_7789,N_8246);
or U11308 (N_11308,N_9325,N_5014);
xor U11309 (N_11309,N_9984,N_5046);
and U11310 (N_11310,N_5314,N_5950);
nand U11311 (N_11311,N_5121,N_9168);
xor U11312 (N_11312,N_5263,N_6137);
nor U11313 (N_11313,N_5775,N_6660);
and U11314 (N_11314,N_7776,N_8490);
nor U11315 (N_11315,N_9102,N_5500);
nor U11316 (N_11316,N_9125,N_8502);
nor U11317 (N_11317,N_5393,N_8837);
nor U11318 (N_11318,N_9524,N_5467);
nand U11319 (N_11319,N_9735,N_7419);
xor U11320 (N_11320,N_9196,N_8117);
xor U11321 (N_11321,N_7649,N_5743);
nand U11322 (N_11322,N_9862,N_6513);
xnor U11323 (N_11323,N_6861,N_9612);
nand U11324 (N_11324,N_6470,N_7780);
and U11325 (N_11325,N_9272,N_5789);
xor U11326 (N_11326,N_8406,N_6457);
nor U11327 (N_11327,N_7602,N_7339);
nor U11328 (N_11328,N_9069,N_9778);
nor U11329 (N_11329,N_6495,N_6009);
and U11330 (N_11330,N_9402,N_9048);
or U11331 (N_11331,N_6515,N_6743);
nand U11332 (N_11332,N_9183,N_9194);
and U11333 (N_11333,N_8327,N_9514);
nand U11334 (N_11334,N_8328,N_7386);
nand U11335 (N_11335,N_6460,N_7879);
or U11336 (N_11336,N_9905,N_9702);
or U11337 (N_11337,N_7300,N_7798);
nand U11338 (N_11338,N_7617,N_8888);
nand U11339 (N_11339,N_8223,N_5718);
nor U11340 (N_11340,N_6280,N_8941);
nand U11341 (N_11341,N_7455,N_7793);
nor U11342 (N_11342,N_6771,N_6115);
nand U11343 (N_11343,N_6480,N_5041);
or U11344 (N_11344,N_5432,N_8402);
and U11345 (N_11345,N_9446,N_7053);
nor U11346 (N_11346,N_9602,N_5502);
nor U11347 (N_11347,N_9728,N_5331);
xor U11348 (N_11348,N_7725,N_6446);
nor U11349 (N_11349,N_8086,N_9814);
nand U11350 (N_11350,N_5107,N_7002);
or U11351 (N_11351,N_5917,N_8162);
or U11352 (N_11352,N_5520,N_5261);
nand U11353 (N_11353,N_6812,N_8147);
or U11354 (N_11354,N_9388,N_7716);
nand U11355 (N_11355,N_6443,N_5629);
or U11356 (N_11356,N_6073,N_6811);
nor U11357 (N_11357,N_9764,N_9659);
nand U11358 (N_11358,N_6617,N_7683);
or U11359 (N_11359,N_6927,N_6312);
nand U11360 (N_11360,N_8244,N_9615);
or U11361 (N_11361,N_6210,N_5465);
nor U11362 (N_11362,N_9528,N_8131);
or U11363 (N_11363,N_7097,N_6413);
and U11364 (N_11364,N_8266,N_9114);
or U11365 (N_11365,N_9228,N_9085);
or U11366 (N_11366,N_6189,N_8192);
and U11367 (N_11367,N_9266,N_6200);
xor U11368 (N_11368,N_9777,N_5406);
xnor U11369 (N_11369,N_7642,N_6874);
nor U11370 (N_11370,N_9928,N_5807);
nand U11371 (N_11371,N_5009,N_5088);
nor U11372 (N_11372,N_7280,N_8656);
xor U11373 (N_11373,N_7066,N_6622);
and U11374 (N_11374,N_9050,N_7174);
nand U11375 (N_11375,N_7456,N_7830);
and U11376 (N_11376,N_5790,N_8604);
or U11377 (N_11377,N_8668,N_9427);
xnor U11378 (N_11378,N_6785,N_9667);
xnor U11379 (N_11379,N_6745,N_5192);
nor U11380 (N_11380,N_5707,N_6763);
or U11381 (N_11381,N_5537,N_7585);
or U11382 (N_11382,N_6385,N_7796);
or U11383 (N_11383,N_7277,N_9726);
xnor U11384 (N_11384,N_9733,N_8480);
nand U11385 (N_11385,N_7973,N_7630);
nand U11386 (N_11386,N_9559,N_8754);
nor U11387 (N_11387,N_6509,N_9173);
nor U11388 (N_11388,N_8667,N_6500);
or U11389 (N_11389,N_9538,N_7815);
and U11390 (N_11390,N_6846,N_6068);
nand U11391 (N_11391,N_5549,N_7850);
and U11392 (N_11392,N_7301,N_7117);
nand U11393 (N_11393,N_8161,N_7537);
or U11394 (N_11394,N_7104,N_8546);
or U11395 (N_11395,N_7098,N_6618);
nand U11396 (N_11396,N_5410,N_6132);
nor U11397 (N_11397,N_9875,N_8361);
nand U11398 (N_11398,N_5231,N_7371);
xnor U11399 (N_11399,N_7444,N_5448);
or U11400 (N_11400,N_7416,N_7693);
nor U11401 (N_11401,N_9829,N_5662);
or U11402 (N_11402,N_6971,N_9312);
or U11403 (N_11403,N_5761,N_8285);
and U11404 (N_11404,N_6097,N_9395);
or U11405 (N_11405,N_8025,N_6796);
or U11406 (N_11406,N_8433,N_7034);
and U11407 (N_11407,N_9478,N_6063);
and U11408 (N_11408,N_5754,N_7601);
nor U11409 (N_11409,N_8168,N_9472);
nand U11410 (N_11410,N_7508,N_7225);
and U11411 (N_11411,N_7551,N_7739);
and U11412 (N_11412,N_8221,N_6002);
nor U11413 (N_11413,N_5222,N_7461);
and U11414 (N_11414,N_9153,N_6547);
or U11415 (N_11415,N_7352,N_6628);
or U11416 (N_11416,N_5622,N_6702);
or U11417 (N_11417,N_6350,N_6040);
nand U11418 (N_11418,N_6048,N_5990);
xor U11419 (N_11419,N_6420,N_7958);
and U11420 (N_11420,N_7990,N_8484);
nor U11421 (N_11421,N_8173,N_6274);
or U11422 (N_11422,N_6085,N_7292);
nor U11423 (N_11423,N_9648,N_6232);
nand U11424 (N_11424,N_9851,N_7013);
or U11425 (N_11425,N_6802,N_8506);
and U11426 (N_11426,N_6016,N_7568);
xor U11427 (N_11427,N_9797,N_6859);
or U11428 (N_11428,N_5898,N_5388);
nand U11429 (N_11429,N_6868,N_6728);
and U11430 (N_11430,N_8498,N_7401);
and U11431 (N_11431,N_8704,N_9333);
xor U11432 (N_11432,N_9475,N_7762);
or U11433 (N_11433,N_8409,N_9430);
xor U11434 (N_11434,N_8407,N_7696);
and U11435 (N_11435,N_9569,N_9959);
nand U11436 (N_11436,N_7893,N_8957);
xnor U11437 (N_11437,N_9588,N_6089);
nand U11438 (N_11438,N_8038,N_5336);
nor U11439 (N_11439,N_7719,N_6264);
nand U11440 (N_11440,N_6196,N_5864);
and U11441 (N_11441,N_8666,N_5787);
nand U11442 (N_11442,N_5450,N_8998);
or U11443 (N_11443,N_8864,N_9917);
nor U11444 (N_11444,N_5526,N_8029);
nand U11445 (N_11445,N_9192,N_5693);
and U11446 (N_11446,N_9240,N_7190);
nor U11447 (N_11447,N_9253,N_9591);
or U11448 (N_11448,N_6658,N_9772);
and U11449 (N_11449,N_6185,N_5971);
nor U11450 (N_11450,N_9315,N_6970);
or U11451 (N_11451,N_5524,N_5540);
xnor U11452 (N_11452,N_8232,N_6220);
nand U11453 (N_11453,N_6199,N_9457);
nand U11454 (N_11454,N_6655,N_5007);
nor U11455 (N_11455,N_9499,N_8525);
and U11456 (N_11456,N_9159,N_5854);
or U11457 (N_11457,N_5564,N_9557);
nor U11458 (N_11458,N_9799,N_5073);
nor U11459 (N_11459,N_6339,N_7184);
nand U11460 (N_11460,N_6602,N_6749);
or U11461 (N_11461,N_9423,N_6095);
nand U11462 (N_11462,N_9677,N_6595);
nand U11463 (N_11463,N_6422,N_5721);
nand U11464 (N_11464,N_5136,N_9024);
or U11465 (N_11465,N_5771,N_6636);
and U11466 (N_11466,N_8354,N_6697);
nor U11467 (N_11467,N_5886,N_6433);
and U11468 (N_11468,N_9028,N_6560);
and U11469 (N_11469,N_7640,N_5000);
or U11470 (N_11470,N_5735,N_6754);
or U11471 (N_11471,N_8587,N_5533);
or U11472 (N_11472,N_8732,N_7345);
xnor U11473 (N_11473,N_6467,N_8593);
or U11474 (N_11474,N_6390,N_9785);
and U11475 (N_11475,N_7701,N_9358);
nor U11476 (N_11476,N_9236,N_9790);
or U11477 (N_11477,N_9081,N_8645);
and U11478 (N_11478,N_6317,N_5104);
nand U11479 (N_11479,N_8006,N_9564);
and U11480 (N_11480,N_7832,N_6284);
nand U11481 (N_11481,N_6151,N_5529);
xor U11482 (N_11482,N_7535,N_5522);
and U11483 (N_11483,N_8472,N_7514);
or U11484 (N_11484,N_8790,N_7178);
nor U11485 (N_11485,N_9517,N_8841);
nand U11486 (N_11486,N_7849,N_8831);
nand U11487 (N_11487,N_6612,N_7033);
nand U11488 (N_11488,N_6365,N_5759);
nor U11489 (N_11489,N_6588,N_8932);
nor U11490 (N_11490,N_9335,N_6112);
xor U11491 (N_11491,N_8314,N_8927);
nor U11492 (N_11492,N_5374,N_7131);
nand U11493 (N_11493,N_8555,N_9768);
nor U11494 (N_11494,N_7878,N_5493);
or U11495 (N_11495,N_9172,N_6254);
or U11496 (N_11496,N_7515,N_9165);
xor U11497 (N_11497,N_5696,N_7387);
xnor U11498 (N_11498,N_5068,N_8769);
nor U11499 (N_11499,N_7443,N_7686);
xor U11500 (N_11500,N_5563,N_7118);
xnor U11501 (N_11501,N_5150,N_6125);
xnor U11502 (N_11502,N_6669,N_6473);
and U11503 (N_11503,N_8031,N_8991);
and U11504 (N_11504,N_8287,N_9941);
or U11505 (N_11505,N_6852,N_9370);
xor U11506 (N_11506,N_6565,N_7273);
and U11507 (N_11507,N_5868,N_7479);
xnor U11508 (N_11508,N_6051,N_6139);
and U11509 (N_11509,N_5719,N_5262);
nand U11510 (N_11510,N_8271,N_9981);
and U11511 (N_11511,N_6556,N_6217);
nand U11512 (N_11512,N_8664,N_8622);
or U11513 (N_11513,N_8558,N_9622);
xor U11514 (N_11514,N_5006,N_7348);
nor U11515 (N_11515,N_7432,N_6102);
and U11516 (N_11516,N_7459,N_6166);
xor U11517 (N_11517,N_5928,N_9220);
xor U11518 (N_11518,N_6975,N_6850);
or U11519 (N_11519,N_9217,N_5963);
and U11520 (N_11520,N_5816,N_6104);
and U11521 (N_11521,N_8224,N_5047);
or U11522 (N_11522,N_6392,N_5827);
nand U11523 (N_11523,N_8208,N_6977);
xor U11524 (N_11524,N_6408,N_5590);
nand U11525 (N_11525,N_5988,N_7763);
xnor U11526 (N_11526,N_9704,N_7186);
xnor U11527 (N_11527,N_6570,N_7538);
xor U11528 (N_11528,N_8291,N_5095);
or U11529 (N_11529,N_7729,N_9497);
or U11530 (N_11530,N_5866,N_9720);
xor U11531 (N_11531,N_6043,N_7547);
nor U11532 (N_11532,N_7148,N_5847);
and U11533 (N_11533,N_9495,N_5836);
and U11534 (N_11534,N_6230,N_8430);
or U11535 (N_11535,N_9392,N_9348);
or U11536 (N_11536,N_8107,N_5456);
xnor U11537 (N_11537,N_8895,N_8436);
and U11538 (N_11538,N_7723,N_7556);
nor U11539 (N_11539,N_5220,N_9998);
xnor U11540 (N_11540,N_7374,N_9097);
nor U11541 (N_11541,N_8282,N_8370);
nor U11542 (N_11542,N_5186,N_8923);
nor U11543 (N_11543,N_7862,N_5409);
nand U11544 (N_11544,N_6150,N_7599);
xnor U11545 (N_11545,N_8865,N_8950);
or U11546 (N_11546,N_7609,N_7275);
and U11547 (N_11547,N_6742,N_9744);
nor U11548 (N_11548,N_9860,N_6571);
nor U11549 (N_11549,N_5844,N_8341);
nand U11550 (N_11550,N_7799,N_6544);
nand U11551 (N_11551,N_6174,N_8078);
nand U11552 (N_11552,N_5413,N_8024);
nand U11553 (N_11553,N_7437,N_8544);
and U11554 (N_11554,N_6677,N_5239);
xor U11555 (N_11555,N_8844,N_5091);
or U11556 (N_11556,N_5001,N_8961);
nor U11557 (N_11557,N_9575,N_5593);
nand U11558 (N_11558,N_9760,N_6080);
xor U11559 (N_11559,N_8103,N_5332);
and U11560 (N_11560,N_6155,N_9013);
nand U11561 (N_11561,N_7106,N_5468);
or U11562 (N_11562,N_7102,N_6266);
nor U11563 (N_11563,N_9131,N_8432);
xor U11564 (N_11564,N_8766,N_7675);
nor U11565 (N_11565,N_6581,N_9697);
or U11566 (N_11566,N_8240,N_7303);
nor U11567 (N_11567,N_6000,N_7756);
nor U11568 (N_11568,N_6322,N_6416);
nand U11569 (N_11569,N_7820,N_9261);
nor U11570 (N_11570,N_6691,N_8550);
xor U11571 (N_11571,N_6613,N_7951);
xnor U11572 (N_11572,N_8630,N_5664);
and U11573 (N_11573,N_8643,N_8922);
or U11574 (N_11574,N_8122,N_9148);
nand U11575 (N_11575,N_5992,N_9724);
nor U11576 (N_11576,N_6106,N_9930);
or U11577 (N_11577,N_6646,N_5487);
nand U11578 (N_11578,N_6360,N_5270);
nor U11579 (N_11579,N_8421,N_9017);
xor U11580 (N_11580,N_6321,N_9580);
xor U11581 (N_11581,N_8258,N_5850);
or U11582 (N_11582,N_6634,N_6478);
or U11583 (N_11583,N_7235,N_9227);
nor U11584 (N_11584,N_8697,N_8716);
and U11585 (N_11585,N_9124,N_5818);
nand U11586 (N_11586,N_8699,N_6531);
nor U11587 (N_11587,N_9966,N_9185);
nand U11588 (N_11588,N_8174,N_5837);
and U11589 (N_11589,N_6074,N_7502);
nand U11590 (N_11590,N_9010,N_9161);
and U11591 (N_11591,N_6344,N_6735);
xor U11592 (N_11592,N_5361,N_8206);
and U11593 (N_11593,N_8631,N_8115);
or U11594 (N_11594,N_5635,N_7646);
nor U11595 (N_11595,N_5208,N_7577);
nand U11596 (N_11596,N_5553,N_7623);
nand U11597 (N_11597,N_9958,N_5244);
and U11598 (N_11598,N_7250,N_8278);
xor U11599 (N_11599,N_7898,N_5170);
nand U11600 (N_11600,N_9737,N_6028);
or U11601 (N_11601,N_5131,N_9471);
nand U11602 (N_11602,N_5475,N_9297);
nor U11603 (N_11603,N_5893,N_6789);
xor U11604 (N_11604,N_6412,N_8916);
nand U11605 (N_11605,N_6561,N_7811);
or U11606 (N_11606,N_7848,N_7740);
and U11607 (N_11607,N_5360,N_7937);
or U11608 (N_11608,N_5373,N_9577);
and U11609 (N_11609,N_7873,N_6782);
and U11610 (N_11610,N_7470,N_9286);
nand U11611 (N_11611,N_5316,N_6598);
nand U11612 (N_11612,N_8048,N_8709);
or U11613 (N_11613,N_9633,N_5157);
xnor U11614 (N_11614,N_8079,N_8508);
and U11615 (N_11615,N_8655,N_5644);
nand U11616 (N_11616,N_5013,N_5446);
nor U11617 (N_11617,N_6411,N_6399);
and U11618 (N_11618,N_9488,N_5350);
nor U11619 (N_11619,N_9820,N_8209);
xor U11620 (N_11620,N_5085,N_6294);
and U11621 (N_11621,N_9736,N_8211);
and U11622 (N_11622,N_6404,N_7071);
or U11623 (N_11623,N_6918,N_7205);
nand U11624 (N_11624,N_8571,N_8004);
nand U11625 (N_11625,N_8469,N_7357);
xnor U11626 (N_11626,N_5182,N_5838);
xor U11627 (N_11627,N_7037,N_8076);
and U11628 (N_11628,N_7889,N_5392);
and U11629 (N_11629,N_7367,N_7666);
nand U11630 (N_11630,N_7772,N_6149);
xor U11631 (N_11631,N_8563,N_5257);
or U11632 (N_11632,N_6920,N_6799);
or U11633 (N_11633,N_6397,N_8913);
or U11634 (N_11634,N_5902,N_6512);
nand U11635 (N_11635,N_5808,N_5581);
or U11636 (N_11636,N_6278,N_5212);
nand U11637 (N_11637,N_9270,N_7202);
nor U11638 (N_11638,N_8216,N_8770);
xor U11639 (N_11639,N_9065,N_5060);
xor U11640 (N_11640,N_7349,N_8448);
nor U11641 (N_11641,N_7315,N_9301);
or U11642 (N_11642,N_9974,N_9122);
nand U11643 (N_11643,N_9310,N_9101);
xnor U11644 (N_11644,N_5059,N_9004);
nor U11645 (N_11645,N_9158,N_9450);
nand U11646 (N_11646,N_8970,N_7625);
or U11647 (N_11647,N_8099,N_5213);
nand U11648 (N_11648,N_6774,N_9911);
nor U11649 (N_11649,N_7674,N_8512);
or U11650 (N_11650,N_8347,N_8966);
nor U11651 (N_11651,N_9645,N_8554);
xnor U11652 (N_11652,N_8995,N_7533);
or U11653 (N_11653,N_8152,N_8785);
nand U11654 (N_11654,N_6133,N_5927);
and U11655 (N_11655,N_7963,N_9498);
and U11656 (N_11656,N_8479,N_5680);
or U11657 (N_11657,N_5799,N_8925);
or U11658 (N_11658,N_9897,N_7650);
nand U11659 (N_11659,N_8636,N_8789);
nand U11660 (N_11660,N_9177,N_6738);
or U11661 (N_11661,N_9749,N_6827);
nor U11662 (N_11662,N_6770,N_6529);
nor U11663 (N_11663,N_6144,N_6471);
and U11664 (N_11664,N_5904,N_9924);
nor U11665 (N_11665,N_7835,N_9418);
or U11666 (N_11666,N_5938,N_6519);
xnor U11667 (N_11667,N_9506,N_6843);
xnor U11668 (N_11668,N_7978,N_8541);
nand U11669 (N_11669,N_6219,N_5479);
xnor U11670 (N_11670,N_6229,N_7305);
and U11671 (N_11671,N_6862,N_8329);
and U11672 (N_11672,N_7029,N_5685);
nor U11673 (N_11673,N_6465,N_7265);
or U11674 (N_11674,N_9515,N_7399);
or U11675 (N_11675,N_9578,N_5690);
or U11676 (N_11676,N_5045,N_5339);
nor U11677 (N_11677,N_7735,N_9119);
and U11678 (N_11678,N_6725,N_6018);
and U11679 (N_11679,N_9086,N_9802);
and U11680 (N_11680,N_5794,N_8902);
nor U11681 (N_11681,N_9881,N_9529);
and U11682 (N_11682,N_8600,N_9856);
and U11683 (N_11683,N_8632,N_9150);
nor U11684 (N_11684,N_8357,N_6760);
nor U11685 (N_11685,N_9411,N_7206);
or U11686 (N_11686,N_8737,N_7209);
or U11687 (N_11687,N_9782,N_8355);
xnor U11688 (N_11688,N_9803,N_5989);
or U11689 (N_11689,N_9649,N_6054);
xor U11690 (N_11690,N_6551,N_9581);
xor U11691 (N_11691,N_9214,N_5463);
and U11692 (N_11692,N_8268,N_5185);
nand U11693 (N_11693,N_8100,N_8017);
xnor U11694 (N_11694,N_8729,N_8128);
nand U11695 (N_11695,N_6610,N_5098);
xor U11696 (N_11696,N_9269,N_7751);
nand U11697 (N_11697,N_9200,N_5656);
nand U11698 (N_11698,N_7024,N_9352);
nand U11699 (N_11699,N_9996,N_8784);
nor U11700 (N_11700,N_5665,N_8030);
and U11701 (N_11701,N_6901,N_8782);
nor U11702 (N_11702,N_6393,N_7372);
or U11703 (N_11703,N_5678,N_5511);
or U11704 (N_11704,N_9181,N_7613);
nor U11705 (N_11705,N_5398,N_9216);
xnor U11706 (N_11706,N_7896,N_7628);
nor U11707 (N_11707,N_9861,N_6221);
and U11708 (N_11708,N_5086,N_5377);
and U11709 (N_11709,N_7194,N_9128);
nor U11710 (N_11710,N_6686,N_6990);
and U11711 (N_11711,N_5958,N_9383);
nor U11712 (N_11712,N_6704,N_6179);
or U11713 (N_11713,N_5924,N_5043);
and U11714 (N_11714,N_7690,N_6315);
xor U11715 (N_11715,N_5044,N_9417);
nand U11716 (N_11716,N_5523,N_8127);
nor U11717 (N_11717,N_7385,N_7008);
or U11718 (N_11718,N_9160,N_8462);
or U11719 (N_11719,N_8960,N_8452);
nor U11720 (N_11720,N_7076,N_6163);
nor U11721 (N_11721,N_5290,N_5282);
nor U11722 (N_11722,N_6651,N_6642);
nor U11723 (N_11723,N_6662,N_5625);
and U11724 (N_11724,N_6003,N_5940);
nor U11725 (N_11725,N_8935,N_8316);
nand U11726 (N_11726,N_8825,N_6730);
or U11727 (N_11727,N_9977,N_5441);
and U11728 (N_11728,N_7633,N_9147);
xnor U11729 (N_11729,N_5211,N_7154);
nor U11730 (N_11730,N_7201,N_5246);
and U11731 (N_11731,N_6521,N_5054);
nand U11732 (N_11732,N_7773,N_7691);
xnor U11733 (N_11733,N_9115,N_9490);
nor U11734 (N_11734,N_7496,N_8556);
nor U11735 (N_11735,N_7614,N_6235);
nor U11736 (N_11736,N_6034,N_5368);
nand U11737 (N_11737,N_8626,N_8334);
or U11738 (N_11738,N_5561,N_7948);
nand U11739 (N_11739,N_9604,N_9926);
xnor U11740 (N_11740,N_5679,N_7940);
nand U11741 (N_11741,N_5825,N_5604);
xnor U11742 (N_11742,N_9218,N_6178);
and U11743 (N_11743,N_9442,N_5137);
nor U11744 (N_11744,N_6299,N_6246);
and U11745 (N_11745,N_8589,N_6171);
and U11746 (N_11746,N_5066,N_6647);
xor U11747 (N_11747,N_9693,N_5312);
or U11748 (N_11748,N_6824,N_6295);
nor U11749 (N_11749,N_5518,N_7475);
or U11750 (N_11750,N_5036,N_5805);
and U11751 (N_11751,N_6442,N_5652);
nand U11752 (N_11752,N_5586,N_6236);
nand U11753 (N_11753,N_8530,N_6286);
nor U11754 (N_11754,N_5733,N_5308);
or U11755 (N_11755,N_9954,N_7018);
and U11756 (N_11756,N_9186,N_9053);
or U11757 (N_11757,N_7052,N_7810);
and U11758 (N_11758,N_8603,N_6205);
and U11759 (N_11759,N_7438,N_9769);
xor U11760 (N_11760,N_7777,N_8396);
nor U11761 (N_11761,N_5736,N_6814);
nor U11762 (N_11762,N_7364,N_7445);
or U11763 (N_11763,N_6320,N_8832);
or U11764 (N_11764,N_8182,N_6053);
nor U11765 (N_11765,N_8538,N_6716);
and U11766 (N_11766,N_5498,N_9121);
nor U11767 (N_11767,N_6514,N_7705);
or U11768 (N_11768,N_7091,N_7458);
and U11769 (N_11769,N_6527,N_5532);
nand U11770 (N_11770,N_5772,N_9546);
xor U11771 (N_11771,N_7095,N_8640);
and U11772 (N_11772,N_8684,N_5822);
nor U11773 (N_11773,N_8047,N_7157);
and U11774 (N_11774,N_6238,N_6123);
xor U11775 (N_11775,N_6657,N_8336);
and U11776 (N_11776,N_6942,N_9088);
xnor U11777 (N_11777,N_6938,N_6481);
or U11778 (N_11778,N_7680,N_8808);
or U11779 (N_11779,N_5640,N_7258);
or U11780 (N_11780,N_7779,N_6759);
or U11781 (N_11781,N_8573,N_5556);
nor U11782 (N_11782,N_6197,N_7383);
nand U11783 (N_11783,N_7911,N_7607);
xnor U11784 (N_11784,N_7304,N_9940);
or U11785 (N_11785,N_8504,N_9701);
or U11786 (N_11786,N_7860,N_7185);
nand U11787 (N_11787,N_8394,N_7610);
xnor U11788 (N_11788,N_5770,N_9380);
and U11789 (N_11789,N_7775,N_8658);
xor U11790 (N_11790,N_6407,N_7541);
or U11791 (N_11791,N_9304,N_6094);
nor U11792 (N_11792,N_5110,N_8193);
or U11793 (N_11793,N_8145,N_7233);
and U11794 (N_11794,N_6228,N_7945);
nor U11795 (N_11795,N_7289,N_7546);
nor U11796 (N_11796,N_5639,N_9742);
or U11797 (N_11797,N_8583,N_8280);
xor U11798 (N_11798,N_8930,N_9850);
and U11799 (N_11799,N_5682,N_5210);
xor U11800 (N_11800,N_9205,N_5663);
xnor U11801 (N_11801,N_5438,N_7545);
nor U11802 (N_11802,N_6965,N_6426);
or U11803 (N_11803,N_6858,N_5488);
nand U11804 (N_11804,N_9385,N_7145);
or U11805 (N_11805,N_6534,N_9327);
xor U11806 (N_11806,N_7757,N_8522);
and U11807 (N_11807,N_9103,N_8876);
or U11808 (N_11808,N_8176,N_8761);
nor U11809 (N_11809,N_9877,N_6353);
nor U11810 (N_11810,N_8718,N_5845);
nor U11811 (N_11811,N_5168,N_6568);
xnor U11812 (N_11812,N_8797,N_8340);
nand U11813 (N_11813,N_5289,N_6621);
nor U11814 (N_11814,N_9651,N_9331);
and U11815 (N_11815,N_7991,N_8787);
nor U11816 (N_11816,N_7015,N_6688);
and U11817 (N_11817,N_8588,N_7003);
nand U11818 (N_11818,N_8678,N_8517);
nor U11819 (N_11819,N_9118,N_7807);
or U11820 (N_11820,N_7704,N_8113);
nand U11821 (N_11821,N_6558,N_7522);
nand U11822 (N_11822,N_8195,N_5268);
nor U11823 (N_11823,N_8330,N_5998);
or U11824 (N_11824,N_8713,N_8568);
and U11825 (N_11825,N_5328,N_9549);
or U11826 (N_11826,N_8918,N_6099);
and U11827 (N_11827,N_6523,N_9923);
nand U11828 (N_11828,N_6816,N_5594);
or U11829 (N_11829,N_8188,N_9329);
or U11830 (N_11830,N_7051,N_6756);
nor U11831 (N_11831,N_7665,N_5288);
xor U11832 (N_11832,N_5547,N_7328);
and U11833 (N_11833,N_7869,N_8774);
xor U11834 (N_11834,N_7022,N_8398);
xnor U11835 (N_11835,N_7510,N_5892);
nor U11836 (N_11836,N_7580,N_8317);
and U11837 (N_11837,N_5959,N_7405);
or U11838 (N_11838,N_9208,N_9000);
xnor U11839 (N_11839,N_5359,N_8456);
or U11840 (N_11840,N_5610,N_6548);
and U11841 (N_11841,N_8714,N_5323);
nand U11842 (N_11842,N_5565,N_5961);
nand U11843 (N_11843,N_8476,N_7253);
nor U11844 (N_11844,N_9489,N_9291);
and U11845 (N_11845,N_5173,N_7516);
nand U11846 (N_11846,N_9611,N_7662);
nor U11847 (N_11847,N_5280,N_5461);
or U11848 (N_11848,N_5449,N_7100);
nand U11849 (N_11849,N_5920,N_7362);
nor U11850 (N_11850,N_8595,N_8060);
or U11851 (N_11851,N_7748,N_9555);
and U11852 (N_11852,N_5147,N_7214);
or U11853 (N_11853,N_6969,N_7094);
xor U11854 (N_11854,N_7626,N_6479);
nand U11855 (N_11855,N_9699,N_9532);
xor U11856 (N_11856,N_9311,N_5309);
xor U11857 (N_11857,N_8395,N_7124);
xor U11858 (N_11858,N_5919,N_9106);
xor U11859 (N_11859,N_8281,N_7509);
xor U11860 (N_11860,N_9821,N_7841);
or U11861 (N_11861,N_7787,N_9454);
or U11862 (N_11862,N_8203,N_8880);
xnor U11863 (N_11863,N_6878,N_6522);
xor U11864 (N_11864,N_9094,N_6552);
xor U11865 (N_11865,N_9326,N_6964);
nand U11866 (N_11866,N_6914,N_5582);
nand U11867 (N_11867,N_5758,N_5329);
nand U11868 (N_11868,N_6082,N_9635);
and U11869 (N_11869,N_5369,N_8241);
nor U11870 (N_11870,N_7931,N_7920);
or U11871 (N_11871,N_8151,N_9077);
or U11872 (N_11872,N_9169,N_5600);
nor U11873 (N_11873,N_5615,N_5253);
nor U11874 (N_11874,N_5571,N_9394);
or U11875 (N_11875,N_5149,N_6808);
nand U11876 (N_11876,N_9502,N_9123);
or U11877 (N_11877,N_6333,N_5637);
and U11878 (N_11878,N_9563,N_9873);
xnor U11879 (N_11879,N_5008,N_9167);
nor U11880 (N_11880,N_9691,N_7128);
nand U11881 (N_11881,N_5801,N_5327);
nor U11882 (N_11882,N_7734,N_6271);
nor U11883 (N_11883,N_5191,N_8875);
or U11884 (N_11884,N_8083,N_6518);
or U11885 (N_11885,N_5861,N_5161);
or U11886 (N_11886,N_8756,N_6654);
or U11887 (N_11887,N_8458,N_5667);
or U11888 (N_11888,N_5143,N_8267);
xnor U11889 (N_11889,N_6242,N_6060);
nor U11890 (N_11890,N_9992,N_7256);
nor U11891 (N_11891,N_5216,N_5153);
and U11892 (N_11892,N_9255,N_9629);
xnor U11893 (N_11893,N_8830,N_6912);
nor U11894 (N_11894,N_8892,N_5869);
nand U11895 (N_11895,N_7410,N_7493);
nand U11896 (N_11896,N_6991,N_8986);
xnor U11897 (N_11897,N_9824,N_5631);
nor U11898 (N_11898,N_8408,N_8276);
nor U11899 (N_11899,N_8890,N_7165);
nand U11900 (N_11900,N_6382,N_9351);
nor U11901 (N_11901,N_8489,N_6764);
nand U11902 (N_11902,N_6502,N_8118);
xnor U11903 (N_11903,N_8043,N_5485);
nand U11904 (N_11904,N_9746,N_6988);
nor U11905 (N_11905,N_7582,N_9662);
and U11906 (N_11906,N_8557,N_7412);
nand U11907 (N_11907,N_8414,N_6694);
nand U11908 (N_11908,N_7228,N_8157);
nand U11909 (N_11909,N_9511,N_6195);
or U11910 (N_11910,N_7158,N_7957);
xnor U11911 (N_11911,N_6381,N_9910);
and U11912 (N_11912,N_8520,N_8940);
xnor U11913 (N_11913,N_5245,N_9858);
nand U11914 (N_11914,N_6611,N_5732);
xnor U11915 (N_11915,N_5768,N_6681);
xnor U11916 (N_11916,N_7550,N_6324);
and U11917 (N_11917,N_5199,N_8531);
nand U11918 (N_11918,N_5371,N_8065);
and U11919 (N_11919,N_8799,N_7946);
and U11920 (N_11920,N_6757,N_8838);
or U11921 (N_11921,N_9864,N_7271);
nor U11922 (N_11922,N_9033,N_5358);
and U11923 (N_11923,N_5981,N_9957);
and U11924 (N_11924,N_6855,N_9567);
xnor U11925 (N_11925,N_8064,N_8342);
nand U11926 (N_11926,N_9830,N_8570);
and U11927 (N_11927,N_6307,N_7749);
or U11928 (N_11928,N_7565,N_7042);
and U11929 (N_11929,N_9280,N_6146);
and U11930 (N_11930,N_5932,N_9287);
and U11931 (N_11931,N_9298,N_7135);
and U11932 (N_11932,N_6817,N_9052);
or U11933 (N_11933,N_5408,N_7113);
or U11934 (N_11934,N_8343,N_7781);
and U11935 (N_11935,N_8228,N_7274);
or U11936 (N_11936,N_8850,N_9283);
xor U11937 (N_11937,N_7771,N_8549);
xor U11938 (N_11938,N_9758,N_6543);
xnor U11939 (N_11939,N_5543,N_8501);
nor U11940 (N_11940,N_7553,N_5266);
nand U11941 (N_11941,N_5120,N_8742);
nor U11942 (N_11942,N_5183,N_5913);
nand U11943 (N_11943,N_8920,N_7361);
nor U11944 (N_11944,N_8883,N_9950);
and U11945 (N_11945,N_8420,N_6626);
xor U11946 (N_11946,N_7995,N_6314);
or U11947 (N_11947,N_6630,N_9919);
or U11948 (N_11948,N_6592,N_7792);
nand U11949 (N_11949,N_6793,N_9433);
nor U11950 (N_11950,N_7040,N_7494);
xnor U11951 (N_11951,N_9483,N_9307);
nor U11952 (N_11952,N_7267,N_5896);
nor U11953 (N_11953,N_7467,N_5764);
nand U11954 (N_11954,N_8628,N_8164);
nor U11955 (N_11955,N_9142,N_7836);
or U11956 (N_11956,N_6832,N_6004);
or U11957 (N_11957,N_6836,N_6805);
and U11958 (N_11958,N_7404,N_9987);
nand U11959 (N_11959,N_7211,N_9835);
nand U11960 (N_11960,N_9305,N_7056);
xor U11961 (N_11961,N_5433,N_7358);
or U11962 (N_11962,N_7231,N_7694);
nor U11963 (N_11963,N_8945,N_8521);
or U11964 (N_11964,N_7518,N_7400);
or U11965 (N_11965,N_8110,N_8415);
nor U11966 (N_11966,N_8013,N_9654);
nor U11967 (N_11967,N_7079,N_9753);
nand U11968 (N_11968,N_7105,N_8015);
nor U11969 (N_11969,N_8416,N_9098);
xor U11970 (N_11970,N_5788,N_8386);
and U11971 (N_11971,N_7293,N_8437);
nand U11972 (N_11972,N_5072,N_5203);
nand U11973 (N_11973,N_5420,N_8819);
xnor U11974 (N_11974,N_9900,N_5163);
nand U11975 (N_11975,N_7954,N_8682);
nor U11976 (N_11976,N_8323,N_9314);
nor U11977 (N_11977,N_7593,N_6872);
nor U11978 (N_11978,N_5067,N_9801);
nor U11979 (N_11979,N_6036,N_9752);
or U11980 (N_11980,N_5267,N_8717);
or U11981 (N_11981,N_9073,N_6113);
and U11982 (N_11982,N_8067,N_7302);
and U11983 (N_11983,N_8978,N_8220);
nor U11984 (N_11984,N_8377,N_5910);
and U11985 (N_11985,N_9090,N_8413);
or U11986 (N_11986,N_5258,N_6375);
nand U11987 (N_11987,N_8175,N_5411);
or U11988 (N_11988,N_8320,N_5684);
nand U11989 (N_11989,N_6775,N_8358);
and U11990 (N_11990,N_6584,N_7232);
or U11991 (N_11991,N_7700,N_7120);
and U11992 (N_11992,N_9199,N_8366);
nand U11993 (N_11993,N_8676,N_7791);
nor U11994 (N_11994,N_8262,N_9247);
and U11995 (N_11995,N_5689,N_6601);
or U11996 (N_11996,N_5084,N_5002);
nand U11997 (N_11997,N_6313,N_9561);
xnor U11998 (N_11998,N_9624,N_9639);
nor U11999 (N_11999,N_8299,N_5412);
or U12000 (N_12000,N_5978,N_5803);
and U12001 (N_12001,N_8496,N_6347);
nand U12002 (N_12002,N_6895,N_8049);
nor U12003 (N_12003,N_9582,N_6899);
and U12004 (N_12004,N_6538,N_7794);
xnor U12005 (N_12005,N_7985,N_6882);
xnor U12006 (N_12006,N_9002,N_6296);
nor U12007 (N_12007,N_8745,N_9231);
and U12008 (N_12008,N_8277,N_6429);
nand U12009 (N_12009,N_6924,N_7490);
nor U12010 (N_12010,N_6695,N_9809);
xor U12011 (N_12011,N_7702,N_8434);
nor U12012 (N_12012,N_7619,N_5930);
or U12013 (N_12013,N_9937,N_7153);
or U12014 (N_12014,N_8980,N_6419);
xnor U12015 (N_12015,N_7485,N_7884);
nand U12016 (N_12016,N_8021,N_9672);
or U12017 (N_12017,N_9359,N_7826);
nor U12018 (N_12018,N_9175,N_6447);
or U12019 (N_12019,N_7440,N_6364);
xnor U12020 (N_12020,N_6915,N_6243);
or U12021 (N_12021,N_7947,N_7672);
nand U12022 (N_12022,N_7965,N_5390);
nor U12023 (N_12023,N_6152,N_6615);
and U12024 (N_12024,N_9713,N_7718);
xor U12025 (N_12025,N_9539,N_5612);
nor U12026 (N_12026,N_5688,N_5675);
or U12027 (N_12027,N_9260,N_7325);
or U12028 (N_12028,N_6889,N_6701);
xnor U12029 (N_12029,N_6898,N_9039);
or U12030 (N_12030,N_6589,N_9571);
nand U12031 (N_12031,N_5428,N_5080);
nor U12032 (N_12032,N_8050,N_7786);
nor U12033 (N_12033,N_5671,N_8040);
or U12034 (N_12034,N_6136,N_5588);
nand U12035 (N_12035,N_5158,N_7909);
nand U12036 (N_12036,N_5784,N_6039);
xnor U12037 (N_12037,N_5922,N_7376);
or U12038 (N_12038,N_5851,N_6906);
nor U12039 (N_12039,N_5626,N_9317);
xor U12040 (N_12040,N_7353,N_5514);
or U12041 (N_12041,N_9918,N_5852);
or U12042 (N_12042,N_6436,N_5109);
or U12043 (N_12043,N_8870,N_6825);
nor U12044 (N_12044,N_9786,N_8928);
nor U12045 (N_12045,N_9847,N_6643);
xnor U12046 (N_12046,N_7121,N_6828);
nand U12047 (N_12047,N_5260,N_9171);
nand U12048 (N_12048,N_8775,N_5776);
nor U12049 (N_12049,N_8859,N_5015);
nand U12050 (N_12050,N_6579,N_7101);
nand U12051 (N_12051,N_8350,N_9723);
nor U12052 (N_12052,N_9091,N_5584);
nand U12053 (N_12053,N_5941,N_9295);
nand U12054 (N_12054,N_5884,N_6856);
and U12055 (N_12055,N_6768,N_8765);
nor U12056 (N_12056,N_5702,N_8601);
and U12057 (N_12057,N_9586,N_5040);
nor U12058 (N_12058,N_7561,N_5247);
xor U12059 (N_12059,N_6116,N_6989);
nor U12060 (N_12060,N_5737,N_8715);
nand U12061 (N_12061,N_6731,N_8899);
nor U12062 (N_12062,N_7355,N_6624);
xor U12063 (N_12063,N_8551,N_5476);
or U12064 (N_12064,N_9234,N_6923);
xor U12065 (N_12065,N_6665,N_5112);
nand U12066 (N_12066,N_7972,N_8236);
or U12067 (N_12067,N_6941,N_5012);
xor U12068 (N_12068,N_9589,N_7637);
nor U12069 (N_12069,N_5455,N_6093);
and U12070 (N_12070,N_6154,N_9705);
xor U12071 (N_12071,N_8798,N_8644);
and U12072 (N_12072,N_5598,N_6475);
and U12073 (N_12073,N_9276,N_6169);
nor U12074 (N_12074,N_5090,N_9934);
and U12075 (N_12075,N_5781,N_5809);
and U12076 (N_12076,N_7212,N_8284);
and U12077 (N_12077,N_5949,N_6903);
and U12078 (N_12078,N_9678,N_5815);
or U12079 (N_12079,N_8417,N_5575);
xnor U12080 (N_12080,N_6675,N_8695);
and U12081 (N_12081,N_6715,N_8424);
xor U12082 (N_12082,N_7007,N_8777);
and U12083 (N_12083,N_6506,N_8475);
and U12084 (N_12084,N_8092,N_9330);
xnor U12085 (N_12085,N_5760,N_5240);
or U12086 (N_12086,N_6995,N_6308);
and U12087 (N_12087,N_7758,N_8942);
or U12088 (N_12088,N_6837,N_5999);
nand U12089 (N_12089,N_5769,N_9379);
or U12090 (N_12090,N_9643,N_8063);
xor U12091 (N_12091,N_8908,N_5102);
nand U12092 (N_12092,N_5548,N_6183);
nand U12093 (N_12093,N_7643,N_5042);
nor U12094 (N_12094,N_8075,N_8529);
nand U12095 (N_12095,N_5076,N_6037);
and U12096 (N_12096,N_7571,N_8623);
nand U12097 (N_12097,N_6854,N_6950);
and U12098 (N_12098,N_8483,N_8312);
nand U12099 (N_12099,N_5839,N_9034);
xnor U12100 (N_12100,N_8901,N_8084);
nand U12101 (N_12101,N_7351,N_8561);
xor U12102 (N_12102,N_6902,N_6260);
xnor U12103 (N_12103,N_7975,N_9057);
nand U12104 (N_12104,N_7208,N_5531);
xor U12105 (N_12105,N_5344,N_8752);
and U12106 (N_12106,N_6966,N_6259);
or U12107 (N_12107,N_7706,N_7724);
and U12108 (N_12108,N_7688,N_9837);
nand U12109 (N_12109,N_9943,N_7843);
nand U12110 (N_12110,N_5401,N_9891);
or U12111 (N_12111,N_9983,N_6087);
nor U12112 (N_12112,N_9566,N_9606);
nor U12113 (N_12113,N_7714,N_5348);
or U12114 (N_12114,N_6306,N_8375);
or U12115 (N_12115,N_7618,N_8811);
and U12116 (N_12116,N_6765,N_9465);
nand U12117 (N_12117,N_9376,N_5826);
nand U12118 (N_12118,N_9481,N_9238);
or U12119 (N_12119,N_9130,N_9817);
nor U12120 (N_12120,N_5340,N_9558);
and U12121 (N_12121,N_5856,N_6753);
nand U12122 (N_12122,N_5491,N_6919);
nor U12123 (N_12123,N_5385,N_8190);
xor U12124 (N_12124,N_5028,N_8428);
nor U12125 (N_12125,N_6932,N_8385);
or U12126 (N_12126,N_9893,N_5889);
nand U12127 (N_12127,N_7962,N_5027);
nor U12128 (N_12128,N_6917,N_6718);
or U12129 (N_12129,N_7413,N_7746);
nor U12130 (N_12130,N_9844,N_7436);
xor U12131 (N_12131,N_6948,N_7075);
and U12132 (N_12132,N_8439,N_5380);
nor U12133 (N_12133,N_6801,N_8012);
nor U12134 (N_12134,N_9663,N_9145);
nand U12135 (N_12135,N_6389,N_7017);
or U12136 (N_12136,N_8247,N_6554);
or U12137 (N_12137,N_6083,N_8349);
and U12138 (N_12138,N_9706,N_9725);
and U12139 (N_12139,N_8612,N_7393);
nand U12140 (N_12140,N_6261,N_9188);
nand U12141 (N_12141,N_5517,N_7021);
nand U12142 (N_12142,N_6790,N_8552);
nor U12143 (N_12143,N_7600,N_7210);
xnor U12144 (N_12144,N_6180,N_5083);
xnor U12145 (N_12145,N_9732,N_7872);
or U12146 (N_12146,N_5954,N_5996);
nor U12147 (N_12147,N_8810,N_9191);
or U12148 (N_12148,N_7760,N_7298);
nand U12149 (N_12149,N_6879,N_6240);
or U12150 (N_12150,N_6377,N_8166);
nor U12151 (N_12151,N_9484,N_7435);
xor U12152 (N_12152,N_5142,N_8042);
or U12153 (N_12153,N_8653,N_5241);
xor U12154 (N_12154,N_8962,N_9328);
and U12155 (N_12155,N_8625,N_6107);
nor U12156 (N_12156,N_5179,N_9852);
and U12157 (N_12157,N_5873,N_5111);
and U12158 (N_12158,N_6371,N_5224);
or U12159 (N_12159,N_7959,N_5730);
nand U12160 (N_12160,N_7488,N_5567);
or U12161 (N_12161,N_8070,N_6035);
nand U12162 (N_12162,N_8856,N_5538);
xor U12163 (N_12163,N_6550,N_6772);
nor U12164 (N_12164,N_5672,N_6204);
xnor U12165 (N_12165,N_7657,N_6398);
or U12166 (N_12166,N_5552,N_6394);
nand U12167 (N_12167,N_6114,N_5135);
xnor U12168 (N_12168,N_9684,N_8647);
and U12169 (N_12169,N_6524,N_9068);
nand U12170 (N_12170,N_9133,N_8133);
or U12171 (N_12171,N_8360,N_6239);
nand U12172 (N_12172,N_8707,N_9007);
xnor U12173 (N_12173,N_8077,N_7864);
xnor U12174 (N_12174,N_6059,N_6750);
xnor U12175 (N_12175,N_9717,N_6563);
nand U12176 (N_12176,N_9823,N_9832);
and U12177 (N_12177,N_5486,N_6866);
or U12178 (N_12178,N_8900,N_7517);
and U12179 (N_12179,N_7685,N_8105);
nand U12180 (N_12180,N_5880,N_6380);
or U12181 (N_12181,N_5724,N_7859);
and U12182 (N_12182,N_9920,N_5322);
and U12183 (N_12183,N_7414,N_7870);
nand U12184 (N_12184,N_8088,N_9781);
nand U12185 (N_12185,N_7663,N_8227);
and U12186 (N_12186,N_8095,N_8988);
or U12187 (N_12187,N_9530,N_7499);
xnor U12188 (N_12188,N_9590,N_9364);
or U12189 (N_12189,N_5668,N_9095);
nand U12190 (N_12190,N_9703,N_7426);
nor U12191 (N_12191,N_8906,N_5232);
nor U12192 (N_12192,N_8548,N_7918);
or U12193 (N_12193,N_7970,N_9252);
or U12194 (N_12194,N_7495,N_6092);
nor U12195 (N_12195,N_6128,N_8665);
or U12196 (N_12196,N_8915,N_8687);
or U12197 (N_12197,N_6499,N_8793);
or U12198 (N_12198,N_7844,N_9550);
nor U12199 (N_12199,N_7336,N_9224);
or U12200 (N_12200,N_5248,N_6921);
nor U12201 (N_12201,N_5597,N_9666);
nand U12202 (N_12202,N_7407,N_9136);
xnor U12203 (N_12203,N_6276,N_5670);
xnor U12204 (N_12204,N_9070,N_7132);
nand U12205 (N_12205,N_5397,N_5614);
nor U12206 (N_12206,N_5562,N_5783);
or U12207 (N_12207,N_8245,N_6431);
or U12208 (N_12208,N_7155,N_9032);
or U12209 (N_12209,N_9390,N_7442);
xor U12210 (N_12210,N_7744,N_6453);
nand U12211 (N_12211,N_8074,N_8981);
nand U12212 (N_12212,N_6664,N_9982);
and U12213 (N_12213,N_8747,N_7434);
or U12214 (N_12214,N_9014,N_6142);
nand U12215 (N_12215,N_9107,N_7366);
and U12216 (N_12216,N_6269,N_7109);
or U12217 (N_12217,N_9036,N_5471);
or U12218 (N_12218,N_8743,N_5035);
nand U12219 (N_12219,N_6692,N_7941);
xor U12220 (N_12220,N_9949,N_5895);
and U12221 (N_12221,N_9426,N_7612);
nor U12222 (N_12222,N_6316,N_8760);
xor U12223 (N_12223,N_9156,N_9078);
xnor U12224 (N_12224,N_8463,N_6486);
nand U12225 (N_12225,N_6255,N_7243);
xor U12226 (N_12226,N_9750,N_5074);
or U12227 (N_12227,N_8829,N_8749);
xnor U12228 (N_12228,N_6030,N_6319);
nand U12229 (N_12229,N_7238,N_7140);
nand U12230 (N_12230,N_5154,N_9229);
nor U12231 (N_12231,N_5744,N_9863);
nor U12232 (N_12232,N_5926,N_5599);
or U12233 (N_12233,N_5037,N_8696);
nand U12234 (N_12234,N_8540,N_5674);
nand U12235 (N_12235,N_5421,N_5310);
and U12236 (N_12236,N_8939,N_5774);
nand U12237 (N_12237,N_9757,N_8973);
and U12238 (N_12238,N_9341,N_9771);
nor U12239 (N_12239,N_8748,N_5123);
nor U12240 (N_12240,N_8639,N_8591);
and U12241 (N_12241,N_8993,N_8814);
nand U12242 (N_12242,N_8565,N_5472);
nand U12243 (N_12243,N_8457,N_5714);
nand U12244 (N_12244,N_9831,N_6949);
nor U12245 (N_12245,N_9176,N_7573);
or U12246 (N_12246,N_9323,N_7259);
nand U12247 (N_12247,N_7687,N_5568);
nor U12248 (N_12248,N_7226,N_5252);
xnor U12249 (N_12249,N_8621,N_9690);
xor U12250 (N_12250,N_8710,N_5661);
nand U12251 (N_12251,N_7028,N_8686);
xnor U12252 (N_12252,N_5030,N_5021);
nor U12253 (N_12253,N_9698,N_6346);
xor U12254 (N_12254,N_7019,N_7635);
and U12255 (N_12255,N_7766,N_5883);
nor U12256 (N_12256,N_8823,N_9585);
nor U12257 (N_12257,N_5504,N_6343);
and U12258 (N_12258,N_9278,N_8274);
xor U12259 (N_12259,N_5293,N_6211);
xor U12260 (N_12260,N_7525,N_5681);
nor U12261 (N_12261,N_7139,N_8404);
and U12262 (N_12262,N_9636,N_7294);
nand U12263 (N_12263,N_9338,N_5929);
nor U12264 (N_12264,N_6177,N_5402);
xor U12265 (N_12265,N_7450,N_9458);
xor U12266 (N_12266,N_7576,N_5145);
nand U12267 (N_12267,N_7449,N_7755);
or U12268 (N_12268,N_8239,N_7195);
or U12269 (N_12269,N_9978,N_9275);
nor U12270 (N_12270,N_6190,N_9715);
xnor U12271 (N_12271,N_9673,N_6953);
xor U12272 (N_12272,N_9139,N_6976);
and U12273 (N_12273,N_9354,N_7876);
or U12274 (N_12274,N_9641,N_9460);
xnor U12275 (N_12275,N_9991,N_7641);
nand U12276 (N_12276,N_9277,N_5100);
or U12277 (N_12277,N_6987,N_7707);
nand U12278 (N_12278,N_7555,N_9780);
or U12279 (N_12279,N_6337,N_7130);
and U12280 (N_12280,N_9384,N_8884);
and U12281 (N_12281,N_8721,N_9047);
or U12282 (N_12282,N_5576,N_6637);
and U12283 (N_12283,N_7005,N_7804);
or U12284 (N_12284,N_6720,N_7334);
nand U12285 (N_12285,N_5492,N_5738);
nand U12286 (N_12286,N_5276,N_9734);
or U12287 (N_12287,N_6810,N_8662);
nor U12288 (N_12288,N_8009,N_9129);
nand U12289 (N_12289,N_5431,N_6913);
nor U12290 (N_12290,N_9686,N_9482);
and U12291 (N_12291,N_6340,N_7592);
nor U12292 (N_12292,N_8764,N_7747);
or U12293 (N_12293,N_9976,N_5489);
nor U12294 (N_12294,N_9134,N_7581);
nor U12295 (N_12295,N_6909,N_9038);
and U12296 (N_12296,N_8313,N_5077);
and U12297 (N_12297,N_8441,N_9045);
nand U12298 (N_12298,N_6138,N_5642);
nor U12299 (N_12299,N_7992,N_6955);
nand U12300 (N_12300,N_6126,N_5630);
nor U12301 (N_12301,N_6367,N_8675);
or U12302 (N_12302,N_5301,N_8315);
and U12303 (N_12303,N_5650,N_5507);
or U12304 (N_12304,N_9387,N_8150);
xnor U12305 (N_12305,N_6430,N_8680);
and U12306 (N_12306,N_7615,N_5676);
or U12307 (N_12307,N_9444,N_9299);
nand U12308 (N_12308,N_9420,N_9035);
nand U12309 (N_12309,N_9761,N_7333);
or U12310 (N_12310,N_6362,N_8477);
nor U12311 (N_12311,N_9120,N_7439);
or U12312 (N_12312,N_5577,N_9108);
xnor U12313 (N_12313,N_5855,N_5101);
and U12314 (N_12314,N_9692,N_8326);
or U12315 (N_12315,N_7783,N_6982);
nand U12316 (N_12316,N_6289,N_6031);
xor U12317 (N_12317,N_7377,N_5660);
xnor U12318 (N_12318,N_9445,N_8418);
nor U12319 (N_12319,N_6461,N_9369);
nand U12320 (N_12320,N_5196,N_7689);
nor U12321 (N_12321,N_5513,N_9062);
nand U12322 (N_12322,N_8002,N_8778);
or U12323 (N_12323,N_8652,N_5829);
or U12324 (N_12324,N_8367,N_6454);
and U12325 (N_12325,N_7813,N_5284);
xnor U12326 (N_12326,N_8791,N_7136);
xnor U12327 (N_12327,N_6057,N_9373);
xnor U12328 (N_12328,N_9242,N_9929);
nor U12329 (N_12329,N_7323,N_5870);
nor U12330 (N_12330,N_7147,N_5250);
xor U12331 (N_12331,N_8982,N_5055);
nand U12332 (N_12332,N_7897,N_6585);
and U12333 (N_12333,N_5334,N_9398);
or U12334 (N_12334,N_9399,N_6599);
and U12335 (N_12335,N_6440,N_6670);
nand U12336 (N_12336,N_9795,N_5200);
nand U12337 (N_12337,N_9970,N_6108);
and U12338 (N_12338,N_5911,N_7409);
or U12339 (N_12339,N_7753,N_8581);
or U12340 (N_12340,N_9074,N_9637);
or U12341 (N_12341,N_7382,N_5830);
nor U12342 (N_12342,N_6644,N_6069);
nand U12343 (N_12343,N_8910,N_9212);
nor U12344 (N_12344,N_7611,N_6052);
xnor U12345 (N_12345,N_5351,N_8346);
nand U12346 (N_12346,N_8701,N_6871);
xnor U12347 (N_12347,N_9839,N_6733);
or U12348 (N_12348,N_6762,N_9848);
xor U12349 (N_12349,N_7890,N_8146);
or U12350 (N_12350,N_9759,N_9041);
xnor U12351 (N_12351,N_5372,N_5400);
nor U12352 (N_12352,N_7661,N_7181);
or U12353 (N_12353,N_5207,N_5643);
nand U12354 (N_12354,N_5587,N_8897);
nand U12355 (N_12355,N_9547,N_9207);
or U12356 (N_12356,N_9367,N_9952);
or U12357 (N_12357,N_8453,N_6290);
nor U12358 (N_12358,N_5271,N_7354);
nor U12359 (N_12359,N_9623,N_9876);
and U12360 (N_12360,N_8302,N_6709);
xnor U12361 (N_12361,N_6297,N_7306);
and U12362 (N_12362,N_5249,N_6121);
nand U12363 (N_12363,N_8608,N_5727);
nand U12364 (N_12364,N_5177,N_9787);
nand U12365 (N_12365,N_8494,N_7840);
or U12366 (N_12366,N_8403,N_5478);
nand U12367 (N_12367,N_6452,N_5508);
or U12368 (N_12368,N_5710,N_5503);
and U12369 (N_12369,N_8574,N_6777);
xor U12370 (N_12370,N_5991,N_7587);
nand U12371 (N_12371,N_7498,N_7648);
nand U12372 (N_12372,N_6300,N_5381);
nand U12373 (N_12373,N_6873,N_8840);
nand U12374 (N_12374,N_7645,N_5976);
nor U12375 (N_12375,N_5105,N_9441);
or U12376 (N_12376,N_8461,N_7431);
nand U12377 (N_12377,N_7934,N_7487);
or U12378 (N_12378,N_6714,N_9059);
or U12379 (N_12379,N_6943,N_8251);
nand U12380 (N_12380,N_6839,N_5470);
nor U12381 (N_12381,N_5125,N_6586);
nand U12382 (N_12382,N_7369,N_5791);
and U12383 (N_12383,N_7603,N_6445);
nor U12384 (N_12384,N_9461,N_6001);
and U12385 (N_12385,N_8733,N_9412);
nor U12386 (N_12386,N_7310,N_6252);
nor U12387 (N_12387,N_8672,N_8362);
nand U12388 (N_12388,N_6800,N_5605);
and U12389 (N_12389,N_8308,N_6739);
and U12390 (N_12390,N_8473,N_5613);
and U12391 (N_12391,N_7322,N_9671);
or U12392 (N_12392,N_9679,N_9084);
or U12393 (N_12393,N_7938,N_5287);
or U12394 (N_12394,N_8014,N_5343);
or U12395 (N_12395,N_5189,N_9343);
nand U12396 (N_12396,N_9695,N_7192);
xnor U12397 (N_12397,N_9360,N_7054);
nor U12398 (N_12398,N_7819,N_5019);
nand U12399 (N_12399,N_8242,N_5057);
xor U12400 (N_12400,N_7481,N_8953);
and U12401 (N_12401,N_7803,N_7221);
or U12402 (N_12402,N_5307,N_7732);
or U12403 (N_12403,N_6356,N_8792);
nand U12404 (N_12404,N_8126,N_9302);
or U12405 (N_12405,N_8478,N_8909);
or U12406 (N_12406,N_8249,N_5705);
nand U12407 (N_12407,N_9904,N_5300);
xor U12408 (N_12408,N_9607,N_8364);
nor U12409 (N_12409,N_6826,N_6201);
nor U12410 (N_12410,N_8804,N_5387);
or U12411 (N_12411,N_5792,N_6727);
xnor U12412 (N_12412,N_6079,N_9040);
nand U12413 (N_12413,N_6635,N_7542);
and U12414 (N_12414,N_7183,N_5403);
or U12415 (N_12415,N_9046,N_6956);
xnor U12416 (N_12416,N_7634,N_5591);
nor U12417 (N_12417,N_7468,N_5324);
xnor U12418 (N_12418,N_5357,N_7741);
xor U12419 (N_12419,N_8339,N_9334);
and U12420 (N_12420,N_8698,N_7847);
and U12421 (N_12421,N_7272,N_9350);
and U12422 (N_12422,N_8154,N_9993);
and U12423 (N_12423,N_8380,N_8321);
xor U12424 (N_12424,N_5139,N_5099);
nand U12425 (N_12425,N_9522,N_6822);
nand U12426 (N_12426,N_7244,N_7073);
nor U12427 (N_12427,N_5506,N_8513);
or U12428 (N_12428,N_7998,N_6723);
nand U12429 (N_12429,N_5481,N_7126);
or U12430 (N_12430,N_5190,N_7875);
xnor U12431 (N_12431,N_8212,N_5653);
xnor U12432 (N_12432,N_5187,N_9432);
nand U12433 (N_12433,N_6505,N_9190);
nor U12434 (N_12434,N_9545,N_8651);
and U12435 (N_12435,N_6532,N_9249);
nand U12436 (N_12436,N_5356,N_5933);
and U12437 (N_12437,N_9798,N_7906);
and U12438 (N_12438,N_9290,N_8990);
nor U12439 (N_12439,N_9416,N_8979);
nor U12440 (N_12440,N_5078,N_9816);
or U12441 (N_12441,N_8868,N_6726);
nand U12442 (N_12442,N_5171,N_8934);
nor U12443 (N_12443,N_7032,N_6961);
nand U12444 (N_12444,N_8351,N_8780);
or U12445 (N_12445,N_6885,N_6794);
xnor U12446 (N_12446,N_7078,N_6705);
nor U12447 (N_12447,N_9909,N_6233);
nor U12448 (N_12448,N_8958,N_5834);
or U12449 (N_12449,N_8149,N_5890);
nand U12450 (N_12450,N_6740,N_7708);
nor U12451 (N_12451,N_7463,N_5061);
xor U12452 (N_12452,N_8028,N_9079);
nor U12453 (N_12453,N_7150,N_8036);
or U12454 (N_12454,N_6567,N_9404);
nor U12455 (N_12455,N_9111,N_7584);
or U12456 (N_12456,N_6576,N_7347);
or U12457 (N_12457,N_7311,N_7472);
nand U12458 (N_12458,N_9344,N_5215);
xnor U12459 (N_12459,N_9003,N_5071);
or U12460 (N_12460,N_7229,N_7567);
and U12461 (N_12461,N_7230,N_8425);
nand U12462 (N_12462,N_5165,N_8053);
and U12463 (N_12463,N_5907,N_8388);
nand U12464 (N_12464,N_6510,N_9990);
or U12465 (N_12465,N_8290,N_7240);
and U12466 (N_12466,N_8537,N_5010);
xor U12467 (N_12467,N_8989,N_6222);
nor U12468 (N_12468,N_9211,N_5956);
xor U12469 (N_12469,N_9281,N_9707);
nor U12470 (N_12470,N_5256,N_6809);
xor U12471 (N_12471,N_5863,N_9826);
and U12472 (N_12472,N_5952,N_8863);
or U12473 (N_12473,N_6352,N_5264);
and U12474 (N_12474,N_8611,N_5669);
nand U12475 (N_12475,N_7482,N_6578);
nand U12476 (N_12476,N_9274,N_8057);
or U12477 (N_12477,N_5146,N_7774);
nand U12478 (N_12478,N_9874,N_9366);
and U12479 (N_12479,N_9754,N_9608);
and U12480 (N_12480,N_8771,N_8659);
xor U12481 (N_12481,N_5651,N_6332);
nor U12482 (N_12482,N_6143,N_5214);
nor U12483 (N_12483,N_9154,N_9355);
or U12484 (N_12484,N_6298,N_8929);
xnor U12485 (N_12485,N_5535,N_9485);
nand U12486 (N_12486,N_6546,N_6071);
nand U12487 (N_12487,N_9548,N_5648);
nand U12488 (N_12488,N_7886,N_7866);
and U12489 (N_12489,N_9292,N_6840);
or U12490 (N_12490,N_6159,N_8087);
and U12491 (N_12491,N_8515,N_9285);
nand U12492 (N_12492,N_8310,N_8708);
nand U12493 (N_12493,N_5132,N_5124);
nand U12494 (N_12494,N_8392,N_6535);
nor U12495 (N_12495,N_5634,N_8230);
nand U12496 (N_12496,N_6311,N_8488);
or U12497 (N_12497,N_6134,N_6088);
nor U12498 (N_12498,N_7782,N_5029);
or U12499 (N_12499,N_7143,N_5659);
nand U12500 (N_12500,N_5116,N_9992);
and U12501 (N_12501,N_9201,N_5291);
nand U12502 (N_12502,N_8311,N_9581);
xor U12503 (N_12503,N_9876,N_9050);
or U12504 (N_12504,N_5379,N_9513);
nand U12505 (N_12505,N_9011,N_7531);
nand U12506 (N_12506,N_7036,N_8587);
xnor U12507 (N_12507,N_5909,N_7463);
xnor U12508 (N_12508,N_9732,N_6389);
or U12509 (N_12509,N_7940,N_5567);
and U12510 (N_12510,N_7844,N_5688);
and U12511 (N_12511,N_7270,N_9141);
nor U12512 (N_12512,N_9506,N_8084);
xor U12513 (N_12513,N_6536,N_8584);
nor U12514 (N_12514,N_8195,N_9148);
nor U12515 (N_12515,N_6586,N_6029);
xnor U12516 (N_12516,N_7686,N_5493);
nand U12517 (N_12517,N_8372,N_6482);
and U12518 (N_12518,N_8951,N_7850);
xnor U12519 (N_12519,N_5811,N_5506);
xnor U12520 (N_12520,N_6482,N_8793);
xnor U12521 (N_12521,N_8156,N_6574);
and U12522 (N_12522,N_9653,N_9926);
xnor U12523 (N_12523,N_8894,N_5129);
xor U12524 (N_12524,N_5513,N_7728);
nand U12525 (N_12525,N_7072,N_8396);
and U12526 (N_12526,N_5199,N_7900);
nand U12527 (N_12527,N_6866,N_5336);
nand U12528 (N_12528,N_8252,N_7483);
and U12529 (N_12529,N_5340,N_6978);
or U12530 (N_12530,N_6466,N_7152);
or U12531 (N_12531,N_6744,N_8660);
or U12532 (N_12532,N_6458,N_6827);
nor U12533 (N_12533,N_5183,N_5407);
and U12534 (N_12534,N_8987,N_8901);
nor U12535 (N_12535,N_9079,N_9463);
nor U12536 (N_12536,N_6817,N_9793);
xor U12537 (N_12537,N_8131,N_7888);
or U12538 (N_12538,N_9378,N_8013);
nor U12539 (N_12539,N_7922,N_9193);
and U12540 (N_12540,N_7026,N_9369);
or U12541 (N_12541,N_8350,N_7934);
or U12542 (N_12542,N_9232,N_8855);
nand U12543 (N_12543,N_6137,N_7686);
or U12544 (N_12544,N_7640,N_5092);
xor U12545 (N_12545,N_7460,N_8321);
and U12546 (N_12546,N_9090,N_9348);
nor U12547 (N_12547,N_8333,N_7754);
nand U12548 (N_12548,N_9909,N_7073);
xnor U12549 (N_12549,N_9989,N_5743);
xor U12550 (N_12550,N_6466,N_5404);
nor U12551 (N_12551,N_7041,N_8464);
xnor U12552 (N_12552,N_7902,N_7822);
or U12553 (N_12553,N_6043,N_8143);
xor U12554 (N_12554,N_9602,N_7178);
and U12555 (N_12555,N_9552,N_7104);
nand U12556 (N_12556,N_5157,N_9017);
nand U12557 (N_12557,N_7324,N_6459);
nor U12558 (N_12558,N_5670,N_5860);
xnor U12559 (N_12559,N_8726,N_6771);
nor U12560 (N_12560,N_9837,N_5510);
nand U12561 (N_12561,N_7647,N_7659);
and U12562 (N_12562,N_6609,N_6589);
xnor U12563 (N_12563,N_8099,N_6943);
nor U12564 (N_12564,N_8926,N_7486);
nand U12565 (N_12565,N_5365,N_6809);
nand U12566 (N_12566,N_6525,N_9456);
and U12567 (N_12567,N_7269,N_9466);
nor U12568 (N_12568,N_9557,N_9762);
xor U12569 (N_12569,N_9514,N_5064);
and U12570 (N_12570,N_6896,N_8495);
nor U12571 (N_12571,N_5326,N_7370);
or U12572 (N_12572,N_5776,N_8322);
and U12573 (N_12573,N_7867,N_5297);
xnor U12574 (N_12574,N_9167,N_8668);
nand U12575 (N_12575,N_7379,N_6533);
nor U12576 (N_12576,N_9225,N_7073);
nand U12577 (N_12577,N_5175,N_9633);
nor U12578 (N_12578,N_5340,N_9585);
nand U12579 (N_12579,N_9814,N_9975);
nand U12580 (N_12580,N_8693,N_6629);
nand U12581 (N_12581,N_5024,N_7174);
and U12582 (N_12582,N_5239,N_5506);
and U12583 (N_12583,N_8747,N_5349);
or U12584 (N_12584,N_6224,N_9957);
and U12585 (N_12585,N_8032,N_7688);
and U12586 (N_12586,N_6283,N_7627);
xnor U12587 (N_12587,N_5360,N_9611);
and U12588 (N_12588,N_8762,N_8468);
and U12589 (N_12589,N_9756,N_6641);
nand U12590 (N_12590,N_8602,N_5316);
nand U12591 (N_12591,N_5684,N_9379);
or U12592 (N_12592,N_9545,N_8333);
nand U12593 (N_12593,N_7748,N_6101);
nor U12594 (N_12594,N_9871,N_6908);
and U12595 (N_12595,N_5709,N_8618);
xor U12596 (N_12596,N_5001,N_5952);
and U12597 (N_12597,N_8043,N_6154);
xor U12598 (N_12598,N_5133,N_5640);
and U12599 (N_12599,N_6268,N_8757);
nor U12600 (N_12600,N_5153,N_6329);
xor U12601 (N_12601,N_6190,N_8995);
or U12602 (N_12602,N_7080,N_6646);
or U12603 (N_12603,N_8050,N_9961);
or U12604 (N_12604,N_8992,N_9659);
or U12605 (N_12605,N_9203,N_8435);
or U12606 (N_12606,N_7026,N_7897);
xor U12607 (N_12607,N_7193,N_6930);
nor U12608 (N_12608,N_6685,N_7813);
nor U12609 (N_12609,N_8167,N_9039);
nor U12610 (N_12610,N_5305,N_6644);
nand U12611 (N_12611,N_8448,N_7775);
or U12612 (N_12612,N_7527,N_7870);
nor U12613 (N_12613,N_6748,N_7620);
nand U12614 (N_12614,N_8664,N_9691);
nor U12615 (N_12615,N_9484,N_8020);
nand U12616 (N_12616,N_9716,N_6822);
xor U12617 (N_12617,N_7887,N_9045);
xnor U12618 (N_12618,N_5090,N_8511);
or U12619 (N_12619,N_5306,N_5138);
and U12620 (N_12620,N_7990,N_7113);
nor U12621 (N_12621,N_8936,N_5995);
or U12622 (N_12622,N_9177,N_6278);
or U12623 (N_12623,N_8831,N_6255);
xor U12624 (N_12624,N_5893,N_8462);
xnor U12625 (N_12625,N_8526,N_9565);
nand U12626 (N_12626,N_8079,N_7607);
nand U12627 (N_12627,N_5466,N_8760);
nor U12628 (N_12628,N_9186,N_8947);
and U12629 (N_12629,N_7333,N_7992);
and U12630 (N_12630,N_6539,N_6835);
and U12631 (N_12631,N_7215,N_7225);
or U12632 (N_12632,N_5499,N_7074);
or U12633 (N_12633,N_9828,N_9553);
xnor U12634 (N_12634,N_7503,N_9629);
and U12635 (N_12635,N_6288,N_9321);
or U12636 (N_12636,N_8063,N_5257);
and U12637 (N_12637,N_7599,N_9429);
xor U12638 (N_12638,N_9613,N_5357);
xnor U12639 (N_12639,N_8928,N_8145);
and U12640 (N_12640,N_7827,N_7911);
xnor U12641 (N_12641,N_8198,N_7989);
xnor U12642 (N_12642,N_8623,N_6572);
or U12643 (N_12643,N_6510,N_6749);
nand U12644 (N_12644,N_9423,N_7430);
and U12645 (N_12645,N_5292,N_8824);
nand U12646 (N_12646,N_5581,N_9136);
nand U12647 (N_12647,N_6528,N_5152);
nor U12648 (N_12648,N_9860,N_6975);
or U12649 (N_12649,N_8851,N_9805);
and U12650 (N_12650,N_9615,N_8155);
xnor U12651 (N_12651,N_8156,N_6011);
xor U12652 (N_12652,N_7687,N_7252);
xor U12653 (N_12653,N_5037,N_7903);
nor U12654 (N_12654,N_7058,N_8470);
or U12655 (N_12655,N_8199,N_6877);
and U12656 (N_12656,N_6473,N_7447);
and U12657 (N_12657,N_5884,N_7158);
and U12658 (N_12658,N_7471,N_5135);
nand U12659 (N_12659,N_9583,N_5994);
and U12660 (N_12660,N_5329,N_9026);
xor U12661 (N_12661,N_8688,N_5136);
or U12662 (N_12662,N_8909,N_7497);
or U12663 (N_12663,N_9250,N_6332);
and U12664 (N_12664,N_8804,N_9541);
nor U12665 (N_12665,N_6978,N_7271);
nor U12666 (N_12666,N_7490,N_5736);
or U12667 (N_12667,N_9842,N_9146);
nand U12668 (N_12668,N_5135,N_9850);
xor U12669 (N_12669,N_5645,N_8438);
nand U12670 (N_12670,N_7116,N_6391);
nand U12671 (N_12671,N_7136,N_6403);
xor U12672 (N_12672,N_9463,N_9004);
and U12673 (N_12673,N_8046,N_6227);
xnor U12674 (N_12674,N_9218,N_6683);
or U12675 (N_12675,N_8320,N_8283);
and U12676 (N_12676,N_9422,N_8064);
nand U12677 (N_12677,N_5171,N_7816);
nor U12678 (N_12678,N_6936,N_9881);
or U12679 (N_12679,N_7721,N_6421);
or U12680 (N_12680,N_7317,N_5648);
and U12681 (N_12681,N_7960,N_7850);
and U12682 (N_12682,N_9346,N_9795);
nand U12683 (N_12683,N_7380,N_5468);
or U12684 (N_12684,N_8762,N_7984);
or U12685 (N_12685,N_5934,N_9751);
nor U12686 (N_12686,N_6766,N_5347);
nor U12687 (N_12687,N_8336,N_8611);
nand U12688 (N_12688,N_7403,N_5349);
nand U12689 (N_12689,N_8024,N_7078);
nand U12690 (N_12690,N_9111,N_9539);
xor U12691 (N_12691,N_8602,N_5634);
or U12692 (N_12692,N_8450,N_5794);
or U12693 (N_12693,N_8525,N_8139);
nand U12694 (N_12694,N_6813,N_7944);
nand U12695 (N_12695,N_6831,N_7445);
or U12696 (N_12696,N_8461,N_8066);
nand U12697 (N_12697,N_5583,N_9730);
nand U12698 (N_12698,N_9775,N_6097);
or U12699 (N_12699,N_7252,N_5914);
nor U12700 (N_12700,N_7632,N_6687);
nor U12701 (N_12701,N_6899,N_5529);
nand U12702 (N_12702,N_9901,N_5691);
xnor U12703 (N_12703,N_6453,N_8456);
xnor U12704 (N_12704,N_8745,N_6068);
xor U12705 (N_12705,N_5665,N_7183);
nor U12706 (N_12706,N_9035,N_9563);
nand U12707 (N_12707,N_8584,N_8416);
nand U12708 (N_12708,N_7160,N_7179);
nor U12709 (N_12709,N_5995,N_6176);
nand U12710 (N_12710,N_9544,N_8811);
or U12711 (N_12711,N_9050,N_5018);
nor U12712 (N_12712,N_7723,N_8667);
nor U12713 (N_12713,N_6475,N_5222);
xnor U12714 (N_12714,N_9717,N_5312);
xnor U12715 (N_12715,N_8729,N_6308);
xnor U12716 (N_12716,N_6274,N_7611);
nand U12717 (N_12717,N_9575,N_5844);
and U12718 (N_12718,N_9426,N_9722);
xnor U12719 (N_12719,N_6649,N_7436);
xnor U12720 (N_12720,N_6441,N_5767);
and U12721 (N_12721,N_5903,N_6050);
or U12722 (N_12722,N_6621,N_9132);
nor U12723 (N_12723,N_7942,N_8734);
nand U12724 (N_12724,N_9864,N_8175);
nand U12725 (N_12725,N_9707,N_9368);
or U12726 (N_12726,N_9360,N_8250);
nor U12727 (N_12727,N_6371,N_7188);
xor U12728 (N_12728,N_7208,N_7970);
and U12729 (N_12729,N_7277,N_8140);
or U12730 (N_12730,N_6577,N_7118);
and U12731 (N_12731,N_9334,N_7534);
and U12732 (N_12732,N_5956,N_6891);
nor U12733 (N_12733,N_7614,N_7061);
nand U12734 (N_12734,N_5199,N_5848);
or U12735 (N_12735,N_6148,N_7421);
xnor U12736 (N_12736,N_6387,N_9925);
and U12737 (N_12737,N_8748,N_5328);
nor U12738 (N_12738,N_7456,N_8860);
xor U12739 (N_12739,N_6286,N_7937);
xor U12740 (N_12740,N_7974,N_8306);
and U12741 (N_12741,N_7080,N_5993);
and U12742 (N_12742,N_8382,N_6045);
or U12743 (N_12743,N_9164,N_5900);
and U12744 (N_12744,N_9168,N_7287);
or U12745 (N_12745,N_8916,N_6322);
nand U12746 (N_12746,N_7063,N_7659);
and U12747 (N_12747,N_6991,N_9405);
nor U12748 (N_12748,N_8607,N_7845);
nor U12749 (N_12749,N_8533,N_7268);
or U12750 (N_12750,N_6454,N_6508);
nand U12751 (N_12751,N_5113,N_5311);
or U12752 (N_12752,N_7514,N_6948);
and U12753 (N_12753,N_9795,N_6713);
nor U12754 (N_12754,N_6775,N_9780);
and U12755 (N_12755,N_5456,N_5013);
nand U12756 (N_12756,N_5708,N_5698);
nand U12757 (N_12757,N_5400,N_8246);
xor U12758 (N_12758,N_9176,N_7273);
xor U12759 (N_12759,N_7932,N_8009);
and U12760 (N_12760,N_7579,N_9656);
and U12761 (N_12761,N_6995,N_5559);
nor U12762 (N_12762,N_5417,N_8349);
xor U12763 (N_12763,N_6645,N_7771);
nor U12764 (N_12764,N_5949,N_6957);
and U12765 (N_12765,N_9260,N_7508);
and U12766 (N_12766,N_6756,N_9985);
nand U12767 (N_12767,N_9429,N_8854);
or U12768 (N_12768,N_7812,N_8196);
and U12769 (N_12769,N_5341,N_9270);
nand U12770 (N_12770,N_8038,N_9098);
xor U12771 (N_12771,N_6667,N_9917);
nor U12772 (N_12772,N_9209,N_8039);
nor U12773 (N_12773,N_8307,N_9944);
xor U12774 (N_12774,N_8816,N_5117);
xor U12775 (N_12775,N_8101,N_9058);
xnor U12776 (N_12776,N_9736,N_8902);
xor U12777 (N_12777,N_6165,N_6302);
and U12778 (N_12778,N_6220,N_9538);
xnor U12779 (N_12779,N_5576,N_9101);
or U12780 (N_12780,N_5126,N_9374);
xor U12781 (N_12781,N_6718,N_5196);
and U12782 (N_12782,N_7582,N_7221);
xor U12783 (N_12783,N_8252,N_8003);
and U12784 (N_12784,N_7336,N_9931);
nor U12785 (N_12785,N_5281,N_9482);
or U12786 (N_12786,N_9985,N_9259);
nor U12787 (N_12787,N_8330,N_8568);
and U12788 (N_12788,N_6003,N_7480);
nand U12789 (N_12789,N_9337,N_9314);
or U12790 (N_12790,N_9861,N_7754);
xnor U12791 (N_12791,N_7277,N_8241);
xnor U12792 (N_12792,N_7698,N_7455);
and U12793 (N_12793,N_5626,N_7703);
or U12794 (N_12794,N_6553,N_6629);
and U12795 (N_12795,N_8755,N_5007);
or U12796 (N_12796,N_8488,N_8355);
nand U12797 (N_12797,N_5752,N_7823);
nand U12798 (N_12798,N_5429,N_8445);
xnor U12799 (N_12799,N_7114,N_9896);
nand U12800 (N_12800,N_5723,N_6581);
nand U12801 (N_12801,N_9665,N_6614);
and U12802 (N_12802,N_7942,N_5390);
nor U12803 (N_12803,N_6044,N_9293);
xnor U12804 (N_12804,N_9006,N_9371);
xnor U12805 (N_12805,N_9687,N_5259);
nor U12806 (N_12806,N_8361,N_9700);
nand U12807 (N_12807,N_9690,N_5393);
or U12808 (N_12808,N_5408,N_8435);
and U12809 (N_12809,N_9123,N_6413);
or U12810 (N_12810,N_8835,N_6890);
nand U12811 (N_12811,N_9348,N_8701);
or U12812 (N_12812,N_8722,N_9762);
nand U12813 (N_12813,N_9209,N_5104);
nor U12814 (N_12814,N_5908,N_7478);
nand U12815 (N_12815,N_6687,N_5340);
xnor U12816 (N_12816,N_9785,N_9671);
and U12817 (N_12817,N_7974,N_6338);
nand U12818 (N_12818,N_7411,N_5977);
nand U12819 (N_12819,N_7617,N_8299);
nand U12820 (N_12820,N_8284,N_8600);
nor U12821 (N_12821,N_8778,N_7384);
nand U12822 (N_12822,N_5201,N_5168);
or U12823 (N_12823,N_8750,N_6924);
xnor U12824 (N_12824,N_9807,N_9804);
xor U12825 (N_12825,N_7375,N_5606);
and U12826 (N_12826,N_6238,N_7120);
nand U12827 (N_12827,N_9593,N_9741);
xnor U12828 (N_12828,N_7460,N_8240);
nand U12829 (N_12829,N_6754,N_5745);
xor U12830 (N_12830,N_8071,N_9223);
and U12831 (N_12831,N_5309,N_8170);
or U12832 (N_12832,N_5197,N_8961);
nor U12833 (N_12833,N_7191,N_8518);
xnor U12834 (N_12834,N_7011,N_8131);
and U12835 (N_12835,N_8145,N_8820);
or U12836 (N_12836,N_6972,N_8803);
or U12837 (N_12837,N_7811,N_5368);
nand U12838 (N_12838,N_7827,N_6385);
and U12839 (N_12839,N_9671,N_7126);
or U12840 (N_12840,N_6843,N_9563);
nand U12841 (N_12841,N_7730,N_6516);
xnor U12842 (N_12842,N_7875,N_7210);
and U12843 (N_12843,N_9730,N_7480);
xnor U12844 (N_12844,N_8378,N_7505);
or U12845 (N_12845,N_6692,N_9091);
nor U12846 (N_12846,N_9272,N_5249);
or U12847 (N_12847,N_7124,N_5819);
and U12848 (N_12848,N_7011,N_7390);
xnor U12849 (N_12849,N_7027,N_6674);
or U12850 (N_12850,N_8414,N_7281);
nor U12851 (N_12851,N_8900,N_5445);
and U12852 (N_12852,N_9376,N_9649);
and U12853 (N_12853,N_9383,N_7479);
nand U12854 (N_12854,N_5421,N_6488);
xor U12855 (N_12855,N_5870,N_8539);
xor U12856 (N_12856,N_9731,N_8617);
xnor U12857 (N_12857,N_8513,N_8653);
and U12858 (N_12858,N_8432,N_6847);
and U12859 (N_12859,N_9058,N_9665);
xnor U12860 (N_12860,N_7477,N_7009);
nand U12861 (N_12861,N_7196,N_7098);
or U12862 (N_12862,N_9921,N_9464);
and U12863 (N_12863,N_9474,N_6842);
xor U12864 (N_12864,N_7864,N_6360);
nand U12865 (N_12865,N_8507,N_5874);
or U12866 (N_12866,N_8453,N_8886);
xnor U12867 (N_12867,N_7193,N_6706);
xnor U12868 (N_12868,N_6189,N_7723);
or U12869 (N_12869,N_5585,N_6661);
nand U12870 (N_12870,N_8453,N_9717);
and U12871 (N_12871,N_8813,N_9947);
or U12872 (N_12872,N_9192,N_8607);
or U12873 (N_12873,N_5664,N_5147);
or U12874 (N_12874,N_8148,N_6183);
or U12875 (N_12875,N_9074,N_9728);
nand U12876 (N_12876,N_9124,N_9756);
nor U12877 (N_12877,N_9936,N_7457);
nor U12878 (N_12878,N_5376,N_5846);
or U12879 (N_12879,N_7558,N_7838);
xnor U12880 (N_12880,N_5597,N_5598);
or U12881 (N_12881,N_5586,N_6581);
nor U12882 (N_12882,N_8008,N_9198);
nor U12883 (N_12883,N_8356,N_6247);
and U12884 (N_12884,N_7440,N_9459);
xnor U12885 (N_12885,N_9864,N_6168);
nor U12886 (N_12886,N_6648,N_8836);
and U12887 (N_12887,N_6013,N_5866);
or U12888 (N_12888,N_9250,N_6688);
and U12889 (N_12889,N_6055,N_8592);
nor U12890 (N_12890,N_7922,N_5187);
nor U12891 (N_12891,N_5238,N_6846);
or U12892 (N_12892,N_7698,N_8221);
nor U12893 (N_12893,N_8500,N_6831);
nand U12894 (N_12894,N_7886,N_7229);
or U12895 (N_12895,N_8350,N_7519);
nand U12896 (N_12896,N_9509,N_5822);
nor U12897 (N_12897,N_6933,N_7746);
xor U12898 (N_12898,N_9539,N_7834);
nand U12899 (N_12899,N_5675,N_6109);
nand U12900 (N_12900,N_7490,N_8994);
and U12901 (N_12901,N_5505,N_7694);
or U12902 (N_12902,N_5063,N_9811);
and U12903 (N_12903,N_5927,N_6474);
xor U12904 (N_12904,N_6485,N_8575);
nand U12905 (N_12905,N_6924,N_5189);
and U12906 (N_12906,N_8895,N_6774);
and U12907 (N_12907,N_6818,N_6519);
nand U12908 (N_12908,N_7446,N_7849);
xnor U12909 (N_12909,N_9159,N_5462);
nand U12910 (N_12910,N_8518,N_5512);
or U12911 (N_12911,N_5170,N_8810);
and U12912 (N_12912,N_9839,N_9181);
nor U12913 (N_12913,N_9849,N_9094);
or U12914 (N_12914,N_9979,N_6790);
nor U12915 (N_12915,N_8967,N_9818);
and U12916 (N_12916,N_9645,N_5788);
nand U12917 (N_12917,N_6393,N_9214);
and U12918 (N_12918,N_5667,N_5215);
nand U12919 (N_12919,N_8605,N_7879);
or U12920 (N_12920,N_5179,N_9469);
nor U12921 (N_12921,N_8186,N_5515);
nor U12922 (N_12922,N_6861,N_5181);
nand U12923 (N_12923,N_6495,N_7232);
and U12924 (N_12924,N_5555,N_8585);
or U12925 (N_12925,N_7054,N_8606);
or U12926 (N_12926,N_6808,N_9915);
nand U12927 (N_12927,N_6419,N_6367);
and U12928 (N_12928,N_7034,N_5590);
nand U12929 (N_12929,N_7819,N_6681);
or U12930 (N_12930,N_7029,N_6179);
xnor U12931 (N_12931,N_5865,N_7812);
xnor U12932 (N_12932,N_6150,N_6399);
and U12933 (N_12933,N_5223,N_6600);
and U12934 (N_12934,N_6110,N_9383);
nor U12935 (N_12935,N_7568,N_6835);
nor U12936 (N_12936,N_6069,N_6297);
and U12937 (N_12937,N_5400,N_9957);
nor U12938 (N_12938,N_8076,N_8849);
or U12939 (N_12939,N_7110,N_5538);
and U12940 (N_12940,N_5837,N_5370);
or U12941 (N_12941,N_9438,N_9919);
xor U12942 (N_12942,N_7244,N_7205);
xnor U12943 (N_12943,N_8478,N_5584);
nor U12944 (N_12944,N_9388,N_8001);
nand U12945 (N_12945,N_7337,N_7842);
nand U12946 (N_12946,N_6241,N_5176);
and U12947 (N_12947,N_8813,N_6096);
or U12948 (N_12948,N_5759,N_5083);
nor U12949 (N_12949,N_8683,N_8308);
and U12950 (N_12950,N_5677,N_8850);
and U12951 (N_12951,N_5987,N_7504);
xnor U12952 (N_12952,N_7865,N_6370);
nor U12953 (N_12953,N_9230,N_7919);
xnor U12954 (N_12954,N_9503,N_5232);
nand U12955 (N_12955,N_5200,N_5173);
xnor U12956 (N_12956,N_7118,N_6064);
xnor U12957 (N_12957,N_5327,N_7977);
xor U12958 (N_12958,N_6018,N_6749);
or U12959 (N_12959,N_8827,N_6309);
xor U12960 (N_12960,N_6033,N_9835);
and U12961 (N_12961,N_8835,N_5936);
nor U12962 (N_12962,N_6692,N_6965);
nor U12963 (N_12963,N_6060,N_9861);
nand U12964 (N_12964,N_5192,N_7926);
xor U12965 (N_12965,N_9970,N_6348);
or U12966 (N_12966,N_6643,N_9398);
nor U12967 (N_12967,N_8270,N_7715);
and U12968 (N_12968,N_8074,N_7892);
and U12969 (N_12969,N_9051,N_5326);
and U12970 (N_12970,N_7160,N_7551);
and U12971 (N_12971,N_5812,N_9930);
nor U12972 (N_12972,N_9061,N_7960);
and U12973 (N_12973,N_7621,N_8296);
nor U12974 (N_12974,N_6612,N_5812);
xor U12975 (N_12975,N_6464,N_5558);
nand U12976 (N_12976,N_9930,N_9118);
or U12977 (N_12977,N_8357,N_7857);
or U12978 (N_12978,N_8921,N_9389);
nand U12979 (N_12979,N_8395,N_5080);
xnor U12980 (N_12980,N_6454,N_5635);
and U12981 (N_12981,N_7967,N_5588);
nor U12982 (N_12982,N_5935,N_9224);
nand U12983 (N_12983,N_9519,N_8181);
and U12984 (N_12984,N_8280,N_6587);
nand U12985 (N_12985,N_8535,N_6506);
xor U12986 (N_12986,N_6256,N_8947);
nand U12987 (N_12987,N_7087,N_5492);
or U12988 (N_12988,N_6423,N_5702);
or U12989 (N_12989,N_5232,N_9253);
or U12990 (N_12990,N_6422,N_6054);
and U12991 (N_12991,N_9952,N_8733);
and U12992 (N_12992,N_7202,N_6695);
nor U12993 (N_12993,N_9977,N_5257);
and U12994 (N_12994,N_7070,N_9947);
and U12995 (N_12995,N_6654,N_7601);
nor U12996 (N_12996,N_8690,N_9494);
nand U12997 (N_12997,N_8282,N_6616);
nor U12998 (N_12998,N_5837,N_7466);
or U12999 (N_12999,N_8771,N_5128);
nand U13000 (N_13000,N_7586,N_9236);
and U13001 (N_13001,N_7319,N_8790);
nor U13002 (N_13002,N_5895,N_5456);
xnor U13003 (N_13003,N_9646,N_7296);
nor U13004 (N_13004,N_7685,N_5001);
and U13005 (N_13005,N_6841,N_8691);
or U13006 (N_13006,N_5549,N_6076);
or U13007 (N_13007,N_7927,N_9913);
nor U13008 (N_13008,N_6543,N_7739);
nand U13009 (N_13009,N_9492,N_9822);
and U13010 (N_13010,N_9568,N_5930);
nor U13011 (N_13011,N_9078,N_6282);
nand U13012 (N_13012,N_9732,N_7300);
or U13013 (N_13013,N_7097,N_5910);
and U13014 (N_13014,N_8938,N_7224);
and U13015 (N_13015,N_5558,N_5918);
nand U13016 (N_13016,N_7221,N_6397);
and U13017 (N_13017,N_8941,N_7981);
and U13018 (N_13018,N_6059,N_8186);
and U13019 (N_13019,N_8040,N_7569);
xor U13020 (N_13020,N_6157,N_9269);
nor U13021 (N_13021,N_5477,N_5126);
xnor U13022 (N_13022,N_8479,N_5873);
and U13023 (N_13023,N_7351,N_5671);
xnor U13024 (N_13024,N_7701,N_9356);
or U13025 (N_13025,N_8137,N_6308);
nor U13026 (N_13026,N_8263,N_7968);
or U13027 (N_13027,N_5351,N_5300);
nor U13028 (N_13028,N_6768,N_6846);
nor U13029 (N_13029,N_9235,N_8984);
xor U13030 (N_13030,N_8069,N_6706);
xnor U13031 (N_13031,N_8821,N_5966);
nor U13032 (N_13032,N_5709,N_7529);
xnor U13033 (N_13033,N_7369,N_7101);
nor U13034 (N_13034,N_6138,N_9674);
nor U13035 (N_13035,N_5989,N_9030);
and U13036 (N_13036,N_6100,N_6476);
or U13037 (N_13037,N_9959,N_9245);
or U13038 (N_13038,N_9913,N_6593);
nand U13039 (N_13039,N_5164,N_8130);
or U13040 (N_13040,N_6361,N_7584);
nand U13041 (N_13041,N_5919,N_6365);
or U13042 (N_13042,N_8704,N_5188);
xnor U13043 (N_13043,N_5832,N_8068);
and U13044 (N_13044,N_6516,N_7715);
nand U13045 (N_13045,N_8522,N_7306);
nor U13046 (N_13046,N_5499,N_7600);
and U13047 (N_13047,N_5839,N_5481);
nand U13048 (N_13048,N_9121,N_5722);
xnor U13049 (N_13049,N_8867,N_8534);
or U13050 (N_13050,N_8887,N_7146);
and U13051 (N_13051,N_6112,N_9402);
nor U13052 (N_13052,N_8959,N_7959);
xnor U13053 (N_13053,N_5868,N_6556);
or U13054 (N_13054,N_5074,N_6372);
and U13055 (N_13055,N_6627,N_7055);
xnor U13056 (N_13056,N_8473,N_8974);
xnor U13057 (N_13057,N_9937,N_7633);
nand U13058 (N_13058,N_6851,N_9569);
xor U13059 (N_13059,N_5099,N_7510);
or U13060 (N_13060,N_9200,N_9471);
nand U13061 (N_13061,N_8848,N_8442);
nand U13062 (N_13062,N_6625,N_5598);
nand U13063 (N_13063,N_7678,N_5291);
nand U13064 (N_13064,N_6315,N_8193);
and U13065 (N_13065,N_6157,N_9550);
or U13066 (N_13066,N_9548,N_7120);
xor U13067 (N_13067,N_8762,N_6172);
or U13068 (N_13068,N_5951,N_8166);
xor U13069 (N_13069,N_7210,N_8746);
nand U13070 (N_13070,N_6606,N_7782);
xnor U13071 (N_13071,N_7287,N_7515);
nor U13072 (N_13072,N_6985,N_5182);
nand U13073 (N_13073,N_6062,N_5281);
xnor U13074 (N_13074,N_6878,N_5988);
and U13075 (N_13075,N_9074,N_7501);
and U13076 (N_13076,N_5668,N_6921);
nor U13077 (N_13077,N_6589,N_6678);
and U13078 (N_13078,N_6736,N_9065);
nand U13079 (N_13079,N_9357,N_6526);
and U13080 (N_13080,N_5390,N_5939);
nand U13081 (N_13081,N_8020,N_8363);
nand U13082 (N_13082,N_8412,N_7692);
xor U13083 (N_13083,N_7815,N_5707);
nand U13084 (N_13084,N_7320,N_8087);
and U13085 (N_13085,N_5499,N_8277);
xnor U13086 (N_13086,N_9904,N_9887);
and U13087 (N_13087,N_7924,N_7816);
or U13088 (N_13088,N_8254,N_6930);
xor U13089 (N_13089,N_9459,N_7388);
or U13090 (N_13090,N_9085,N_9130);
and U13091 (N_13091,N_6631,N_6637);
nor U13092 (N_13092,N_7611,N_9692);
nor U13093 (N_13093,N_9987,N_8573);
and U13094 (N_13094,N_8741,N_5656);
or U13095 (N_13095,N_6227,N_5813);
or U13096 (N_13096,N_7463,N_9384);
or U13097 (N_13097,N_5872,N_9960);
xnor U13098 (N_13098,N_6118,N_8327);
nor U13099 (N_13099,N_7615,N_6464);
nor U13100 (N_13100,N_5337,N_6397);
nand U13101 (N_13101,N_6338,N_9834);
and U13102 (N_13102,N_9160,N_6438);
nand U13103 (N_13103,N_5061,N_7923);
nor U13104 (N_13104,N_9403,N_7434);
or U13105 (N_13105,N_9829,N_6162);
or U13106 (N_13106,N_5674,N_5168);
and U13107 (N_13107,N_8914,N_5012);
or U13108 (N_13108,N_9278,N_6235);
nand U13109 (N_13109,N_6575,N_5151);
nor U13110 (N_13110,N_9270,N_8617);
xnor U13111 (N_13111,N_7265,N_5162);
xor U13112 (N_13112,N_8938,N_9142);
nor U13113 (N_13113,N_7933,N_5657);
or U13114 (N_13114,N_6261,N_8107);
nand U13115 (N_13115,N_5586,N_8926);
and U13116 (N_13116,N_5634,N_8370);
and U13117 (N_13117,N_8307,N_7053);
nor U13118 (N_13118,N_9064,N_6487);
nand U13119 (N_13119,N_7017,N_8768);
nor U13120 (N_13120,N_8590,N_5219);
xor U13121 (N_13121,N_8203,N_5029);
or U13122 (N_13122,N_6353,N_5960);
and U13123 (N_13123,N_6465,N_7203);
nand U13124 (N_13124,N_5893,N_5885);
and U13125 (N_13125,N_6199,N_6487);
nand U13126 (N_13126,N_9707,N_7799);
nor U13127 (N_13127,N_5279,N_8668);
xor U13128 (N_13128,N_7389,N_7293);
nand U13129 (N_13129,N_8966,N_9293);
nor U13130 (N_13130,N_8950,N_6333);
nand U13131 (N_13131,N_7119,N_5813);
or U13132 (N_13132,N_9966,N_8533);
nor U13133 (N_13133,N_6448,N_7792);
or U13134 (N_13134,N_7877,N_6150);
nand U13135 (N_13135,N_6599,N_8853);
nor U13136 (N_13136,N_6900,N_9407);
or U13137 (N_13137,N_5986,N_5110);
or U13138 (N_13138,N_7667,N_8799);
or U13139 (N_13139,N_5216,N_9060);
nand U13140 (N_13140,N_9510,N_8442);
nor U13141 (N_13141,N_7760,N_7887);
nand U13142 (N_13142,N_9613,N_8641);
and U13143 (N_13143,N_8895,N_6457);
nor U13144 (N_13144,N_8717,N_5241);
nor U13145 (N_13145,N_6437,N_8334);
nor U13146 (N_13146,N_8382,N_9209);
nor U13147 (N_13147,N_6584,N_7120);
nor U13148 (N_13148,N_9831,N_5516);
nand U13149 (N_13149,N_9959,N_8263);
xnor U13150 (N_13150,N_9448,N_5105);
nor U13151 (N_13151,N_6903,N_6038);
or U13152 (N_13152,N_6873,N_7095);
nor U13153 (N_13153,N_7001,N_9027);
nand U13154 (N_13154,N_7556,N_7592);
or U13155 (N_13155,N_8026,N_7839);
nor U13156 (N_13156,N_5062,N_5258);
nor U13157 (N_13157,N_7563,N_8395);
nor U13158 (N_13158,N_6759,N_6213);
nor U13159 (N_13159,N_5926,N_7867);
nand U13160 (N_13160,N_5762,N_9055);
xor U13161 (N_13161,N_9451,N_5371);
or U13162 (N_13162,N_6717,N_8765);
nand U13163 (N_13163,N_9140,N_9709);
or U13164 (N_13164,N_7106,N_7792);
xnor U13165 (N_13165,N_6249,N_6009);
nand U13166 (N_13166,N_5701,N_9166);
xor U13167 (N_13167,N_7046,N_5425);
nor U13168 (N_13168,N_6603,N_6840);
and U13169 (N_13169,N_6191,N_7877);
nand U13170 (N_13170,N_8044,N_6336);
nand U13171 (N_13171,N_7898,N_5246);
or U13172 (N_13172,N_8202,N_6539);
nor U13173 (N_13173,N_5462,N_5416);
and U13174 (N_13174,N_7900,N_7753);
nor U13175 (N_13175,N_6169,N_9979);
or U13176 (N_13176,N_8579,N_7829);
nor U13177 (N_13177,N_9195,N_8177);
nor U13178 (N_13178,N_6170,N_7455);
and U13179 (N_13179,N_8983,N_9235);
nand U13180 (N_13180,N_6350,N_5371);
xnor U13181 (N_13181,N_6173,N_7356);
and U13182 (N_13182,N_5484,N_7615);
or U13183 (N_13183,N_7001,N_9476);
xor U13184 (N_13184,N_6272,N_6203);
nor U13185 (N_13185,N_5990,N_6399);
and U13186 (N_13186,N_9555,N_9569);
nor U13187 (N_13187,N_5752,N_6681);
nor U13188 (N_13188,N_8870,N_7270);
nand U13189 (N_13189,N_7737,N_5334);
xor U13190 (N_13190,N_6227,N_8188);
nor U13191 (N_13191,N_9292,N_5196);
xor U13192 (N_13192,N_6999,N_8259);
nor U13193 (N_13193,N_7969,N_5907);
xnor U13194 (N_13194,N_5452,N_5119);
or U13195 (N_13195,N_5184,N_5399);
nor U13196 (N_13196,N_5839,N_8112);
nand U13197 (N_13197,N_8303,N_8012);
and U13198 (N_13198,N_6703,N_7283);
and U13199 (N_13199,N_8427,N_8163);
nand U13200 (N_13200,N_7722,N_6684);
or U13201 (N_13201,N_9021,N_5600);
nor U13202 (N_13202,N_6334,N_9273);
xor U13203 (N_13203,N_7549,N_5512);
nand U13204 (N_13204,N_6433,N_5776);
nand U13205 (N_13205,N_6006,N_9765);
xor U13206 (N_13206,N_7739,N_7846);
or U13207 (N_13207,N_8582,N_8898);
nor U13208 (N_13208,N_7695,N_9750);
and U13209 (N_13209,N_6512,N_5370);
nor U13210 (N_13210,N_7989,N_5693);
nor U13211 (N_13211,N_9611,N_6405);
or U13212 (N_13212,N_5773,N_5492);
xnor U13213 (N_13213,N_8856,N_6629);
and U13214 (N_13214,N_6724,N_9050);
and U13215 (N_13215,N_7819,N_9224);
xnor U13216 (N_13216,N_7906,N_5160);
or U13217 (N_13217,N_5559,N_8994);
nor U13218 (N_13218,N_5616,N_9734);
or U13219 (N_13219,N_9812,N_8152);
xor U13220 (N_13220,N_7636,N_9800);
or U13221 (N_13221,N_8034,N_8313);
nor U13222 (N_13222,N_6400,N_9505);
or U13223 (N_13223,N_5227,N_8394);
and U13224 (N_13224,N_9264,N_6310);
or U13225 (N_13225,N_8284,N_8490);
and U13226 (N_13226,N_7079,N_9357);
or U13227 (N_13227,N_9908,N_8064);
xor U13228 (N_13228,N_9387,N_7457);
or U13229 (N_13229,N_5202,N_5897);
nand U13230 (N_13230,N_6522,N_8515);
nor U13231 (N_13231,N_9850,N_8533);
and U13232 (N_13232,N_6172,N_7589);
nand U13233 (N_13233,N_7728,N_5648);
nor U13234 (N_13234,N_9130,N_5328);
xor U13235 (N_13235,N_7665,N_9066);
or U13236 (N_13236,N_9566,N_9828);
or U13237 (N_13237,N_6076,N_8396);
or U13238 (N_13238,N_5878,N_6761);
or U13239 (N_13239,N_9861,N_9356);
xnor U13240 (N_13240,N_5120,N_5596);
nand U13241 (N_13241,N_6875,N_9445);
nand U13242 (N_13242,N_6886,N_9813);
xnor U13243 (N_13243,N_9270,N_7371);
nor U13244 (N_13244,N_7670,N_9435);
and U13245 (N_13245,N_5270,N_5307);
nand U13246 (N_13246,N_6148,N_9771);
or U13247 (N_13247,N_6195,N_7968);
xnor U13248 (N_13248,N_5120,N_6973);
nor U13249 (N_13249,N_7682,N_5939);
nand U13250 (N_13250,N_6789,N_9441);
nor U13251 (N_13251,N_7835,N_5225);
nand U13252 (N_13252,N_5609,N_8139);
xor U13253 (N_13253,N_7225,N_6836);
xnor U13254 (N_13254,N_8732,N_8176);
nand U13255 (N_13255,N_8730,N_7405);
and U13256 (N_13256,N_8148,N_9239);
nand U13257 (N_13257,N_5425,N_8989);
or U13258 (N_13258,N_9421,N_8193);
and U13259 (N_13259,N_5350,N_8280);
and U13260 (N_13260,N_5001,N_8468);
xnor U13261 (N_13261,N_5168,N_8541);
xor U13262 (N_13262,N_8230,N_7412);
and U13263 (N_13263,N_8366,N_5416);
nand U13264 (N_13264,N_6600,N_9273);
and U13265 (N_13265,N_9376,N_6279);
nand U13266 (N_13266,N_5513,N_8749);
xnor U13267 (N_13267,N_5513,N_8235);
or U13268 (N_13268,N_9770,N_9711);
nor U13269 (N_13269,N_9241,N_6785);
or U13270 (N_13270,N_9970,N_5245);
xnor U13271 (N_13271,N_9108,N_8489);
xor U13272 (N_13272,N_8330,N_6892);
and U13273 (N_13273,N_8346,N_9831);
nor U13274 (N_13274,N_8850,N_8070);
or U13275 (N_13275,N_6712,N_5179);
nand U13276 (N_13276,N_8333,N_6997);
and U13277 (N_13277,N_5739,N_8711);
and U13278 (N_13278,N_8109,N_9984);
nand U13279 (N_13279,N_8362,N_6798);
nand U13280 (N_13280,N_8134,N_9177);
and U13281 (N_13281,N_5642,N_9220);
and U13282 (N_13282,N_6303,N_8741);
nor U13283 (N_13283,N_7363,N_5932);
nor U13284 (N_13284,N_7239,N_6178);
or U13285 (N_13285,N_6638,N_7255);
nor U13286 (N_13286,N_7471,N_9370);
nor U13287 (N_13287,N_9991,N_7956);
nand U13288 (N_13288,N_9249,N_7142);
xor U13289 (N_13289,N_6047,N_7674);
and U13290 (N_13290,N_7106,N_6137);
nand U13291 (N_13291,N_5170,N_9243);
and U13292 (N_13292,N_7867,N_8570);
nand U13293 (N_13293,N_5624,N_6344);
or U13294 (N_13294,N_7520,N_7451);
xnor U13295 (N_13295,N_9937,N_5915);
and U13296 (N_13296,N_6226,N_7080);
nand U13297 (N_13297,N_9521,N_7742);
and U13298 (N_13298,N_6098,N_5573);
or U13299 (N_13299,N_8808,N_5600);
or U13300 (N_13300,N_6922,N_5228);
xnor U13301 (N_13301,N_9523,N_7288);
xor U13302 (N_13302,N_5325,N_7862);
and U13303 (N_13303,N_9517,N_9614);
xor U13304 (N_13304,N_6408,N_9246);
nor U13305 (N_13305,N_8004,N_8817);
and U13306 (N_13306,N_9929,N_6534);
nand U13307 (N_13307,N_8051,N_8347);
nand U13308 (N_13308,N_5859,N_9396);
and U13309 (N_13309,N_6440,N_5160);
nand U13310 (N_13310,N_7328,N_5143);
nor U13311 (N_13311,N_8386,N_9573);
xor U13312 (N_13312,N_8799,N_5643);
nand U13313 (N_13313,N_6676,N_7844);
nor U13314 (N_13314,N_8875,N_9389);
nor U13315 (N_13315,N_7702,N_9496);
and U13316 (N_13316,N_8900,N_5086);
and U13317 (N_13317,N_8924,N_9983);
nand U13318 (N_13318,N_9908,N_8862);
and U13319 (N_13319,N_9966,N_9703);
nor U13320 (N_13320,N_8145,N_5474);
or U13321 (N_13321,N_6469,N_5560);
nor U13322 (N_13322,N_9800,N_5869);
nand U13323 (N_13323,N_5131,N_9026);
xnor U13324 (N_13324,N_5712,N_9820);
and U13325 (N_13325,N_8683,N_9747);
nor U13326 (N_13326,N_7865,N_8815);
nand U13327 (N_13327,N_9440,N_6532);
and U13328 (N_13328,N_5974,N_5397);
nor U13329 (N_13329,N_8330,N_6092);
xnor U13330 (N_13330,N_7984,N_6409);
and U13331 (N_13331,N_8695,N_9436);
or U13332 (N_13332,N_7830,N_6828);
xor U13333 (N_13333,N_5485,N_6970);
nor U13334 (N_13334,N_7144,N_6964);
nor U13335 (N_13335,N_5506,N_8273);
nor U13336 (N_13336,N_5438,N_9144);
nor U13337 (N_13337,N_7367,N_9093);
xnor U13338 (N_13338,N_6070,N_6872);
xor U13339 (N_13339,N_6012,N_7319);
nand U13340 (N_13340,N_8518,N_6174);
nand U13341 (N_13341,N_8340,N_6803);
and U13342 (N_13342,N_5330,N_5097);
xnor U13343 (N_13343,N_9536,N_5961);
or U13344 (N_13344,N_5777,N_7088);
nor U13345 (N_13345,N_6962,N_7448);
and U13346 (N_13346,N_8523,N_6545);
nand U13347 (N_13347,N_7201,N_8026);
nor U13348 (N_13348,N_7898,N_9740);
xor U13349 (N_13349,N_8303,N_7350);
nor U13350 (N_13350,N_5608,N_9347);
xor U13351 (N_13351,N_5007,N_5097);
nand U13352 (N_13352,N_6178,N_5272);
xor U13353 (N_13353,N_7637,N_6731);
and U13354 (N_13354,N_7310,N_7444);
xor U13355 (N_13355,N_6639,N_7378);
xor U13356 (N_13356,N_9405,N_6143);
or U13357 (N_13357,N_6720,N_6055);
nand U13358 (N_13358,N_8205,N_5547);
nor U13359 (N_13359,N_6550,N_6026);
nand U13360 (N_13360,N_9740,N_5573);
and U13361 (N_13361,N_7697,N_9882);
nor U13362 (N_13362,N_7621,N_9270);
xor U13363 (N_13363,N_6253,N_7777);
xor U13364 (N_13364,N_5563,N_8903);
nand U13365 (N_13365,N_6726,N_9323);
or U13366 (N_13366,N_5513,N_7842);
nand U13367 (N_13367,N_7329,N_6048);
nor U13368 (N_13368,N_7361,N_5979);
xnor U13369 (N_13369,N_7823,N_6124);
nand U13370 (N_13370,N_6107,N_5030);
xnor U13371 (N_13371,N_7837,N_8398);
nand U13372 (N_13372,N_9424,N_5609);
xnor U13373 (N_13373,N_5557,N_5690);
xor U13374 (N_13374,N_9418,N_9439);
nand U13375 (N_13375,N_6443,N_8720);
xnor U13376 (N_13376,N_7502,N_6023);
nand U13377 (N_13377,N_9167,N_7124);
nand U13378 (N_13378,N_6671,N_5662);
nor U13379 (N_13379,N_9449,N_5248);
xor U13380 (N_13380,N_7833,N_7844);
xor U13381 (N_13381,N_5660,N_6236);
nand U13382 (N_13382,N_5826,N_9825);
nor U13383 (N_13383,N_7746,N_7953);
xor U13384 (N_13384,N_7003,N_9633);
xor U13385 (N_13385,N_6415,N_7492);
or U13386 (N_13386,N_9338,N_9345);
nand U13387 (N_13387,N_5584,N_8650);
or U13388 (N_13388,N_6591,N_6488);
and U13389 (N_13389,N_8989,N_9150);
nand U13390 (N_13390,N_7118,N_9056);
xor U13391 (N_13391,N_6477,N_8634);
xor U13392 (N_13392,N_6612,N_5323);
or U13393 (N_13393,N_6193,N_9608);
or U13394 (N_13394,N_7469,N_9597);
and U13395 (N_13395,N_7321,N_9327);
and U13396 (N_13396,N_6507,N_8883);
nand U13397 (N_13397,N_5440,N_9255);
and U13398 (N_13398,N_5698,N_7083);
and U13399 (N_13399,N_8719,N_8311);
nand U13400 (N_13400,N_5748,N_8915);
xnor U13401 (N_13401,N_7346,N_7922);
nand U13402 (N_13402,N_8389,N_6997);
nand U13403 (N_13403,N_7190,N_8963);
and U13404 (N_13404,N_5719,N_9914);
or U13405 (N_13405,N_9603,N_9029);
or U13406 (N_13406,N_8202,N_7075);
or U13407 (N_13407,N_5639,N_9497);
nand U13408 (N_13408,N_7731,N_6851);
or U13409 (N_13409,N_9919,N_9835);
nor U13410 (N_13410,N_9155,N_8561);
and U13411 (N_13411,N_9217,N_8591);
xor U13412 (N_13412,N_5728,N_6069);
and U13413 (N_13413,N_6429,N_8853);
nor U13414 (N_13414,N_8748,N_9360);
nand U13415 (N_13415,N_6422,N_9459);
nand U13416 (N_13416,N_5978,N_8768);
xor U13417 (N_13417,N_7866,N_5463);
nand U13418 (N_13418,N_9052,N_5373);
xnor U13419 (N_13419,N_5331,N_7185);
or U13420 (N_13420,N_7098,N_9303);
nand U13421 (N_13421,N_7626,N_6702);
and U13422 (N_13422,N_6150,N_6550);
and U13423 (N_13423,N_9876,N_8483);
or U13424 (N_13424,N_5055,N_7504);
nand U13425 (N_13425,N_5517,N_7200);
and U13426 (N_13426,N_7065,N_8471);
nor U13427 (N_13427,N_9515,N_9032);
nor U13428 (N_13428,N_8226,N_5676);
nand U13429 (N_13429,N_6931,N_7998);
nor U13430 (N_13430,N_6468,N_5168);
xor U13431 (N_13431,N_8301,N_5287);
nand U13432 (N_13432,N_7556,N_9204);
or U13433 (N_13433,N_7258,N_7017);
xor U13434 (N_13434,N_7499,N_9315);
nand U13435 (N_13435,N_7701,N_5450);
nor U13436 (N_13436,N_8267,N_9490);
nor U13437 (N_13437,N_7077,N_8257);
and U13438 (N_13438,N_5438,N_8598);
nor U13439 (N_13439,N_5243,N_7007);
xor U13440 (N_13440,N_7362,N_6892);
nor U13441 (N_13441,N_9562,N_7440);
nand U13442 (N_13442,N_5145,N_8812);
nor U13443 (N_13443,N_9838,N_8237);
nand U13444 (N_13444,N_8217,N_5971);
nor U13445 (N_13445,N_9664,N_5597);
or U13446 (N_13446,N_8599,N_8359);
nand U13447 (N_13447,N_7153,N_8629);
nand U13448 (N_13448,N_7274,N_7862);
nand U13449 (N_13449,N_5505,N_9090);
nor U13450 (N_13450,N_5369,N_9092);
nor U13451 (N_13451,N_9988,N_5152);
nand U13452 (N_13452,N_6177,N_5884);
and U13453 (N_13453,N_5502,N_7616);
nor U13454 (N_13454,N_8026,N_5651);
nand U13455 (N_13455,N_5669,N_5087);
or U13456 (N_13456,N_8388,N_6182);
and U13457 (N_13457,N_8162,N_7474);
xor U13458 (N_13458,N_8262,N_6014);
xnor U13459 (N_13459,N_6950,N_6553);
and U13460 (N_13460,N_5577,N_8062);
nor U13461 (N_13461,N_8470,N_5067);
nand U13462 (N_13462,N_8554,N_5500);
and U13463 (N_13463,N_6642,N_8443);
and U13464 (N_13464,N_8263,N_7491);
nor U13465 (N_13465,N_6779,N_7738);
xor U13466 (N_13466,N_6473,N_7680);
nor U13467 (N_13467,N_6075,N_8992);
or U13468 (N_13468,N_8924,N_8219);
xor U13469 (N_13469,N_6173,N_7056);
xor U13470 (N_13470,N_7328,N_7203);
or U13471 (N_13471,N_8739,N_7133);
nor U13472 (N_13472,N_9949,N_9063);
or U13473 (N_13473,N_9024,N_5951);
nand U13474 (N_13474,N_7120,N_7799);
or U13475 (N_13475,N_9692,N_6307);
nor U13476 (N_13476,N_6516,N_7170);
nand U13477 (N_13477,N_7041,N_7335);
and U13478 (N_13478,N_7853,N_9450);
nand U13479 (N_13479,N_9949,N_8551);
nand U13480 (N_13480,N_7066,N_5092);
xor U13481 (N_13481,N_5135,N_7781);
or U13482 (N_13482,N_8882,N_7267);
xnor U13483 (N_13483,N_7324,N_7716);
xor U13484 (N_13484,N_9149,N_8367);
nand U13485 (N_13485,N_7239,N_5391);
and U13486 (N_13486,N_9061,N_5150);
and U13487 (N_13487,N_8973,N_9227);
and U13488 (N_13488,N_8783,N_5791);
or U13489 (N_13489,N_6961,N_9142);
and U13490 (N_13490,N_7368,N_7888);
xor U13491 (N_13491,N_6334,N_5308);
nor U13492 (N_13492,N_7987,N_7233);
or U13493 (N_13493,N_5809,N_7737);
xnor U13494 (N_13494,N_8134,N_6072);
and U13495 (N_13495,N_5830,N_5594);
or U13496 (N_13496,N_8715,N_9892);
xor U13497 (N_13497,N_6853,N_9869);
nor U13498 (N_13498,N_9627,N_6826);
and U13499 (N_13499,N_9754,N_5801);
xor U13500 (N_13500,N_5949,N_6779);
nor U13501 (N_13501,N_6778,N_8887);
nand U13502 (N_13502,N_9765,N_5174);
nand U13503 (N_13503,N_5005,N_7523);
xnor U13504 (N_13504,N_9760,N_6976);
or U13505 (N_13505,N_9259,N_5099);
nor U13506 (N_13506,N_6563,N_9967);
nor U13507 (N_13507,N_7917,N_5092);
nor U13508 (N_13508,N_6486,N_9619);
xor U13509 (N_13509,N_5352,N_9420);
and U13510 (N_13510,N_8952,N_7645);
or U13511 (N_13511,N_9032,N_7407);
or U13512 (N_13512,N_9449,N_9381);
nor U13513 (N_13513,N_5039,N_9834);
and U13514 (N_13514,N_8454,N_6010);
or U13515 (N_13515,N_7895,N_5906);
or U13516 (N_13516,N_8022,N_7926);
or U13517 (N_13517,N_6761,N_7254);
nand U13518 (N_13518,N_7226,N_5164);
or U13519 (N_13519,N_6350,N_6332);
nand U13520 (N_13520,N_9328,N_8077);
and U13521 (N_13521,N_8725,N_9310);
or U13522 (N_13522,N_5464,N_5391);
nand U13523 (N_13523,N_9802,N_6077);
nor U13524 (N_13524,N_9218,N_9759);
nor U13525 (N_13525,N_9168,N_7654);
and U13526 (N_13526,N_9882,N_6926);
and U13527 (N_13527,N_9058,N_6710);
and U13528 (N_13528,N_5423,N_6219);
xor U13529 (N_13529,N_6705,N_6523);
nand U13530 (N_13530,N_5386,N_6027);
nand U13531 (N_13531,N_9881,N_9000);
nand U13532 (N_13532,N_6527,N_9045);
xor U13533 (N_13533,N_7665,N_6461);
nor U13534 (N_13534,N_8832,N_8667);
xor U13535 (N_13535,N_5629,N_9615);
nor U13536 (N_13536,N_8050,N_7344);
nor U13537 (N_13537,N_6755,N_6872);
or U13538 (N_13538,N_6950,N_8662);
xnor U13539 (N_13539,N_7893,N_9657);
or U13540 (N_13540,N_5029,N_5172);
nand U13541 (N_13541,N_8905,N_8195);
xor U13542 (N_13542,N_6728,N_8455);
xnor U13543 (N_13543,N_5538,N_9890);
xor U13544 (N_13544,N_6370,N_9473);
nor U13545 (N_13545,N_6418,N_5638);
nand U13546 (N_13546,N_8816,N_8567);
nand U13547 (N_13547,N_8628,N_9892);
xnor U13548 (N_13548,N_7863,N_9232);
nor U13549 (N_13549,N_6530,N_9014);
and U13550 (N_13550,N_6084,N_7578);
xor U13551 (N_13551,N_5056,N_5136);
nor U13552 (N_13552,N_7450,N_6698);
or U13553 (N_13553,N_5881,N_8929);
xor U13554 (N_13554,N_7446,N_8434);
and U13555 (N_13555,N_8332,N_8278);
nor U13556 (N_13556,N_8067,N_9840);
nor U13557 (N_13557,N_9262,N_5081);
and U13558 (N_13558,N_9354,N_6547);
or U13559 (N_13559,N_5792,N_7793);
and U13560 (N_13560,N_6955,N_5007);
or U13561 (N_13561,N_6906,N_9407);
nand U13562 (N_13562,N_9781,N_6896);
nor U13563 (N_13563,N_8633,N_9484);
nand U13564 (N_13564,N_6681,N_9097);
and U13565 (N_13565,N_8879,N_5504);
nor U13566 (N_13566,N_5042,N_8136);
nor U13567 (N_13567,N_6705,N_8183);
and U13568 (N_13568,N_5136,N_6875);
nand U13569 (N_13569,N_6184,N_5088);
and U13570 (N_13570,N_9810,N_7217);
and U13571 (N_13571,N_7522,N_5518);
nor U13572 (N_13572,N_8088,N_8876);
xnor U13573 (N_13573,N_9008,N_9444);
and U13574 (N_13574,N_7633,N_8971);
or U13575 (N_13575,N_8310,N_8468);
and U13576 (N_13576,N_5816,N_9727);
nand U13577 (N_13577,N_9781,N_5067);
nand U13578 (N_13578,N_8518,N_8695);
or U13579 (N_13579,N_9248,N_5825);
xnor U13580 (N_13580,N_6903,N_6181);
and U13581 (N_13581,N_5450,N_6897);
nor U13582 (N_13582,N_5271,N_6635);
nand U13583 (N_13583,N_7474,N_7020);
or U13584 (N_13584,N_7738,N_8736);
and U13585 (N_13585,N_6664,N_5953);
xnor U13586 (N_13586,N_8855,N_8658);
nor U13587 (N_13587,N_9951,N_8715);
nand U13588 (N_13588,N_6405,N_9896);
nand U13589 (N_13589,N_6736,N_8184);
nor U13590 (N_13590,N_7342,N_8910);
nand U13591 (N_13591,N_7968,N_7667);
nand U13592 (N_13592,N_9610,N_8314);
and U13593 (N_13593,N_8164,N_5573);
or U13594 (N_13594,N_5543,N_9830);
nor U13595 (N_13595,N_7409,N_9791);
xnor U13596 (N_13596,N_8642,N_8543);
and U13597 (N_13597,N_9556,N_9061);
and U13598 (N_13598,N_7195,N_8775);
or U13599 (N_13599,N_6861,N_9361);
nor U13600 (N_13600,N_6973,N_5965);
nand U13601 (N_13601,N_7964,N_6370);
nand U13602 (N_13602,N_5154,N_7692);
nor U13603 (N_13603,N_6320,N_9605);
xor U13604 (N_13604,N_6787,N_9442);
nor U13605 (N_13605,N_8435,N_7740);
or U13606 (N_13606,N_8060,N_5118);
nand U13607 (N_13607,N_6210,N_9028);
xnor U13608 (N_13608,N_5038,N_5856);
nor U13609 (N_13609,N_9373,N_5194);
nor U13610 (N_13610,N_8176,N_6145);
or U13611 (N_13611,N_6218,N_5625);
or U13612 (N_13612,N_5498,N_6645);
and U13613 (N_13613,N_9485,N_7904);
nor U13614 (N_13614,N_9833,N_8589);
nor U13615 (N_13615,N_6561,N_8728);
and U13616 (N_13616,N_6753,N_5560);
and U13617 (N_13617,N_5637,N_7726);
and U13618 (N_13618,N_9998,N_5116);
nand U13619 (N_13619,N_9431,N_5906);
xnor U13620 (N_13620,N_5284,N_7994);
xor U13621 (N_13621,N_5542,N_7031);
or U13622 (N_13622,N_7150,N_6932);
nand U13623 (N_13623,N_9045,N_5788);
nand U13624 (N_13624,N_7139,N_5036);
and U13625 (N_13625,N_8234,N_8117);
xnor U13626 (N_13626,N_5477,N_6709);
nor U13627 (N_13627,N_6952,N_6677);
and U13628 (N_13628,N_5136,N_7347);
or U13629 (N_13629,N_6112,N_8954);
xnor U13630 (N_13630,N_6613,N_7330);
or U13631 (N_13631,N_9805,N_9371);
xor U13632 (N_13632,N_8296,N_7177);
and U13633 (N_13633,N_7129,N_6925);
or U13634 (N_13634,N_7887,N_7950);
nand U13635 (N_13635,N_7447,N_5365);
and U13636 (N_13636,N_5941,N_5304);
or U13637 (N_13637,N_9814,N_8859);
nand U13638 (N_13638,N_9438,N_9432);
nand U13639 (N_13639,N_8346,N_5925);
or U13640 (N_13640,N_8381,N_7500);
nand U13641 (N_13641,N_8946,N_6698);
nand U13642 (N_13642,N_5501,N_6874);
nand U13643 (N_13643,N_8285,N_5979);
and U13644 (N_13644,N_6855,N_6951);
nor U13645 (N_13645,N_5741,N_7031);
xnor U13646 (N_13646,N_6687,N_9628);
xnor U13647 (N_13647,N_7297,N_9787);
and U13648 (N_13648,N_9060,N_6991);
nand U13649 (N_13649,N_8463,N_5828);
and U13650 (N_13650,N_6984,N_9194);
or U13651 (N_13651,N_7174,N_5394);
nand U13652 (N_13652,N_6382,N_7404);
xnor U13653 (N_13653,N_6435,N_8142);
and U13654 (N_13654,N_6806,N_9571);
and U13655 (N_13655,N_6978,N_9497);
and U13656 (N_13656,N_5117,N_7182);
xor U13657 (N_13657,N_5895,N_5823);
or U13658 (N_13658,N_8330,N_5960);
xnor U13659 (N_13659,N_8203,N_6582);
nor U13660 (N_13660,N_8386,N_5207);
xnor U13661 (N_13661,N_5652,N_6678);
and U13662 (N_13662,N_6980,N_5565);
or U13663 (N_13663,N_7097,N_7796);
or U13664 (N_13664,N_9827,N_9146);
nand U13665 (N_13665,N_6108,N_7501);
and U13666 (N_13666,N_7942,N_7971);
nand U13667 (N_13667,N_5979,N_8147);
nor U13668 (N_13668,N_7844,N_5406);
nand U13669 (N_13669,N_6074,N_9182);
nand U13670 (N_13670,N_6676,N_6897);
nor U13671 (N_13671,N_6102,N_5697);
nand U13672 (N_13672,N_7347,N_6010);
and U13673 (N_13673,N_7354,N_7356);
nor U13674 (N_13674,N_9223,N_5832);
or U13675 (N_13675,N_8772,N_8863);
and U13676 (N_13676,N_6688,N_8413);
or U13677 (N_13677,N_5090,N_9732);
or U13678 (N_13678,N_9139,N_8411);
nand U13679 (N_13679,N_6029,N_6280);
or U13680 (N_13680,N_7992,N_7706);
nor U13681 (N_13681,N_7029,N_5954);
or U13682 (N_13682,N_9334,N_9191);
nor U13683 (N_13683,N_5814,N_9765);
or U13684 (N_13684,N_5470,N_8348);
or U13685 (N_13685,N_6242,N_6814);
or U13686 (N_13686,N_7195,N_8272);
xnor U13687 (N_13687,N_9762,N_9038);
and U13688 (N_13688,N_8648,N_8790);
nor U13689 (N_13689,N_9897,N_5912);
nor U13690 (N_13690,N_9858,N_7186);
nand U13691 (N_13691,N_6465,N_9923);
or U13692 (N_13692,N_8383,N_6899);
nor U13693 (N_13693,N_5384,N_8501);
nor U13694 (N_13694,N_5158,N_7043);
nor U13695 (N_13695,N_5897,N_7525);
nand U13696 (N_13696,N_6994,N_8947);
nor U13697 (N_13697,N_9026,N_8530);
xor U13698 (N_13698,N_5638,N_8876);
or U13699 (N_13699,N_9156,N_5817);
and U13700 (N_13700,N_7222,N_5085);
or U13701 (N_13701,N_8052,N_6343);
nor U13702 (N_13702,N_8014,N_9954);
nor U13703 (N_13703,N_7586,N_9260);
or U13704 (N_13704,N_6540,N_8676);
and U13705 (N_13705,N_6603,N_5471);
xor U13706 (N_13706,N_8953,N_8070);
nand U13707 (N_13707,N_5877,N_7811);
nand U13708 (N_13708,N_7271,N_6695);
or U13709 (N_13709,N_9685,N_5116);
or U13710 (N_13710,N_7831,N_7154);
or U13711 (N_13711,N_7486,N_7754);
xnor U13712 (N_13712,N_5727,N_9619);
and U13713 (N_13713,N_5859,N_9246);
and U13714 (N_13714,N_9374,N_6596);
and U13715 (N_13715,N_7900,N_7337);
nor U13716 (N_13716,N_8915,N_6296);
xnor U13717 (N_13717,N_7260,N_9795);
xnor U13718 (N_13718,N_9527,N_8934);
nand U13719 (N_13719,N_6652,N_8385);
xor U13720 (N_13720,N_5524,N_8331);
and U13721 (N_13721,N_5681,N_5286);
xor U13722 (N_13722,N_9413,N_6953);
nand U13723 (N_13723,N_6671,N_7793);
or U13724 (N_13724,N_5676,N_8899);
nand U13725 (N_13725,N_9000,N_6648);
nor U13726 (N_13726,N_5961,N_5805);
or U13727 (N_13727,N_5654,N_5027);
nor U13728 (N_13728,N_8215,N_5865);
or U13729 (N_13729,N_6848,N_9908);
nand U13730 (N_13730,N_9736,N_7041);
or U13731 (N_13731,N_7335,N_9485);
or U13732 (N_13732,N_6645,N_8479);
or U13733 (N_13733,N_8629,N_7426);
nand U13734 (N_13734,N_5759,N_9458);
and U13735 (N_13735,N_5948,N_7787);
xor U13736 (N_13736,N_8263,N_5949);
xor U13737 (N_13737,N_5002,N_6606);
xnor U13738 (N_13738,N_6439,N_9929);
xnor U13739 (N_13739,N_5308,N_5751);
or U13740 (N_13740,N_8384,N_5004);
nor U13741 (N_13741,N_5192,N_7325);
xnor U13742 (N_13742,N_9911,N_8294);
nand U13743 (N_13743,N_9421,N_6032);
or U13744 (N_13744,N_9898,N_8885);
nand U13745 (N_13745,N_8616,N_6190);
nor U13746 (N_13746,N_9470,N_6308);
nor U13747 (N_13747,N_8556,N_6454);
nand U13748 (N_13748,N_6017,N_9608);
or U13749 (N_13749,N_9400,N_8903);
nor U13750 (N_13750,N_6531,N_8768);
xnor U13751 (N_13751,N_9089,N_8081);
xnor U13752 (N_13752,N_7413,N_5235);
or U13753 (N_13753,N_9492,N_5197);
xor U13754 (N_13754,N_7499,N_9165);
nor U13755 (N_13755,N_7310,N_5491);
and U13756 (N_13756,N_9949,N_9373);
xor U13757 (N_13757,N_8450,N_6826);
xor U13758 (N_13758,N_7717,N_6496);
nand U13759 (N_13759,N_8398,N_6700);
nand U13760 (N_13760,N_8114,N_9609);
nand U13761 (N_13761,N_8706,N_7530);
xor U13762 (N_13762,N_7031,N_7072);
xor U13763 (N_13763,N_5377,N_9187);
or U13764 (N_13764,N_9693,N_6140);
or U13765 (N_13765,N_9964,N_9254);
and U13766 (N_13766,N_7062,N_6945);
nor U13767 (N_13767,N_6643,N_9924);
and U13768 (N_13768,N_5848,N_9863);
or U13769 (N_13769,N_6545,N_7083);
xnor U13770 (N_13770,N_8322,N_5494);
and U13771 (N_13771,N_9256,N_7545);
xnor U13772 (N_13772,N_8353,N_6424);
nor U13773 (N_13773,N_8293,N_5478);
nand U13774 (N_13774,N_8703,N_6023);
nand U13775 (N_13775,N_8036,N_9353);
or U13776 (N_13776,N_5043,N_8788);
xnor U13777 (N_13777,N_9866,N_8226);
and U13778 (N_13778,N_6227,N_5502);
nor U13779 (N_13779,N_7043,N_5635);
or U13780 (N_13780,N_8797,N_6460);
or U13781 (N_13781,N_7762,N_6512);
or U13782 (N_13782,N_8134,N_8410);
nor U13783 (N_13783,N_6991,N_6762);
or U13784 (N_13784,N_5066,N_8033);
nand U13785 (N_13785,N_6353,N_6970);
nand U13786 (N_13786,N_9682,N_8721);
nand U13787 (N_13787,N_8509,N_8242);
xor U13788 (N_13788,N_7345,N_9076);
or U13789 (N_13789,N_5562,N_5498);
nand U13790 (N_13790,N_6035,N_8446);
xnor U13791 (N_13791,N_9392,N_7497);
and U13792 (N_13792,N_6660,N_6012);
nor U13793 (N_13793,N_8325,N_7571);
or U13794 (N_13794,N_9602,N_7848);
and U13795 (N_13795,N_8070,N_5662);
nand U13796 (N_13796,N_6083,N_5265);
nand U13797 (N_13797,N_5584,N_8543);
and U13798 (N_13798,N_7035,N_8111);
nor U13799 (N_13799,N_9993,N_8954);
or U13800 (N_13800,N_6133,N_7222);
nor U13801 (N_13801,N_8271,N_5635);
xor U13802 (N_13802,N_7006,N_7760);
or U13803 (N_13803,N_5777,N_9108);
nor U13804 (N_13804,N_6535,N_7135);
nand U13805 (N_13805,N_6277,N_8991);
or U13806 (N_13806,N_9922,N_5086);
xnor U13807 (N_13807,N_6606,N_9363);
nand U13808 (N_13808,N_5694,N_9202);
or U13809 (N_13809,N_7698,N_9775);
nand U13810 (N_13810,N_7925,N_5274);
nand U13811 (N_13811,N_6167,N_9323);
xor U13812 (N_13812,N_9202,N_9472);
nand U13813 (N_13813,N_6573,N_5492);
or U13814 (N_13814,N_8224,N_6039);
and U13815 (N_13815,N_5472,N_5685);
nor U13816 (N_13816,N_7110,N_5623);
xnor U13817 (N_13817,N_7202,N_7203);
and U13818 (N_13818,N_5080,N_6721);
or U13819 (N_13819,N_9885,N_6962);
xor U13820 (N_13820,N_9410,N_6749);
xnor U13821 (N_13821,N_7359,N_9756);
or U13822 (N_13822,N_5822,N_5023);
nor U13823 (N_13823,N_8033,N_7801);
and U13824 (N_13824,N_9590,N_6910);
or U13825 (N_13825,N_5137,N_5800);
nand U13826 (N_13826,N_6639,N_6079);
or U13827 (N_13827,N_5631,N_5858);
xor U13828 (N_13828,N_8250,N_6246);
xor U13829 (N_13829,N_7414,N_7059);
and U13830 (N_13830,N_6074,N_5939);
xnor U13831 (N_13831,N_7079,N_7224);
xnor U13832 (N_13832,N_6771,N_6437);
or U13833 (N_13833,N_7862,N_7575);
or U13834 (N_13834,N_5503,N_7253);
xor U13835 (N_13835,N_5122,N_5704);
and U13836 (N_13836,N_8050,N_6276);
nor U13837 (N_13837,N_8379,N_7369);
nand U13838 (N_13838,N_8188,N_6412);
xor U13839 (N_13839,N_5625,N_9779);
nor U13840 (N_13840,N_5816,N_9366);
nor U13841 (N_13841,N_7930,N_6023);
or U13842 (N_13842,N_6319,N_9771);
and U13843 (N_13843,N_5413,N_9417);
nor U13844 (N_13844,N_6076,N_5753);
nand U13845 (N_13845,N_8177,N_6931);
and U13846 (N_13846,N_6158,N_8766);
xnor U13847 (N_13847,N_9863,N_7341);
nand U13848 (N_13848,N_5999,N_9320);
or U13849 (N_13849,N_7237,N_7752);
or U13850 (N_13850,N_5702,N_5568);
or U13851 (N_13851,N_9071,N_7848);
and U13852 (N_13852,N_5435,N_9547);
or U13853 (N_13853,N_5760,N_8326);
and U13854 (N_13854,N_7739,N_7182);
nand U13855 (N_13855,N_5107,N_9480);
and U13856 (N_13856,N_5228,N_7891);
nor U13857 (N_13857,N_6562,N_6252);
nor U13858 (N_13858,N_9770,N_8394);
or U13859 (N_13859,N_9515,N_7645);
xor U13860 (N_13860,N_8561,N_8057);
or U13861 (N_13861,N_6244,N_8157);
xor U13862 (N_13862,N_5114,N_6769);
nand U13863 (N_13863,N_5256,N_6314);
nand U13864 (N_13864,N_7717,N_7214);
nand U13865 (N_13865,N_8800,N_8650);
nor U13866 (N_13866,N_8782,N_6165);
xnor U13867 (N_13867,N_7488,N_7972);
nor U13868 (N_13868,N_6977,N_8065);
or U13869 (N_13869,N_9723,N_7860);
nor U13870 (N_13870,N_8679,N_5598);
and U13871 (N_13871,N_6729,N_9318);
nand U13872 (N_13872,N_9857,N_9257);
or U13873 (N_13873,N_6631,N_6443);
nor U13874 (N_13874,N_9194,N_6554);
nor U13875 (N_13875,N_7940,N_8042);
or U13876 (N_13876,N_5464,N_9358);
nor U13877 (N_13877,N_8250,N_7387);
or U13878 (N_13878,N_6252,N_8796);
and U13879 (N_13879,N_5535,N_6636);
nand U13880 (N_13880,N_7084,N_6834);
and U13881 (N_13881,N_9056,N_6491);
nor U13882 (N_13882,N_6985,N_5168);
nand U13883 (N_13883,N_7894,N_8363);
nand U13884 (N_13884,N_8335,N_8095);
nand U13885 (N_13885,N_5110,N_6168);
nand U13886 (N_13886,N_9740,N_8141);
or U13887 (N_13887,N_6681,N_6342);
or U13888 (N_13888,N_6727,N_5229);
nor U13889 (N_13889,N_8866,N_9199);
nor U13890 (N_13890,N_9810,N_6642);
and U13891 (N_13891,N_8204,N_9668);
xor U13892 (N_13892,N_6567,N_6412);
or U13893 (N_13893,N_6652,N_6975);
nor U13894 (N_13894,N_8091,N_5645);
or U13895 (N_13895,N_6517,N_5718);
xor U13896 (N_13896,N_5929,N_9469);
nor U13897 (N_13897,N_9011,N_6879);
or U13898 (N_13898,N_8849,N_5394);
and U13899 (N_13899,N_6259,N_6454);
xor U13900 (N_13900,N_7975,N_8401);
and U13901 (N_13901,N_5087,N_7395);
and U13902 (N_13902,N_8171,N_7265);
xnor U13903 (N_13903,N_7946,N_7481);
nand U13904 (N_13904,N_7949,N_8594);
nor U13905 (N_13905,N_9317,N_5760);
nand U13906 (N_13906,N_5483,N_7884);
and U13907 (N_13907,N_5971,N_5347);
or U13908 (N_13908,N_7644,N_9443);
nand U13909 (N_13909,N_9674,N_5278);
xor U13910 (N_13910,N_6849,N_9573);
nand U13911 (N_13911,N_7376,N_8827);
nand U13912 (N_13912,N_8807,N_7658);
xnor U13913 (N_13913,N_9924,N_7894);
xnor U13914 (N_13914,N_8649,N_6138);
nor U13915 (N_13915,N_9278,N_5159);
nor U13916 (N_13916,N_8931,N_5498);
or U13917 (N_13917,N_5433,N_8336);
nand U13918 (N_13918,N_7627,N_5574);
nor U13919 (N_13919,N_8810,N_8062);
and U13920 (N_13920,N_8614,N_6009);
nor U13921 (N_13921,N_8069,N_6123);
and U13922 (N_13922,N_8864,N_7854);
and U13923 (N_13923,N_5106,N_8564);
xor U13924 (N_13924,N_8671,N_7869);
xnor U13925 (N_13925,N_9443,N_9128);
and U13926 (N_13926,N_6264,N_6299);
nor U13927 (N_13927,N_9641,N_8062);
and U13928 (N_13928,N_6569,N_8711);
and U13929 (N_13929,N_6719,N_5181);
or U13930 (N_13930,N_6840,N_5125);
nor U13931 (N_13931,N_9275,N_7180);
or U13932 (N_13932,N_5796,N_6256);
or U13933 (N_13933,N_7640,N_8080);
and U13934 (N_13934,N_8420,N_5803);
xor U13935 (N_13935,N_8111,N_9091);
and U13936 (N_13936,N_7688,N_5296);
and U13937 (N_13937,N_7193,N_5529);
or U13938 (N_13938,N_6166,N_6295);
and U13939 (N_13939,N_6663,N_5991);
xor U13940 (N_13940,N_6718,N_6111);
nor U13941 (N_13941,N_7428,N_6588);
nor U13942 (N_13942,N_6418,N_5161);
xor U13943 (N_13943,N_6187,N_6763);
nor U13944 (N_13944,N_9267,N_7464);
nor U13945 (N_13945,N_9038,N_6149);
nor U13946 (N_13946,N_7101,N_9184);
or U13947 (N_13947,N_5454,N_9587);
nand U13948 (N_13948,N_9836,N_9145);
xor U13949 (N_13949,N_5685,N_9826);
xnor U13950 (N_13950,N_5074,N_8152);
nand U13951 (N_13951,N_5708,N_8942);
and U13952 (N_13952,N_9970,N_9023);
and U13953 (N_13953,N_9215,N_9840);
nor U13954 (N_13954,N_5388,N_5588);
nand U13955 (N_13955,N_6428,N_6572);
nand U13956 (N_13956,N_7754,N_7847);
nor U13957 (N_13957,N_6290,N_9691);
and U13958 (N_13958,N_6946,N_8790);
xnor U13959 (N_13959,N_9911,N_5998);
nand U13960 (N_13960,N_5134,N_9897);
or U13961 (N_13961,N_9769,N_5982);
nand U13962 (N_13962,N_5359,N_8040);
xor U13963 (N_13963,N_5924,N_7587);
or U13964 (N_13964,N_8830,N_7839);
nand U13965 (N_13965,N_7807,N_9077);
or U13966 (N_13966,N_9216,N_9488);
and U13967 (N_13967,N_6239,N_5449);
xnor U13968 (N_13968,N_5070,N_7953);
or U13969 (N_13969,N_8603,N_7780);
or U13970 (N_13970,N_5741,N_8449);
or U13971 (N_13971,N_9102,N_8291);
xor U13972 (N_13972,N_5266,N_5230);
xor U13973 (N_13973,N_9131,N_9702);
nand U13974 (N_13974,N_8231,N_6938);
nor U13975 (N_13975,N_6151,N_6212);
xor U13976 (N_13976,N_8928,N_9877);
or U13977 (N_13977,N_6626,N_7107);
or U13978 (N_13978,N_9844,N_6587);
or U13979 (N_13979,N_5890,N_6762);
nor U13980 (N_13980,N_7206,N_9976);
nor U13981 (N_13981,N_8514,N_7070);
xor U13982 (N_13982,N_5338,N_6597);
or U13983 (N_13983,N_7274,N_7893);
or U13984 (N_13984,N_8376,N_9949);
and U13985 (N_13985,N_8047,N_6181);
or U13986 (N_13986,N_8956,N_9492);
nor U13987 (N_13987,N_7043,N_9785);
and U13988 (N_13988,N_6337,N_5632);
nor U13989 (N_13989,N_8341,N_9446);
nand U13990 (N_13990,N_5708,N_5050);
or U13991 (N_13991,N_5406,N_6115);
xor U13992 (N_13992,N_8324,N_7053);
or U13993 (N_13993,N_7611,N_9131);
nand U13994 (N_13994,N_7969,N_6352);
or U13995 (N_13995,N_6298,N_9625);
nor U13996 (N_13996,N_9052,N_6188);
nand U13997 (N_13997,N_7118,N_6176);
xnor U13998 (N_13998,N_7264,N_5775);
xor U13999 (N_13999,N_8649,N_8071);
xnor U14000 (N_14000,N_6101,N_8826);
nor U14001 (N_14001,N_7216,N_8595);
nand U14002 (N_14002,N_5912,N_9870);
or U14003 (N_14003,N_6111,N_9589);
or U14004 (N_14004,N_9113,N_5363);
xor U14005 (N_14005,N_8397,N_9781);
or U14006 (N_14006,N_9676,N_9318);
nand U14007 (N_14007,N_6459,N_8692);
and U14008 (N_14008,N_9560,N_6615);
and U14009 (N_14009,N_6291,N_5675);
and U14010 (N_14010,N_5374,N_6729);
xnor U14011 (N_14011,N_9407,N_8054);
or U14012 (N_14012,N_6921,N_5690);
nor U14013 (N_14013,N_8946,N_5049);
nor U14014 (N_14014,N_6055,N_9782);
nand U14015 (N_14015,N_9781,N_8129);
xnor U14016 (N_14016,N_7445,N_9117);
nand U14017 (N_14017,N_9064,N_8870);
nand U14018 (N_14018,N_7247,N_7177);
nand U14019 (N_14019,N_8280,N_9934);
nor U14020 (N_14020,N_8581,N_7275);
nor U14021 (N_14021,N_8209,N_8775);
xnor U14022 (N_14022,N_5480,N_5523);
and U14023 (N_14023,N_8327,N_8817);
and U14024 (N_14024,N_8050,N_6367);
xor U14025 (N_14025,N_6058,N_9617);
nor U14026 (N_14026,N_7258,N_7716);
xnor U14027 (N_14027,N_6230,N_7033);
nor U14028 (N_14028,N_6683,N_6122);
nor U14029 (N_14029,N_7032,N_9099);
nor U14030 (N_14030,N_8106,N_8456);
nand U14031 (N_14031,N_7035,N_5587);
and U14032 (N_14032,N_8966,N_7212);
nand U14033 (N_14033,N_6662,N_6236);
or U14034 (N_14034,N_8313,N_9806);
or U14035 (N_14035,N_7786,N_6631);
and U14036 (N_14036,N_8908,N_5399);
or U14037 (N_14037,N_7214,N_6247);
or U14038 (N_14038,N_8273,N_5834);
xor U14039 (N_14039,N_8381,N_9345);
xnor U14040 (N_14040,N_5581,N_5481);
and U14041 (N_14041,N_7396,N_9674);
nand U14042 (N_14042,N_9077,N_8243);
and U14043 (N_14043,N_7660,N_9857);
nand U14044 (N_14044,N_9279,N_7750);
nand U14045 (N_14045,N_9674,N_6154);
nand U14046 (N_14046,N_9148,N_5770);
xor U14047 (N_14047,N_7748,N_6021);
nor U14048 (N_14048,N_9490,N_5666);
nor U14049 (N_14049,N_7965,N_7834);
and U14050 (N_14050,N_8395,N_7224);
or U14051 (N_14051,N_7588,N_6568);
and U14052 (N_14052,N_6418,N_5605);
or U14053 (N_14053,N_5990,N_5904);
nor U14054 (N_14054,N_9628,N_9417);
and U14055 (N_14055,N_9623,N_8981);
nand U14056 (N_14056,N_7149,N_6914);
nor U14057 (N_14057,N_9817,N_9184);
xnor U14058 (N_14058,N_7173,N_5275);
nor U14059 (N_14059,N_6502,N_5712);
nand U14060 (N_14060,N_9921,N_8720);
nor U14061 (N_14061,N_8860,N_9802);
nand U14062 (N_14062,N_5992,N_8423);
nand U14063 (N_14063,N_9244,N_7784);
xnor U14064 (N_14064,N_9569,N_6790);
nor U14065 (N_14065,N_8431,N_6283);
xor U14066 (N_14066,N_5340,N_6159);
and U14067 (N_14067,N_8630,N_5468);
xor U14068 (N_14068,N_5939,N_7517);
xor U14069 (N_14069,N_8545,N_8724);
nor U14070 (N_14070,N_6131,N_6335);
xnor U14071 (N_14071,N_6391,N_5211);
nor U14072 (N_14072,N_8260,N_5532);
nor U14073 (N_14073,N_8072,N_5778);
nand U14074 (N_14074,N_8017,N_6305);
or U14075 (N_14075,N_9345,N_8281);
xor U14076 (N_14076,N_5194,N_9184);
nand U14077 (N_14077,N_9388,N_9389);
xor U14078 (N_14078,N_9997,N_8586);
and U14079 (N_14079,N_7645,N_5369);
and U14080 (N_14080,N_7403,N_6120);
or U14081 (N_14081,N_8425,N_8683);
nor U14082 (N_14082,N_6354,N_6536);
nor U14083 (N_14083,N_5298,N_8464);
nand U14084 (N_14084,N_6657,N_7511);
nand U14085 (N_14085,N_7001,N_8674);
xor U14086 (N_14086,N_8338,N_5277);
or U14087 (N_14087,N_7475,N_8428);
nor U14088 (N_14088,N_9949,N_7060);
nand U14089 (N_14089,N_6046,N_5001);
or U14090 (N_14090,N_9942,N_9919);
or U14091 (N_14091,N_8975,N_9598);
nand U14092 (N_14092,N_8877,N_7867);
or U14093 (N_14093,N_5192,N_7014);
xnor U14094 (N_14094,N_8286,N_7762);
nand U14095 (N_14095,N_8304,N_6698);
nor U14096 (N_14096,N_6641,N_5984);
xor U14097 (N_14097,N_9282,N_8204);
and U14098 (N_14098,N_5020,N_9158);
nand U14099 (N_14099,N_9799,N_7907);
nand U14100 (N_14100,N_9492,N_9988);
nand U14101 (N_14101,N_7684,N_9466);
nor U14102 (N_14102,N_8793,N_5295);
and U14103 (N_14103,N_7174,N_5417);
xnor U14104 (N_14104,N_6904,N_9046);
nor U14105 (N_14105,N_8942,N_5879);
and U14106 (N_14106,N_6260,N_6499);
xnor U14107 (N_14107,N_6458,N_6545);
or U14108 (N_14108,N_8315,N_6231);
and U14109 (N_14109,N_5704,N_5877);
nand U14110 (N_14110,N_9635,N_6608);
or U14111 (N_14111,N_5969,N_7722);
xnor U14112 (N_14112,N_8956,N_5184);
or U14113 (N_14113,N_8699,N_7738);
or U14114 (N_14114,N_9836,N_7507);
nor U14115 (N_14115,N_9114,N_5243);
and U14116 (N_14116,N_5361,N_6795);
or U14117 (N_14117,N_8819,N_8512);
or U14118 (N_14118,N_8199,N_9003);
and U14119 (N_14119,N_5605,N_5593);
or U14120 (N_14120,N_9407,N_7178);
nor U14121 (N_14121,N_5117,N_8417);
nand U14122 (N_14122,N_8256,N_5803);
and U14123 (N_14123,N_8234,N_5549);
or U14124 (N_14124,N_7586,N_8477);
or U14125 (N_14125,N_6399,N_5870);
nand U14126 (N_14126,N_6559,N_8415);
or U14127 (N_14127,N_5316,N_5596);
nand U14128 (N_14128,N_6029,N_7982);
nand U14129 (N_14129,N_8051,N_9294);
nor U14130 (N_14130,N_9312,N_7797);
nor U14131 (N_14131,N_8921,N_8614);
xnor U14132 (N_14132,N_8531,N_9879);
nor U14133 (N_14133,N_7578,N_6167);
nand U14134 (N_14134,N_9466,N_7558);
or U14135 (N_14135,N_8825,N_5612);
nor U14136 (N_14136,N_8964,N_5518);
nor U14137 (N_14137,N_9305,N_6410);
or U14138 (N_14138,N_8978,N_6142);
and U14139 (N_14139,N_8014,N_6877);
xor U14140 (N_14140,N_5148,N_6863);
or U14141 (N_14141,N_7112,N_8901);
nand U14142 (N_14142,N_5561,N_6710);
or U14143 (N_14143,N_5641,N_5629);
and U14144 (N_14144,N_9437,N_7837);
xor U14145 (N_14145,N_8661,N_7290);
xnor U14146 (N_14146,N_9336,N_6054);
or U14147 (N_14147,N_9356,N_7180);
nand U14148 (N_14148,N_6991,N_7871);
or U14149 (N_14149,N_5210,N_7529);
or U14150 (N_14150,N_8635,N_9408);
xor U14151 (N_14151,N_5169,N_9894);
and U14152 (N_14152,N_6601,N_6830);
nand U14153 (N_14153,N_8460,N_6359);
and U14154 (N_14154,N_6631,N_7391);
and U14155 (N_14155,N_8268,N_6809);
and U14156 (N_14156,N_7279,N_6475);
xnor U14157 (N_14157,N_8384,N_9644);
nand U14158 (N_14158,N_6990,N_5993);
nor U14159 (N_14159,N_5810,N_6884);
and U14160 (N_14160,N_7639,N_5035);
and U14161 (N_14161,N_7198,N_8291);
nand U14162 (N_14162,N_5749,N_5661);
and U14163 (N_14163,N_8914,N_8422);
xor U14164 (N_14164,N_7611,N_7240);
nand U14165 (N_14165,N_7357,N_9477);
nand U14166 (N_14166,N_5717,N_9004);
or U14167 (N_14167,N_6201,N_8870);
nor U14168 (N_14168,N_7599,N_6786);
or U14169 (N_14169,N_9748,N_6850);
xnor U14170 (N_14170,N_9703,N_8189);
xor U14171 (N_14171,N_5741,N_9923);
nor U14172 (N_14172,N_6329,N_9149);
and U14173 (N_14173,N_9839,N_8417);
nand U14174 (N_14174,N_5818,N_9894);
xor U14175 (N_14175,N_6751,N_5758);
or U14176 (N_14176,N_9974,N_6950);
or U14177 (N_14177,N_6589,N_7093);
and U14178 (N_14178,N_6912,N_8500);
xnor U14179 (N_14179,N_8342,N_5946);
or U14180 (N_14180,N_7244,N_5762);
or U14181 (N_14181,N_5561,N_7464);
nor U14182 (N_14182,N_6931,N_5059);
nor U14183 (N_14183,N_9435,N_6146);
nor U14184 (N_14184,N_5622,N_8003);
xnor U14185 (N_14185,N_5972,N_7585);
xor U14186 (N_14186,N_9861,N_5859);
nand U14187 (N_14187,N_7546,N_8301);
and U14188 (N_14188,N_8172,N_9024);
or U14189 (N_14189,N_9682,N_7682);
nor U14190 (N_14190,N_8375,N_7766);
nor U14191 (N_14191,N_7252,N_5399);
and U14192 (N_14192,N_9889,N_6472);
xor U14193 (N_14193,N_5310,N_5988);
or U14194 (N_14194,N_5691,N_7937);
nand U14195 (N_14195,N_7199,N_9527);
nor U14196 (N_14196,N_8659,N_7795);
or U14197 (N_14197,N_9986,N_9116);
nand U14198 (N_14198,N_9410,N_8839);
nor U14199 (N_14199,N_6959,N_7764);
nor U14200 (N_14200,N_8835,N_5886);
nand U14201 (N_14201,N_8318,N_8725);
and U14202 (N_14202,N_8618,N_7133);
xnor U14203 (N_14203,N_7135,N_6917);
nand U14204 (N_14204,N_9605,N_6117);
xnor U14205 (N_14205,N_5529,N_7162);
nor U14206 (N_14206,N_5734,N_8193);
nor U14207 (N_14207,N_8221,N_6404);
nor U14208 (N_14208,N_6660,N_8741);
nor U14209 (N_14209,N_5871,N_5926);
xor U14210 (N_14210,N_7017,N_6245);
or U14211 (N_14211,N_7979,N_9439);
and U14212 (N_14212,N_8576,N_9023);
xnor U14213 (N_14213,N_9305,N_6998);
or U14214 (N_14214,N_7894,N_9235);
nor U14215 (N_14215,N_6690,N_5518);
and U14216 (N_14216,N_5904,N_9518);
nand U14217 (N_14217,N_7926,N_7103);
nand U14218 (N_14218,N_7050,N_9851);
nor U14219 (N_14219,N_8463,N_7339);
nand U14220 (N_14220,N_8075,N_9311);
and U14221 (N_14221,N_7047,N_7920);
nand U14222 (N_14222,N_7084,N_6166);
xnor U14223 (N_14223,N_6339,N_9807);
or U14224 (N_14224,N_6269,N_5780);
nor U14225 (N_14225,N_8544,N_8365);
nand U14226 (N_14226,N_8917,N_9748);
nor U14227 (N_14227,N_5226,N_9096);
xnor U14228 (N_14228,N_7291,N_9351);
xor U14229 (N_14229,N_9520,N_7500);
or U14230 (N_14230,N_6938,N_8896);
and U14231 (N_14231,N_6150,N_6183);
nor U14232 (N_14232,N_6047,N_8776);
xnor U14233 (N_14233,N_7903,N_5393);
and U14234 (N_14234,N_7674,N_9641);
and U14235 (N_14235,N_9944,N_9024);
nand U14236 (N_14236,N_7445,N_8149);
xnor U14237 (N_14237,N_7664,N_7913);
xor U14238 (N_14238,N_8635,N_8096);
or U14239 (N_14239,N_8115,N_6862);
nand U14240 (N_14240,N_8138,N_6126);
xor U14241 (N_14241,N_8189,N_8905);
and U14242 (N_14242,N_9698,N_7315);
nor U14243 (N_14243,N_5712,N_5959);
nor U14244 (N_14244,N_7610,N_8633);
nor U14245 (N_14245,N_6476,N_5286);
nand U14246 (N_14246,N_5981,N_5900);
xor U14247 (N_14247,N_5350,N_7598);
nand U14248 (N_14248,N_7212,N_5324);
nand U14249 (N_14249,N_7214,N_9215);
or U14250 (N_14250,N_8852,N_6198);
nor U14251 (N_14251,N_7783,N_8589);
xnor U14252 (N_14252,N_5781,N_9268);
and U14253 (N_14253,N_7738,N_5316);
xnor U14254 (N_14254,N_5862,N_6857);
and U14255 (N_14255,N_5694,N_8323);
nor U14256 (N_14256,N_7615,N_5050);
nor U14257 (N_14257,N_8208,N_7670);
xor U14258 (N_14258,N_8695,N_5322);
and U14259 (N_14259,N_5835,N_9303);
nand U14260 (N_14260,N_9597,N_5661);
xnor U14261 (N_14261,N_5779,N_9160);
nand U14262 (N_14262,N_5908,N_5137);
xnor U14263 (N_14263,N_9101,N_9267);
nor U14264 (N_14264,N_5474,N_6553);
or U14265 (N_14265,N_6603,N_9895);
nand U14266 (N_14266,N_6520,N_7909);
xnor U14267 (N_14267,N_6114,N_7790);
nor U14268 (N_14268,N_6675,N_7819);
nor U14269 (N_14269,N_7484,N_8942);
nor U14270 (N_14270,N_9874,N_8274);
and U14271 (N_14271,N_7374,N_6296);
and U14272 (N_14272,N_8407,N_8410);
and U14273 (N_14273,N_6874,N_9607);
and U14274 (N_14274,N_9021,N_8451);
or U14275 (N_14275,N_6245,N_8234);
or U14276 (N_14276,N_6871,N_9250);
nand U14277 (N_14277,N_9916,N_9522);
nor U14278 (N_14278,N_7713,N_6373);
nor U14279 (N_14279,N_7879,N_7354);
nor U14280 (N_14280,N_6925,N_7032);
nand U14281 (N_14281,N_6102,N_5893);
nor U14282 (N_14282,N_5261,N_8276);
xor U14283 (N_14283,N_6743,N_6053);
and U14284 (N_14284,N_8682,N_9384);
xnor U14285 (N_14285,N_8131,N_7895);
nor U14286 (N_14286,N_6067,N_9651);
and U14287 (N_14287,N_7853,N_6298);
and U14288 (N_14288,N_9577,N_6598);
xor U14289 (N_14289,N_7457,N_8047);
or U14290 (N_14290,N_8873,N_7836);
and U14291 (N_14291,N_8504,N_6371);
and U14292 (N_14292,N_5120,N_9005);
nand U14293 (N_14293,N_7807,N_6746);
or U14294 (N_14294,N_6530,N_9587);
and U14295 (N_14295,N_7259,N_6721);
nor U14296 (N_14296,N_5610,N_5178);
nand U14297 (N_14297,N_8741,N_7924);
xor U14298 (N_14298,N_6217,N_9270);
xnor U14299 (N_14299,N_7986,N_8513);
nand U14300 (N_14300,N_6535,N_7360);
nor U14301 (N_14301,N_7549,N_5167);
or U14302 (N_14302,N_6268,N_8715);
or U14303 (N_14303,N_8730,N_7876);
or U14304 (N_14304,N_7513,N_6854);
nor U14305 (N_14305,N_9521,N_8343);
nand U14306 (N_14306,N_5077,N_6014);
or U14307 (N_14307,N_5328,N_8816);
xor U14308 (N_14308,N_7976,N_5955);
nor U14309 (N_14309,N_6376,N_8860);
nor U14310 (N_14310,N_6410,N_7651);
and U14311 (N_14311,N_5101,N_9069);
and U14312 (N_14312,N_6283,N_8602);
nor U14313 (N_14313,N_6757,N_6130);
and U14314 (N_14314,N_9013,N_6067);
nor U14315 (N_14315,N_5843,N_7747);
and U14316 (N_14316,N_6931,N_5185);
nand U14317 (N_14317,N_6745,N_9039);
nor U14318 (N_14318,N_9557,N_5885);
and U14319 (N_14319,N_7107,N_8661);
xnor U14320 (N_14320,N_5363,N_7299);
and U14321 (N_14321,N_5702,N_8259);
nand U14322 (N_14322,N_7028,N_6363);
and U14323 (N_14323,N_9764,N_5106);
nand U14324 (N_14324,N_9333,N_7720);
nand U14325 (N_14325,N_8954,N_6215);
nor U14326 (N_14326,N_9478,N_6952);
nand U14327 (N_14327,N_7366,N_8296);
nor U14328 (N_14328,N_9731,N_5675);
and U14329 (N_14329,N_6295,N_8546);
and U14330 (N_14330,N_6907,N_6326);
xor U14331 (N_14331,N_5461,N_8248);
xor U14332 (N_14332,N_7890,N_5996);
and U14333 (N_14333,N_5649,N_5660);
or U14334 (N_14334,N_8337,N_6293);
nor U14335 (N_14335,N_9051,N_9599);
nor U14336 (N_14336,N_5757,N_8535);
xor U14337 (N_14337,N_7180,N_6161);
or U14338 (N_14338,N_6787,N_8033);
xnor U14339 (N_14339,N_9879,N_6343);
and U14340 (N_14340,N_5484,N_5837);
and U14341 (N_14341,N_8729,N_6344);
or U14342 (N_14342,N_6425,N_8870);
nand U14343 (N_14343,N_8259,N_9295);
nand U14344 (N_14344,N_7184,N_6499);
xor U14345 (N_14345,N_7483,N_6318);
nand U14346 (N_14346,N_5964,N_5437);
nand U14347 (N_14347,N_6117,N_6178);
nand U14348 (N_14348,N_6135,N_6882);
nor U14349 (N_14349,N_5465,N_9880);
nand U14350 (N_14350,N_6876,N_7949);
and U14351 (N_14351,N_8525,N_8043);
and U14352 (N_14352,N_8345,N_9929);
xnor U14353 (N_14353,N_9157,N_5385);
nor U14354 (N_14354,N_8919,N_9244);
nand U14355 (N_14355,N_8310,N_6011);
nand U14356 (N_14356,N_7576,N_6129);
nand U14357 (N_14357,N_6107,N_8949);
or U14358 (N_14358,N_7288,N_9579);
nand U14359 (N_14359,N_8390,N_9032);
nand U14360 (N_14360,N_7182,N_5771);
or U14361 (N_14361,N_9134,N_5535);
nor U14362 (N_14362,N_5759,N_7669);
nor U14363 (N_14363,N_8120,N_8863);
xnor U14364 (N_14364,N_5152,N_9761);
nand U14365 (N_14365,N_5936,N_8683);
nor U14366 (N_14366,N_8062,N_8669);
xnor U14367 (N_14367,N_9831,N_5472);
or U14368 (N_14368,N_5155,N_6898);
nand U14369 (N_14369,N_6630,N_7073);
xnor U14370 (N_14370,N_9009,N_9085);
nand U14371 (N_14371,N_7943,N_8291);
nor U14372 (N_14372,N_6775,N_5200);
nand U14373 (N_14373,N_8590,N_9141);
xnor U14374 (N_14374,N_8043,N_5151);
nand U14375 (N_14375,N_8868,N_9092);
xor U14376 (N_14376,N_9901,N_5205);
nor U14377 (N_14377,N_7140,N_5426);
xnor U14378 (N_14378,N_5554,N_5071);
and U14379 (N_14379,N_6991,N_9450);
xnor U14380 (N_14380,N_5433,N_9192);
or U14381 (N_14381,N_7375,N_8345);
nand U14382 (N_14382,N_8458,N_8897);
or U14383 (N_14383,N_8705,N_9731);
xnor U14384 (N_14384,N_5975,N_7345);
xnor U14385 (N_14385,N_7252,N_5045);
xnor U14386 (N_14386,N_5897,N_5289);
nand U14387 (N_14387,N_7713,N_6836);
or U14388 (N_14388,N_6303,N_8090);
xnor U14389 (N_14389,N_8404,N_5517);
nor U14390 (N_14390,N_6336,N_7045);
and U14391 (N_14391,N_6235,N_6468);
xnor U14392 (N_14392,N_8114,N_6895);
or U14393 (N_14393,N_8904,N_8022);
and U14394 (N_14394,N_5320,N_8442);
nor U14395 (N_14395,N_6550,N_5854);
and U14396 (N_14396,N_9134,N_9010);
nor U14397 (N_14397,N_9635,N_9192);
nor U14398 (N_14398,N_8057,N_7749);
nand U14399 (N_14399,N_5199,N_7574);
nor U14400 (N_14400,N_6328,N_7767);
xnor U14401 (N_14401,N_5643,N_7145);
nand U14402 (N_14402,N_7295,N_8240);
xnor U14403 (N_14403,N_9220,N_7104);
nand U14404 (N_14404,N_7443,N_6970);
nand U14405 (N_14405,N_9180,N_6585);
xnor U14406 (N_14406,N_7181,N_8905);
xor U14407 (N_14407,N_6717,N_6589);
xor U14408 (N_14408,N_8672,N_6309);
and U14409 (N_14409,N_6716,N_7578);
nor U14410 (N_14410,N_7855,N_9868);
nand U14411 (N_14411,N_5907,N_7287);
xor U14412 (N_14412,N_6912,N_8871);
xor U14413 (N_14413,N_7108,N_6260);
nor U14414 (N_14414,N_5088,N_6123);
nand U14415 (N_14415,N_6489,N_8252);
nor U14416 (N_14416,N_5012,N_9112);
xor U14417 (N_14417,N_5773,N_9172);
nand U14418 (N_14418,N_7338,N_7807);
or U14419 (N_14419,N_6567,N_6583);
nor U14420 (N_14420,N_5873,N_8430);
and U14421 (N_14421,N_9052,N_9645);
nor U14422 (N_14422,N_9981,N_8803);
and U14423 (N_14423,N_6497,N_8275);
or U14424 (N_14424,N_6095,N_9287);
and U14425 (N_14425,N_8781,N_6294);
or U14426 (N_14426,N_5292,N_6075);
or U14427 (N_14427,N_9327,N_7006);
and U14428 (N_14428,N_9655,N_5256);
nand U14429 (N_14429,N_6742,N_8263);
and U14430 (N_14430,N_5577,N_9125);
and U14431 (N_14431,N_6907,N_7676);
xnor U14432 (N_14432,N_7303,N_5011);
xnor U14433 (N_14433,N_7659,N_7446);
nor U14434 (N_14434,N_8816,N_6562);
xnor U14435 (N_14435,N_9311,N_9317);
xor U14436 (N_14436,N_5950,N_6876);
nand U14437 (N_14437,N_9001,N_7470);
xor U14438 (N_14438,N_8482,N_8782);
and U14439 (N_14439,N_6837,N_7679);
or U14440 (N_14440,N_5234,N_6192);
nor U14441 (N_14441,N_5799,N_5505);
xnor U14442 (N_14442,N_5089,N_8198);
and U14443 (N_14443,N_5447,N_9206);
and U14444 (N_14444,N_8301,N_6618);
or U14445 (N_14445,N_7020,N_9491);
xor U14446 (N_14446,N_5209,N_8438);
xor U14447 (N_14447,N_9509,N_7559);
nor U14448 (N_14448,N_6257,N_5386);
xnor U14449 (N_14449,N_5555,N_9672);
and U14450 (N_14450,N_8083,N_6908);
and U14451 (N_14451,N_8118,N_7296);
or U14452 (N_14452,N_8299,N_5610);
xnor U14453 (N_14453,N_8045,N_9839);
and U14454 (N_14454,N_7173,N_9782);
nor U14455 (N_14455,N_9722,N_6065);
and U14456 (N_14456,N_8668,N_8183);
xor U14457 (N_14457,N_5277,N_7695);
nand U14458 (N_14458,N_6838,N_9673);
nand U14459 (N_14459,N_9698,N_8741);
or U14460 (N_14460,N_8750,N_8312);
xor U14461 (N_14461,N_8862,N_6413);
nor U14462 (N_14462,N_9733,N_5424);
xor U14463 (N_14463,N_8683,N_7301);
nor U14464 (N_14464,N_6810,N_5363);
and U14465 (N_14465,N_7558,N_7432);
nor U14466 (N_14466,N_8267,N_8409);
nor U14467 (N_14467,N_7831,N_8183);
or U14468 (N_14468,N_8761,N_5196);
nand U14469 (N_14469,N_8211,N_7501);
or U14470 (N_14470,N_7226,N_5648);
nor U14471 (N_14471,N_6672,N_7177);
nor U14472 (N_14472,N_8233,N_8126);
nand U14473 (N_14473,N_5874,N_6987);
nor U14474 (N_14474,N_7113,N_5327);
xor U14475 (N_14475,N_9143,N_7735);
nand U14476 (N_14476,N_5191,N_8710);
nand U14477 (N_14477,N_5100,N_6331);
xor U14478 (N_14478,N_5621,N_9955);
nand U14479 (N_14479,N_6757,N_8327);
nor U14480 (N_14480,N_8544,N_7590);
and U14481 (N_14481,N_6326,N_8109);
nand U14482 (N_14482,N_8452,N_7570);
nand U14483 (N_14483,N_8077,N_7737);
nor U14484 (N_14484,N_7743,N_9751);
nor U14485 (N_14485,N_8183,N_6040);
nand U14486 (N_14486,N_7497,N_8030);
and U14487 (N_14487,N_7742,N_7381);
nand U14488 (N_14488,N_8299,N_8084);
or U14489 (N_14489,N_6168,N_6856);
and U14490 (N_14490,N_6258,N_5478);
nand U14491 (N_14491,N_5037,N_6220);
or U14492 (N_14492,N_9884,N_5813);
nand U14493 (N_14493,N_7315,N_5859);
nand U14494 (N_14494,N_7394,N_6763);
xor U14495 (N_14495,N_5265,N_9268);
nand U14496 (N_14496,N_6052,N_9801);
and U14497 (N_14497,N_6360,N_8522);
xnor U14498 (N_14498,N_9399,N_5750);
xor U14499 (N_14499,N_8433,N_5973);
nand U14500 (N_14500,N_5506,N_5823);
and U14501 (N_14501,N_8933,N_5211);
or U14502 (N_14502,N_5767,N_9164);
nor U14503 (N_14503,N_8145,N_8017);
xor U14504 (N_14504,N_9318,N_8723);
xor U14505 (N_14505,N_8094,N_5016);
or U14506 (N_14506,N_8341,N_9450);
and U14507 (N_14507,N_5561,N_6861);
xnor U14508 (N_14508,N_6567,N_5177);
and U14509 (N_14509,N_9243,N_5598);
nor U14510 (N_14510,N_7733,N_7439);
or U14511 (N_14511,N_6287,N_8300);
or U14512 (N_14512,N_8362,N_5338);
or U14513 (N_14513,N_5017,N_5242);
or U14514 (N_14514,N_7351,N_8735);
nand U14515 (N_14515,N_6323,N_6356);
or U14516 (N_14516,N_7648,N_5578);
or U14517 (N_14517,N_5253,N_5984);
nor U14518 (N_14518,N_9022,N_7016);
or U14519 (N_14519,N_5627,N_8184);
and U14520 (N_14520,N_7432,N_5148);
nor U14521 (N_14521,N_9076,N_5334);
nand U14522 (N_14522,N_7697,N_6165);
and U14523 (N_14523,N_5614,N_6336);
or U14524 (N_14524,N_7307,N_7544);
or U14525 (N_14525,N_9289,N_7069);
and U14526 (N_14526,N_7708,N_6459);
and U14527 (N_14527,N_9189,N_8665);
xnor U14528 (N_14528,N_7477,N_6573);
nand U14529 (N_14529,N_9150,N_5773);
and U14530 (N_14530,N_8453,N_5363);
nor U14531 (N_14531,N_7048,N_6411);
nor U14532 (N_14532,N_9866,N_7688);
xnor U14533 (N_14533,N_7927,N_9314);
xnor U14534 (N_14534,N_7278,N_9435);
and U14535 (N_14535,N_5613,N_7369);
nand U14536 (N_14536,N_7368,N_7557);
or U14537 (N_14537,N_7412,N_7625);
xnor U14538 (N_14538,N_7637,N_9991);
or U14539 (N_14539,N_6651,N_6092);
nor U14540 (N_14540,N_7147,N_7263);
nor U14541 (N_14541,N_6556,N_8229);
or U14542 (N_14542,N_8153,N_6096);
nand U14543 (N_14543,N_9075,N_7327);
and U14544 (N_14544,N_7555,N_8287);
nand U14545 (N_14545,N_9922,N_8800);
nand U14546 (N_14546,N_5683,N_6500);
or U14547 (N_14547,N_9384,N_9343);
xnor U14548 (N_14548,N_7693,N_6110);
and U14549 (N_14549,N_8735,N_7986);
or U14550 (N_14550,N_8062,N_6176);
or U14551 (N_14551,N_8368,N_8851);
and U14552 (N_14552,N_5111,N_8873);
and U14553 (N_14553,N_8961,N_6852);
or U14554 (N_14554,N_8619,N_9645);
xor U14555 (N_14555,N_9787,N_8115);
xor U14556 (N_14556,N_7416,N_7581);
or U14557 (N_14557,N_6630,N_5622);
nor U14558 (N_14558,N_7494,N_8921);
and U14559 (N_14559,N_6622,N_7865);
or U14560 (N_14560,N_6943,N_8847);
nor U14561 (N_14561,N_6057,N_8192);
xnor U14562 (N_14562,N_8449,N_7637);
nand U14563 (N_14563,N_6870,N_6405);
xor U14564 (N_14564,N_7356,N_7968);
and U14565 (N_14565,N_5087,N_6851);
and U14566 (N_14566,N_8710,N_5535);
xnor U14567 (N_14567,N_8798,N_7865);
nand U14568 (N_14568,N_7176,N_5606);
xnor U14569 (N_14569,N_7935,N_7673);
nand U14570 (N_14570,N_6736,N_8359);
nand U14571 (N_14571,N_6124,N_7504);
nor U14572 (N_14572,N_8196,N_6656);
xnor U14573 (N_14573,N_9536,N_8995);
or U14574 (N_14574,N_8727,N_6907);
and U14575 (N_14575,N_8088,N_7083);
nand U14576 (N_14576,N_8648,N_6904);
nand U14577 (N_14577,N_9128,N_7324);
xor U14578 (N_14578,N_6012,N_8494);
nand U14579 (N_14579,N_6489,N_9497);
xor U14580 (N_14580,N_7709,N_6015);
nand U14581 (N_14581,N_5532,N_7652);
and U14582 (N_14582,N_6181,N_8162);
nor U14583 (N_14583,N_7471,N_6075);
or U14584 (N_14584,N_5882,N_6359);
nand U14585 (N_14585,N_8738,N_5962);
and U14586 (N_14586,N_9756,N_5964);
and U14587 (N_14587,N_9140,N_6963);
nand U14588 (N_14588,N_7649,N_8013);
nor U14589 (N_14589,N_8588,N_8382);
and U14590 (N_14590,N_9973,N_6960);
xnor U14591 (N_14591,N_6367,N_8795);
nor U14592 (N_14592,N_8645,N_5656);
xnor U14593 (N_14593,N_5462,N_8648);
xor U14594 (N_14594,N_9391,N_6040);
nand U14595 (N_14595,N_8195,N_9983);
and U14596 (N_14596,N_6637,N_5588);
nor U14597 (N_14597,N_7407,N_8129);
xnor U14598 (N_14598,N_9840,N_6272);
nor U14599 (N_14599,N_5555,N_6508);
and U14600 (N_14600,N_6289,N_6049);
xor U14601 (N_14601,N_7088,N_6111);
and U14602 (N_14602,N_9496,N_5297);
xnor U14603 (N_14603,N_6984,N_9541);
nand U14604 (N_14604,N_8593,N_7761);
and U14605 (N_14605,N_7821,N_7698);
or U14606 (N_14606,N_5921,N_9273);
nor U14607 (N_14607,N_9560,N_9153);
or U14608 (N_14608,N_5251,N_9651);
and U14609 (N_14609,N_5151,N_5237);
or U14610 (N_14610,N_9437,N_7273);
xnor U14611 (N_14611,N_8007,N_6574);
xor U14612 (N_14612,N_5895,N_8113);
or U14613 (N_14613,N_5870,N_8619);
nor U14614 (N_14614,N_7864,N_7128);
nor U14615 (N_14615,N_6323,N_9318);
xnor U14616 (N_14616,N_9367,N_8425);
and U14617 (N_14617,N_7588,N_8913);
and U14618 (N_14618,N_5524,N_6287);
nor U14619 (N_14619,N_5843,N_9579);
xor U14620 (N_14620,N_7150,N_7551);
xnor U14621 (N_14621,N_7368,N_7391);
xnor U14622 (N_14622,N_6643,N_6455);
or U14623 (N_14623,N_5070,N_9695);
nand U14624 (N_14624,N_6488,N_9375);
nand U14625 (N_14625,N_5007,N_7664);
nand U14626 (N_14626,N_8237,N_9558);
nand U14627 (N_14627,N_5237,N_8245);
xor U14628 (N_14628,N_9681,N_6539);
nor U14629 (N_14629,N_5799,N_7566);
xnor U14630 (N_14630,N_7354,N_5433);
and U14631 (N_14631,N_5245,N_5653);
xor U14632 (N_14632,N_8178,N_9466);
xnor U14633 (N_14633,N_6955,N_7439);
and U14634 (N_14634,N_7511,N_8240);
or U14635 (N_14635,N_9338,N_5097);
and U14636 (N_14636,N_7510,N_6820);
xor U14637 (N_14637,N_7237,N_9296);
or U14638 (N_14638,N_8585,N_7083);
or U14639 (N_14639,N_9986,N_6866);
and U14640 (N_14640,N_9080,N_9785);
and U14641 (N_14641,N_6975,N_7185);
and U14642 (N_14642,N_7155,N_5181);
nand U14643 (N_14643,N_8407,N_5337);
or U14644 (N_14644,N_9498,N_6621);
or U14645 (N_14645,N_5160,N_7347);
nand U14646 (N_14646,N_5081,N_6353);
and U14647 (N_14647,N_5361,N_5227);
and U14648 (N_14648,N_6636,N_6156);
and U14649 (N_14649,N_5055,N_5537);
and U14650 (N_14650,N_5198,N_8875);
nand U14651 (N_14651,N_9080,N_6909);
and U14652 (N_14652,N_7132,N_8975);
and U14653 (N_14653,N_9019,N_8702);
or U14654 (N_14654,N_6527,N_7210);
xnor U14655 (N_14655,N_8447,N_7141);
xor U14656 (N_14656,N_6133,N_8060);
and U14657 (N_14657,N_6234,N_9313);
nor U14658 (N_14658,N_9763,N_8442);
nor U14659 (N_14659,N_9320,N_8553);
nand U14660 (N_14660,N_9234,N_8115);
xnor U14661 (N_14661,N_5792,N_5180);
and U14662 (N_14662,N_8621,N_6794);
xnor U14663 (N_14663,N_8439,N_7037);
or U14664 (N_14664,N_5213,N_5054);
xor U14665 (N_14665,N_8740,N_6773);
xnor U14666 (N_14666,N_6211,N_5147);
and U14667 (N_14667,N_8030,N_8568);
or U14668 (N_14668,N_5639,N_6282);
and U14669 (N_14669,N_5171,N_5527);
nand U14670 (N_14670,N_7068,N_5250);
or U14671 (N_14671,N_9997,N_7361);
and U14672 (N_14672,N_9470,N_7538);
or U14673 (N_14673,N_6777,N_9637);
and U14674 (N_14674,N_9988,N_8221);
nand U14675 (N_14675,N_5961,N_6409);
nand U14676 (N_14676,N_5094,N_8186);
and U14677 (N_14677,N_6558,N_9139);
xnor U14678 (N_14678,N_6191,N_9588);
nand U14679 (N_14679,N_6521,N_8982);
or U14680 (N_14680,N_8571,N_6591);
nand U14681 (N_14681,N_9409,N_7629);
or U14682 (N_14682,N_6056,N_9269);
xnor U14683 (N_14683,N_6028,N_8891);
and U14684 (N_14684,N_7846,N_9588);
or U14685 (N_14685,N_7702,N_9874);
and U14686 (N_14686,N_7470,N_5596);
xnor U14687 (N_14687,N_6229,N_6499);
nand U14688 (N_14688,N_5838,N_8251);
nand U14689 (N_14689,N_9676,N_5596);
or U14690 (N_14690,N_9375,N_6386);
and U14691 (N_14691,N_8170,N_8696);
nand U14692 (N_14692,N_7004,N_9601);
xor U14693 (N_14693,N_8544,N_8699);
nor U14694 (N_14694,N_6142,N_7040);
xnor U14695 (N_14695,N_7737,N_9400);
xnor U14696 (N_14696,N_8220,N_7188);
or U14697 (N_14697,N_9131,N_5449);
and U14698 (N_14698,N_6719,N_8592);
and U14699 (N_14699,N_7229,N_5058);
or U14700 (N_14700,N_9581,N_5993);
and U14701 (N_14701,N_5681,N_5079);
and U14702 (N_14702,N_5660,N_5294);
or U14703 (N_14703,N_6105,N_9589);
and U14704 (N_14704,N_5951,N_7832);
nor U14705 (N_14705,N_6177,N_9983);
xor U14706 (N_14706,N_7207,N_9501);
nor U14707 (N_14707,N_7672,N_9772);
nor U14708 (N_14708,N_5541,N_6808);
nor U14709 (N_14709,N_8008,N_9633);
nand U14710 (N_14710,N_8141,N_6877);
and U14711 (N_14711,N_5535,N_8304);
and U14712 (N_14712,N_9087,N_7914);
nand U14713 (N_14713,N_9330,N_6333);
and U14714 (N_14714,N_9513,N_8069);
nor U14715 (N_14715,N_8872,N_9817);
and U14716 (N_14716,N_8611,N_5002);
xor U14717 (N_14717,N_7800,N_6279);
or U14718 (N_14718,N_8458,N_7726);
xor U14719 (N_14719,N_7481,N_5574);
nand U14720 (N_14720,N_8765,N_7315);
and U14721 (N_14721,N_8940,N_6880);
or U14722 (N_14722,N_9766,N_7465);
or U14723 (N_14723,N_7825,N_7355);
and U14724 (N_14724,N_5131,N_8232);
and U14725 (N_14725,N_8604,N_5253);
nor U14726 (N_14726,N_7617,N_7509);
nor U14727 (N_14727,N_5818,N_5870);
nor U14728 (N_14728,N_7342,N_5830);
and U14729 (N_14729,N_8749,N_7980);
and U14730 (N_14730,N_6096,N_5464);
nor U14731 (N_14731,N_9024,N_6534);
or U14732 (N_14732,N_7250,N_9014);
and U14733 (N_14733,N_9796,N_8637);
and U14734 (N_14734,N_6086,N_5257);
nor U14735 (N_14735,N_8696,N_5256);
xor U14736 (N_14736,N_9023,N_8259);
nor U14737 (N_14737,N_6297,N_9025);
nor U14738 (N_14738,N_9922,N_6668);
nor U14739 (N_14739,N_6010,N_5136);
nor U14740 (N_14740,N_8598,N_7703);
xnor U14741 (N_14741,N_6661,N_8648);
xnor U14742 (N_14742,N_8518,N_6018);
and U14743 (N_14743,N_9817,N_8029);
or U14744 (N_14744,N_6340,N_5483);
and U14745 (N_14745,N_9640,N_9553);
nor U14746 (N_14746,N_5872,N_9294);
nand U14747 (N_14747,N_9826,N_7351);
nor U14748 (N_14748,N_6622,N_6902);
nor U14749 (N_14749,N_6125,N_8817);
nor U14750 (N_14750,N_5582,N_7746);
nand U14751 (N_14751,N_6749,N_9184);
xor U14752 (N_14752,N_7049,N_9094);
xor U14753 (N_14753,N_8929,N_7981);
xnor U14754 (N_14754,N_7370,N_6402);
nand U14755 (N_14755,N_7061,N_5956);
nand U14756 (N_14756,N_7129,N_6945);
and U14757 (N_14757,N_6908,N_7090);
and U14758 (N_14758,N_8094,N_6000);
nor U14759 (N_14759,N_5955,N_5579);
nor U14760 (N_14760,N_5570,N_6596);
xor U14761 (N_14761,N_5477,N_8031);
nand U14762 (N_14762,N_7008,N_8847);
nor U14763 (N_14763,N_7928,N_9422);
and U14764 (N_14764,N_8920,N_5418);
nand U14765 (N_14765,N_5402,N_7624);
and U14766 (N_14766,N_7617,N_5279);
nor U14767 (N_14767,N_7810,N_8889);
xor U14768 (N_14768,N_9791,N_6981);
nand U14769 (N_14769,N_8886,N_6967);
nor U14770 (N_14770,N_7997,N_6673);
nor U14771 (N_14771,N_5538,N_8939);
xor U14772 (N_14772,N_5603,N_7760);
nand U14773 (N_14773,N_7272,N_8326);
nor U14774 (N_14774,N_6686,N_5269);
nand U14775 (N_14775,N_9060,N_7630);
or U14776 (N_14776,N_9616,N_8921);
nor U14777 (N_14777,N_9409,N_9407);
and U14778 (N_14778,N_6199,N_9755);
nand U14779 (N_14779,N_8569,N_9118);
nand U14780 (N_14780,N_9264,N_8363);
and U14781 (N_14781,N_9915,N_8739);
nand U14782 (N_14782,N_7080,N_6893);
and U14783 (N_14783,N_6019,N_8294);
and U14784 (N_14784,N_9588,N_7495);
nor U14785 (N_14785,N_7697,N_8616);
xnor U14786 (N_14786,N_5810,N_9776);
xor U14787 (N_14787,N_5474,N_9689);
nand U14788 (N_14788,N_6551,N_5656);
nor U14789 (N_14789,N_7414,N_7796);
nand U14790 (N_14790,N_8719,N_9464);
xnor U14791 (N_14791,N_9340,N_5650);
and U14792 (N_14792,N_5381,N_7967);
or U14793 (N_14793,N_7015,N_8672);
nand U14794 (N_14794,N_7020,N_9854);
and U14795 (N_14795,N_6039,N_8180);
and U14796 (N_14796,N_9515,N_5926);
and U14797 (N_14797,N_5924,N_7375);
nand U14798 (N_14798,N_7097,N_8805);
nor U14799 (N_14799,N_6977,N_9081);
nand U14800 (N_14800,N_5053,N_7335);
nor U14801 (N_14801,N_7563,N_8360);
xnor U14802 (N_14802,N_8716,N_7572);
or U14803 (N_14803,N_7893,N_9771);
xor U14804 (N_14804,N_7268,N_5848);
nand U14805 (N_14805,N_5202,N_8277);
xor U14806 (N_14806,N_9017,N_7521);
nor U14807 (N_14807,N_8820,N_6216);
nand U14808 (N_14808,N_6797,N_9659);
and U14809 (N_14809,N_9192,N_6343);
nor U14810 (N_14810,N_6076,N_8116);
nand U14811 (N_14811,N_9767,N_8718);
and U14812 (N_14812,N_6011,N_9487);
nand U14813 (N_14813,N_5144,N_8200);
nor U14814 (N_14814,N_5718,N_8517);
nand U14815 (N_14815,N_5328,N_8277);
or U14816 (N_14816,N_9646,N_5604);
nor U14817 (N_14817,N_7529,N_7966);
nand U14818 (N_14818,N_7587,N_8585);
and U14819 (N_14819,N_9128,N_7020);
xor U14820 (N_14820,N_9683,N_6684);
nand U14821 (N_14821,N_6391,N_8135);
xor U14822 (N_14822,N_7972,N_5207);
nand U14823 (N_14823,N_5696,N_8639);
xnor U14824 (N_14824,N_7727,N_9043);
xor U14825 (N_14825,N_5633,N_6308);
or U14826 (N_14826,N_7654,N_6028);
and U14827 (N_14827,N_7796,N_7710);
or U14828 (N_14828,N_8497,N_7360);
nor U14829 (N_14829,N_7267,N_5489);
xor U14830 (N_14830,N_6405,N_6927);
nor U14831 (N_14831,N_7622,N_8113);
and U14832 (N_14832,N_5170,N_9585);
and U14833 (N_14833,N_5781,N_7684);
xor U14834 (N_14834,N_6133,N_6899);
nor U14835 (N_14835,N_5381,N_9725);
xnor U14836 (N_14836,N_7384,N_9046);
nand U14837 (N_14837,N_7044,N_8373);
and U14838 (N_14838,N_8679,N_5278);
or U14839 (N_14839,N_8143,N_9941);
or U14840 (N_14840,N_8512,N_8296);
and U14841 (N_14841,N_8844,N_6271);
or U14842 (N_14842,N_5850,N_9948);
or U14843 (N_14843,N_9146,N_6749);
or U14844 (N_14844,N_9179,N_6968);
or U14845 (N_14845,N_5479,N_5173);
nand U14846 (N_14846,N_9099,N_6504);
nor U14847 (N_14847,N_5673,N_7816);
nand U14848 (N_14848,N_5283,N_5161);
xnor U14849 (N_14849,N_7087,N_8253);
nor U14850 (N_14850,N_6357,N_7804);
nand U14851 (N_14851,N_6314,N_8829);
nand U14852 (N_14852,N_5613,N_5105);
nor U14853 (N_14853,N_6357,N_9529);
nor U14854 (N_14854,N_7835,N_7913);
xor U14855 (N_14855,N_7934,N_5331);
xor U14856 (N_14856,N_6066,N_5291);
nand U14857 (N_14857,N_7554,N_6163);
or U14858 (N_14858,N_9238,N_9815);
nand U14859 (N_14859,N_6898,N_6675);
xnor U14860 (N_14860,N_6183,N_9087);
xor U14861 (N_14861,N_9874,N_5284);
and U14862 (N_14862,N_6376,N_5476);
or U14863 (N_14863,N_9018,N_5273);
nand U14864 (N_14864,N_5338,N_9016);
and U14865 (N_14865,N_8503,N_9035);
or U14866 (N_14866,N_5382,N_6359);
or U14867 (N_14867,N_6979,N_7137);
nor U14868 (N_14868,N_6382,N_7371);
xnor U14869 (N_14869,N_6572,N_5201);
nand U14870 (N_14870,N_6927,N_9649);
or U14871 (N_14871,N_9508,N_5388);
nor U14872 (N_14872,N_8807,N_6583);
nor U14873 (N_14873,N_5230,N_5257);
nor U14874 (N_14874,N_6580,N_7642);
and U14875 (N_14875,N_5294,N_8011);
or U14876 (N_14876,N_6092,N_9502);
nor U14877 (N_14877,N_6429,N_5124);
and U14878 (N_14878,N_6754,N_9863);
nand U14879 (N_14879,N_8594,N_8418);
nor U14880 (N_14880,N_5428,N_5043);
xnor U14881 (N_14881,N_8664,N_9767);
and U14882 (N_14882,N_8537,N_6317);
nor U14883 (N_14883,N_6891,N_8054);
xor U14884 (N_14884,N_9859,N_8179);
and U14885 (N_14885,N_9100,N_5810);
xor U14886 (N_14886,N_5601,N_9494);
xnor U14887 (N_14887,N_9745,N_5003);
or U14888 (N_14888,N_9576,N_6438);
nand U14889 (N_14889,N_6213,N_5140);
nor U14890 (N_14890,N_5209,N_9392);
or U14891 (N_14891,N_7511,N_6482);
nor U14892 (N_14892,N_6360,N_8770);
or U14893 (N_14893,N_6834,N_7696);
nand U14894 (N_14894,N_6317,N_9392);
nand U14895 (N_14895,N_7396,N_8269);
and U14896 (N_14896,N_8933,N_8299);
nand U14897 (N_14897,N_6872,N_7425);
xor U14898 (N_14898,N_6476,N_5231);
nor U14899 (N_14899,N_8171,N_6686);
and U14900 (N_14900,N_8677,N_8908);
nor U14901 (N_14901,N_6408,N_7770);
and U14902 (N_14902,N_8484,N_8936);
xor U14903 (N_14903,N_8847,N_7513);
xnor U14904 (N_14904,N_7672,N_5825);
xnor U14905 (N_14905,N_9138,N_7073);
or U14906 (N_14906,N_8580,N_6619);
xnor U14907 (N_14907,N_5105,N_8249);
and U14908 (N_14908,N_6806,N_6424);
or U14909 (N_14909,N_7556,N_5617);
and U14910 (N_14910,N_8195,N_8749);
nand U14911 (N_14911,N_8358,N_6699);
xnor U14912 (N_14912,N_9252,N_5607);
nand U14913 (N_14913,N_9868,N_6225);
xnor U14914 (N_14914,N_9952,N_5897);
nand U14915 (N_14915,N_8453,N_8293);
or U14916 (N_14916,N_9681,N_6163);
and U14917 (N_14917,N_9319,N_9993);
or U14918 (N_14918,N_7549,N_9466);
nand U14919 (N_14919,N_5458,N_6948);
nor U14920 (N_14920,N_8002,N_7429);
and U14921 (N_14921,N_8051,N_8586);
xor U14922 (N_14922,N_9284,N_8260);
nand U14923 (N_14923,N_6028,N_8203);
and U14924 (N_14924,N_7497,N_8213);
and U14925 (N_14925,N_7633,N_9586);
and U14926 (N_14926,N_6989,N_6159);
and U14927 (N_14927,N_8684,N_5650);
or U14928 (N_14928,N_6985,N_5285);
nand U14929 (N_14929,N_7283,N_9709);
or U14930 (N_14930,N_5772,N_6637);
xnor U14931 (N_14931,N_5608,N_8489);
nand U14932 (N_14932,N_9983,N_6146);
xor U14933 (N_14933,N_5048,N_6605);
nand U14934 (N_14934,N_7609,N_8420);
nor U14935 (N_14935,N_6928,N_7425);
nand U14936 (N_14936,N_9410,N_7212);
xor U14937 (N_14937,N_5241,N_5287);
nor U14938 (N_14938,N_5699,N_8956);
nand U14939 (N_14939,N_5057,N_5822);
nand U14940 (N_14940,N_5010,N_7546);
xor U14941 (N_14941,N_5503,N_9345);
nor U14942 (N_14942,N_8831,N_7889);
nand U14943 (N_14943,N_9079,N_7800);
or U14944 (N_14944,N_6336,N_5568);
nand U14945 (N_14945,N_7561,N_5518);
xor U14946 (N_14946,N_7103,N_8793);
or U14947 (N_14947,N_5394,N_6329);
nand U14948 (N_14948,N_9151,N_8343);
nor U14949 (N_14949,N_7889,N_8590);
and U14950 (N_14950,N_6256,N_9311);
nand U14951 (N_14951,N_7202,N_5601);
or U14952 (N_14952,N_8787,N_8755);
or U14953 (N_14953,N_6667,N_6644);
and U14954 (N_14954,N_5700,N_8306);
nor U14955 (N_14955,N_6101,N_8993);
and U14956 (N_14956,N_8335,N_9822);
or U14957 (N_14957,N_8849,N_9691);
nand U14958 (N_14958,N_9485,N_7211);
or U14959 (N_14959,N_9003,N_6390);
nor U14960 (N_14960,N_6951,N_7099);
nor U14961 (N_14961,N_5118,N_8685);
nor U14962 (N_14962,N_8567,N_8244);
and U14963 (N_14963,N_7455,N_6509);
or U14964 (N_14964,N_8899,N_8730);
and U14965 (N_14965,N_8729,N_8275);
xnor U14966 (N_14966,N_6152,N_9002);
nand U14967 (N_14967,N_8217,N_6206);
nor U14968 (N_14968,N_8512,N_7978);
and U14969 (N_14969,N_8144,N_9065);
xor U14970 (N_14970,N_9015,N_5243);
or U14971 (N_14971,N_7347,N_5208);
and U14972 (N_14972,N_6276,N_5212);
nand U14973 (N_14973,N_6745,N_9408);
or U14974 (N_14974,N_6845,N_5610);
nor U14975 (N_14975,N_7233,N_6836);
nor U14976 (N_14976,N_9068,N_9374);
nor U14977 (N_14977,N_9293,N_6006);
or U14978 (N_14978,N_7048,N_6934);
or U14979 (N_14979,N_5858,N_6234);
or U14980 (N_14980,N_6058,N_6451);
nor U14981 (N_14981,N_6404,N_5888);
and U14982 (N_14982,N_7713,N_9533);
and U14983 (N_14983,N_6526,N_9338);
nand U14984 (N_14984,N_5360,N_9278);
nor U14985 (N_14985,N_9341,N_7027);
nand U14986 (N_14986,N_7649,N_9738);
xor U14987 (N_14987,N_7410,N_6466);
xor U14988 (N_14988,N_9905,N_8321);
or U14989 (N_14989,N_5765,N_7829);
nor U14990 (N_14990,N_6509,N_7685);
and U14991 (N_14991,N_7705,N_9806);
nor U14992 (N_14992,N_8709,N_9921);
or U14993 (N_14993,N_8818,N_7579);
xnor U14994 (N_14994,N_7257,N_8218);
nor U14995 (N_14995,N_7966,N_5283);
and U14996 (N_14996,N_8880,N_9565);
nor U14997 (N_14997,N_9301,N_5358);
nor U14998 (N_14998,N_7761,N_9961);
nand U14999 (N_14999,N_6030,N_7514);
xor U15000 (N_15000,N_10527,N_12351);
and U15001 (N_15001,N_12341,N_11467);
xor U15002 (N_15002,N_14244,N_13261);
and U15003 (N_15003,N_14005,N_14819);
nand U15004 (N_15004,N_10280,N_14956);
or U15005 (N_15005,N_12765,N_12720);
nor U15006 (N_15006,N_11611,N_13866);
xnor U15007 (N_15007,N_10849,N_11164);
nand U15008 (N_15008,N_10069,N_13985);
xor U15009 (N_15009,N_10377,N_12870);
and U15010 (N_15010,N_10437,N_12953);
nand U15011 (N_15011,N_10734,N_14303);
or U15012 (N_15012,N_11753,N_10468);
xor U15013 (N_15013,N_11483,N_11718);
or U15014 (N_15014,N_10400,N_12163);
and U15015 (N_15015,N_12108,N_13542);
xor U15016 (N_15016,N_10754,N_12338);
or U15017 (N_15017,N_10108,N_10550);
or U15018 (N_15018,N_13804,N_12919);
nand U15019 (N_15019,N_14578,N_14935);
or U15020 (N_15020,N_11955,N_12233);
xnor U15021 (N_15021,N_13802,N_13943);
nor U15022 (N_15022,N_14734,N_14473);
and U15023 (N_15023,N_13235,N_12181);
nand U15024 (N_15024,N_11821,N_12121);
nand U15025 (N_15025,N_12712,N_13563);
xor U15026 (N_15026,N_14988,N_11680);
and U15027 (N_15027,N_14326,N_11002);
or U15028 (N_15028,N_11339,N_13726);
and U15029 (N_15029,N_13275,N_11288);
or U15030 (N_15030,N_12867,N_10884);
xor U15031 (N_15031,N_13553,N_13256);
and U15032 (N_15032,N_13383,N_14368);
or U15033 (N_15033,N_12826,N_12923);
nand U15034 (N_15034,N_14875,N_14806);
and U15035 (N_15035,N_11970,N_13351);
nand U15036 (N_15036,N_13225,N_10154);
nand U15037 (N_15037,N_10781,N_13783);
and U15038 (N_15038,N_12392,N_14438);
xor U15039 (N_15039,N_14260,N_14727);
xor U15040 (N_15040,N_13741,N_13897);
nor U15041 (N_15041,N_11953,N_13703);
nor U15042 (N_15042,N_10014,N_14736);
or U15043 (N_15043,N_11185,N_12489);
or U15044 (N_15044,N_10023,N_13872);
xnor U15045 (N_15045,N_11171,N_12693);
nor U15046 (N_15046,N_12795,N_12492);
or U15047 (N_15047,N_12323,N_10887);
nor U15048 (N_15048,N_10399,N_11292);
xor U15049 (N_15049,N_12902,N_10316);
nand U15050 (N_15050,N_10523,N_14812);
nor U15051 (N_15051,N_11357,N_10963);
nor U15052 (N_15052,N_10463,N_13270);
nand U15053 (N_15053,N_13458,N_13240);
nand U15054 (N_15054,N_11628,N_10715);
or U15055 (N_15055,N_12397,N_10691);
or U15056 (N_15056,N_10586,N_12628);
nand U15057 (N_15057,N_10984,N_11617);
or U15058 (N_15058,N_12822,N_13020);
nor U15059 (N_15059,N_13330,N_10766);
nand U15060 (N_15060,N_14279,N_13909);
and U15061 (N_15061,N_10825,N_10495);
nand U15062 (N_15062,N_11222,N_13205);
xnor U15063 (N_15063,N_13614,N_14141);
xor U15064 (N_15064,N_11360,N_14766);
nor U15065 (N_15065,N_12992,N_10322);
or U15066 (N_15066,N_11771,N_14485);
and U15067 (N_15067,N_14525,N_13878);
nand U15068 (N_15068,N_14721,N_12728);
nand U15069 (N_15069,N_10654,N_11275);
nor U15070 (N_15070,N_13396,N_12428);
xnor U15071 (N_15071,N_14581,N_12624);
and U15072 (N_15072,N_12709,N_10513);
nor U15073 (N_15073,N_12276,N_10676);
nor U15074 (N_15074,N_14767,N_13829);
and U15075 (N_15075,N_10137,N_14362);
nor U15076 (N_15076,N_10829,N_12914);
and U15077 (N_15077,N_10362,N_10904);
and U15078 (N_15078,N_12944,N_14732);
nand U15079 (N_15079,N_12139,N_13486);
nor U15080 (N_15080,N_10896,N_11077);
or U15081 (N_15081,N_11717,N_11981);
xnor U15082 (N_15082,N_14940,N_11957);
xor U15083 (N_15083,N_11911,N_13352);
xnor U15084 (N_15084,N_14207,N_13737);
and U15085 (N_15085,N_12807,N_14064);
and U15086 (N_15086,N_13833,N_13013);
nor U15087 (N_15087,N_10445,N_14430);
or U15088 (N_15088,N_13095,N_14567);
nor U15089 (N_15089,N_10290,N_14807);
or U15090 (N_15090,N_10001,N_13090);
xnor U15091 (N_15091,N_11330,N_10057);
xnor U15092 (N_15092,N_12474,N_11128);
or U15093 (N_15093,N_12223,N_14523);
and U15094 (N_15094,N_12009,N_12898);
nand U15095 (N_15095,N_10058,N_13334);
xnor U15096 (N_15096,N_12660,N_12295);
nand U15097 (N_15097,N_12639,N_14038);
nand U15098 (N_15098,N_14809,N_14881);
nand U15099 (N_15099,N_10927,N_10041);
or U15100 (N_15100,N_14841,N_13271);
nand U15101 (N_15101,N_12806,N_12935);
and U15102 (N_15102,N_11367,N_11010);
or U15103 (N_15103,N_11337,N_11472);
nand U15104 (N_15104,N_12832,N_10009);
nor U15105 (N_15105,N_14185,N_12472);
xnor U15106 (N_15106,N_10130,N_13962);
xor U15107 (N_15107,N_14879,N_12705);
or U15108 (N_15108,N_10895,N_13107);
or U15109 (N_15109,N_10354,N_13482);
xor U15110 (N_15110,N_13129,N_11057);
nor U15111 (N_15111,N_14846,N_12852);
xor U15112 (N_15112,N_11751,N_12873);
nand U15113 (N_15113,N_14212,N_14001);
nand U15114 (N_15114,N_12636,N_11258);
and U15115 (N_15115,N_12547,N_10350);
xnor U15116 (N_15116,N_10355,N_12941);
and U15117 (N_15117,N_13559,N_14650);
and U15118 (N_15118,N_14288,N_13036);
nand U15119 (N_15119,N_12597,N_14811);
xnor U15120 (N_15120,N_10481,N_13864);
xor U15121 (N_15121,N_10277,N_14059);
nor U15122 (N_15122,N_14883,N_10585);
or U15123 (N_15123,N_11815,N_12051);
nor U15124 (N_15124,N_10040,N_14179);
and U15125 (N_15125,N_12371,N_11789);
or U15126 (N_15126,N_11799,N_11690);
and U15127 (N_15127,N_13386,N_11481);
nand U15128 (N_15128,N_14055,N_14825);
nand U15129 (N_15129,N_14254,N_14393);
xor U15130 (N_15130,N_13638,N_12741);
and U15131 (N_15131,N_12420,N_12286);
nand U15132 (N_15132,N_13886,N_10665);
or U15133 (N_15133,N_11384,N_11712);
nand U15134 (N_15134,N_13997,N_14345);
or U15135 (N_15135,N_14715,N_10753);
or U15136 (N_15136,N_11013,N_14320);
or U15137 (N_15137,N_10480,N_14124);
nand U15138 (N_15138,N_14286,N_10938);
nand U15139 (N_15139,N_10744,N_13565);
xnor U15140 (N_15140,N_11852,N_14389);
and U15141 (N_15141,N_10060,N_11172);
nand U15142 (N_15142,N_13100,N_14927);
nor U15143 (N_15143,N_13440,N_14192);
and U15144 (N_15144,N_14187,N_10484);
or U15145 (N_15145,N_12643,N_11791);
nor U15146 (N_15146,N_11266,N_10006);
and U15147 (N_15147,N_13582,N_14941);
xor U15148 (N_15148,N_10148,N_12389);
or U15149 (N_15149,N_11140,N_11933);
xnor U15150 (N_15150,N_12846,N_13282);
xnor U15151 (N_15151,N_10308,N_14224);
xor U15152 (N_15152,N_14028,N_10250);
xnor U15153 (N_15153,N_12706,N_13471);
nor U15154 (N_15154,N_11301,N_14171);
nor U15155 (N_15155,N_13716,N_10637);
xnor U15156 (N_15156,N_11592,N_14282);
nand U15157 (N_15157,N_10470,N_13195);
nand U15158 (N_15158,N_13697,N_10748);
nor U15159 (N_15159,N_14667,N_13319);
and U15160 (N_15160,N_14090,N_13549);
and U15161 (N_15161,N_10440,N_11640);
and U15162 (N_15162,N_14822,N_10672);
or U15163 (N_15163,N_14067,N_11631);
xnor U15164 (N_15164,N_11543,N_11445);
and U15165 (N_15165,N_12932,N_12861);
and U15166 (N_15166,N_10363,N_13687);
nor U15167 (N_15167,N_10318,N_13644);
nor U15168 (N_15168,N_14772,N_14234);
or U15169 (N_15169,N_12101,N_14200);
xor U15170 (N_15170,N_14016,N_11584);
nor U15171 (N_15171,N_13893,N_10779);
nand U15172 (N_15172,N_14645,N_14552);
or U15173 (N_15173,N_13402,N_13349);
and U15174 (N_15174,N_12685,N_13144);
or U15175 (N_15175,N_10537,N_10692);
and U15176 (N_15176,N_11734,N_12525);
nor U15177 (N_15177,N_10084,N_10852);
nor U15178 (N_15178,N_10155,N_13372);
or U15179 (N_15179,N_13409,N_14503);
or U15180 (N_15180,N_10858,N_11954);
or U15181 (N_15181,N_12933,N_13010);
xnor U15182 (N_15182,N_13841,N_14607);
or U15183 (N_15183,N_11961,N_14747);
nand U15184 (N_15184,N_13541,N_13269);
or U15185 (N_15185,N_12137,N_12752);
and U15186 (N_15186,N_12251,N_10421);
xor U15187 (N_15187,N_12533,N_10908);
nand U15188 (N_15188,N_10985,N_10086);
or U15189 (N_15189,N_10374,N_12230);
nor U15190 (N_15190,N_13785,N_10799);
xnor U15191 (N_15191,N_14256,N_13747);
or U15192 (N_15192,N_11050,N_14551);
nor U15193 (N_15193,N_14031,N_12893);
nor U15194 (N_15194,N_13288,N_10539);
nand U15195 (N_15195,N_12847,N_10420);
xnor U15196 (N_15196,N_10732,N_14202);
and U15197 (N_15197,N_14040,N_11693);
nor U15198 (N_15198,N_10589,N_12042);
nor U15199 (N_15199,N_11987,N_10172);
and U15200 (N_15200,N_14112,N_13685);
xor U15201 (N_15201,N_13593,N_12481);
and U15202 (N_15202,N_10590,N_14538);
xnor U15203 (N_15203,N_11232,N_11676);
nand U15204 (N_15204,N_12616,N_10689);
and U15205 (N_15205,N_14239,N_14189);
nor U15206 (N_15206,N_14061,N_10169);
nand U15207 (N_15207,N_10945,N_10405);
nor U15208 (N_15208,N_13949,N_13053);
and U15209 (N_15209,N_11532,N_14198);
xnor U15210 (N_15210,N_11219,N_11972);
nand U15211 (N_15211,N_12446,N_10558);
nand U15212 (N_15212,N_13260,N_11353);
nand U15213 (N_15213,N_14768,N_11423);
or U15214 (N_15214,N_10446,N_14412);
xor U15215 (N_15215,N_14564,N_13366);
xnor U15216 (N_15216,N_13336,N_14818);
and U15217 (N_15217,N_14101,N_12577);
and U15218 (N_15218,N_12048,N_14268);
xor U15219 (N_15219,N_12094,N_13576);
or U15220 (N_15220,N_14114,N_11215);
and U15221 (N_15221,N_14103,N_13989);
and U15222 (N_15222,N_11835,N_13736);
and U15223 (N_15223,N_14745,N_11395);
and U15224 (N_15224,N_10150,N_12566);
xnor U15225 (N_15225,N_14878,N_13973);
nor U15226 (N_15226,N_10901,N_11929);
or U15227 (N_15227,N_12247,N_11218);
or U15228 (N_15228,N_13203,N_10635);
or U15229 (N_15229,N_14088,N_12776);
or U15230 (N_15230,N_11999,N_10509);
xor U15231 (N_15231,N_14131,N_11873);
or U15232 (N_15232,N_11444,N_11843);
xor U15233 (N_15233,N_10663,N_14197);
or U15234 (N_15234,N_11985,N_13964);
and U15235 (N_15235,N_11525,N_10430);
xor U15236 (N_15236,N_11126,N_11660);
and U15237 (N_15237,N_14446,N_13339);
xnor U15238 (N_15238,N_10479,N_12751);
nor U15239 (N_15239,N_14252,N_12904);
xnor U15240 (N_15240,N_13656,N_12991);
xnor U15241 (N_15241,N_14774,N_11029);
and U15242 (N_15242,N_12391,N_12975);
nand U15243 (N_15243,N_10571,N_13792);
or U15244 (N_15244,N_11283,N_12204);
and U15245 (N_15245,N_13231,N_13572);
nor U15246 (N_15246,N_12329,N_14025);
xnor U15247 (N_15247,N_11786,N_14639);
xor U15248 (N_15248,N_13201,N_13185);
nor U15249 (N_15249,N_13031,N_10203);
or U15250 (N_15250,N_11148,N_12239);
nand U15251 (N_15251,N_10990,N_11465);
xor U15252 (N_15252,N_13934,N_13573);
and U15253 (N_15253,N_14281,N_13627);
or U15254 (N_15254,N_12172,N_14802);
nand U15255 (N_15255,N_11784,N_14494);
nor U15256 (N_15256,N_13557,N_12862);
or U15257 (N_15257,N_14902,N_12655);
xor U15258 (N_15258,N_10013,N_11073);
nand U15259 (N_15259,N_10360,N_13771);
and U15260 (N_15260,N_13450,N_11143);
and U15261 (N_15261,N_11274,N_13818);
or U15262 (N_15262,N_13923,N_12138);
and U15263 (N_15263,N_10534,N_10288);
xor U15264 (N_15264,N_14582,N_12425);
nor U15265 (N_15265,N_10687,N_14621);
xor U15266 (N_15266,N_11839,N_13534);
nand U15267 (N_15267,N_13150,N_10449);
xor U15268 (N_15268,N_13320,N_10969);
and U15269 (N_15269,N_13710,N_12416);
nand U15270 (N_15270,N_14756,N_11198);
xor U15271 (N_15271,N_10098,N_12294);
or U15272 (N_15272,N_11897,N_14991);
or U15273 (N_15273,N_13170,N_11313);
nor U15274 (N_15274,N_11428,N_14539);
nand U15275 (N_15275,N_12015,N_10876);
and U15276 (N_15276,N_13359,N_11342);
or U15277 (N_15277,N_11358,N_13300);
nor U15278 (N_15278,N_10580,N_10928);
xor U15279 (N_15279,N_12354,N_12766);
nand U15280 (N_15280,N_14405,N_14882);
nand U15281 (N_15281,N_13158,N_12538);
xor U15282 (N_15282,N_14793,N_13143);
nor U15283 (N_15283,N_10533,N_12155);
nor U15284 (N_15284,N_11094,N_11881);
or U15285 (N_15285,N_12005,N_11036);
or U15286 (N_15286,N_13731,N_11382);
xor U15287 (N_15287,N_12197,N_13212);
nand U15288 (N_15288,N_13507,N_11776);
or U15289 (N_15289,N_12558,N_13561);
and U15290 (N_15290,N_13718,N_14985);
nand U15291 (N_15291,N_12789,N_14643);
nor U15292 (N_15292,N_13532,N_12322);
nand U15293 (N_15293,N_10338,N_13154);
nand U15294 (N_15294,N_12673,N_11832);
xnor U15295 (N_15295,N_13418,N_10543);
or U15296 (N_15296,N_13827,N_10349);
nor U15297 (N_15297,N_10147,N_12549);
nand U15298 (N_15298,N_11149,N_11325);
nor U15299 (N_15299,N_10679,N_14009);
and U15300 (N_15300,N_10071,N_14333);
nor U15301 (N_15301,N_12092,N_12278);
xor U15302 (N_15302,N_14466,N_14419);
and U15303 (N_15303,N_13437,N_11421);
xnor U15304 (N_15304,N_10903,N_12955);
and U15305 (N_15305,N_11937,N_12308);
and U15306 (N_15306,N_13654,N_11931);
xor U15307 (N_15307,N_14426,N_12262);
and U15308 (N_15308,N_14498,N_14140);
or U15309 (N_15309,N_14614,N_11847);
nand U15310 (N_15310,N_13925,N_13536);
nor U15311 (N_15311,N_13057,N_13972);
and U15312 (N_15312,N_12460,N_14855);
nand U15313 (N_15313,N_11888,N_14153);
nor U15314 (N_15314,N_12764,N_12754);
nand U15315 (N_15315,N_14442,N_11643);
nor U15316 (N_15316,N_10462,N_12109);
xor U15317 (N_15317,N_11397,N_10961);
nand U15318 (N_15318,N_14905,N_11404);
and U15319 (N_15319,N_14535,N_13114);
and U15320 (N_15320,N_10145,N_13752);
nor U15321 (N_15321,N_13890,N_12373);
and U15322 (N_15322,N_13018,N_14449);
and U15323 (N_15323,N_12250,N_14157);
nand U15324 (N_15324,N_11299,N_14337);
xor U15325 (N_15325,N_10820,N_12997);
and U15326 (N_15326,N_12833,N_14835);
xor U15327 (N_15327,N_10972,N_11539);
and U15328 (N_15328,N_14454,N_12622);
or U15329 (N_15329,N_10500,N_14801);
and U15330 (N_15330,N_13246,N_12993);
or U15331 (N_15331,N_10854,N_11066);
or U15332 (N_15332,N_12114,N_13005);
or U15333 (N_15333,N_12951,N_12856);
and U15334 (N_15334,N_11666,N_12340);
nand U15335 (N_15335,N_13904,N_10043);
or U15336 (N_15336,N_14482,N_14886);
or U15337 (N_15337,N_10999,N_11677);
nand U15338 (N_15338,N_11665,N_14250);
nor U15339 (N_15339,N_10407,N_14218);
or U15340 (N_15340,N_14152,N_10565);
nand U15341 (N_15341,N_12488,N_13938);
nand U15342 (N_15342,N_10140,N_12604);
and U15343 (N_15343,N_14850,N_14929);
nand U15344 (N_15344,N_11567,N_10240);
nor U15345 (N_15345,N_13043,N_13634);
or U15346 (N_15346,N_10074,N_14472);
xnor U15347 (N_15347,N_13564,N_14050);
nor U15348 (N_15348,N_10604,N_11398);
and U15349 (N_15349,N_13297,N_13773);
or U15350 (N_15350,N_10486,N_13473);
or U15351 (N_15351,N_12285,N_10202);
and U15352 (N_15352,N_13377,N_10456);
and U15353 (N_15353,N_11440,N_10222);
nor U15354 (N_15354,N_12125,N_14936);
xnor U15355 (N_15355,N_14743,N_14508);
xor U15356 (N_15356,N_11540,N_11189);
nor U15357 (N_15357,N_13676,N_11755);
nor U15358 (N_15358,N_14257,N_11829);
or U15359 (N_15359,N_11635,N_10770);
and U15360 (N_15360,N_14297,N_14360);
nor U15361 (N_15361,N_10656,N_14020);
and U15362 (N_15362,N_13173,N_12543);
nor U15363 (N_15363,N_11757,N_10844);
nor U15364 (N_15364,N_12699,N_14838);
nor U15365 (N_15365,N_13007,N_11741);
and U15366 (N_15366,N_13867,N_11427);
and U15367 (N_15367,N_10883,N_10158);
nand U15368 (N_15368,N_12788,N_11262);
nand U15369 (N_15369,N_13488,N_14617);
xor U15370 (N_15370,N_14366,N_11515);
nand U15371 (N_15371,N_12206,N_10015);
xor U15372 (N_15372,N_14350,N_14945);
or U15373 (N_15373,N_14355,N_12288);
or U15374 (N_15374,N_11716,N_12606);
or U15375 (N_15375,N_13219,N_13509);
nor U15376 (N_15376,N_11583,N_10957);
or U15377 (N_15377,N_11458,N_14019);
nand U15378 (N_15378,N_12877,N_14738);
nor U15379 (N_15379,N_10409,N_10746);
and U15380 (N_15380,N_14572,N_12056);
nand U15381 (N_15381,N_10011,N_10593);
nor U15382 (N_15382,N_10392,N_11302);
or U15383 (N_15383,N_11728,N_11890);
xor U15384 (N_15384,N_13861,N_11141);
xor U15385 (N_15385,N_11912,N_12696);
nand U15386 (N_15386,N_10906,N_14637);
nor U15387 (N_15387,N_14527,N_12773);
or U15388 (N_15388,N_14713,N_10309);
xor U15389 (N_15389,N_14497,N_11824);
nor U15390 (N_15390,N_12656,N_14866);
nor U15391 (N_15391,N_11098,N_14555);
nand U15392 (N_15392,N_13842,N_11920);
or U15393 (N_15393,N_13957,N_14893);
or U15394 (N_15394,N_13424,N_13119);
or U15395 (N_15395,N_12845,N_10971);
and U15396 (N_15396,N_14587,N_12621);
xor U15397 (N_15397,N_10067,N_11502);
nand U15398 (N_15398,N_11706,N_14222);
nor U15399 (N_15399,N_13375,N_13296);
and U15400 (N_15400,N_11116,N_12364);
nand U15401 (N_15401,N_14773,N_12212);
nand U15402 (N_15402,N_13592,N_11963);
nor U15403 (N_15403,N_10707,N_14294);
xor U15404 (N_15404,N_11979,N_13127);
or U15405 (N_15405,N_14459,N_13454);
xnor U15406 (N_15406,N_12080,N_12333);
nand U15407 (N_15407,N_12670,N_14383);
or U15408 (N_15408,N_13786,N_10866);
or U15409 (N_15409,N_14335,N_13419);
nand U15410 (N_15410,N_14007,N_14477);
or U15411 (N_15411,N_13629,N_10369);
and U15412 (N_15412,N_14432,N_13503);
nand U15413 (N_15413,N_13528,N_12190);
and U15414 (N_15414,N_12073,N_12229);
and U15415 (N_15415,N_11346,N_13817);
or U15416 (N_15416,N_14741,N_13669);
nor U15417 (N_15417,N_12189,N_13538);
and U15418 (N_15418,N_12309,N_13781);
nor U15419 (N_15419,N_12762,N_11740);
nor U15420 (N_15420,N_12700,N_13215);
or U15421 (N_15421,N_14313,N_13226);
nand U15422 (N_15422,N_10919,N_14012);
nand U15423 (N_15423,N_14820,N_13208);
nor U15424 (N_15424,N_13157,N_10598);
xor U15425 (N_15425,N_10167,N_14467);
nor U15426 (N_15426,N_11874,N_11366);
or U15427 (N_15427,N_11595,N_11183);
nor U15428 (N_15428,N_11156,N_12086);
nor U15429 (N_15429,N_14947,N_13798);
xnor U15430 (N_15430,N_13527,N_13796);
nor U15431 (N_15431,N_14828,N_10767);
nor U15432 (N_15432,N_13019,N_10302);
nand U15433 (N_15433,N_12062,N_12217);
and U15434 (N_15434,N_14182,N_11329);
xor U15435 (N_15435,N_12046,N_13524);
xor U15436 (N_15436,N_14908,N_11271);
and U15437 (N_15437,N_12735,N_10012);
or U15438 (N_15438,N_10246,N_13530);
nand U15439 (N_15439,N_10375,N_14147);
xnor U15440 (N_15440,N_14990,N_10299);
nand U15441 (N_15441,N_11615,N_14106);
nor U15442 (N_15442,N_11780,N_13717);
or U15443 (N_15443,N_13394,N_14054);
xnor U15444 (N_15444,N_14394,N_12055);
or U15445 (N_15445,N_12120,N_11766);
nor U15446 (N_15446,N_14409,N_11737);
and U15447 (N_15447,N_14896,N_12858);
and U15448 (N_15448,N_12544,N_12891);
xnor U15449 (N_15449,N_13317,N_13001);
nor U15450 (N_15450,N_12718,N_14762);
nand U15451 (N_15451,N_12698,N_10930);
and U15452 (N_15452,N_12519,N_11343);
or U15453 (N_15453,N_13956,N_13560);
and U15454 (N_15454,N_13663,N_14563);
xor U15455 (N_15455,N_12282,N_14674);
or U15456 (N_15456,N_11831,N_10822);
and U15457 (N_15457,N_11240,N_12300);
and U15458 (N_15458,N_10986,N_12482);
and U15459 (N_15459,N_14327,N_11768);
or U15460 (N_15460,N_10410,N_13596);
nand U15461 (N_15461,N_14378,N_12067);
nor U15462 (N_15462,N_14813,N_14652);
xnor U15463 (N_15463,N_11949,N_13191);
and U15464 (N_15464,N_12730,N_10877);
nor U15465 (N_15465,N_10815,N_14986);
nand U15466 (N_15466,N_12814,N_14119);
and U15467 (N_15467,N_11752,N_14964);
or U15468 (N_15468,N_11811,N_14373);
nor U15469 (N_15469,N_14511,N_13908);
nand U15470 (N_15470,N_10346,N_13689);
and U15471 (N_15471,N_14792,N_11093);
xnor U15472 (N_15472,N_12084,N_12447);
nand U15473 (N_15473,N_12287,N_12458);
and U15474 (N_15474,N_13218,N_10152);
nand U15475 (N_15475,N_12952,N_14399);
nand U15476 (N_15476,N_13599,N_11800);
xnor U15477 (N_15477,N_14249,N_11188);
nor U15478 (N_15478,N_13969,N_14190);
nand U15479 (N_15479,N_12794,N_13373);
nand U15480 (N_15480,N_14330,N_12224);
xnor U15481 (N_15481,N_10343,N_10136);
nor U15482 (N_15482,N_14663,N_14966);
and U15483 (N_15483,N_12792,N_11169);
nor U15484 (N_15484,N_14862,N_10287);
nand U15485 (N_15485,N_11469,N_11909);
xnor U15486 (N_15486,N_10646,N_12855);
xnor U15487 (N_15487,N_10133,N_13978);
or U15488 (N_15488,N_14478,N_10457);
or U15489 (N_15489,N_14853,N_13840);
and U15490 (N_15490,N_14684,N_13705);
xor U15491 (N_15491,N_12343,N_11151);
nand U15492 (N_15492,N_13584,N_11005);
nand U15493 (N_15493,N_10819,N_14410);
and U15494 (N_15494,N_12771,N_13164);
or U15495 (N_15495,N_10621,N_13683);
and U15496 (N_15496,N_14894,N_10776);
or U15497 (N_15497,N_11359,N_13006);
nor U15498 (N_15498,N_10588,N_10454);
or U15499 (N_15499,N_11416,N_13302);
or U15500 (N_15500,N_13673,N_14136);
and U15501 (N_15501,N_11808,N_12469);
nand U15502 (N_15502,N_14686,N_14094);
nand U15503 (N_15503,N_11935,N_14557);
nand U15504 (N_15504,N_10115,N_11180);
xnor U15505 (N_15505,N_10891,N_11297);
nand U15506 (N_15506,N_11788,N_12584);
and U15507 (N_15507,N_11074,N_11162);
or U15508 (N_15508,N_14787,N_12203);
or U15509 (N_15509,N_10282,N_13766);
or U15510 (N_15510,N_10982,N_11088);
nor U15511 (N_15511,N_11580,N_11704);
nor U15512 (N_15512,N_11489,N_12804);
nor U15513 (N_15513,N_12401,N_13678);
xor U15514 (N_15514,N_14474,N_10076);
nand U15515 (N_15515,N_14354,N_11739);
xor U15516 (N_15516,N_12298,N_13285);
and U15517 (N_15517,N_12559,N_12746);
nand U15518 (N_15518,N_13052,N_10391);
or U15519 (N_15519,N_12240,N_10900);
or U15520 (N_15520,N_10857,N_10226);
nand U15521 (N_15521,N_10636,N_13954);
nor U15522 (N_15522,N_11659,N_12913);
and U15523 (N_15523,N_10038,N_14417);
or U15524 (N_15524,N_11105,N_10960);
xnor U15525 (N_15525,N_13589,N_14702);
nor U15526 (N_15526,N_13287,N_13074);
or U15527 (N_15527,N_11109,N_14951);
and U15528 (N_15528,N_11927,N_12557);
nor U15529 (N_15529,N_11461,N_11474);
or U15530 (N_15530,N_13788,N_12014);
and U15531 (N_15531,N_13476,N_13876);
nand U15532 (N_15532,N_10219,N_12595);
nor U15533 (N_15533,N_13868,N_11528);
nor U15534 (N_15534,N_10907,N_12651);
xnor U15535 (N_15535,N_11490,N_13124);
or U15536 (N_15536,N_11682,N_12742);
and U15537 (N_15537,N_10089,N_12423);
nor U15538 (N_15538,N_14403,N_12964);
xnor U15539 (N_15539,N_13623,N_10261);
xnor U15540 (N_15540,N_13784,N_10688);
nand U15541 (N_15541,N_12611,N_11983);
nand U15542 (N_15542,N_13380,N_13042);
or U15543 (N_15543,N_12648,N_14944);
xnor U15544 (N_15544,N_11125,N_11177);
xnor U15545 (N_15545,N_12328,N_11411);
nand U15546 (N_15546,N_14544,N_14556);
or U15547 (N_15547,N_13233,N_10652);
nand U15548 (N_15548,N_13649,N_14406);
and U15549 (N_15549,N_10438,N_13066);
and U15550 (N_15550,N_12967,N_12226);
nor U15551 (N_15551,N_10267,N_14673);
or U15552 (N_15552,N_11235,N_11376);
or U15553 (N_15553,N_13603,N_12678);
nor U15554 (N_15554,N_13775,N_13912);
and U15555 (N_15555,N_10054,N_10867);
or U15556 (N_15556,N_12219,N_10326);
nor U15557 (N_15557,N_14679,N_10105);
or U15558 (N_15558,N_13675,N_11224);
nor U15559 (N_15559,N_12111,N_13657);
nand U15560 (N_15560,N_12860,N_10244);
nor U15561 (N_15561,N_14634,N_11208);
xor U15562 (N_15562,N_14460,N_10220);
or U15563 (N_15563,N_13499,N_11229);
nor U15564 (N_15564,N_12812,N_13739);
or U15565 (N_15565,N_10572,N_10805);
xor U15566 (N_15566,N_10991,N_11804);
and U15567 (N_15567,N_13602,N_12380);
or U15568 (N_15568,N_13984,N_14471);
nor U15569 (N_15569,N_10893,N_13738);
and U15570 (N_15570,N_13193,N_13082);
nand U15571 (N_15571,N_14204,N_13055);
or U15572 (N_15572,N_11834,N_10499);
or U15573 (N_15573,N_14369,N_14687);
nand U15574 (N_15574,N_14913,N_12183);
xnor U15575 (N_15575,N_14962,N_13166);
xnor U15576 (N_15576,N_14380,N_12161);
or U15577 (N_15577,N_14598,N_12357);
nor U15578 (N_15578,N_12938,N_11585);
or U15579 (N_15579,N_14411,N_14719);
nand U15580 (N_15580,N_13358,N_14586);
nand U15581 (N_15581,N_13748,N_13812);
and U15582 (N_15582,N_12457,N_13456);
or U15583 (N_15583,N_11389,N_14909);
xor U15584 (N_15584,N_13674,N_11966);
nand U15585 (N_15585,N_11312,N_14829);
or U15586 (N_15586,N_12803,N_13898);
or U15587 (N_15587,N_13955,N_12963);
and U15588 (N_15588,N_13648,N_10774);
nor U15589 (N_15589,N_13910,N_11577);
xnor U15590 (N_15590,N_12390,N_14181);
and U15591 (N_15591,N_14566,N_10185);
and U15592 (N_15592,N_11875,N_13677);
nor U15593 (N_15593,N_10874,N_13243);
or U15594 (N_15594,N_12269,N_10289);
nor U15595 (N_15595,N_14876,N_10127);
nand U15596 (N_15596,N_12571,N_14992);
xor U15597 (N_15597,N_10125,N_10498);
nand U15598 (N_15598,N_11899,N_13836);
and U15599 (N_15599,N_14423,N_12756);
nand U15600 (N_15600,N_14895,N_11760);
and U15601 (N_15601,N_13051,N_14517);
or U15602 (N_15602,N_11498,N_11928);
nand U15603 (N_15603,N_11364,N_10268);
or U15604 (N_15604,N_14761,N_13077);
nor U15605 (N_15605,N_14151,N_12827);
nor U15606 (N_15606,N_13624,N_11403);
or U15607 (N_15607,N_13617,N_13408);
xor U15608 (N_15608,N_11626,N_13023);
or U15609 (N_15609,N_10601,N_12324);
nand U15610 (N_15610,N_10995,N_13998);
and U15611 (N_15611,N_12451,N_14897);
and U15612 (N_15612,N_12296,N_10847);
or U15613 (N_15613,N_11893,N_14892);
nor U15614 (N_15614,N_11306,N_11076);
and U15615 (N_15615,N_14796,N_13690);
nand U15616 (N_15616,N_12507,N_13828);
and U15617 (N_15617,N_12727,N_12502);
nor U15618 (N_15618,N_14826,N_13940);
and U15619 (N_15619,N_11158,N_14359);
or U15620 (N_15620,N_10521,N_13307);
xnor U15621 (N_15621,N_14000,N_11068);
nor U15622 (N_15622,N_10817,N_13126);
and U15623 (N_15623,N_11405,N_12917);
and U15624 (N_15624,N_12588,N_11394);
nor U15625 (N_15625,N_14946,N_10000);
and U15626 (N_15626,N_13278,N_14798);
xor U15627 (N_15627,N_13782,N_12205);
nor U15628 (N_15628,N_13284,N_12920);
nor U15629 (N_15629,N_13498,N_14255);
nand U15630 (N_15630,N_12277,N_13682);
nand U15631 (N_15631,N_14208,N_14970);
and U15632 (N_15632,N_10976,N_11494);
nor U15633 (N_15633,N_13884,N_11549);
nand U15634 (N_15634,N_10525,N_12940);
nand U15635 (N_15635,N_10120,N_14830);
or U15636 (N_15636,N_13038,N_14044);
nand U15637 (N_15637,N_11634,N_10795);
or U15638 (N_15638,N_12816,N_14868);
nand U15639 (N_15639,N_11513,N_10758);
nand U15640 (N_15640,N_14270,N_10541);
nor U15641 (N_15641,N_11655,N_13298);
and U15642 (N_15642,N_12851,N_13725);
nor U15643 (N_15643,N_10826,N_11946);
nand U15644 (N_15644,N_10745,N_14512);
xor U15645 (N_15645,N_13911,N_10929);
nand U15646 (N_15646,N_12602,N_11586);
or U15647 (N_15647,N_13971,N_11167);
or U15648 (N_15648,N_10083,N_11062);
or U15649 (N_15649,N_11316,N_12180);
or U15650 (N_15650,N_13483,N_11134);
nor U15651 (N_15651,N_13381,N_10488);
nand U15652 (N_15652,N_11310,N_13293);
and U15653 (N_15653,N_14717,N_10394);
or U15654 (N_15654,N_12066,N_13546);
or U15655 (N_15655,N_10649,N_14641);
nor U15656 (N_15656,N_11984,N_11255);
nor U15657 (N_15657,N_13734,N_11907);
or U15658 (N_15658,N_13655,N_11363);
nand U15659 (N_15659,N_12440,N_10804);
and U15660 (N_15660,N_10764,N_13044);
or U15661 (N_15661,N_13839,N_12103);
nor U15662 (N_15662,N_11708,N_10889);
nand U15663 (N_15663,N_13210,N_12045);
xor U15664 (N_15664,N_13120,N_12291);
nor U15665 (N_15665,N_14311,N_10317);
and U15666 (N_15666,N_10021,N_10017);
nor U15667 (N_15667,N_10393,N_14034);
xor U15668 (N_15668,N_13000,N_11697);
nand U15669 (N_15669,N_11825,N_11600);
or U15670 (N_15670,N_13264,N_13751);
nor U15671 (N_15671,N_13831,N_12159);
and U15672 (N_15672,N_10843,N_11372);
nor U15673 (N_15673,N_13601,N_12072);
nand U15674 (N_15674,N_12667,N_12411);
nor U15675 (N_15675,N_11259,N_11812);
xnor U15676 (N_15676,N_10755,N_12242);
nand U15677 (N_15677,N_13214,N_12388);
xnor U15678 (N_15678,N_14594,N_10913);
or U15679 (N_15679,N_13891,N_10518);
xor U15680 (N_15680,N_12631,N_11940);
nor U15681 (N_15681,N_12041,N_10295);
xor U15682 (N_15682,N_11083,N_13996);
or U15683 (N_15683,N_11182,N_14126);
nor U15684 (N_15684,N_10863,N_12743);
xnor U15685 (N_15685,N_13443,N_14654);
nor U15686 (N_15686,N_13301,N_14023);
or U15687 (N_15687,N_14008,N_13887);
xnor U15688 (N_15688,N_14760,N_14857);
and U15689 (N_15689,N_10485,N_12249);
and U15690 (N_15690,N_11419,N_14770);
nand U15691 (N_15691,N_14248,N_11850);
nor U15692 (N_15692,N_11747,N_12647);
xnor U15693 (N_15693,N_12409,N_13496);
and U15694 (N_15694,N_11967,N_14500);
xnor U15695 (N_15695,N_13417,N_12976);
nor U15696 (N_15696,N_13937,N_12899);
or U15697 (N_15697,N_13303,N_14553);
nand U15698 (N_15698,N_11335,N_14261);
nor U15699 (N_15699,N_13730,N_12442);
nand U15700 (N_15700,N_12707,N_13490);
or U15701 (N_15701,N_10283,N_12657);
or U15702 (N_15702,N_12471,N_14493);
xor U15703 (N_15703,N_11123,N_13354);
nand U15704 (N_15704,N_14264,N_12593);
and U15705 (N_15705,N_14521,N_11767);
xor U15706 (N_15706,N_13459,N_11978);
nand U15707 (N_15707,N_11137,N_11736);
xor U15708 (N_15708,N_11443,N_12290);
nand U15709 (N_15709,N_14914,N_14993);
and U15710 (N_15710,N_11206,N_14163);
nor U15711 (N_15711,N_11155,N_13980);
or U15712 (N_15712,N_10242,N_10677);
or U15713 (N_15713,N_11025,N_14245);
and U15714 (N_15714,N_12417,N_11826);
nor U15715 (N_15715,N_12927,N_10583);
and U15716 (N_15716,N_10107,N_13160);
and U15717 (N_15717,N_14575,N_12237);
and U15718 (N_15718,N_12868,N_12578);
xnor U15719 (N_15719,N_11432,N_12615);
xor U15720 (N_15720,N_12010,N_12671);
or U15721 (N_15721,N_13029,N_12116);
or U15722 (N_15722,N_10157,N_10304);
or U15723 (N_15723,N_14125,N_11015);
or U15724 (N_15724,N_13147,N_10497);
and U15725 (N_15725,N_12107,N_12126);
nand U15726 (N_15726,N_12626,N_14541);
or U15727 (N_15727,N_14532,N_11892);
nor U15728 (N_15728,N_10594,N_14976);
xor U15729 (N_15729,N_13508,N_10914);
nor U15730 (N_15730,N_12869,N_11048);
or U15731 (N_15731,N_13174,N_12065);
or U15732 (N_15732,N_12808,N_11522);
and U15733 (N_15733,N_12630,N_12077);
nand U15734 (N_15734,N_11043,N_13117);
xor U15735 (N_15735,N_10717,N_11355);
and U15736 (N_15736,N_13765,N_11544);
nor U15737 (N_15737,N_14416,N_12536);
and U15738 (N_15738,N_11209,N_14849);
nand U15739 (N_15739,N_13039,N_13385);
or U15740 (N_15740,N_13753,N_11377);
or U15741 (N_15741,N_14074,N_14998);
nor U15742 (N_15742,N_12801,N_13034);
or U15743 (N_15743,N_12838,N_11067);
or U15744 (N_15744,N_10808,N_11194);
nor U15745 (N_15745,N_14085,N_10714);
or U15746 (N_15746,N_13196,N_13586);
and U15747 (N_15747,N_14974,N_11533);
or U15748 (N_15748,N_11478,N_10181);
xor U15749 (N_15749,N_12949,N_14357);
nor U15750 (N_15750,N_12337,N_13387);
or U15751 (N_15751,N_13382,N_11318);
or U15752 (N_15752,N_11721,N_12866);
nor U15753 (N_15753,N_11894,N_14305);
xnor U15754 (N_15754,N_10342,N_13290);
xor U15755 (N_15755,N_13209,N_10785);
nand U15756 (N_15756,N_13763,N_10933);
xor U15757 (N_15757,N_10494,N_14549);
or U15758 (N_15758,N_13384,N_13684);
xnor U15759 (N_15759,N_14274,N_14138);
xor U15760 (N_15760,N_10018,N_14280);
or U15761 (N_15761,N_14922,N_12321);
nand U15762 (N_15762,N_12527,N_14904);
xor U15763 (N_15763,N_12311,N_13457);
xnor U15764 (N_15764,N_11569,N_10793);
nand U15765 (N_15765,N_11032,N_13525);
nor U15766 (N_15766,N_14027,N_14431);
nor U15767 (N_15767,N_14568,N_11506);
and U15768 (N_15768,N_11018,N_14194);
and U15769 (N_15769,N_14758,N_11186);
or U15770 (N_15770,N_11558,N_12158);
and U15771 (N_15771,N_14920,N_10207);
nand U15772 (N_15772,N_14919,N_12837);
xor U15773 (N_15773,N_13640,N_12880);
and U15774 (N_15774,N_14509,N_12688);
nor U15775 (N_15775,N_11724,N_10081);
nor U15776 (N_15776,N_10048,N_14167);
and U15777 (N_15777,N_13583,N_12270);
xnor U15778 (N_15778,N_10653,N_13744);
and U15779 (N_15779,N_12924,N_13360);
nand U15780 (N_15780,N_14601,N_11244);
nor U15781 (N_15781,N_13446,N_12091);
or U15782 (N_15782,N_10164,N_12129);
xnor U15783 (N_15783,N_12254,N_14884);
and U15784 (N_15784,N_12510,N_10078);
xnor U15785 (N_15785,N_14132,N_12036);
nor U15786 (N_15786,N_11883,N_11742);
or U15787 (N_15787,N_10542,N_10591);
nor U15788 (N_15788,N_12444,N_12115);
or U15789 (N_15789,N_12185,N_10979);
nand U15790 (N_15790,N_13658,N_10294);
nand U15791 (N_15791,N_13847,N_14488);
or U15792 (N_15792,N_12785,N_13016);
or U15793 (N_15793,N_13723,N_10227);
nor U15794 (N_15794,N_14097,N_11779);
and U15795 (N_15795,N_13668,N_12132);
and U15796 (N_15796,N_12740,N_10905);
nand U15797 (N_15797,N_14491,N_12382);
and U15798 (N_15798,N_11249,N_13445);
and U15799 (N_15799,N_12459,N_14971);
nand U15800 (N_15800,N_12884,N_10987);
nand U15801 (N_15801,N_13850,N_14166);
xor U15802 (N_15802,N_12995,N_13213);
or U15803 (N_15803,N_11925,N_12970);
or U15804 (N_15804,N_11070,N_13277);
or U15805 (N_15805,N_13720,N_12214);
xor U15806 (N_15806,N_11251,N_13050);
xor U15807 (N_15807,N_12818,N_14469);
and U15808 (N_15808,N_11857,N_12347);
xnor U15809 (N_15809,N_10735,N_13578);
and U15810 (N_15810,N_13379,N_13406);
xor U15811 (N_15811,N_13709,N_11564);
or U15812 (N_15812,N_11959,N_14953);
xnor U15813 (N_15813,N_11199,N_12130);
nor U15814 (N_15814,N_14695,N_11977);
or U15815 (N_15815,N_10293,N_12922);
or U15816 (N_15816,N_12252,N_13838);
nor U15817 (N_15817,N_10460,N_11236);
and U15818 (N_15818,N_11618,N_12499);
and U15819 (N_15819,N_12609,N_10639);
and U15820 (N_15820,N_10567,N_10123);
nor U15821 (N_15821,N_11192,N_11060);
and U15822 (N_15822,N_10345,N_13961);
nor U15823 (N_15823,N_12026,N_11340);
or U15824 (N_15824,N_11726,N_11166);
or U15825 (N_15825,N_10366,N_10070);
nor U15826 (N_15826,N_10216,N_11414);
and U15827 (N_15827,N_10812,N_13073);
xor U15828 (N_15828,N_12516,N_13309);
nand U15829 (N_15829,N_14206,N_10373);
and U15830 (N_15830,N_14242,N_14630);
nor U15831 (N_15831,N_14371,N_10441);
xnor U15832 (N_15832,N_13182,N_10631);
and U15833 (N_15833,N_13568,N_11848);
or U15834 (N_15834,N_14092,N_14603);
xnor U15835 (N_15835,N_13948,N_12642);
xor U15836 (N_15836,N_11459,N_13965);
nor U15837 (N_15837,N_10619,N_11114);
and U15838 (N_15838,N_12675,N_10121);
or U15839 (N_15839,N_14874,N_12767);
nand U15840 (N_15840,N_14616,N_10536);
nor U15841 (N_15841,N_10046,N_11644);
nor U15842 (N_15842,N_13764,N_14422);
nand U15843 (N_15843,N_11059,N_12724);
nand U15844 (N_15844,N_14595,N_12750);
nor U15845 (N_15845,N_14424,N_10401);
or U15846 (N_15846,N_13577,N_12225);
nor U15847 (N_15847,N_10153,N_12452);
and U15848 (N_15848,N_13825,N_13625);
nor U15849 (N_15849,N_11499,N_11027);
and U15850 (N_15850,N_12144,N_14045);
or U15851 (N_15851,N_12843,N_10728);
or U15852 (N_15852,N_10188,N_10175);
or U15853 (N_15853,N_11647,N_14624);
and U15854 (N_15854,N_13922,N_14742);
nor U15855 (N_15855,N_12307,N_14340);
nand U15856 (N_15856,N_13493,N_13813);
nor U15857 (N_15857,N_11948,N_10413);
and U15858 (N_15858,N_13612,N_10260);
nand U15859 (N_15859,N_10696,N_14324);
xor U15860 (N_15860,N_11527,N_11696);
xor U15861 (N_15861,N_13249,N_13939);
nand U15862 (N_15862,N_10578,N_12087);
nand U15863 (N_15863,N_12059,N_14217);
and U15864 (N_15864,N_10853,N_11152);
nor U15865 (N_15865,N_14089,N_10111);
nand U15866 (N_15866,N_13421,N_11713);
xnor U15867 (N_15867,N_10996,N_12708);
nor U15868 (N_15868,N_11797,N_13291);
or U15869 (N_15869,N_14385,N_10200);
and U15870 (N_15870,N_11160,N_11869);
or U15871 (N_15871,N_10699,N_11727);
nor U15872 (N_15872,N_10917,N_12495);
nor U15873 (N_15873,N_13745,N_14891);
xor U15874 (N_15874,N_11345,N_12016);
or U15875 (N_15875,N_14047,N_11645);
or U15876 (N_15876,N_13464,N_14933);
nor U15877 (N_15877,N_11971,N_12758);
nand U15878 (N_15878,N_12395,N_12148);
and U15879 (N_15879,N_12582,N_10209);
nand U15880 (N_15880,N_12537,N_14386);
nand U15881 (N_15881,N_14604,N_10331);
nand U15882 (N_15882,N_11153,N_12334);
nor U15883 (N_15883,N_14699,N_11511);
nand U15884 (N_15884,N_14292,N_11352);
xnor U15885 (N_15885,N_13787,N_14611);
and U15886 (N_15886,N_14858,N_14455);
nand U15887 (N_15887,N_12601,N_12053);
and U15888 (N_15888,N_13635,N_14547);
xnor U15889 (N_15889,N_10482,N_13686);
or U15890 (N_15890,N_14075,N_13853);
nand U15891 (N_15891,N_11065,N_11891);
nand U15892 (N_15892,N_10129,N_11058);
nor U15893 (N_15893,N_14636,N_11714);
or U15894 (N_15894,N_11594,N_14296);
nand U15895 (N_15895,N_11793,N_10415);
nand U15896 (N_15896,N_10340,N_13048);
and U15897 (N_15897,N_12532,N_14791);
nand U15898 (N_15898,N_13345,N_11576);
nand U15899 (N_15899,N_12836,N_12479);
or U15900 (N_15900,N_14869,N_11441);
or U15901 (N_15901,N_13701,N_13809);
or U15902 (N_15902,N_10501,N_12315);
nand U15903 (N_15903,N_12633,N_14465);
nor U15904 (N_15904,N_13338,N_11919);
xor U15905 (N_15905,N_14571,N_10694);
or U15906 (N_15906,N_11175,N_12503);
nor U15907 (N_15907,N_13047,N_12037);
nor U15908 (N_15908,N_13181,N_10718);
nor U15909 (N_15909,N_11968,N_10119);
nand U15910 (N_15910,N_14427,N_10313);
xnor U15911 (N_15911,N_11482,N_12534);
xnor U15912 (N_15912,N_12744,N_14515);
nor U15913 (N_15913,N_13451,N_12775);
nand U15914 (N_15914,N_12184,N_10684);
nand U15915 (N_15915,N_12717,N_10099);
nor U15916 (N_15916,N_14058,N_10697);
nand U15917 (N_15917,N_11625,N_14010);
and U15918 (N_15918,N_11849,N_12666);
xnor U15919 (N_15919,N_11276,N_14628);
and U15920 (N_15920,N_10506,N_13979);
nand U15921 (N_15921,N_11264,N_14718);
and U15922 (N_15922,N_13332,N_10842);
xor U15923 (N_15923,N_13777,N_11989);
xor U15924 (N_15924,N_14546,N_11268);
xnor U15925 (N_15925,N_12432,N_12890);
xnor U15926 (N_15926,N_13435,N_13945);
nand U15927 (N_15927,N_12236,N_13035);
xnor U15928 (N_15928,N_11038,N_14816);
nor U15929 (N_15929,N_10861,N_11331);
and U15930 (N_15930,N_14984,N_13704);
or U15931 (N_15931,N_13848,N_14480);
and U15932 (N_15932,N_13959,N_10659);
or U15933 (N_15933,N_10235,N_12320);
nor U15934 (N_15934,N_13378,N_11723);
nand U15935 (N_15935,N_11455,N_11260);
or U15936 (N_15936,N_12632,N_10620);
nand U15937 (N_15937,N_11460,N_10712);
and U15938 (N_15938,N_14276,N_14203);
or U15939 (N_15939,N_12231,N_14158);
nand U15940 (N_15940,N_13229,N_11632);
or U15941 (N_15941,N_12683,N_14965);
nor U15942 (N_15942,N_12520,N_11994);
nor U15943 (N_15943,N_10025,N_11636);
or U15944 (N_15944,N_10778,N_14172);
or U15945 (N_15945,N_10379,N_11962);
xnor U15946 (N_15946,N_13273,N_14086);
or U15947 (N_15947,N_14155,N_13981);
nor U15948 (N_15948,N_10114,N_13670);
xnor U15949 (N_15949,N_12317,N_10737);
nor U15950 (N_15950,N_14492,N_10773);
or U15951 (N_15951,N_10416,N_11082);
nor U15952 (N_15952,N_12119,N_14562);
xnor U15953 (N_15953,N_14435,N_13982);
nand U15954 (N_15954,N_14445,N_13449);
or U15955 (N_15955,N_10554,N_12984);
xor U15956 (N_15956,N_12165,N_12802);
xnor U15957 (N_15957,N_14180,N_13580);
nor U15958 (N_15958,N_10894,N_13846);
nor U15959 (N_15959,N_14588,N_14322);
or U15960 (N_15960,N_14087,N_13376);
and U15961 (N_15961,N_10865,N_12694);
xor U15962 (N_15962,N_10942,N_11486);
and U15963 (N_15963,N_14174,N_11765);
xor U15964 (N_15964,N_14880,N_13305);
xnor U15965 (N_15965,N_13845,N_12028);
or U15966 (N_15966,N_12674,N_13632);
xnor U15967 (N_15967,N_12003,N_12448);
nor U15968 (N_15968,N_11895,N_12907);
nor U15969 (N_15969,N_10547,N_11551);
or U15970 (N_15970,N_13025,N_14642);
and U15971 (N_15971,N_14994,N_14127);
and U15972 (N_15972,N_12526,N_12258);
and U15973 (N_15973,N_12954,N_10729);
and U15974 (N_15974,N_14444,N_12823);
xnor U15975 (N_15975,N_10918,N_12177);
or U15976 (N_15976,N_10595,N_11099);
nor U15977 (N_15977,N_11165,N_14213);
xnor U15978 (N_15978,N_10909,N_14068);
or U15979 (N_15979,N_14827,N_11572);
xnor U15980 (N_15980,N_13466,N_10073);
and U15981 (N_15981,N_13228,N_11537);
nor U15982 (N_15982,N_12345,N_11684);
xnor U15983 (N_15983,N_13187,N_10532);
nand U15984 (N_15984,N_12406,N_14569);
nor U15985 (N_15985,N_14302,N_10810);
and U15986 (N_15986,N_12484,N_11668);
or U15987 (N_15987,N_13340,N_10837);
nand U15988 (N_15988,N_10045,N_14821);
and U15989 (N_15989,N_10897,N_12259);
xnor U15990 (N_15990,N_11896,N_11866);
and U15991 (N_15991,N_10833,N_14262);
xnor U15992 (N_15992,N_11656,N_12088);
nand U15993 (N_15993,N_10841,N_13312);
xor U15994 (N_15994,N_12906,N_13136);
nor U15995 (N_15995,N_13310,N_13914);
or U15996 (N_15996,N_11604,N_10024);
nor U15997 (N_15997,N_13698,N_12198);
nand U15998 (N_15998,N_14219,N_11031);
or U15999 (N_15999,N_10189,N_12824);
nand U16000 (N_16000,N_11542,N_10613);
nor U16001 (N_16001,N_11009,N_12905);
and U16002 (N_16002,N_14754,N_11196);
or U16003 (N_16003,N_11853,N_13768);
nand U16004 (N_16004,N_10870,N_13562);
nand U16005 (N_16005,N_10934,N_11449);
nand U16006 (N_16006,N_13543,N_13975);
or U16007 (N_16007,N_14030,N_12052);
and U16008 (N_16008,N_10705,N_13167);
nand U16009 (N_16009,N_12734,N_11534);
xor U16010 (N_16010,N_11496,N_13433);
nor U16011 (N_16011,N_14644,N_12179);
nand U16012 (N_16012,N_10587,N_14843);
xor U16013 (N_16013,N_13272,N_11493);
and U16014 (N_16014,N_14196,N_12805);
nor U16015 (N_16015,N_11884,N_14076);
xnor U16016 (N_16016,N_14267,N_12859);
or U16017 (N_16017,N_11621,N_13636);
and U16018 (N_16018,N_12480,N_11733);
and U16019 (N_16019,N_14317,N_14915);
nor U16020 (N_16020,N_10881,N_10165);
nand U16021 (N_16021,N_13361,N_11004);
nor U16022 (N_16022,N_12178,N_13571);
and U16023 (N_16023,N_14247,N_13370);
nand U16024 (N_16024,N_11000,N_10256);
nand U16025 (N_16025,N_13590,N_12921);
or U16026 (N_16026,N_14156,N_14082);
or U16027 (N_16027,N_13924,N_10824);
or U16028 (N_16028,N_12063,N_12883);
and U16029 (N_16029,N_12506,N_13362);
xor U16030 (N_16030,N_11448,N_11293);
nor U16031 (N_16031,N_12719,N_14273);
nor U16032 (N_16032,N_11778,N_11488);
or U16033 (N_16033,N_12449,N_10711);
or U16034 (N_16034,N_11021,N_13145);
or U16035 (N_16035,N_12672,N_12878);
and U16036 (N_16036,N_14982,N_11154);
nor U16037 (N_16037,N_11601,N_13033);
or U16038 (N_16038,N_11409,N_12372);
nor U16039 (N_16039,N_10270,N_12738);
and U16040 (N_16040,N_13097,N_11619);
nand U16041 (N_16041,N_14649,N_14233);
nand U16042 (N_16042,N_11921,N_13223);
or U16043 (N_16043,N_12649,N_10834);
nor U16044 (N_16044,N_10212,N_13333);
nor U16045 (N_16045,N_13068,N_10258);
xor U16046 (N_16046,N_14149,N_12676);
xor U16047 (N_16047,N_11550,N_13027);
nor U16048 (N_16048,N_10080,N_14483);
or U16049 (N_16049,N_11593,N_10757);
or U16050 (N_16050,N_12829,N_13063);
nand U16051 (N_16051,N_11320,N_10628);
nand U16052 (N_16052,N_14854,N_12521);
and U16053 (N_16053,N_10634,N_14379);
and U16054 (N_16054,N_10756,N_14698);
nand U16055 (N_16055,N_10703,N_13628);
xor U16056 (N_16056,N_10075,N_11356);
and U16057 (N_16057,N_11227,N_12043);
and U16058 (N_16058,N_11011,N_12303);
nand U16059 (N_16059,N_11091,N_12098);
nor U16060 (N_16060,N_12942,N_13211);
and U16061 (N_16061,N_12564,N_14640);
nor U16062 (N_16062,N_13594,N_14903);
nor U16063 (N_16063,N_12702,N_12478);
or U16064 (N_16064,N_14154,N_10278);
nor U16065 (N_16065,N_13587,N_10149);
and U16066 (N_16066,N_12950,N_14709);
nand U16067 (N_16067,N_12413,N_14887);
xor U16068 (N_16068,N_14015,N_14696);
nand U16069 (N_16069,N_10466,N_10178);
xor U16070 (N_16070,N_14524,N_12844);
nand U16071 (N_16071,N_13515,N_12625);
nor U16072 (N_16072,N_12079,N_14671);
or U16073 (N_16073,N_13830,N_14115);
nor U16074 (N_16074,N_11798,N_12514);
or U16075 (N_16075,N_13517,N_10180);
xor U16076 (N_16076,N_14958,N_11915);
or U16077 (N_16077,N_11650,N_14954);
nor U16078 (N_16078,N_10388,N_11947);
nand U16079 (N_16079,N_14496,N_14889);
and U16080 (N_16080,N_13263,N_10848);
xor U16081 (N_16081,N_13505,N_11686);
and U16082 (N_16082,N_10949,N_11090);
nor U16083 (N_16083,N_11334,N_14229);
and U16084 (N_16084,N_13609,N_14706);
nor U16085 (N_16085,N_10487,N_10680);
nand U16086 (N_16086,N_13719,N_12335);
and U16087 (N_16087,N_14782,N_11950);
and U16088 (N_16088,N_13148,N_12191);
xor U16089 (N_16089,N_14786,N_12591);
nand U16090 (N_16090,N_10491,N_12722);
xor U16091 (N_16091,N_10265,N_12418);
nand U16092 (N_16092,N_13616,N_14980);
nor U16093 (N_16093,N_11161,N_11247);
nor U16094 (N_16094,N_10103,N_13974);
xnor U16095 (N_16095,N_11379,N_10708);
and U16096 (N_16096,N_10030,N_10618);
or U16097 (N_16097,N_10932,N_12590);
nor U16098 (N_16098,N_14540,N_11311);
nand U16099 (N_16099,N_11484,N_12594);
nand U16100 (N_16100,N_10693,N_14856);
nor U16101 (N_16101,N_12305,N_12462);
nor U16102 (N_16102,N_12035,N_14672);
nand U16103 (N_16103,N_10784,N_14703);
nand U16104 (N_16104,N_14918,N_10428);
xnor U16105 (N_16105,N_13030,N_11485);
and U16106 (N_16106,N_11055,N_10997);
nand U16107 (N_16107,N_11840,N_14823);
nor U16108 (N_16108,N_13061,N_13976);
and U16109 (N_16109,N_10062,N_10221);
or U16110 (N_16110,N_14259,N_13328);
nor U16111 (N_16111,N_14499,N_11579);
nand U16112 (N_16112,N_11942,N_11622);
xor U16113 (N_16113,N_11017,N_13900);
and U16114 (N_16114,N_10576,N_14216);
nand U16115 (N_16115,N_14522,N_11307);
nor U16116 (N_16116,N_13236,N_13795);
nor U16117 (N_16117,N_13465,N_10031);
or U16118 (N_16118,N_10436,N_11900);
xnor U16119 (N_16119,N_11370,N_11842);
or U16120 (N_16120,N_10947,N_13420);
or U16121 (N_16121,N_14284,N_12703);
nor U16122 (N_16122,N_13991,N_13863);
xnor U16123 (N_16123,N_10952,N_10455);
and U16124 (N_16124,N_13012,N_11012);
or U16125 (N_16125,N_12979,N_14657);
or U16126 (N_16126,N_11863,N_14318);
nand U16127 (N_16127,N_13645,N_12358);
and U16128 (N_16128,N_11195,N_10332);
xor U16129 (N_16129,N_10850,N_11020);
xnor U16130 (N_16130,N_10271,N_14906);
xnor U16131 (N_16131,N_12466,N_12221);
xor U16132 (N_16132,N_11877,N_13299);
nand U16133 (N_16133,N_12136,N_10439);
and U16134 (N_16134,N_14026,N_11212);
nor U16135 (N_16135,N_13882,N_11980);
and U16136 (N_16136,N_13369,N_10469);
nor U16137 (N_16137,N_10386,N_14241);
and U16138 (N_16138,N_14057,N_14004);
nand U16139 (N_16139,N_14968,N_13441);
nand U16140 (N_16140,N_11879,N_11654);
nor U16141 (N_16141,N_12068,N_10396);
or U16142 (N_16142,N_14220,N_12810);
or U16143 (N_16143,N_10403,N_11790);
nand U16144 (N_16144,N_14374,N_11801);
nand U16145 (N_16145,N_10275,N_12882);
or U16146 (N_16146,N_11362,N_12528);
xor U16147 (N_16147,N_11633,N_14429);
nor U16148 (N_16148,N_13889,N_14618);
xor U16149 (N_16149,N_11252,N_13661);
xnor U16150 (N_16150,N_11092,N_11658);
or U16151 (N_16151,N_10088,N_11328);
or U16152 (N_16152,N_13142,N_10759);
nand U16153 (N_16153,N_10638,N_12496);
xnor U16154 (N_16154,N_14315,N_14739);
and U16155 (N_16155,N_13279,N_13113);
and U16156 (N_16156,N_11226,N_10101);
nor U16157 (N_16157,N_10994,N_10049);
and U16158 (N_16158,N_13059,N_11267);
xnor U16159 (N_16159,N_14135,N_11319);
or U16160 (N_16160,N_10236,N_12760);
nand U16161 (N_16161,N_14078,N_11147);
or U16162 (N_16162,N_13216,N_12176);
nor U16163 (N_16163,N_11295,N_14073);
nor U16164 (N_16164,N_12908,N_13823);
xnor U16165 (N_16165,N_11992,N_11936);
or U16166 (N_16166,N_13165,N_11882);
nand U16167 (N_16167,N_12398,N_10683);
xor U16168 (N_16168,N_11918,N_12122);
xnor U16169 (N_16169,N_11545,N_10704);
and U16170 (N_16170,N_14447,N_11715);
nor U16171 (N_16171,N_11436,N_14590);
nand U16172 (N_16172,N_12187,N_10378);
and U16173 (N_16173,N_13192,N_11034);
xnor U16174 (N_16174,N_13414,N_12336);
xor U16175 (N_16175,N_11938,N_10615);
nand U16176 (N_16176,N_12790,N_14312);
or U16177 (N_16177,N_13929,N_10739);
and U16178 (N_16178,N_12024,N_14402);
nor U16179 (N_16179,N_12375,N_10406);
and U16180 (N_16180,N_11559,N_13902);
nand U16181 (N_16181,N_13916,N_14720);
or U16182 (N_16182,N_13247,N_14425);
or U16183 (N_16183,N_11517,N_10916);
xnor U16184 (N_16184,N_10898,N_13992);
or U16185 (N_16185,N_13761,N_12895);
nor U16186 (N_16186,N_13315,N_14839);
xor U16187 (N_16187,N_14108,N_14613);
xnor U16188 (N_16188,N_10020,N_12061);
or U16189 (N_16189,N_13122,N_11749);
nor U16190 (N_16190,N_11904,N_11986);
xnor U16191 (N_16191,N_12228,N_12297);
nand U16192 (N_16192,N_10596,N_14343);
and U16193 (N_16193,N_13472,N_13462);
nor U16194 (N_16194,N_12424,N_11273);
nor U16195 (N_16195,N_10353,N_14865);
nand U16196 (N_16196,N_12433,N_12265);
nand U16197 (N_16197,N_11323,N_12608);
or U16198 (N_16198,N_10072,N_10471);
nand U16199 (N_16199,N_10561,N_13774);
nand U16200 (N_16200,N_11287,N_11243);
nand U16201 (N_16201,N_11956,N_12326);
or U16202 (N_16202,N_13058,N_14271);
xnor U16203 (N_16203,N_14441,N_14486);
nand U16204 (N_16204,N_14997,N_12113);
nand U16205 (N_16205,N_11976,N_13570);
nor U16206 (N_16206,N_14580,N_11401);
xor U16207 (N_16207,N_14697,N_10551);
xnor U16208 (N_16208,N_13133,N_10606);
or U16209 (N_16209,N_13259,N_10800);
xor U16210 (N_16210,N_11187,N_12280);
nor U16211 (N_16211,N_10037,N_11127);
nor U16212 (N_16212,N_11278,N_13041);
nand U16213 (N_16213,N_14808,N_10033);
nand U16214 (N_16214,N_12599,N_10489);
or U16215 (N_16215,N_14353,N_13179);
and U16216 (N_16216,N_13368,N_12665);
or U16217 (N_16217,N_12173,N_12004);
nor U16218 (N_16218,N_11475,N_11672);
or U16219 (N_16219,N_12517,N_12407);
nor U16220 (N_16220,N_13918,N_12542);
xor U16221 (N_16221,N_10423,N_13397);
xnor U16222 (N_16222,N_11535,N_13631);
or U16223 (N_16223,N_13102,N_10490);
or U16224 (N_16224,N_14145,N_10056);
nand U16225 (N_16225,N_11435,N_10139);
nand U16226 (N_16226,N_11072,N_12029);
or U16227 (N_16227,N_11121,N_10749);
and U16228 (N_16228,N_13659,N_12974);
nor U16229 (N_16229,N_11738,N_13688);
nand U16230 (N_16230,N_10871,N_13680);
or U16231 (N_16231,N_10052,N_10556);
nor U16232 (N_16232,N_12264,N_14795);
and U16233 (N_16233,N_12778,N_12901);
xnor U16234 (N_16234,N_13754,N_14646);
nand U16235 (N_16235,N_12485,N_14323);
xor U16236 (N_16236,N_12617,N_11599);
or U16237 (N_16237,N_10783,N_14143);
nor U16238 (N_16238,N_12931,N_10723);
xnor U16239 (N_16239,N_12075,N_11468);
nor U16240 (N_16240,N_10022,N_10102);
or U16241 (N_16241,N_12574,N_14888);
xor U16242 (N_16242,N_12875,N_14864);
and U16243 (N_16243,N_12936,N_11113);
or U16244 (N_16244,N_13919,N_11385);
nor U16245 (N_16245,N_14408,N_12193);
nand U16246 (N_16246,N_11282,N_11591);
or U16247 (N_16247,N_14771,N_14332);
or U16248 (N_16248,N_14170,N_14824);
nand U16249 (N_16249,N_11581,N_12095);
xnor U16250 (N_16250,N_11383,N_10528);
nand U16251 (N_16251,N_14093,N_14148);
nand U16252 (N_16252,N_11885,N_10726);
or U16253 (N_16253,N_12483,N_13481);
xnor U16254 (N_16254,N_11699,N_11652);
and U16255 (N_16255,N_11916,N_13968);
xnor U16256 (N_16256,N_13755,N_13639);
or U16257 (N_16257,N_11446,N_13484);
nor U16258 (N_16258,N_14711,N_12194);
nor U16259 (N_16259,N_11476,N_10003);
nand U16260 (N_16260,N_11692,N_13611);
or U16261 (N_16261,N_10027,N_11523);
or U16262 (N_16262,N_14765,N_13797);
nand U16263 (N_16263,N_13917,N_13502);
or U16264 (N_16264,N_11806,N_12874);
and U16265 (N_16265,N_10570,N_13091);
nor U16266 (N_16266,N_12691,N_10142);
nand U16267 (N_16267,N_14121,N_12268);
nand U16268 (N_16268,N_13140,N_10760);
nand U16269 (N_16269,N_12218,N_11047);
or U16270 (N_16270,N_10300,N_12679);
nand U16271 (N_16271,N_12008,N_10474);
or U16272 (N_16272,N_14495,N_14193);
nor U16273 (N_16273,N_10787,N_14937);
and U16274 (N_16274,N_10650,N_11859);
nand U16275 (N_16275,N_11336,N_13161);
and U16276 (N_16276,N_14134,N_12710);
nand U16277 (N_16277,N_12266,N_11639);
nor U16278 (N_16278,N_11056,N_10965);
nand U16279 (N_16279,N_10176,N_11053);
or U16280 (N_16280,N_13186,N_13815);
and U16281 (N_16281,N_10065,N_14665);
and U16282 (N_16282,N_10141,N_11590);
nand U16283 (N_16283,N_12112,N_14710);
or U16284 (N_16284,N_10303,N_13115);
or U16285 (N_16285,N_14232,N_13742);
nor U16286 (N_16286,N_13987,N_11042);
xnor U16287 (N_16287,N_11103,N_13003);
and U16288 (N_16288,N_12220,N_12151);
nor U16289 (N_16289,N_13963,N_13575);
nand U16290 (N_16290,N_11190,N_11663);
or U16291 (N_16291,N_13343,N_14275);
xnor U16292 (N_16292,N_10284,N_10845);
nand U16293 (N_16293,N_14077,N_13156);
and U16294 (N_16294,N_14056,N_11819);
and U16295 (N_16295,N_13808,N_12962);
or U16296 (N_16296,N_12222,N_13960);
xnor U16297 (N_16297,N_11390,N_13200);
nand U16298 (N_16298,N_14414,N_11146);
nor U16299 (N_16299,N_11315,N_11969);
nand U16300 (N_16300,N_10197,N_14520);
or U16301 (N_16301,N_10584,N_13951);
and U16302 (N_16302,N_13544,N_11609);
xor U16303 (N_16303,N_11304,N_12629);
nor U16304 (N_16304,N_14533,N_10791);
or U16305 (N_16305,N_12403,N_11095);
or U16306 (N_16306,N_12579,N_13901);
and U16307 (N_16307,N_12256,N_12208);
nor U16308 (N_16308,N_14209,N_14413);
nand U16309 (N_16309,N_12813,N_10798);
or U16310 (N_16310,N_10182,N_14404);
nor U16311 (N_16311,N_14448,N_14287);
or U16312 (N_16312,N_11795,N_11867);
nand U16313 (N_16313,N_12721,N_10879);
xor U16314 (N_16314,N_12786,N_12141);
nor U16315 (N_16315,N_14769,N_11872);
nand U16316 (N_16316,N_12662,N_13128);
xnor U16317 (N_16317,N_12968,N_14033);
and U16318 (N_16318,N_10545,N_11388);
nor U16319 (N_16319,N_10633,N_11844);
nand U16320 (N_16320,N_12260,N_12040);
or U16321 (N_16321,N_11097,N_12128);
nand U16322 (N_16322,N_12216,N_12487);
nand U16323 (N_16323,N_11735,N_12463);
xor U16324 (N_16324,N_14836,N_14356);
nand U16325 (N_16325,N_14817,N_12568);
xor U16326 (N_16326,N_11807,N_11245);
xnor U16327 (N_16327,N_14785,N_13190);
or U16328 (N_16328,N_11637,N_13990);
nand U16329 (N_16329,N_10291,N_14367);
nor U16330 (N_16330,N_10183,N_12490);
nor U16331 (N_16331,N_13494,N_14128);
nor U16332 (N_16332,N_10229,N_12289);
nor U16333 (N_16333,N_10361,N_12529);
and U16334 (N_16334,N_13130,N_12374);
nor U16335 (N_16335,N_13986,N_12658);
nor U16336 (N_16336,N_11833,N_14877);
or U16337 (N_16337,N_11413,N_10771);
nor U16338 (N_16338,N_10004,N_12070);
or U16339 (N_16339,N_10035,N_14781);
and U16340 (N_16340,N_13926,N_12349);
nand U16341 (N_16341,N_12819,N_13807);
xnor U16342 (N_16342,N_11557,N_11378);
and U16343 (N_16343,N_14342,N_11453);
and U16344 (N_16344,N_10859,N_11203);
nor U16345 (N_16345,N_13743,N_12355);
and U16346 (N_16346,N_14104,N_10166);
nand U16347 (N_16347,N_10968,N_14955);
nand U16348 (N_16348,N_11993,N_14625);
or U16349 (N_16349,N_10980,N_10002);
and U16350 (N_16350,N_12497,N_10008);
or U16351 (N_16351,N_11191,N_14682);
xnor U16352 (N_16352,N_13469,N_14885);
nand U16353 (N_16353,N_10029,N_11348);
nor U16354 (N_16354,N_10097,N_10940);
and U16355 (N_16355,N_13642,N_10955);
nor U16356 (N_16356,N_10511,N_14859);
or U16357 (N_16357,N_11492,N_12664);
and U16358 (N_16358,N_13325,N_10138);
nor U16359 (N_16359,N_12124,N_13491);
or U16360 (N_16360,N_11707,N_11285);
nor U16361 (N_16361,N_14724,N_10389);
xor U16362 (N_16362,N_12811,N_10186);
or U16363 (N_16363,N_10724,N_14443);
nor U16364 (N_16364,N_12896,N_10811);
nor U16365 (N_16365,N_10519,N_11828);
and U16366 (N_16366,N_10608,N_13535);
and U16367 (N_16367,N_10297,N_10381);
nor U16368 (N_16368,N_11084,N_10337);
nor U16369 (N_16369,N_14173,N_13694);
and U16370 (N_16370,N_11670,N_10559);
nand U16371 (N_16371,N_12793,N_11439);
nand U16372 (N_16372,N_13064,N_12310);
and U16373 (N_16373,N_10981,N_14983);
xor U16374 (N_16374,N_14610,N_14633);
xnor U16375 (N_16375,N_11106,N_12306);
xor U16376 (N_16376,N_10126,N_11371);
xnor U16377 (N_16377,N_12987,N_12753);
nor U16378 (N_16378,N_12399,N_12147);
nand U16379 (N_16379,N_13715,N_13248);
nor U16380 (N_16380,N_11033,N_11679);
or U16381 (N_16381,N_11974,N_11399);
nor U16382 (N_16382,N_11851,N_14308);
or U16383 (N_16383,N_12032,N_11373);
nor U16384 (N_16384,N_13388,N_14063);
nand U16385 (N_16385,N_14648,N_13447);
nand U16386 (N_16386,N_10607,N_14609);
nor U16387 (N_16387,N_12999,N_13106);
and U16388 (N_16388,N_14669,N_14489);
and U16389 (N_16389,N_11861,N_14907);
nor U16390 (N_16390,N_11415,N_14339);
nand U16391 (N_16391,N_10873,N_12586);
nand U16392 (N_16392,N_10128,N_10862);
nor U16393 (N_16393,N_14870,N_12565);
nand U16394 (N_16394,N_13054,N_10796);
and U16395 (N_16395,N_11023,N_11040);
nor U16396 (N_16396,N_12243,N_14949);
nand U16397 (N_16397,N_12248,N_14957);
nor U16398 (N_16398,N_13920,N_13999);
and U16399 (N_16399,N_11136,N_14840);
or U16400 (N_16400,N_11437,N_13239);
xor U16401 (N_16401,N_13477,N_12695);
and U16402 (N_16402,N_12563,N_14740);
nor U16403 (N_16403,N_10998,N_11231);
and U16404 (N_16404,N_14931,N_13531);
xor U16405 (N_16405,N_10371,N_13163);
nand U16406 (N_16406,N_12779,N_12825);
xor U16407 (N_16407,N_12293,N_11814);
or U16408 (N_16408,N_13389,N_12175);
nor U16409 (N_16409,N_12925,N_11623);
nand U16410 (N_16410,N_14502,N_13252);
or U16411 (N_16411,N_10762,N_14363);
and U16412 (N_16412,N_10557,N_10702);
nor U16413 (N_16413,N_14924,N_14221);
nand U16414 (N_16414,N_11351,N_11234);
nor U16415 (N_16415,N_10765,N_14246);
nor U16416 (N_16416,N_13870,N_10026);
nand U16417 (N_16417,N_12605,N_13337);
nor U16418 (N_16418,N_10674,N_10892);
nor U16419 (N_16419,N_10179,N_14737);
and U16420 (N_16420,N_12284,N_12798);
or U16421 (N_16421,N_12684,N_11582);
nor U16422 (N_16422,N_11118,N_14168);
nand U16423 (N_16423,N_11613,N_13037);
nor U16424 (N_16424,N_12958,N_11597);
nand U16425 (N_16425,N_12455,N_14692);
and U16426 (N_16426,N_12319,N_10269);
nand U16427 (N_16427,N_11197,N_11810);
or U16428 (N_16428,N_12909,N_14479);
and U16429 (N_16429,N_12404,N_12253);
nand U16430 (N_16430,N_13605,N_14691);
nor U16431 (N_16431,N_10993,N_14775);
nor U16432 (N_16432,N_14381,N_11573);
nand U16433 (N_16433,N_14752,N_14506);
and U16434 (N_16434,N_11754,N_11748);
nor U16435 (N_16435,N_13630,N_12551);
nand U16436 (N_16436,N_13060,N_13197);
nand U16437 (N_16437,N_10973,N_10467);
xnor U16438 (N_16438,N_11286,N_11424);
nand U16439 (N_16439,N_10132,N_13832);
or U16440 (N_16440,N_12716,N_11629);
or U16441 (N_16441,N_12437,N_13526);
or U16442 (N_16442,N_11179,N_13588);
nand U16443 (N_16443,N_12381,N_10273);
or U16444 (N_16444,N_12415,N_12835);
nor U16445 (N_16445,N_13110,N_13556);
nor U16446 (N_16446,N_12209,N_13222);
nor U16447 (N_16447,N_13393,N_11045);
nor U16448 (N_16448,N_12644,N_12476);
nor U16449 (N_16449,N_10645,N_13121);
xnor U16450 (N_16450,N_10382,N_12244);
nor U16451 (N_16451,N_10344,N_12486);
nor U16452 (N_16452,N_13619,N_11225);
nand U16453 (N_16453,N_13873,N_13692);
xor U16454 (N_16454,N_13118,N_14011);
and U16455 (N_16455,N_14837,N_12562);
nand U16456 (N_16456,N_11426,N_13146);
nor U16457 (N_16457,N_12638,N_11321);
and U16458 (N_16458,N_11512,N_12021);
xnor U16459 (N_16459,N_14722,N_10044);
and U16460 (N_16460,N_10162,N_13183);
nor U16461 (N_16461,N_11711,N_12555);
or U16462 (N_16462,N_11939,N_14797);
and U16463 (N_16463,N_13672,N_14600);
or U16464 (N_16464,N_12560,N_11028);
nor U16465 (N_16465,N_10335,N_14129);
xnor U16466 (N_16466,N_11781,N_13323);
xor U16467 (N_16467,N_11168,N_14690);
or U16468 (N_16468,N_11173,N_13610);
and U16469 (N_16469,N_13921,N_14666);
nand U16470 (N_16470,N_14759,N_12841);
or U16471 (N_16471,N_12467,N_10698);
nor U16472 (N_16472,N_10662,N_12099);
nor U16473 (N_16473,N_12973,N_13567);
nor U16474 (N_16474,N_11019,N_11349);
nor U16475 (N_16475,N_10540,N_10670);
xnor U16476 (N_16476,N_10953,N_14049);
or U16477 (N_16477,N_10685,N_14051);
nor U16478 (N_16478,N_14436,N_11568);
or U16479 (N_16479,N_13652,N_13995);
or U16480 (N_16480,N_11932,N_11332);
or U16481 (N_16481,N_11051,N_13152);
or U16482 (N_16482,N_14146,N_10092);
nand U16483 (N_16483,N_11200,N_13514);
and U16484 (N_16484,N_13155,N_10215);
and U16485 (N_16485,N_12465,N_10535);
nand U16486 (N_16486,N_12654,N_13168);
or U16487 (N_16487,N_14463,N_10019);
nand U16488 (N_16488,N_10851,N_11407);
nor U16489 (N_16489,N_12839,N_14507);
and U16490 (N_16490,N_14358,N_11732);
nor U16491 (N_16491,N_13522,N_13607);
nor U16492 (N_16492,N_14080,N_13810);
and U16493 (N_16493,N_11965,N_10255);
xor U16494 (N_16494,N_12600,N_12635);
nand U16495 (N_16495,N_11117,N_10365);
nand U16496 (N_16496,N_14948,N_10159);
or U16497 (N_16497,N_11087,N_11616);
nor U16498 (N_16498,N_10061,N_12524);
and U16499 (N_16499,N_13262,N_11035);
or U16500 (N_16500,N_13112,N_10251);
and U16501 (N_16501,N_13316,N_12412);
and U16502 (N_16502,N_11201,N_13932);
or U16503 (N_16503,N_11926,N_10673);
and U16504 (N_16504,N_12201,N_11603);
nand U16505 (N_16505,N_14066,N_14400);
xnor U16506 (N_16506,N_10790,N_12828);
or U16507 (N_16507,N_12791,N_11674);
or U16508 (N_16508,N_12339,N_14475);
nand U16509 (N_16509,N_10951,N_13487);
xor U16510 (N_16510,N_14597,N_10742);
and U16511 (N_16511,N_13237,N_11291);
or U16512 (N_16512,N_11773,N_14139);
nand U16513 (N_16513,N_14748,N_13930);
and U16514 (N_16514,N_11281,N_13400);
nor U16515 (N_16515,N_14678,N_10701);
xor U16516 (N_16516,N_12234,N_14391);
and U16517 (N_16517,N_14161,N_13407);
nand U16518 (N_16518,N_13801,N_13626);
or U16519 (N_16519,N_10869,N_10364);
nor U16520 (N_16520,N_14397,N_10882);
or U16521 (N_16521,N_10305,N_13885);
and U16522 (N_16522,N_13858,N_14842);
or U16523 (N_16523,N_13879,N_13518);
or U16524 (N_16524,N_14178,N_11254);
or U16525 (N_16525,N_13501,N_10974);
or U16526 (N_16526,N_12238,N_14231);
and U16527 (N_16527,N_13497,N_10681);
nor U16528 (N_16528,N_12149,N_12800);
nand U16529 (N_16529,N_12535,N_13109);
xor U16530 (N_16530,N_10367,N_14120);
xnor U16531 (N_16531,N_10324,N_10730);
or U16532 (N_16532,N_13461,N_10828);
or U16533 (N_16533,N_12996,N_10736);
or U16534 (N_16534,N_13722,N_11864);
nand U16535 (N_16535,N_13342,N_13566);
or U16536 (N_16536,N_10347,N_11089);
nand U16537 (N_16537,N_13094,N_12400);
or U16538 (N_16538,N_14018,N_11574);
or U16539 (N_16539,N_10066,N_11846);
nor U16540 (N_16540,N_12312,N_11447);
and U16541 (N_16541,N_12422,N_13177);
or U16542 (N_16542,N_12945,N_12977);
and U16543 (N_16543,N_12039,N_12772);
nor U16544 (N_16544,N_10124,N_14585);
or U16545 (N_16545,N_10989,N_10775);
or U16546 (N_16546,N_11063,N_13907);
nand U16547 (N_16547,N_10777,N_10926);
or U16548 (N_16548,N_14901,N_14693);
nand U16549 (N_16549,N_13172,N_12232);
and U16550 (N_16550,N_12821,N_12815);
nand U16551 (N_16551,N_11157,N_12689);
or U16552 (N_16552,N_14593,N_14647);
xor U16553 (N_16553,N_14352,N_12570);
xnor U16554 (N_16554,N_12156,N_11284);
xnor U16555 (N_16555,N_12000,N_12182);
xor U16556 (N_16556,N_11142,N_12246);
nand U16557 (N_16557,N_14969,N_11495);
xnor U16558 (N_16558,N_10939,N_11408);
or U16559 (N_16559,N_12352,N_14790);
nand U16560 (N_16560,N_11277,N_11669);
nor U16561 (N_16561,N_11111,N_14627);
nor U16562 (N_16562,N_10418,N_13392);
or U16563 (N_16563,N_11880,N_10356);
or U16564 (N_16564,N_12887,N_10266);
and U16565 (N_16565,N_12211,N_13983);
or U16566 (N_16566,N_10296,N_14852);
xnor U16567 (N_16567,N_10552,N_12386);
and U16568 (N_16568,N_13280,N_11845);
nor U16569 (N_16569,N_11237,N_12508);
and U16570 (N_16570,N_14118,N_10924);
xnor U16571 (N_16571,N_11081,N_14017);
xor U16572 (N_16572,N_13108,N_11958);
nor U16573 (N_16573,N_12589,N_12598);
or U16574 (N_16574,N_10225,N_13579);
xnor U16575 (N_16575,N_14799,N_11520);
nor U16576 (N_16576,N_14291,N_11910);
xor U16577 (N_16577,N_10431,N_14528);
xnor U16578 (N_16578,N_12505,N_12863);
and U16579 (N_16579,N_13913,N_14130);
xnor U16580 (N_16580,N_13510,N_11995);
nand U16581 (N_16581,N_11233,N_13412);
and U16582 (N_16582,N_11817,N_10156);
and U16583 (N_16583,N_10085,N_12074);
nor U16584 (N_16584,N_13967,N_12610);
and U16585 (N_16585,N_14319,N_12273);
and U16586 (N_16586,N_14505,N_11473);
nor U16587 (N_16587,N_12985,N_10118);
nor U16588 (N_16588,N_13621,N_13062);
or U16589 (N_16589,N_13346,N_10546);
xnor U16590 (N_16590,N_12245,N_10720);
nor U16591 (N_16591,N_12049,N_12145);
or U16592 (N_16592,N_10232,N_10763);
or U16593 (N_16593,N_13295,N_13554);
or U16594 (N_16594,N_11239,N_13865);
xnor U16595 (N_16595,N_14053,N_13448);
and U16596 (N_16596,N_12518,N_10211);
and U16597 (N_16597,N_11546,N_13286);
xnor U16598 (N_16598,N_14476,N_13281);
nand U16599 (N_16599,N_12799,N_12044);
xnor U16600 (N_16600,N_10959,N_13004);
and U16601 (N_16601,N_11868,N_10093);
and U16602 (N_16602,N_13516,N_12515);
xor U16603 (N_16603,N_10885,N_13189);
and U16604 (N_16604,N_13606,N_14860);
and U16605 (N_16605,N_12876,N_14606);
nor U16606 (N_16606,N_13727,N_10478);
or U16607 (N_16607,N_11648,N_13915);
and U16608 (N_16608,N_11400,N_12168);
xor U16609 (N_16609,N_10643,N_11975);
nand U16610 (N_16610,N_10641,N_11008);
xor U16611 (N_16611,N_11470,N_10034);
nand U16612 (N_16612,N_11750,N_12131);
xor U16613 (N_16613,N_13857,N_11841);
xor U16614 (N_16614,N_12396,N_14100);
or U16615 (N_16615,N_11688,N_14235);
and U16616 (N_16616,N_13306,N_12681);
xnor U16617 (N_16617,N_10605,N_12550);
or U16618 (N_16618,N_12889,N_11887);
or U16619 (N_16619,N_10792,N_13653);
nand U16620 (N_16620,N_13079,N_14675);
and U16621 (N_16621,N_11997,N_14537);
xnor U16622 (N_16622,N_11479,N_13367);
nand U16623 (N_16623,N_11662,N_10333);
xor U16624 (N_16624,N_12872,N_12780);
or U16625 (N_16625,N_13267,N_12152);
nor U16626 (N_16626,N_12782,N_10950);
or U16627 (N_16627,N_10104,N_12302);
and U16628 (N_16628,N_13242,N_11354);
nand U16629 (N_16629,N_14928,N_11037);
xnor U16630 (N_16630,N_10526,N_10193);
nor U16631 (N_16631,N_11314,N_10948);
and U16632 (N_16632,N_13758,N_12279);
nor U16633 (N_16633,N_10199,N_13520);
and U16634 (N_16634,N_10100,N_14243);
nand U16635 (N_16635,N_10579,N_11054);
xor U16636 (N_16636,N_14632,N_10983);
or U16637 (N_16637,N_14815,N_11220);
xor U16638 (N_16638,N_14230,N_13439);
xnor U16639 (N_16639,N_14712,N_13083);
or U16640 (N_16640,N_14923,N_13153);
nor U16641 (N_16641,N_13395,N_13660);
nor U16642 (N_16642,N_12006,N_10727);
xor U16643 (N_16643,N_10522,N_11505);
xnor U16644 (N_16644,N_13098,N_10146);
nor U16645 (N_16645,N_13022,N_14784);
nand U16646 (N_16646,N_10068,N_10855);
and U16647 (N_16647,N_12934,N_14390);
xnor U16648 (N_16648,N_13671,N_10064);
or U16649 (N_16649,N_12038,N_13254);
nand U16650 (N_16650,N_13096,N_12441);
or U16651 (N_16651,N_13227,N_11001);
xnor U16652 (N_16652,N_13480,N_11772);
or U16653 (N_16653,N_10609,N_12668);
nor U16654 (N_16654,N_13356,N_14205);
xor U16655 (N_16655,N_14300,N_12018);
or U16656 (N_16656,N_11317,N_10334);
and U16657 (N_16657,N_14733,N_12948);
nor U16658 (N_16658,N_10402,N_11462);
or U16659 (N_16659,N_12356,N_12202);
or U16660 (N_16660,N_14728,N_14534);
or U16661 (N_16661,N_13304,N_12645);
nand U16662 (N_16662,N_10234,N_14635);
and U16663 (N_16663,N_10320,N_10272);
or U16664 (N_16664,N_13134,N_12569);
nor U16665 (N_16665,N_12747,N_13733);
and U16666 (N_16666,N_10624,N_14210);
nor U16667 (N_16667,N_10238,N_13289);
xor U16668 (N_16668,N_12769,N_14309);
nand U16669 (N_16669,N_14750,N_14890);
or U16670 (N_16670,N_13724,N_14024);
nor U16671 (N_16671,N_14211,N_14591);
and U16672 (N_16672,N_10517,N_10325);
and U16673 (N_16673,N_11944,N_12272);
or U16674 (N_16674,N_11991,N_11996);
or U16675 (N_16675,N_14764,N_10582);
and U16676 (N_16676,N_10872,N_13266);
or U16677 (N_16677,N_12959,N_13327);
nor U16678 (N_16678,N_10516,N_12620);
xnor U16679 (N_16679,N_10657,N_10922);
or U16680 (N_16680,N_12986,N_12267);
and U16681 (N_16681,N_14638,N_10821);
or U16682 (N_16682,N_12663,N_11519);
or U16683 (N_16683,N_10201,N_14307);
xor U16684 (N_16684,N_12379,N_14452);
xnor U16685 (N_16685,N_13390,N_12690);
nor U16686 (N_16686,N_10629,N_10359);
nor U16687 (N_16687,N_10492,N_11500);
xnor U16688 (N_16688,N_13151,N_14457);
nor U16689 (N_16689,N_11886,N_13455);
and U16690 (N_16690,N_14845,N_13608);
nand U16691 (N_16691,N_11973,N_14468);
nor U16692 (N_16692,N_12960,N_11322);
nand U16693 (N_16693,N_10218,N_12659);
xor U16694 (N_16694,N_12033,N_12002);
and U16695 (N_16695,N_14107,N_12546);
and U16696 (N_16696,N_12939,N_14069);
nor U16697 (N_16697,N_12704,N_14110);
nor U16698 (N_16698,N_10191,N_11856);
or U16699 (N_16699,N_14814,N_12093);
nor U16700 (N_16700,N_11396,N_13806);
xnor U16701 (N_16701,N_14789,N_10890);
and U16702 (N_16702,N_14510,N_14071);
or U16703 (N_16703,N_10453,N_13778);
and U16704 (N_16704,N_10192,N_11694);
nor U16705 (N_16705,N_11794,N_14612);
or U16706 (N_16706,N_12215,N_14659);
nor U16707 (N_16707,N_10886,N_12929);
nand U16708 (N_16708,N_14925,N_12331);
nand U16709 (N_16709,N_11368,N_13093);
and U16710 (N_16710,N_14516,N_12082);
xnor U16711 (N_16711,N_14341,N_12715);
or U16712 (N_16712,N_10690,N_10285);
nor U16713 (N_16713,N_10978,N_11518);
xor U16714 (N_16714,N_14003,N_12434);
nor U16715 (N_16715,N_11170,N_13399);
and U16716 (N_16716,N_13749,N_12972);
xor U16717 (N_16717,N_10328,N_13411);
and U16718 (N_16718,N_11589,N_10450);
nor U16719 (N_16719,N_14744,N_11782);
and U16720 (N_16720,N_11391,N_12301);
nor U16721 (N_16721,N_14735,N_13049);
or U16722 (N_16722,N_10912,N_11341);
nand U16723 (N_16723,N_12102,N_10616);
or U16724 (N_16724,N_12840,N_13791);
xnor U16725 (N_16725,N_13816,N_14348);
xor U16726 (N_16726,N_13790,N_10564);
or U16727 (N_16727,N_11112,N_11547);
or U16728 (N_16728,N_11988,N_10206);
xor U16729 (N_16729,N_13085,N_10452);
nor U16730 (N_16730,N_14298,N_11906);
xnor U16731 (N_16731,N_12383,N_12646);
or U16732 (N_16732,N_12274,N_10856);
and U16733 (N_16733,N_12614,N_10010);
or U16734 (N_16734,N_11101,N_12393);
or U16735 (N_16735,N_12737,N_14458);
nand U16736 (N_16736,N_12001,N_14861);
nand U16737 (N_16737,N_11438,N_12761);
or U16738 (N_16738,N_13432,N_10577);
nor U16739 (N_16739,N_11338,N_14470);
or U16740 (N_16740,N_14456,N_12910);
and U16741 (N_16741,N_14726,N_10053);
and U16742 (N_16742,N_13169,N_10042);
or U16743 (N_16743,N_11638,N_14415);
and U16744 (N_16744,N_14123,N_11624);
nor U16745 (N_16745,N_14975,N_10864);
nor U16746 (N_16746,N_13175,N_11003);
xor U16747 (N_16747,N_14757,N_14215);
and U16748 (N_16748,N_11709,N_12783);
nor U16749 (N_16749,N_14437,N_14081);
xnor U16750 (N_16750,N_10307,N_10549);
nor U16751 (N_16751,N_13702,N_12370);
or U16752 (N_16752,N_12344,N_14299);
and U16753 (N_16753,N_10187,N_11150);
or U16754 (N_16754,N_11129,N_13953);
xor U16755 (N_16755,N_12100,N_13826);
nand U16756 (N_16756,N_14631,N_14169);
nand U16757 (N_16757,N_11380,N_14428);
nor U16758 (N_16758,N_10507,N_12892);
nor U16759 (N_16759,N_10427,N_13641);
nor U16760 (N_16760,N_12548,N_13065);
and U16761 (N_16761,N_13321,N_12154);
and U16762 (N_16762,N_12134,N_12842);
and U16763 (N_16763,N_11309,N_11620);
or U16764 (N_16764,N_13595,N_13008);
nor U16765 (N_16765,N_11902,N_14910);
nand U16766 (N_16766,N_10306,N_11497);
nand U16767 (N_16767,N_14658,N_11216);
and U16768 (N_16768,N_14952,N_14035);
nor U16769 (N_16769,N_13899,N_11176);
xnor U16770 (N_16770,N_12998,N_14851);
nand U16771 (N_16771,N_13941,N_14421);
xor U16772 (N_16772,N_13903,N_12327);
nand U16773 (N_16773,N_12110,N_14763);
xnor U16774 (N_16774,N_14943,N_10977);
nand U16775 (N_16775,N_12607,N_10569);
and U16776 (N_16776,N_11664,N_14096);
xnor U16777 (N_16777,N_14677,N_11228);
and U16778 (N_16778,N_10422,N_13966);
and U16779 (N_16779,N_12857,N_13413);
nor U16780 (N_16780,N_12350,N_13952);
and U16781 (N_16781,N_10710,N_12736);
and U16782 (N_16782,N_11530,N_11642);
nand U16783 (N_16783,N_10512,N_13391);
or U16784 (N_16784,N_12034,N_13851);
xnor U16785 (N_16785,N_13696,N_14225);
nor U16786 (N_16786,N_13474,N_13318);
nor U16787 (N_16787,N_11207,N_13721);
and U16788 (N_16788,N_10741,N_10946);
nand U16789 (N_16789,N_11466,N_12573);
and U16790 (N_16790,N_12552,N_13131);
xor U16791 (N_16791,N_11563,N_10243);
and U16792 (N_16792,N_11745,N_12160);
xor U16793 (N_16793,N_14314,N_11333);
nor U16794 (N_16794,N_10505,N_11661);
nor U16795 (N_16795,N_13811,N_12733);
nor U16796 (N_16796,N_11526,N_11104);
or U16797 (N_16797,N_10135,N_12150);
nor U16798 (N_16798,N_12106,N_12947);
and U16799 (N_16799,N_11830,N_14099);
and U16800 (N_16800,N_13877,N_10095);
nand U16801 (N_16801,N_14084,N_14453);
or U16802 (N_16802,N_14175,N_10666);
and U16803 (N_16803,N_10713,N_12281);
nand U16804 (N_16804,N_13946,N_14384);
and U16805 (N_16805,N_11431,N_14052);
nor U16806 (N_16806,N_10803,N_14401);
xnor U16807 (N_16807,N_10177,N_12493);
and U16808 (N_16808,N_12797,N_12990);
xnor U16809 (N_16809,N_12325,N_13712);
xor U16810 (N_16810,N_10797,N_12263);
or U16811 (N_16811,N_12849,N_14191);
xnor U16812 (N_16812,N_10789,N_12171);
and U16813 (N_16813,N_14266,N_11683);
and U16814 (N_16814,N_10496,N_10610);
nand U16815 (N_16815,N_11096,N_13892);
nor U16816 (N_16816,N_10016,N_12342);
nand U16817 (N_16817,N_12714,N_12157);
or U16818 (N_16818,N_11369,N_12957);
xor U16819 (N_16819,N_12162,N_14701);
or U16820 (N_16820,N_14395,N_13251);
and U16821 (N_16821,N_14306,N_11420);
xor U16822 (N_16822,N_13423,N_10039);
xnor U16823 (N_16823,N_12575,N_13162);
nor U16824 (N_16824,N_12781,N_12085);
xnor U16825 (N_16825,N_10780,N_14749);
nand U16826 (N_16826,N_11744,N_12146);
or U16827 (N_16827,N_12348,N_12313);
nand U16828 (N_16828,N_13888,N_14681);
and U16829 (N_16829,N_11816,N_10050);
xnor U16830 (N_16830,N_13086,N_13364);
and U16831 (N_16831,N_11761,N_11132);
nor U16832 (N_16832,N_10096,N_10695);
and U16833 (N_16833,N_12427,N_12725);
xnor U16834 (N_16834,N_14560,N_12435);
and U16835 (N_16835,N_13452,N_12530);
nand U16836 (N_16836,N_11115,N_14900);
xor U16837 (N_16837,N_13779,N_10311);
and U16838 (N_16838,N_14979,N_13993);
and U16839 (N_16839,N_12912,N_10082);
nor U16840 (N_16840,N_12429,N_11324);
nand U16841 (N_16841,N_13679,N_10248);
or U16842 (N_16842,N_11673,N_13199);
or U16843 (N_16843,N_13024,N_11722);
and U16844 (N_16844,N_12916,N_13555);
or U16845 (N_16845,N_14987,N_12711);
xnor U16846 (N_16846,N_11250,N_13729);
xor U16847 (N_16847,N_11785,N_14977);
nor U16848 (N_16848,N_14950,N_13906);
and U16849 (N_16849,N_14109,N_13326);
xnor U16850 (N_16850,N_14926,N_13762);
xnor U16851 (N_16851,N_14543,N_12627);
and U16852 (N_16852,N_13257,N_13468);
or U16853 (N_16853,N_13711,N_11705);
and U16854 (N_16854,N_11908,N_14912);
or U16855 (N_16855,N_11130,N_13475);
nor U16856 (N_16856,N_11565,N_13224);
and U16857 (N_16857,N_10597,N_11695);
xor U16858 (N_16858,N_10448,N_13548);
nor U16859 (N_16859,N_13067,N_12089);
xnor U16860 (N_16860,N_13511,N_10925);
xor U16861 (N_16861,N_14960,N_14660);
nand U16862 (N_16862,N_14228,N_11144);
nor U16863 (N_16863,N_13207,N_13180);
nand U16864 (N_16864,N_10253,N_13728);
or U16865 (N_16865,N_11653,N_12531);
xnor U16866 (N_16866,N_10109,N_10249);
nor U16867 (N_16867,N_13234,N_13854);
or U16868 (N_16868,N_11607,N_12915);
nand U16869 (N_16869,N_11272,N_10247);
xor U16870 (N_16870,N_13069,N_11730);
nor U16871 (N_16871,N_13819,N_11560);
xor U16872 (N_16872,N_11257,N_13881);
nand U16873 (N_16873,N_14226,N_14176);
and U16874 (N_16874,N_12956,N_10323);
or U16875 (N_16875,N_14137,N_13500);
xor U16876 (N_16876,N_13895,N_12142);
xor U16877 (N_16877,N_14655,N_10264);
nor U16878 (N_16878,N_11303,N_14558);
nor U16879 (N_16879,N_12612,N_14440);
nand U16880 (N_16880,N_14227,N_10134);
nand U16881 (N_16881,N_10806,N_11792);
nand U16882 (N_16882,N_11211,N_13335);
and U16883 (N_16883,N_11344,N_13089);
nand U16884 (N_16884,N_14481,N_12509);
xor U16885 (N_16885,N_10411,N_13651);
and U16886 (N_16886,N_14559,N_14592);
or U16887 (N_16887,N_11818,N_11365);
nand U16888 (N_16888,N_10899,N_14542);
and U16889 (N_16889,N_14573,N_14844);
nor U16890 (N_16890,N_12686,N_10630);
xor U16891 (N_16891,N_11406,N_13849);
nand U16892 (N_16892,N_13427,N_10644);
or U16893 (N_16893,N_10336,N_10880);
xnor U16894 (N_16894,N_11703,N_14626);
nor U16895 (N_16895,N_13371,N_12366);
xor U16896 (N_16896,N_13075,N_12661);
nand U16897 (N_16897,N_13894,N_10213);
xor U16898 (N_16898,N_13880,N_13422);
nor U16899 (N_16899,N_14365,N_10315);
and U16900 (N_16900,N_12763,N_10640);
or U16901 (N_16901,N_13415,N_10395);
xor U16902 (N_16902,N_10443,N_12900);
nand U16903 (N_16903,N_10761,N_10944);
nand U16904 (N_16904,N_11296,N_14032);
and U16905 (N_16905,N_12971,N_12363);
and U16906 (N_16906,N_11510,N_11646);
nand U16907 (N_16907,N_13241,N_11796);
xor U16908 (N_16908,N_11387,N_14916);
nand U16909 (N_16909,N_14388,N_12257);
and U16910 (N_16910,N_13513,N_14872);
and U16911 (N_16911,N_11903,N_14186);
nand U16912 (N_16912,N_10807,N_14490);
nor U16913 (N_16913,N_10743,N_11681);
xor U16914 (N_16914,N_13404,N_13776);
nor U16915 (N_16915,N_13871,N_10622);
xnor U16916 (N_16916,N_13141,N_11913);
xnor U16917 (N_16917,N_10956,N_10493);
nor U16918 (N_16918,N_12701,N_10544);
nor U16919 (N_16919,N_14091,N_13859);
nor U16920 (N_16920,N_13139,N_13665);
or U16921 (N_16921,N_14783,N_11022);
or U16922 (N_16922,N_10830,N_13283);
nor U16923 (N_16923,N_12494,N_12076);
or U16924 (N_16924,N_14265,N_11914);
xor U16925 (N_16925,N_11210,N_13695);
nand U16926 (N_16926,N_13426,N_14995);
nor U16927 (N_16927,N_11425,N_14289);
or U16928 (N_16928,N_12213,N_14867);
or U16929 (N_16929,N_14779,N_10625);
xnor U16930 (N_16930,N_12894,N_10827);
or U16931 (N_16931,N_12983,N_10975);
xor U16932 (N_16932,N_13707,N_14680);
xnor U16933 (N_16933,N_12384,N_12013);
or U16934 (N_16934,N_12834,N_11836);
or U16935 (N_16935,N_10560,N_12123);
and U16936 (N_16936,N_13011,N_14670);
nand U16937 (N_16937,N_11064,N_12755);
nor U16938 (N_16938,N_11687,N_10962);
and U16939 (N_16939,N_10614,N_11702);
nor U16940 (N_16940,N_13374,N_14930);
nor U16941 (N_16941,N_10747,N_14002);
nand U16942 (N_16942,N_11507,N_12966);
xor U16943 (N_16943,N_14105,N_10252);
nand U16944 (N_16944,N_12587,N_14550);
nand U16945 (N_16945,N_10429,N_13014);
or U16946 (N_16946,N_11131,N_10245);
and U16947 (N_16947,N_13104,N_10915);
or U16948 (N_16948,N_11951,N_10079);
and U16949 (N_16949,N_14545,N_13017);
nor U16950 (N_16950,N_12445,N_12408);
xor U16951 (N_16951,N_12541,N_12653);
nor U16952 (N_16952,N_14978,N_10254);
nor U16953 (N_16953,N_10465,N_13485);
xnor U16954 (N_16954,N_10174,N_14251);
xor U16955 (N_16955,N_14370,N_10722);
xnor U16956 (N_16956,N_12820,N_13944);
nand U16957 (N_16957,N_14961,N_11410);
nand U16958 (N_16958,N_13478,N_12652);
and U16959 (N_16959,N_12596,N_11982);
or U16960 (N_16960,N_13852,N_11710);
nand U16961 (N_16961,N_11756,N_10434);
and U16962 (N_16962,N_12911,N_13820);
and U16963 (N_16963,N_14277,N_12513);
nand U16964 (N_16964,N_13708,N_11667);
and U16965 (N_16965,N_12928,N_14602);
and U16966 (N_16966,N_10671,N_14159);
nand U16967 (N_16967,N_12731,N_14536);
and U16968 (N_16968,N_11256,N_10312);
nor U16969 (N_16969,N_11774,N_11014);
nor U16970 (N_16970,N_14777,N_11217);
nor U16971 (N_16971,N_12637,N_11787);
nand U16972 (N_16972,N_11270,N_14661);
or U16973 (N_16973,N_11657,N_10327);
and U16974 (N_16974,N_11429,N_11044);
nor U16975 (N_16975,N_13935,N_13551);
nand U16976 (N_16976,N_13255,N_10160);
and U16977 (N_16977,N_14530,N_11998);
nand U16978 (N_16978,N_11605,N_11374);
nand U16979 (N_16979,N_11561,N_13540);
xnor U16980 (N_16980,N_12097,N_13401);
and U16981 (N_16981,N_14529,N_13431);
and U16982 (N_16982,N_10725,N_11536);
xnor U16983 (N_16983,N_14361,N_14668);
nand U16984 (N_16984,N_13245,N_12454);
nand U16985 (N_16985,N_13159,N_13453);
or U16986 (N_16986,N_12362,N_10194);
nor U16987 (N_16987,N_14651,N_10651);
xnor U16988 (N_16988,N_13620,N_11945);
nand U16989 (N_16989,N_13405,N_10351);
and U16990 (N_16990,N_13026,N_11464);
or U16991 (N_16991,N_11614,N_12854);
and U16992 (N_16992,N_10738,N_14046);
or U16993 (N_16993,N_11361,N_13799);
nand U16994 (N_16994,N_14863,N_12768);
and U16995 (N_16995,N_12853,N_14464);
xnor U16996 (N_16996,N_13078,N_12271);
or U16997 (N_16997,N_12314,N_11080);
nand U16998 (N_16998,N_10515,N_12982);
xnor U16999 (N_16999,N_11078,N_14615);
nand U17000 (N_17000,N_10091,N_11178);
nor U17001 (N_17001,N_14407,N_11862);
xor U17002 (N_17002,N_14514,N_13344);
xor U17003 (N_17003,N_12385,N_11265);
or U17004 (N_17004,N_11375,N_10801);
xnor U17005 (N_17005,N_11290,N_10425);
or U17006 (N_17006,N_14039,N_10520);
nand U17007 (N_17007,N_13101,N_12903);
xnor U17008 (N_17008,N_13132,N_12438);
and U17009 (N_17009,N_13428,N_12511);
and U17010 (N_17010,N_12188,N_13740);
xor U17011 (N_17011,N_11566,N_14072);
or U17012 (N_17012,N_10298,N_12431);
and U17013 (N_17013,N_14664,N_14605);
or U17014 (N_17014,N_13045,N_14921);
xor U17015 (N_17015,N_13434,N_10077);
nand U17016 (N_17016,N_10835,N_12369);
nand U17017 (N_17017,N_13613,N_12619);
and U17018 (N_17018,N_14364,N_12081);
nor U17019 (N_17019,N_13598,N_12030);
and U17020 (N_17020,N_12353,N_12749);
and U17021 (N_17021,N_13355,N_13111);
nand U17022 (N_17022,N_10612,N_13927);
nor U17023 (N_17023,N_11030,N_12879);
and U17024 (N_17024,N_14331,N_12135);
and U17025 (N_17025,N_13217,N_10398);
xnor U17026 (N_17026,N_14165,N_12969);
nor U17027 (N_17027,N_11487,N_13550);
nand U17028 (N_17028,N_12576,N_12453);
nand U17029 (N_17029,N_12227,N_13869);
or U17030 (N_17030,N_11562,N_12143);
nand U17031 (N_17031,N_12186,N_12897);
and U17032 (N_17032,N_10846,N_12640);
nand U17033 (N_17033,N_14518,N_12618);
or U17034 (N_17034,N_11417,N_12980);
or U17035 (N_17035,N_11941,N_13470);
or U17036 (N_17036,N_12170,N_11898);
nand U17037 (N_17037,N_13615,N_12332);
nor U17038 (N_17038,N_10599,N_13780);
xor U17039 (N_17039,N_14751,N_10214);
and U17040 (N_17040,N_10788,N_11181);
nor U17041 (N_17041,N_13253,N_14676);
xnor U17042 (N_17042,N_14574,N_14942);
and U17043 (N_17043,N_12241,N_13767);
or U17044 (N_17044,N_14959,N_10233);
nor U17045 (N_17045,N_10259,N_10911);
or U17046 (N_17046,N_10329,N_12745);
or U17047 (N_17047,N_12020,N_14548);
or U17048 (N_17048,N_13009,N_14608);
xnor U17049 (N_17049,N_12864,N_13537);
nand U17050 (N_17050,N_13504,N_14293);
xnor U17051 (N_17051,N_10113,N_12978);
and U17052 (N_17052,N_10504,N_10447);
and U17053 (N_17053,N_13824,N_13942);
nor U17054 (N_17054,N_13529,N_12064);
nor U17055 (N_17055,N_11689,N_10387);
and U17056 (N_17056,N_10208,N_13803);
xor U17057 (N_17057,N_10875,N_14321);
and U17058 (N_17058,N_13221,N_13206);
nor U17059 (N_17059,N_13977,N_14351);
xnor U17060 (N_17060,N_10530,N_12071);
or U17061 (N_17061,N_13046,N_13539);
or U17062 (N_17062,N_14014,N_13250);
nand U17063 (N_17063,N_13403,N_13874);
nand U17064 (N_17064,N_10195,N_13347);
nor U17065 (N_17065,N_11214,N_11871);
and U17066 (N_17066,N_12117,N_10005);
or U17067 (N_17067,N_13643,N_10627);
and U17068 (N_17068,N_13028,N_10339);
and U17069 (N_17069,N_14272,N_11678);
xnor U17070 (N_17070,N_13600,N_12572);
nand U17071 (N_17071,N_10967,N_12050);
xor U17072 (N_17072,N_10007,N_13834);
xnor U17073 (N_17073,N_10581,N_12926);
xnor U17074 (N_17074,N_10941,N_11463);
nand U17075 (N_17075,N_14329,N_12634);
nor U17076 (N_17076,N_14041,N_12871);
xor U17077 (N_17077,N_12669,N_12019);
xnor U17078 (N_17078,N_13547,N_10281);
and U17079 (N_17079,N_11430,N_10611);
nand U17080 (N_17080,N_12436,N_13691);
and U17081 (N_17081,N_10626,N_12988);
or U17082 (N_17082,N_13444,N_11725);
or U17083 (N_17083,N_13202,N_12153);
or U17084 (N_17084,N_10224,N_10813);
and U17085 (N_17085,N_11878,N_12830);
nand U17086 (N_17086,N_11477,N_14150);
nor U17087 (N_17087,N_14462,N_10823);
xor U17088 (N_17088,N_10330,N_12692);
or U17089 (N_17089,N_10417,N_11770);
nor U17090 (N_17090,N_11422,N_14396);
xor U17091 (N_17091,N_14439,N_10686);
and U17092 (N_17092,N_14344,N_12943);
nor U17093 (N_17093,N_14622,N_14079);
nand U17094 (N_17094,N_11606,N_11248);
or U17095 (N_17095,N_13088,N_13230);
nand U17096 (N_17096,N_14981,N_13805);
nand U17097 (N_17097,N_14375,N_11596);
xnor U17098 (N_17098,N_11006,N_11491);
nor U17099 (N_17099,N_11720,N_11759);
and U17100 (N_17100,N_11531,N_13633);
and U17101 (N_17101,N_13512,N_12981);
or U17102 (N_17102,N_11300,N_13015);
or U17103 (N_17103,N_13770,N_10840);
nor U17104 (N_17104,N_10992,N_10555);
xor U17105 (N_17105,N_12881,N_11193);
nand U17106 (N_17106,N_14095,N_12196);
or U17107 (N_17107,N_13341,N_11503);
xnor U17108 (N_17108,N_14304,N_12831);
and U17109 (N_17109,N_10832,N_11269);
xnor U17110 (N_17110,N_11803,N_12104);
and U17111 (N_17111,N_13410,N_12023);
nor U17112 (N_17112,N_12726,N_14253);
nand U17113 (N_17113,N_10404,N_11238);
xnor U17114 (N_17114,N_14584,N_10433);
nand U17115 (N_17115,N_10964,N_11651);
nand U17116 (N_17116,N_14144,N_11553);
xor U17117 (N_17117,N_14021,N_11280);
or U17118 (N_17118,N_12174,N_13198);
or U17119 (N_17119,N_10786,N_11124);
and U17120 (N_17120,N_10751,N_11764);
or U17121 (N_17121,N_12540,N_11102);
xor U17122 (N_17122,N_10368,N_11024);
xor U17123 (N_17123,N_14484,N_13357);
and U17124 (N_17124,N_14704,N_12360);
or U17125 (N_17125,N_14834,N_10036);
or U17126 (N_17126,N_10818,N_13714);
xnor U17127 (N_17127,N_10831,N_13521);
xor U17128 (N_17128,N_11202,N_12199);
or U17129 (N_17129,N_11860,N_13933);
nand U17130 (N_17130,N_11026,N_11823);
and U17131 (N_17131,N_10196,N_12025);
and U17132 (N_17132,N_12553,N_13931);
or U17133 (N_17133,N_10435,N_10772);
xor U17134 (N_17134,N_11433,N_11777);
nor U17135 (N_17135,N_13232,N_14623);
xor U17136 (N_17136,N_14688,N_11610);
nand U17137 (N_17137,N_13313,N_14685);
nor U17138 (N_17138,N_14805,N_13265);
or U17139 (N_17139,N_11571,N_14346);
nand U17140 (N_17140,N_10660,N_11556);
nand U17141 (N_17141,N_10385,N_12994);
nor U17142 (N_17142,N_14029,N_10143);
nand U17143 (N_17143,N_13294,N_12777);
nand U17144 (N_17144,N_11049,N_10414);
nor U17145 (N_17145,N_11347,N_14729);
nand U17146 (N_17146,N_10563,N_14800);
and U17147 (N_17147,N_12677,N_10719);
and U17148 (N_17148,N_14450,N_10257);
nand U17149 (N_17149,N_11163,N_11729);
and U17150 (N_17150,N_11452,N_14689);
xor U17151 (N_17151,N_10372,N_11381);
nor U17152 (N_17152,N_14102,N_13021);
or U17153 (N_17153,N_14160,N_12561);
or U17154 (N_17154,N_10144,N_10573);
nand U17155 (N_17155,N_12585,N_12613);
or U17156 (N_17156,N_10602,N_11854);
nor U17157 (N_17157,N_10920,N_10168);
xnor U17158 (N_17158,N_11627,N_10575);
nand U17159 (N_17159,N_13238,N_14576);
xnor U17160 (N_17160,N_12426,N_10921);
or U17161 (N_17161,N_10087,N_12759);
nand U17162 (N_17162,N_14098,N_13416);
nor U17163 (N_17163,N_12210,N_10902);
and U17164 (N_17164,N_12169,N_11719);
xor U17165 (N_17165,N_10970,N_10566);
or U17166 (N_17166,N_11085,N_11598);
nand U17167 (N_17167,N_13519,N_14531);
and U17168 (N_17168,N_10473,N_10553);
and U17169 (N_17169,N_14263,N_13681);
xnor U17170 (N_17170,N_13835,N_12192);
nand U17171 (N_17171,N_14022,N_11876);
xor U17172 (N_17172,N_12346,N_10700);
nand U17173 (N_17173,N_11174,N_14487);
xnor U17174 (N_17174,N_11552,N_14513);
nor U17175 (N_17175,N_14434,N_10055);
and U17176 (N_17176,N_11016,N_14973);
nand U17177 (N_17177,N_14778,N_12031);
and U17178 (N_17178,N_10531,N_11641);
nand U17179 (N_17179,N_12167,N_12774);
xor U17180 (N_17180,N_14847,N_11889);
nand U17181 (N_17181,N_12361,N_12378);
xnor U17182 (N_17182,N_11612,N_11294);
nor U17183 (N_17183,N_10301,N_12680);
xor U17184 (N_17184,N_10274,N_10529);
xnor U17185 (N_17185,N_11923,N_13759);
nand U17186 (N_17186,N_14504,N_13591);
and U17187 (N_17187,N_10574,N_14042);
nor U17188 (N_17188,N_10348,N_12498);
xnor U17189 (N_17189,N_13099,N_10459);
or U17190 (N_17190,N_10161,N_12946);
nor U17191 (N_17191,N_11204,N_12567);
or U17192 (N_17192,N_10424,N_10476);
and U17193 (N_17193,N_13793,N_11608);
nand U17194 (N_17194,N_12292,N_13184);
or U17195 (N_17195,N_10426,N_11762);
or U17196 (N_17196,N_14755,N_11434);
and U17197 (N_17197,N_12105,N_11922);
or U17198 (N_17198,N_12770,N_14996);
nor U17199 (N_17199,N_10878,N_14336);
or U17200 (N_17200,N_12027,N_14589);
or U17201 (N_17201,N_13814,N_14338);
nor U17202 (N_17202,N_10310,N_14037);
nand U17203 (N_17203,N_13905,N_14730);
or U17204 (N_17204,N_14725,N_12090);
nor U17205 (N_17205,N_10090,N_13425);
nor U17206 (N_17206,N_10352,N_14392);
and U17207 (N_17207,N_10514,N_14519);
and U17208 (N_17208,N_13800,N_12523);
and U17209 (N_17209,N_10935,N_10131);
xnor U17210 (N_17210,N_11327,N_14269);
nor U17211 (N_17211,N_13092,N_14620);
or U17212 (N_17212,N_12603,N_14583);
nor U17213 (N_17213,N_14070,N_13970);
nor U17214 (N_17214,N_13574,N_11386);
nand U17215 (N_17215,N_10655,N_12368);
nor U17216 (N_17216,N_13769,N_12410);
nand U17217 (N_17217,N_14999,N_10223);
nand U17218 (N_17218,N_14899,N_12318);
and U17219 (N_17219,N_11242,N_11007);
nand U17220 (N_17220,N_12200,N_14387);
or U17221 (N_17221,N_14048,N_13116);
nand U17222 (N_17222,N_13438,N_10868);
nor U17223 (N_17223,N_12047,N_14258);
xnor U17224 (N_17224,N_10592,N_14184);
xor U17225 (N_17225,N_12096,N_10668);
nor U17226 (N_17226,N_11769,N_11541);
nand U17227 (N_17227,N_13436,N_10954);
nand U17228 (N_17228,N_12283,N_11086);
and U17229 (N_17229,N_13569,N_10475);
nand U17230 (N_17230,N_11570,N_13699);
nor U17231 (N_17231,N_12491,N_12739);
and U17232 (N_17232,N_10966,N_11305);
nand U17233 (N_17233,N_10357,N_11071);
and U17234 (N_17234,N_10838,N_14328);
and U17235 (N_17235,N_11521,N_13002);
nor U17236 (N_17236,N_14599,N_10669);
and U17237 (N_17237,N_10241,N_14653);
or U17238 (N_17238,N_12387,N_13244);
or U17239 (N_17239,N_10279,N_13604);
xor U17240 (N_17240,N_12961,N_11504);
xor U17241 (N_17241,N_10508,N_13329);
nor U17242 (N_17242,N_12965,N_14295);
nand U17243 (N_17243,N_13103,N_10600);
nor U17244 (N_17244,N_13348,N_10782);
or U17245 (N_17245,N_12848,N_12545);
or U17246 (N_17246,N_12500,N_10028);
and U17247 (N_17247,N_10032,N_13958);
or U17248 (N_17248,N_10816,N_13084);
xor U17249 (N_17249,N_10116,N_13178);
nor U17250 (N_17250,N_14117,N_11213);
and U17251 (N_17251,N_11046,N_10682);
nand U17252 (N_17252,N_14013,N_11575);
or U17253 (N_17253,N_14237,N_11253);
and U17254 (N_17254,N_12468,N_11763);
xnor U17255 (N_17255,N_11039,N_14656);
xor U17256 (N_17256,N_10432,N_13896);
nand U17257 (N_17257,N_10286,N_14062);
nor U17258 (N_17258,N_12022,N_10276);
or U17259 (N_17259,N_11649,N_14596);
and U17260 (N_17260,N_14382,N_12060);
or U17261 (N_17261,N_13581,N_13647);
nand U17262 (N_17262,N_13928,N_10198);
xor U17263 (N_17263,N_13750,N_14290);
nand U17264 (N_17264,N_14377,N_13666);
nor U17265 (N_17265,N_10461,N_14418);
or U17266 (N_17266,N_10510,N_14334);
nor U17267 (N_17267,N_11261,N_14898);
nor U17268 (N_17268,N_13489,N_12118);
and U17269 (N_17269,N_10860,N_10442);
or U17270 (N_17270,N_14871,N_14911);
and U17271 (N_17271,N_12888,N_13467);
or U17272 (N_17272,N_10444,N_14917);
or U17273 (N_17273,N_11223,N_10262);
xnor U17274 (N_17274,N_10809,N_14873);
nand U17275 (N_17275,N_11069,N_13662);
nor U17276 (N_17276,N_12054,N_14006);
xor U17277 (N_17277,N_12501,N_12592);
and U17278 (N_17278,N_12164,N_12439);
nor U17279 (N_17279,N_12011,N_11827);
nor U17280 (N_17280,N_11456,N_13650);
or U17281 (N_17281,N_13292,N_14972);
nand U17282 (N_17282,N_12729,N_14111);
xor U17283 (N_17283,N_12850,N_11061);
or U17284 (N_17284,N_14065,N_10051);
and U17285 (N_17285,N_14451,N_14810);
xor U17286 (N_17286,N_13533,N_10661);
nor U17287 (N_17287,N_13950,N_12450);
nand U17288 (N_17288,N_11138,N_14939);
nor U17289 (N_17289,N_12207,N_13713);
and U17290 (N_17290,N_11685,N_11960);
or U17291 (N_17291,N_13706,N_13324);
nand U17292 (N_17292,N_14788,N_14932);
or U17293 (N_17293,N_11700,N_12748);
nand U17294 (N_17294,N_11691,N_12885);
or U17295 (N_17295,N_14683,N_10632);
or U17296 (N_17296,N_14832,N_13081);
nand U17297 (N_17297,N_12430,N_11865);
nor U17298 (N_17298,N_10170,N_12058);
or U17299 (N_17299,N_11514,N_14238);
nor U17300 (N_17300,N_10814,N_12083);
nand U17301 (N_17301,N_13545,N_12255);
nand U17302 (N_17302,N_12787,N_10390);
xor U17303 (N_17303,N_13429,N_10464);
nand U17304 (N_17304,N_10292,N_12583);
xnor U17305 (N_17305,N_12930,N_10642);
nor U17306 (N_17306,N_12682,N_13772);
nor U17307 (N_17307,N_11731,N_14201);
xor U17308 (N_17308,N_11837,N_11924);
and U17309 (N_17309,N_11350,N_10603);
xor U17310 (N_17310,N_14433,N_12127);
nor U17311 (N_17311,N_12316,N_13492);
nor U17312 (N_17312,N_13032,N_13821);
nor U17313 (N_17313,N_11952,N_10836);
nand U17314 (N_17314,N_10483,N_13258);
xnor U17315 (N_17315,N_13523,N_12405);
nand U17316 (N_17316,N_13552,N_11508);
nand U17317 (N_17317,N_14619,N_13860);
xnor U17318 (N_17318,N_12713,N_10230);
nor U17319 (N_17319,N_10931,N_11241);
and U17320 (N_17320,N_11870,N_11905);
xnor U17321 (N_17321,N_14122,N_10667);
and U17322 (N_17322,N_14731,N_12732);
and U17323 (N_17323,N_11820,N_14325);
nand U17324 (N_17324,N_13087,N_11442);
xnor U17325 (N_17325,N_11139,N_14376);
or U17326 (N_17326,N_10358,N_11587);
and U17327 (N_17327,N_12817,N_13618);
nand U17328 (N_17328,N_11107,N_11471);
nor U17329 (N_17329,N_11145,N_10752);
nand U17330 (N_17330,N_10376,N_13463);
and U17331 (N_17331,N_11548,N_10063);
xor U17332 (N_17332,N_12539,N_10239);
xnor U17333 (N_17333,N_13149,N_10190);
xor U17334 (N_17334,N_14283,N_12133);
xor U17335 (N_17335,N_13204,N_10888);
nor U17336 (N_17336,N_12697,N_13756);
nand U17337 (N_17337,N_11122,N_13664);
xnor U17338 (N_17338,N_11079,N_11917);
nand U17339 (N_17339,N_14794,N_10794);
and U17340 (N_17340,N_10171,N_12402);
and U17341 (N_17341,N_11279,N_10958);
nand U17342 (N_17342,N_10658,N_10936);
xnor U17343 (N_17343,N_11822,N_13460);
nand U17344 (N_17344,N_11230,N_10769);
or U17345 (N_17345,N_13070,N_12470);
xor U17346 (N_17346,N_12419,N_14723);
xor U17347 (N_17347,N_10341,N_12473);
nand U17348 (N_17348,N_12687,N_10204);
nor U17349 (N_17349,N_10412,N_12623);
nand U17350 (N_17350,N_12809,N_14501);
xnor U17351 (N_17351,N_14083,N_11159);
nand U17352 (N_17352,N_12365,N_10664);
or U17353 (N_17353,N_10451,N_10937);
and U17354 (N_17354,N_12456,N_11454);
xor U17355 (N_17355,N_13495,N_10721);
and U17356 (N_17356,N_14803,N_13274);
and U17357 (N_17357,N_13040,N_11701);
and U17358 (N_17358,N_14967,N_10151);
and U17359 (N_17359,N_12512,N_13171);
and U17360 (N_17360,N_14278,N_11205);
and U17361 (N_17361,N_11524,N_10458);
nor U17362 (N_17362,N_13350,N_14780);
nor U17363 (N_17363,N_14989,N_10568);
nand U17364 (N_17364,N_12477,N_14372);
nor U17365 (N_17365,N_10716,N_13822);
nor U17366 (N_17366,N_13220,N_12078);
or U17367 (N_17367,N_11326,N_14240);
xor U17368 (N_17368,N_10988,N_14236);
or U17369 (N_17369,N_13430,N_12414);
xor U17370 (N_17370,N_12918,N_12641);
nor U17371 (N_17371,N_10617,N_12464);
and U17372 (N_17372,N_11501,N_14570);
or U17373 (N_17373,N_11221,N_10548);
xor U17374 (N_17374,N_14716,N_14662);
or U17375 (N_17375,N_14133,N_10472);
or U17376 (N_17376,N_14963,N_11392);
xor U17377 (N_17377,N_13597,N_13331);
and U17378 (N_17378,N_13138,N_10094);
nand U17379 (N_17379,N_11578,N_14526);
and U17380 (N_17380,N_11602,N_12556);
or U17381 (N_17381,N_12195,N_13735);
xor U17382 (N_17382,N_13760,N_10733);
xnor U17383 (N_17383,N_10562,N_11964);
nor U17384 (N_17384,N_12757,N_11298);
or U17385 (N_17385,N_14183,N_10110);
and U17386 (N_17386,N_12057,N_14707);
nor U17387 (N_17387,N_13875,N_13637);
or U17388 (N_17388,N_11934,N_14398);
xor U17389 (N_17389,N_11930,N_14833);
or U17390 (N_17390,N_13072,N_13883);
nor U17391 (N_17391,N_11802,N_10923);
and U17392 (N_17392,N_11418,N_14700);
or U17393 (N_17393,N_14561,N_14714);
xor U17394 (N_17394,N_11630,N_11783);
or U17395 (N_17395,N_13076,N_10047);
and U17396 (N_17396,N_14214,N_11402);
nor U17397 (N_17397,N_10647,N_13056);
xor U17398 (N_17398,N_14938,N_11393);
nand U17399 (N_17399,N_13365,N_13363);
nor U17400 (N_17400,N_13442,N_14776);
and U17401 (N_17401,N_11675,N_11746);
xor U17402 (N_17402,N_10503,N_10477);
and U17403 (N_17403,N_11538,N_12886);
nor U17404 (N_17404,N_12166,N_10319);
nand U17405 (N_17405,N_12504,N_12299);
nor U17406 (N_17406,N_14554,N_10502);
xnor U17407 (N_17407,N_11108,N_13558);
nor U17408 (N_17408,N_10740,N_13506);
or U17409 (N_17409,N_10408,N_14565);
or U17410 (N_17410,N_13276,N_11943);
nor U17411 (N_17411,N_12522,N_13353);
or U17412 (N_17412,N_10210,N_11743);
and U17413 (N_17413,N_10524,N_12376);
xnor U17414 (N_17414,N_11133,N_12865);
xor U17415 (N_17415,N_11858,N_10228);
xnor U17416 (N_17416,N_10263,N_10163);
nand U17417 (N_17417,N_11516,N_12650);
and U17418 (N_17418,N_12937,N_10384);
nor U17419 (N_17419,N_14188,N_11120);
xor U17420 (N_17420,N_10217,N_11412);
or U17421 (N_17421,N_11838,N_11041);
and U17422 (N_17422,N_14831,N_12421);
nand U17423 (N_17423,N_11457,N_11289);
or U17424 (N_17424,N_13398,N_12461);
or U17425 (N_17425,N_12784,N_10383);
xnor U17426 (N_17426,N_11100,N_12359);
or U17427 (N_17427,N_13794,N_11758);
and U17428 (N_17428,N_12377,N_10802);
or U17429 (N_17429,N_13856,N_12796);
nand U17430 (N_17430,N_11809,N_14629);
or U17431 (N_17431,N_14316,N_13789);
or U17432 (N_17432,N_14043,N_14116);
nor U17433 (N_17433,N_11529,N_13732);
nand U17434 (N_17434,N_13994,N_14301);
or U17435 (N_17435,N_12069,N_14349);
or U17436 (N_17436,N_10910,N_10106);
or U17437 (N_17437,N_11075,N_14177);
or U17438 (N_17438,N_11855,N_13646);
or U17439 (N_17439,N_13071,N_14113);
nor U17440 (N_17440,N_10419,N_13757);
nand U17441 (N_17441,N_13308,N_11990);
and U17442 (N_17442,N_14848,N_14347);
or U17443 (N_17443,N_14746,N_11246);
xnor U17444 (N_17444,N_13988,N_11263);
nor U17445 (N_17445,N_13936,N_13585);
nor U17446 (N_17446,N_13479,N_10122);
and U17447 (N_17447,N_13135,N_14708);
or U17448 (N_17448,N_14579,N_14036);
or U17449 (N_17449,N_13176,N_13268);
nor U17450 (N_17450,N_14142,N_13855);
or U17451 (N_17451,N_14223,N_14934);
and U17452 (N_17452,N_12261,N_10059);
and U17453 (N_17453,N_10380,N_12235);
nor U17454 (N_17454,N_10173,N_14804);
nand U17455 (N_17455,N_10675,N_14577);
nand U17456 (N_17456,N_13862,N_11450);
nor U17457 (N_17457,N_11451,N_11480);
nand U17458 (N_17458,N_10314,N_10623);
nand U17459 (N_17459,N_10750,N_13700);
xor U17460 (N_17460,N_12554,N_11052);
xor U17461 (N_17461,N_10321,N_12304);
and U17462 (N_17462,N_12140,N_13137);
nand U17463 (N_17463,N_14461,N_12581);
and U17464 (N_17464,N_12989,N_13322);
or U17465 (N_17465,N_13844,N_13311);
nor U17466 (N_17466,N_11308,N_13123);
or U17467 (N_17467,N_10184,N_14694);
and U17468 (N_17468,N_12017,N_14753);
or U17469 (N_17469,N_11805,N_11509);
or U17470 (N_17470,N_12012,N_11698);
xor U17471 (N_17471,N_12475,N_11775);
nand U17472 (N_17472,N_13125,N_13837);
xor U17473 (N_17473,N_12275,N_14195);
or U17474 (N_17474,N_10397,N_13746);
xor U17475 (N_17475,N_12394,N_13314);
nand U17476 (N_17476,N_11813,N_13843);
xor U17477 (N_17477,N_13188,N_10943);
nor U17478 (N_17478,N_13947,N_14705);
nor U17479 (N_17479,N_14060,N_10768);
nor U17480 (N_17480,N_14199,N_13080);
xor U17481 (N_17481,N_13667,N_12580);
nor U17482 (N_17482,N_10231,N_10839);
or U17483 (N_17483,N_10538,N_10205);
or U17484 (N_17484,N_13693,N_14420);
or U17485 (N_17485,N_11135,N_10237);
nor U17486 (N_17486,N_10117,N_11554);
and U17487 (N_17487,N_10706,N_14162);
nor U17488 (N_17488,N_10678,N_10648);
xnor U17489 (N_17489,N_11901,N_10370);
or U17490 (N_17490,N_11671,N_12723);
and U17491 (N_17491,N_11110,N_11184);
and U17492 (N_17492,N_11119,N_10112);
xnor U17493 (N_17493,N_13194,N_12330);
xnor U17494 (N_17494,N_14310,N_10731);
xnor U17495 (N_17495,N_10709,N_12007);
and U17496 (N_17496,N_13622,N_11588);
nand U17497 (N_17497,N_11555,N_14285);
xor U17498 (N_17498,N_14164,N_12443);
nand U17499 (N_17499,N_12367,N_13105);
xor U17500 (N_17500,N_13068,N_12756);
xnor U17501 (N_17501,N_13610,N_13645);
and U17502 (N_17502,N_12275,N_11503);
or U17503 (N_17503,N_14483,N_13052);
nand U17504 (N_17504,N_12625,N_13954);
or U17505 (N_17505,N_10992,N_12972);
and U17506 (N_17506,N_12440,N_13105);
nor U17507 (N_17507,N_11326,N_10328);
xnor U17508 (N_17508,N_10188,N_13221);
or U17509 (N_17509,N_13225,N_14806);
xnor U17510 (N_17510,N_11518,N_14254);
nand U17511 (N_17511,N_10659,N_10281);
and U17512 (N_17512,N_12996,N_14824);
nand U17513 (N_17513,N_13384,N_14887);
xor U17514 (N_17514,N_13827,N_11061);
xor U17515 (N_17515,N_10151,N_11596);
or U17516 (N_17516,N_12575,N_14981);
or U17517 (N_17517,N_10448,N_11299);
nor U17518 (N_17518,N_14124,N_12642);
nand U17519 (N_17519,N_14735,N_10568);
and U17520 (N_17520,N_13704,N_14118);
nand U17521 (N_17521,N_14601,N_14325);
xnor U17522 (N_17522,N_11228,N_14640);
or U17523 (N_17523,N_14514,N_10491);
nor U17524 (N_17524,N_13753,N_11926);
or U17525 (N_17525,N_13396,N_12629);
or U17526 (N_17526,N_10711,N_10555);
and U17527 (N_17527,N_10984,N_12385);
nor U17528 (N_17528,N_11242,N_14924);
nand U17529 (N_17529,N_11170,N_10390);
and U17530 (N_17530,N_11561,N_13369);
nor U17531 (N_17531,N_11143,N_11047);
nand U17532 (N_17532,N_14207,N_12738);
xor U17533 (N_17533,N_11117,N_13547);
or U17534 (N_17534,N_10606,N_11764);
nand U17535 (N_17535,N_13537,N_12584);
xor U17536 (N_17536,N_12848,N_10606);
or U17537 (N_17537,N_13795,N_10402);
or U17538 (N_17538,N_14998,N_10338);
xnor U17539 (N_17539,N_13902,N_11387);
or U17540 (N_17540,N_10559,N_11873);
nor U17541 (N_17541,N_14196,N_13012);
nor U17542 (N_17542,N_14285,N_14130);
nand U17543 (N_17543,N_12117,N_13756);
nand U17544 (N_17544,N_14645,N_14482);
and U17545 (N_17545,N_11396,N_10544);
and U17546 (N_17546,N_11705,N_12865);
nor U17547 (N_17547,N_13074,N_11343);
and U17548 (N_17548,N_12735,N_10034);
nor U17549 (N_17549,N_11092,N_14713);
nand U17550 (N_17550,N_12948,N_10708);
and U17551 (N_17551,N_14692,N_14292);
and U17552 (N_17552,N_14357,N_11888);
nor U17553 (N_17553,N_14957,N_10074);
nor U17554 (N_17554,N_13103,N_12657);
and U17555 (N_17555,N_10153,N_12301);
or U17556 (N_17556,N_12431,N_11020);
nor U17557 (N_17557,N_14214,N_10603);
or U17558 (N_17558,N_10638,N_12590);
xor U17559 (N_17559,N_11453,N_13868);
or U17560 (N_17560,N_10150,N_13428);
nor U17561 (N_17561,N_13016,N_14873);
nor U17562 (N_17562,N_12300,N_11374);
nor U17563 (N_17563,N_10915,N_10518);
and U17564 (N_17564,N_14121,N_12291);
and U17565 (N_17565,N_14094,N_12429);
xnor U17566 (N_17566,N_13033,N_12440);
nand U17567 (N_17567,N_13469,N_11910);
nand U17568 (N_17568,N_13260,N_13643);
xnor U17569 (N_17569,N_12336,N_11418);
or U17570 (N_17570,N_10200,N_12324);
nor U17571 (N_17571,N_12230,N_13511);
or U17572 (N_17572,N_13547,N_12605);
xnor U17573 (N_17573,N_13791,N_11242);
and U17574 (N_17574,N_12415,N_13257);
and U17575 (N_17575,N_14986,N_10958);
nor U17576 (N_17576,N_12860,N_14101);
xor U17577 (N_17577,N_11732,N_14841);
nor U17578 (N_17578,N_13741,N_10578);
xor U17579 (N_17579,N_12057,N_11250);
or U17580 (N_17580,N_13614,N_14323);
nor U17581 (N_17581,N_10611,N_13887);
nor U17582 (N_17582,N_12240,N_11711);
or U17583 (N_17583,N_14513,N_10524);
nor U17584 (N_17584,N_14267,N_11808);
nand U17585 (N_17585,N_10965,N_14652);
and U17586 (N_17586,N_11548,N_11110);
xnor U17587 (N_17587,N_10987,N_11831);
or U17588 (N_17588,N_14281,N_10658);
nor U17589 (N_17589,N_14183,N_14358);
or U17590 (N_17590,N_10864,N_14128);
nor U17591 (N_17591,N_11949,N_13041);
xnor U17592 (N_17592,N_10540,N_13488);
xor U17593 (N_17593,N_13686,N_12373);
nor U17594 (N_17594,N_10406,N_10607);
nand U17595 (N_17595,N_13286,N_13626);
xor U17596 (N_17596,N_12148,N_12800);
or U17597 (N_17597,N_13141,N_13288);
xnor U17598 (N_17598,N_14366,N_12196);
xnor U17599 (N_17599,N_10224,N_14825);
or U17600 (N_17600,N_10618,N_14937);
xnor U17601 (N_17601,N_13305,N_13502);
or U17602 (N_17602,N_10151,N_14711);
or U17603 (N_17603,N_11705,N_12431);
nor U17604 (N_17604,N_13470,N_10131);
nand U17605 (N_17605,N_14022,N_12312);
and U17606 (N_17606,N_13345,N_12602);
nand U17607 (N_17607,N_14482,N_12481);
nor U17608 (N_17608,N_11061,N_12879);
nand U17609 (N_17609,N_13682,N_10797);
nor U17610 (N_17610,N_11145,N_10243);
nand U17611 (N_17611,N_11856,N_11538);
and U17612 (N_17612,N_13133,N_13558);
xor U17613 (N_17613,N_12065,N_14177);
nor U17614 (N_17614,N_10075,N_10106);
nand U17615 (N_17615,N_12855,N_12753);
or U17616 (N_17616,N_12952,N_14772);
and U17617 (N_17617,N_11017,N_14297);
nor U17618 (N_17618,N_11260,N_13502);
and U17619 (N_17619,N_14886,N_10840);
xnor U17620 (N_17620,N_13745,N_10920);
nand U17621 (N_17621,N_13884,N_13105);
xnor U17622 (N_17622,N_12402,N_13125);
nand U17623 (N_17623,N_10038,N_11930);
and U17624 (N_17624,N_10042,N_13626);
and U17625 (N_17625,N_11114,N_14325);
and U17626 (N_17626,N_13805,N_14302);
nor U17627 (N_17627,N_10161,N_13151);
nand U17628 (N_17628,N_10505,N_10272);
xnor U17629 (N_17629,N_11526,N_12182);
or U17630 (N_17630,N_10080,N_10754);
or U17631 (N_17631,N_14780,N_14852);
nor U17632 (N_17632,N_14954,N_12821);
nand U17633 (N_17633,N_10871,N_11060);
or U17634 (N_17634,N_13537,N_12162);
nand U17635 (N_17635,N_14659,N_13070);
and U17636 (N_17636,N_12610,N_11552);
nor U17637 (N_17637,N_14661,N_12323);
and U17638 (N_17638,N_14125,N_11959);
nor U17639 (N_17639,N_14683,N_14669);
and U17640 (N_17640,N_14731,N_12281);
xor U17641 (N_17641,N_13841,N_10275);
xnor U17642 (N_17642,N_12777,N_10903);
xor U17643 (N_17643,N_13802,N_10573);
or U17644 (N_17644,N_12771,N_12757);
nor U17645 (N_17645,N_12245,N_10380);
xor U17646 (N_17646,N_14282,N_12364);
nand U17647 (N_17647,N_14743,N_13381);
or U17648 (N_17648,N_13870,N_11882);
or U17649 (N_17649,N_12498,N_14182);
nand U17650 (N_17650,N_12406,N_12292);
or U17651 (N_17651,N_11858,N_13235);
xor U17652 (N_17652,N_13573,N_14696);
nor U17653 (N_17653,N_14107,N_10160);
and U17654 (N_17654,N_12110,N_14434);
and U17655 (N_17655,N_11426,N_12814);
nor U17656 (N_17656,N_13897,N_11071);
nor U17657 (N_17657,N_11046,N_11531);
xor U17658 (N_17658,N_11387,N_13556);
nor U17659 (N_17659,N_14981,N_11018);
nor U17660 (N_17660,N_10637,N_13920);
nand U17661 (N_17661,N_12673,N_12083);
xor U17662 (N_17662,N_10489,N_13901);
nor U17663 (N_17663,N_10680,N_13310);
or U17664 (N_17664,N_11768,N_14542);
xnor U17665 (N_17665,N_11754,N_11142);
nand U17666 (N_17666,N_12164,N_13016);
xnor U17667 (N_17667,N_11287,N_10169);
nand U17668 (N_17668,N_12389,N_12663);
or U17669 (N_17669,N_10574,N_12367);
or U17670 (N_17670,N_12886,N_11235);
nor U17671 (N_17671,N_11622,N_11576);
xor U17672 (N_17672,N_14083,N_13313);
or U17673 (N_17673,N_12077,N_10811);
and U17674 (N_17674,N_11188,N_14714);
or U17675 (N_17675,N_10573,N_14700);
nor U17676 (N_17676,N_11132,N_14564);
or U17677 (N_17677,N_14171,N_12303);
and U17678 (N_17678,N_13222,N_14216);
nor U17679 (N_17679,N_14517,N_11954);
or U17680 (N_17680,N_10436,N_10283);
xnor U17681 (N_17681,N_10986,N_13302);
and U17682 (N_17682,N_10068,N_11912);
xnor U17683 (N_17683,N_13903,N_14869);
nand U17684 (N_17684,N_10459,N_12181);
nor U17685 (N_17685,N_12976,N_12152);
or U17686 (N_17686,N_12981,N_13516);
or U17687 (N_17687,N_10669,N_12631);
nand U17688 (N_17688,N_10895,N_13166);
nor U17689 (N_17689,N_11462,N_10196);
xor U17690 (N_17690,N_13621,N_10058);
xnor U17691 (N_17691,N_14245,N_10444);
or U17692 (N_17692,N_10661,N_11812);
nor U17693 (N_17693,N_11822,N_11933);
or U17694 (N_17694,N_12601,N_12860);
or U17695 (N_17695,N_14581,N_13303);
or U17696 (N_17696,N_12556,N_14005);
or U17697 (N_17697,N_11795,N_13023);
and U17698 (N_17698,N_10009,N_14399);
nand U17699 (N_17699,N_12628,N_11834);
and U17700 (N_17700,N_13143,N_12285);
or U17701 (N_17701,N_10135,N_10173);
nand U17702 (N_17702,N_10076,N_13139);
or U17703 (N_17703,N_10399,N_14681);
and U17704 (N_17704,N_12928,N_12681);
xnor U17705 (N_17705,N_13305,N_14315);
xnor U17706 (N_17706,N_14688,N_12864);
and U17707 (N_17707,N_13431,N_10139);
nor U17708 (N_17708,N_10087,N_12041);
xnor U17709 (N_17709,N_12871,N_12269);
or U17710 (N_17710,N_10936,N_10540);
and U17711 (N_17711,N_13697,N_10155);
nand U17712 (N_17712,N_10405,N_13160);
nand U17713 (N_17713,N_13458,N_12227);
or U17714 (N_17714,N_10623,N_10867);
and U17715 (N_17715,N_11283,N_12109);
xor U17716 (N_17716,N_14619,N_13438);
nor U17717 (N_17717,N_13812,N_11415);
nand U17718 (N_17718,N_13611,N_10268);
nand U17719 (N_17719,N_11115,N_13574);
nor U17720 (N_17720,N_14881,N_13597);
nor U17721 (N_17721,N_12612,N_11283);
nor U17722 (N_17722,N_12287,N_12099);
and U17723 (N_17723,N_10450,N_14304);
or U17724 (N_17724,N_13340,N_14421);
and U17725 (N_17725,N_13724,N_10770);
and U17726 (N_17726,N_10536,N_14715);
nor U17727 (N_17727,N_10383,N_13958);
xnor U17728 (N_17728,N_11848,N_11682);
nand U17729 (N_17729,N_11393,N_12735);
nand U17730 (N_17730,N_11207,N_11285);
or U17731 (N_17731,N_14363,N_14345);
or U17732 (N_17732,N_12682,N_14544);
or U17733 (N_17733,N_12581,N_13262);
and U17734 (N_17734,N_13012,N_13624);
nand U17735 (N_17735,N_11308,N_14079);
or U17736 (N_17736,N_13970,N_10708);
and U17737 (N_17737,N_14472,N_14261);
and U17738 (N_17738,N_12916,N_14823);
and U17739 (N_17739,N_10520,N_10558);
and U17740 (N_17740,N_10480,N_10236);
and U17741 (N_17741,N_14862,N_11883);
nand U17742 (N_17742,N_10793,N_13357);
xnor U17743 (N_17743,N_10192,N_11917);
nor U17744 (N_17744,N_12242,N_14515);
and U17745 (N_17745,N_14151,N_11870);
or U17746 (N_17746,N_14426,N_12192);
nand U17747 (N_17747,N_14715,N_13353);
xor U17748 (N_17748,N_13446,N_12513);
nand U17749 (N_17749,N_13974,N_12798);
nand U17750 (N_17750,N_13788,N_13718);
or U17751 (N_17751,N_11652,N_14108);
xnor U17752 (N_17752,N_10192,N_10708);
xor U17753 (N_17753,N_14387,N_14352);
nand U17754 (N_17754,N_10919,N_11397);
and U17755 (N_17755,N_11873,N_11741);
or U17756 (N_17756,N_11890,N_12485);
nand U17757 (N_17757,N_11968,N_13968);
and U17758 (N_17758,N_14961,N_13641);
and U17759 (N_17759,N_13471,N_14184);
nor U17760 (N_17760,N_10459,N_14890);
xor U17761 (N_17761,N_12921,N_10695);
xor U17762 (N_17762,N_11510,N_12970);
nor U17763 (N_17763,N_10152,N_11904);
and U17764 (N_17764,N_13305,N_14457);
nand U17765 (N_17765,N_12759,N_12315);
nor U17766 (N_17766,N_14777,N_12315);
nand U17767 (N_17767,N_14210,N_12241);
nor U17768 (N_17768,N_11322,N_13711);
and U17769 (N_17769,N_14802,N_10198);
xnor U17770 (N_17770,N_14368,N_10264);
and U17771 (N_17771,N_11563,N_14185);
nor U17772 (N_17772,N_11563,N_14702);
and U17773 (N_17773,N_13857,N_13881);
nor U17774 (N_17774,N_13331,N_11241);
xnor U17775 (N_17775,N_14932,N_11454);
or U17776 (N_17776,N_13739,N_11697);
and U17777 (N_17777,N_12386,N_10792);
xor U17778 (N_17778,N_12909,N_14154);
nand U17779 (N_17779,N_10884,N_11961);
nor U17780 (N_17780,N_12335,N_13429);
xor U17781 (N_17781,N_12380,N_13659);
and U17782 (N_17782,N_10937,N_14366);
or U17783 (N_17783,N_10828,N_13307);
nor U17784 (N_17784,N_14941,N_12857);
xnor U17785 (N_17785,N_11459,N_12767);
or U17786 (N_17786,N_13097,N_11883);
nor U17787 (N_17787,N_12774,N_11658);
or U17788 (N_17788,N_11270,N_14252);
nor U17789 (N_17789,N_13206,N_12476);
nand U17790 (N_17790,N_11678,N_13252);
nor U17791 (N_17791,N_10341,N_10225);
or U17792 (N_17792,N_14550,N_11476);
nor U17793 (N_17793,N_14922,N_10305);
and U17794 (N_17794,N_13286,N_14029);
and U17795 (N_17795,N_14814,N_11941);
or U17796 (N_17796,N_10896,N_10938);
nand U17797 (N_17797,N_10960,N_13383);
and U17798 (N_17798,N_13411,N_14039);
or U17799 (N_17799,N_13805,N_13330);
and U17800 (N_17800,N_13616,N_12749);
xor U17801 (N_17801,N_11490,N_13088);
xnor U17802 (N_17802,N_14046,N_12308);
nand U17803 (N_17803,N_12697,N_14538);
nor U17804 (N_17804,N_13920,N_14759);
nand U17805 (N_17805,N_12138,N_13115);
or U17806 (N_17806,N_10453,N_12386);
or U17807 (N_17807,N_11984,N_14352);
xor U17808 (N_17808,N_14943,N_13685);
or U17809 (N_17809,N_12636,N_11045);
or U17810 (N_17810,N_11773,N_14649);
or U17811 (N_17811,N_13046,N_14365);
and U17812 (N_17812,N_10755,N_11623);
nand U17813 (N_17813,N_14568,N_13769);
nor U17814 (N_17814,N_12895,N_12542);
xor U17815 (N_17815,N_11410,N_10012);
nor U17816 (N_17816,N_13968,N_10278);
or U17817 (N_17817,N_10588,N_13089);
and U17818 (N_17818,N_12570,N_14963);
nand U17819 (N_17819,N_11150,N_14886);
and U17820 (N_17820,N_14570,N_12294);
nor U17821 (N_17821,N_13449,N_12057);
nand U17822 (N_17822,N_10031,N_14157);
and U17823 (N_17823,N_12508,N_10675);
nor U17824 (N_17824,N_12945,N_10138);
nand U17825 (N_17825,N_11983,N_12610);
nand U17826 (N_17826,N_14514,N_11857);
xnor U17827 (N_17827,N_10796,N_11731);
nor U17828 (N_17828,N_10540,N_14142);
xnor U17829 (N_17829,N_12742,N_14607);
nor U17830 (N_17830,N_11604,N_10211);
or U17831 (N_17831,N_14296,N_13659);
nand U17832 (N_17832,N_12319,N_10193);
nand U17833 (N_17833,N_13125,N_14632);
xor U17834 (N_17834,N_10354,N_14419);
nand U17835 (N_17835,N_12617,N_11921);
or U17836 (N_17836,N_12602,N_11737);
or U17837 (N_17837,N_11593,N_10546);
nor U17838 (N_17838,N_14326,N_14660);
or U17839 (N_17839,N_11262,N_11480);
and U17840 (N_17840,N_10745,N_10464);
and U17841 (N_17841,N_12893,N_11255);
or U17842 (N_17842,N_11189,N_12437);
and U17843 (N_17843,N_13397,N_12820);
nand U17844 (N_17844,N_12093,N_14759);
and U17845 (N_17845,N_11876,N_12464);
and U17846 (N_17846,N_14061,N_12622);
nor U17847 (N_17847,N_14165,N_10849);
nand U17848 (N_17848,N_11146,N_13751);
or U17849 (N_17849,N_10382,N_12863);
xnor U17850 (N_17850,N_13033,N_13503);
nand U17851 (N_17851,N_11109,N_12796);
xnor U17852 (N_17852,N_14883,N_13832);
nand U17853 (N_17853,N_14232,N_12651);
xor U17854 (N_17854,N_11183,N_13829);
or U17855 (N_17855,N_13573,N_14971);
nor U17856 (N_17856,N_14004,N_12692);
nand U17857 (N_17857,N_14827,N_13504);
nor U17858 (N_17858,N_13758,N_12987);
nor U17859 (N_17859,N_13266,N_11866);
nand U17860 (N_17860,N_11379,N_11609);
and U17861 (N_17861,N_13410,N_11166);
or U17862 (N_17862,N_12108,N_11247);
and U17863 (N_17863,N_12730,N_10977);
nand U17864 (N_17864,N_11556,N_10404);
xor U17865 (N_17865,N_10574,N_12159);
nand U17866 (N_17866,N_13672,N_10546);
or U17867 (N_17867,N_13803,N_12131);
nor U17868 (N_17868,N_14450,N_13383);
nor U17869 (N_17869,N_12866,N_11474);
or U17870 (N_17870,N_11204,N_10972);
nor U17871 (N_17871,N_13542,N_11279);
xor U17872 (N_17872,N_14990,N_12131);
nand U17873 (N_17873,N_11224,N_12493);
nand U17874 (N_17874,N_14252,N_13829);
xnor U17875 (N_17875,N_10416,N_12169);
xor U17876 (N_17876,N_14450,N_11812);
nor U17877 (N_17877,N_11878,N_11837);
and U17878 (N_17878,N_10642,N_14423);
or U17879 (N_17879,N_10319,N_14579);
xor U17880 (N_17880,N_11626,N_12083);
nand U17881 (N_17881,N_12483,N_12474);
xor U17882 (N_17882,N_13225,N_10862);
and U17883 (N_17883,N_14793,N_12225);
and U17884 (N_17884,N_10760,N_11660);
or U17885 (N_17885,N_13894,N_11965);
and U17886 (N_17886,N_11285,N_14047);
and U17887 (N_17887,N_11328,N_14922);
nor U17888 (N_17888,N_11360,N_10371);
or U17889 (N_17889,N_13865,N_11162);
nor U17890 (N_17890,N_10362,N_14980);
nand U17891 (N_17891,N_10636,N_10981);
or U17892 (N_17892,N_12142,N_14707);
nand U17893 (N_17893,N_12376,N_14919);
xor U17894 (N_17894,N_12416,N_10973);
or U17895 (N_17895,N_12774,N_10554);
nand U17896 (N_17896,N_14930,N_14139);
nand U17897 (N_17897,N_14268,N_10825);
nor U17898 (N_17898,N_12897,N_13813);
xor U17899 (N_17899,N_14704,N_10238);
xor U17900 (N_17900,N_13271,N_14599);
or U17901 (N_17901,N_11547,N_10291);
and U17902 (N_17902,N_11835,N_14753);
nand U17903 (N_17903,N_13461,N_13868);
and U17904 (N_17904,N_10746,N_13633);
xnor U17905 (N_17905,N_12275,N_10643);
or U17906 (N_17906,N_11807,N_10803);
and U17907 (N_17907,N_12998,N_10359);
nand U17908 (N_17908,N_13572,N_10463);
or U17909 (N_17909,N_13895,N_14715);
nor U17910 (N_17910,N_13706,N_11677);
xnor U17911 (N_17911,N_13579,N_14662);
and U17912 (N_17912,N_14394,N_14820);
xnor U17913 (N_17913,N_12406,N_10038);
or U17914 (N_17914,N_11661,N_12988);
xor U17915 (N_17915,N_11909,N_11954);
nand U17916 (N_17916,N_10884,N_11746);
nand U17917 (N_17917,N_10785,N_13144);
and U17918 (N_17918,N_12342,N_13441);
and U17919 (N_17919,N_11179,N_10962);
nor U17920 (N_17920,N_11388,N_13479);
or U17921 (N_17921,N_12241,N_13831);
or U17922 (N_17922,N_12877,N_13042);
nor U17923 (N_17923,N_10798,N_12906);
nor U17924 (N_17924,N_13925,N_10534);
nor U17925 (N_17925,N_13844,N_14340);
or U17926 (N_17926,N_12187,N_13911);
and U17927 (N_17927,N_14597,N_12611);
xnor U17928 (N_17928,N_14073,N_11881);
and U17929 (N_17929,N_13146,N_12031);
or U17930 (N_17930,N_14368,N_14644);
nor U17931 (N_17931,N_12055,N_13152);
and U17932 (N_17932,N_12052,N_12546);
or U17933 (N_17933,N_11768,N_12618);
xor U17934 (N_17934,N_13670,N_12295);
xnor U17935 (N_17935,N_11698,N_14554);
nor U17936 (N_17936,N_12031,N_13215);
nor U17937 (N_17937,N_12451,N_12515);
nand U17938 (N_17938,N_14258,N_10638);
nor U17939 (N_17939,N_13345,N_14521);
or U17940 (N_17940,N_12832,N_14710);
nand U17941 (N_17941,N_11648,N_14176);
or U17942 (N_17942,N_11067,N_14402);
or U17943 (N_17943,N_11723,N_10195);
xnor U17944 (N_17944,N_10960,N_13812);
and U17945 (N_17945,N_12535,N_11108);
nand U17946 (N_17946,N_11831,N_12114);
nand U17947 (N_17947,N_12241,N_13622);
nor U17948 (N_17948,N_13135,N_12400);
nor U17949 (N_17949,N_11856,N_12031);
and U17950 (N_17950,N_10554,N_10940);
or U17951 (N_17951,N_14961,N_12433);
and U17952 (N_17952,N_13854,N_11602);
nand U17953 (N_17953,N_10762,N_12463);
nor U17954 (N_17954,N_12078,N_13329);
xor U17955 (N_17955,N_10192,N_13514);
nand U17956 (N_17956,N_13672,N_13070);
xnor U17957 (N_17957,N_12312,N_11914);
nor U17958 (N_17958,N_10851,N_14305);
nand U17959 (N_17959,N_11379,N_12876);
nor U17960 (N_17960,N_13691,N_14937);
xor U17961 (N_17961,N_10409,N_12260);
and U17962 (N_17962,N_14635,N_13377);
nand U17963 (N_17963,N_13077,N_11421);
nor U17964 (N_17964,N_11523,N_10808);
or U17965 (N_17965,N_12878,N_11616);
nand U17966 (N_17966,N_14854,N_14680);
and U17967 (N_17967,N_11229,N_14836);
or U17968 (N_17968,N_11636,N_12360);
and U17969 (N_17969,N_13527,N_14496);
nand U17970 (N_17970,N_10741,N_12356);
xnor U17971 (N_17971,N_13204,N_11915);
nor U17972 (N_17972,N_10700,N_11999);
and U17973 (N_17973,N_11380,N_14276);
nand U17974 (N_17974,N_13949,N_11811);
and U17975 (N_17975,N_13883,N_10993);
or U17976 (N_17976,N_10171,N_11987);
nor U17977 (N_17977,N_14009,N_12170);
xor U17978 (N_17978,N_12488,N_10744);
xnor U17979 (N_17979,N_10828,N_14377);
nand U17980 (N_17980,N_11237,N_12853);
nor U17981 (N_17981,N_10812,N_12069);
or U17982 (N_17982,N_14739,N_10647);
or U17983 (N_17983,N_11025,N_11763);
nor U17984 (N_17984,N_14602,N_10804);
nand U17985 (N_17985,N_14350,N_13056);
nand U17986 (N_17986,N_10923,N_14685);
and U17987 (N_17987,N_10570,N_10038);
nand U17988 (N_17988,N_12467,N_13613);
and U17989 (N_17989,N_13110,N_14378);
and U17990 (N_17990,N_12046,N_13121);
nand U17991 (N_17991,N_10352,N_10224);
nor U17992 (N_17992,N_10844,N_13088);
and U17993 (N_17993,N_10681,N_13110);
or U17994 (N_17994,N_11917,N_11519);
nor U17995 (N_17995,N_10239,N_13659);
or U17996 (N_17996,N_11870,N_12909);
nand U17997 (N_17997,N_13698,N_12967);
and U17998 (N_17998,N_10030,N_13652);
and U17999 (N_17999,N_12694,N_11515);
and U18000 (N_18000,N_10744,N_12772);
or U18001 (N_18001,N_10559,N_12614);
xor U18002 (N_18002,N_12150,N_13651);
nor U18003 (N_18003,N_11162,N_10806);
or U18004 (N_18004,N_13725,N_12641);
nor U18005 (N_18005,N_14764,N_10133);
or U18006 (N_18006,N_10810,N_13383);
nor U18007 (N_18007,N_13673,N_11175);
nor U18008 (N_18008,N_12963,N_10621);
nand U18009 (N_18009,N_14095,N_11638);
and U18010 (N_18010,N_11422,N_13360);
and U18011 (N_18011,N_14580,N_10900);
nand U18012 (N_18012,N_13560,N_14130);
or U18013 (N_18013,N_11449,N_10796);
xor U18014 (N_18014,N_12888,N_13834);
and U18015 (N_18015,N_13572,N_11205);
and U18016 (N_18016,N_12738,N_11460);
xnor U18017 (N_18017,N_14120,N_13523);
nand U18018 (N_18018,N_14971,N_11091);
nor U18019 (N_18019,N_13531,N_14536);
nand U18020 (N_18020,N_13573,N_11969);
xnor U18021 (N_18021,N_13689,N_12762);
xor U18022 (N_18022,N_14508,N_14632);
and U18023 (N_18023,N_13342,N_14014);
nor U18024 (N_18024,N_13139,N_14526);
nor U18025 (N_18025,N_14912,N_14084);
or U18026 (N_18026,N_11510,N_10492);
xor U18027 (N_18027,N_13661,N_14498);
or U18028 (N_18028,N_11239,N_12825);
nand U18029 (N_18029,N_12651,N_13314);
nor U18030 (N_18030,N_14597,N_13756);
and U18031 (N_18031,N_10667,N_10084);
or U18032 (N_18032,N_13870,N_13200);
xor U18033 (N_18033,N_12426,N_13109);
xor U18034 (N_18034,N_10145,N_12428);
and U18035 (N_18035,N_12680,N_11723);
or U18036 (N_18036,N_11890,N_12652);
xor U18037 (N_18037,N_13974,N_13261);
and U18038 (N_18038,N_14379,N_13439);
nand U18039 (N_18039,N_13731,N_12153);
and U18040 (N_18040,N_11240,N_11262);
or U18041 (N_18041,N_10722,N_11987);
nor U18042 (N_18042,N_14876,N_13702);
xor U18043 (N_18043,N_10894,N_13141);
nand U18044 (N_18044,N_10381,N_11178);
nor U18045 (N_18045,N_13008,N_14101);
nand U18046 (N_18046,N_13990,N_13301);
nand U18047 (N_18047,N_12832,N_13414);
nand U18048 (N_18048,N_10419,N_10492);
nor U18049 (N_18049,N_10155,N_14745);
or U18050 (N_18050,N_12566,N_12623);
and U18051 (N_18051,N_14911,N_11296);
or U18052 (N_18052,N_11762,N_11542);
nand U18053 (N_18053,N_13117,N_13441);
nand U18054 (N_18054,N_13902,N_11055);
and U18055 (N_18055,N_11706,N_11484);
nor U18056 (N_18056,N_10859,N_13769);
nor U18057 (N_18057,N_14675,N_10842);
nand U18058 (N_18058,N_12600,N_14982);
or U18059 (N_18059,N_12222,N_10155);
nor U18060 (N_18060,N_11465,N_11255);
or U18061 (N_18061,N_10998,N_14768);
or U18062 (N_18062,N_13443,N_11926);
and U18063 (N_18063,N_12396,N_10057);
nor U18064 (N_18064,N_12396,N_11449);
nand U18065 (N_18065,N_12275,N_10265);
or U18066 (N_18066,N_11936,N_14617);
nor U18067 (N_18067,N_13794,N_13910);
or U18068 (N_18068,N_10646,N_13618);
nand U18069 (N_18069,N_14174,N_13132);
xor U18070 (N_18070,N_14004,N_11344);
or U18071 (N_18071,N_11117,N_14130);
nor U18072 (N_18072,N_11842,N_12515);
and U18073 (N_18073,N_14103,N_12375);
and U18074 (N_18074,N_13554,N_14864);
or U18075 (N_18075,N_14008,N_13810);
nor U18076 (N_18076,N_13058,N_10187);
nand U18077 (N_18077,N_13143,N_13374);
and U18078 (N_18078,N_12569,N_12031);
nand U18079 (N_18079,N_10926,N_10229);
xnor U18080 (N_18080,N_14181,N_12879);
and U18081 (N_18081,N_13638,N_14638);
and U18082 (N_18082,N_11246,N_13319);
xnor U18083 (N_18083,N_14644,N_12963);
xnor U18084 (N_18084,N_11540,N_12326);
and U18085 (N_18085,N_13878,N_10588);
nor U18086 (N_18086,N_10972,N_14703);
and U18087 (N_18087,N_12559,N_12589);
nand U18088 (N_18088,N_14459,N_11561);
xor U18089 (N_18089,N_12930,N_10166);
nand U18090 (N_18090,N_12038,N_13162);
nand U18091 (N_18091,N_13738,N_11786);
or U18092 (N_18092,N_11931,N_12137);
and U18093 (N_18093,N_14555,N_11411);
nand U18094 (N_18094,N_13187,N_13610);
nor U18095 (N_18095,N_11942,N_14277);
nor U18096 (N_18096,N_12730,N_10582);
nor U18097 (N_18097,N_14036,N_13451);
or U18098 (N_18098,N_12038,N_13457);
and U18099 (N_18099,N_10325,N_14388);
xor U18100 (N_18100,N_13717,N_12545);
nand U18101 (N_18101,N_10078,N_11045);
nand U18102 (N_18102,N_11119,N_12526);
and U18103 (N_18103,N_12310,N_12237);
or U18104 (N_18104,N_10927,N_12725);
xnor U18105 (N_18105,N_13311,N_12408);
nor U18106 (N_18106,N_13138,N_10470);
xnor U18107 (N_18107,N_13977,N_11374);
xor U18108 (N_18108,N_10103,N_11535);
and U18109 (N_18109,N_13812,N_13665);
nor U18110 (N_18110,N_14848,N_14819);
nor U18111 (N_18111,N_14007,N_14690);
nand U18112 (N_18112,N_12144,N_11258);
xnor U18113 (N_18113,N_13038,N_10995);
and U18114 (N_18114,N_13813,N_11081);
nand U18115 (N_18115,N_11530,N_12751);
xor U18116 (N_18116,N_12548,N_14812);
or U18117 (N_18117,N_12293,N_13846);
xor U18118 (N_18118,N_12209,N_12965);
nor U18119 (N_18119,N_10767,N_14668);
and U18120 (N_18120,N_11848,N_12957);
and U18121 (N_18121,N_11911,N_11245);
nor U18122 (N_18122,N_12542,N_14840);
or U18123 (N_18123,N_12563,N_11216);
nor U18124 (N_18124,N_12208,N_13528);
nand U18125 (N_18125,N_14475,N_14301);
and U18126 (N_18126,N_11970,N_10500);
nor U18127 (N_18127,N_10859,N_12530);
xor U18128 (N_18128,N_11200,N_11704);
nor U18129 (N_18129,N_14212,N_11469);
or U18130 (N_18130,N_14192,N_12477);
nand U18131 (N_18131,N_11429,N_13462);
xnor U18132 (N_18132,N_14646,N_13346);
or U18133 (N_18133,N_12445,N_10944);
and U18134 (N_18134,N_12368,N_13685);
or U18135 (N_18135,N_12746,N_13541);
or U18136 (N_18136,N_13848,N_14635);
xnor U18137 (N_18137,N_14243,N_14785);
nor U18138 (N_18138,N_11577,N_11791);
nor U18139 (N_18139,N_10391,N_12352);
or U18140 (N_18140,N_11856,N_11636);
and U18141 (N_18141,N_13097,N_14352);
xor U18142 (N_18142,N_11144,N_14176);
xnor U18143 (N_18143,N_11418,N_12458);
nand U18144 (N_18144,N_14926,N_13089);
and U18145 (N_18145,N_12454,N_14967);
or U18146 (N_18146,N_11244,N_10965);
or U18147 (N_18147,N_11957,N_14479);
and U18148 (N_18148,N_13617,N_13474);
or U18149 (N_18149,N_14868,N_14131);
xor U18150 (N_18150,N_10355,N_12536);
and U18151 (N_18151,N_10183,N_11725);
or U18152 (N_18152,N_12901,N_10834);
or U18153 (N_18153,N_10417,N_10802);
nor U18154 (N_18154,N_11153,N_12539);
nor U18155 (N_18155,N_13013,N_14921);
and U18156 (N_18156,N_13104,N_10737);
and U18157 (N_18157,N_13572,N_14527);
or U18158 (N_18158,N_12496,N_13419);
nand U18159 (N_18159,N_11598,N_13968);
or U18160 (N_18160,N_12090,N_12486);
xor U18161 (N_18161,N_11833,N_12784);
xor U18162 (N_18162,N_13625,N_13424);
xor U18163 (N_18163,N_12274,N_11071);
and U18164 (N_18164,N_10662,N_12341);
nor U18165 (N_18165,N_12905,N_13453);
or U18166 (N_18166,N_12915,N_11602);
nand U18167 (N_18167,N_13087,N_12404);
xnor U18168 (N_18168,N_11539,N_11320);
xnor U18169 (N_18169,N_14719,N_14508);
or U18170 (N_18170,N_14540,N_13012);
and U18171 (N_18171,N_13103,N_11725);
or U18172 (N_18172,N_10450,N_12565);
or U18173 (N_18173,N_14395,N_12625);
nor U18174 (N_18174,N_12821,N_11687);
nand U18175 (N_18175,N_10329,N_12576);
nor U18176 (N_18176,N_11584,N_10296);
nand U18177 (N_18177,N_10179,N_14478);
nor U18178 (N_18178,N_11661,N_10088);
nand U18179 (N_18179,N_14061,N_11010);
or U18180 (N_18180,N_12898,N_11343);
and U18181 (N_18181,N_13792,N_12491);
nand U18182 (N_18182,N_14039,N_14257);
or U18183 (N_18183,N_12399,N_11072);
nor U18184 (N_18184,N_10524,N_14619);
nand U18185 (N_18185,N_13938,N_14525);
or U18186 (N_18186,N_10342,N_10850);
nand U18187 (N_18187,N_10154,N_11004);
nor U18188 (N_18188,N_10179,N_13100);
nor U18189 (N_18189,N_14088,N_11293);
xnor U18190 (N_18190,N_13476,N_10659);
and U18191 (N_18191,N_12712,N_13380);
or U18192 (N_18192,N_11850,N_10362);
nor U18193 (N_18193,N_12577,N_11050);
nor U18194 (N_18194,N_11976,N_12144);
nor U18195 (N_18195,N_13170,N_12432);
or U18196 (N_18196,N_12487,N_11905);
nand U18197 (N_18197,N_12541,N_14517);
nand U18198 (N_18198,N_10305,N_13601);
xnor U18199 (N_18199,N_12493,N_10066);
or U18200 (N_18200,N_12626,N_13029);
xor U18201 (N_18201,N_12062,N_13135);
nor U18202 (N_18202,N_11739,N_14988);
xnor U18203 (N_18203,N_12677,N_12211);
xnor U18204 (N_18204,N_12216,N_11273);
nor U18205 (N_18205,N_14004,N_12986);
nor U18206 (N_18206,N_11195,N_13507);
nand U18207 (N_18207,N_12335,N_10597);
or U18208 (N_18208,N_13951,N_13004);
xor U18209 (N_18209,N_13327,N_12484);
nand U18210 (N_18210,N_11254,N_14591);
or U18211 (N_18211,N_11649,N_14954);
nor U18212 (N_18212,N_11240,N_14459);
nor U18213 (N_18213,N_14038,N_10930);
nand U18214 (N_18214,N_13102,N_12741);
xor U18215 (N_18215,N_10173,N_10103);
xor U18216 (N_18216,N_12859,N_13126);
or U18217 (N_18217,N_10399,N_10385);
or U18218 (N_18218,N_10307,N_12540);
nand U18219 (N_18219,N_11164,N_13303);
nand U18220 (N_18220,N_10738,N_14806);
xnor U18221 (N_18221,N_13727,N_14740);
nand U18222 (N_18222,N_10418,N_10025);
or U18223 (N_18223,N_12352,N_11408);
or U18224 (N_18224,N_14235,N_12988);
or U18225 (N_18225,N_14593,N_12016);
nand U18226 (N_18226,N_10793,N_12651);
or U18227 (N_18227,N_14288,N_11506);
nand U18228 (N_18228,N_13728,N_12338);
and U18229 (N_18229,N_14876,N_11125);
nand U18230 (N_18230,N_14649,N_14517);
nand U18231 (N_18231,N_13888,N_10371);
xor U18232 (N_18232,N_13564,N_11040);
xnor U18233 (N_18233,N_11719,N_14558);
xor U18234 (N_18234,N_14709,N_14967);
and U18235 (N_18235,N_13565,N_13603);
xor U18236 (N_18236,N_11598,N_11091);
xor U18237 (N_18237,N_14598,N_13476);
nor U18238 (N_18238,N_11648,N_10183);
nor U18239 (N_18239,N_10633,N_12828);
and U18240 (N_18240,N_12213,N_13968);
and U18241 (N_18241,N_11102,N_13526);
nor U18242 (N_18242,N_13197,N_14069);
and U18243 (N_18243,N_12417,N_13923);
or U18244 (N_18244,N_12552,N_13914);
and U18245 (N_18245,N_14330,N_11953);
nand U18246 (N_18246,N_11593,N_12164);
or U18247 (N_18247,N_12857,N_10268);
nand U18248 (N_18248,N_14690,N_14516);
or U18249 (N_18249,N_14776,N_10009);
nand U18250 (N_18250,N_13606,N_11112);
nor U18251 (N_18251,N_13040,N_11044);
nor U18252 (N_18252,N_12373,N_12214);
nand U18253 (N_18253,N_13879,N_11550);
nand U18254 (N_18254,N_12575,N_14672);
nand U18255 (N_18255,N_13499,N_10849);
nor U18256 (N_18256,N_13253,N_13098);
nand U18257 (N_18257,N_10454,N_13563);
and U18258 (N_18258,N_10962,N_14064);
and U18259 (N_18259,N_11689,N_10195);
nand U18260 (N_18260,N_11868,N_13559);
and U18261 (N_18261,N_10015,N_10793);
nor U18262 (N_18262,N_14196,N_12198);
or U18263 (N_18263,N_10468,N_12594);
or U18264 (N_18264,N_13687,N_10652);
xor U18265 (N_18265,N_11810,N_11932);
and U18266 (N_18266,N_12430,N_11580);
nand U18267 (N_18267,N_11218,N_10988);
xor U18268 (N_18268,N_10819,N_11274);
and U18269 (N_18269,N_13502,N_14600);
or U18270 (N_18270,N_11058,N_11040);
nand U18271 (N_18271,N_12844,N_11248);
or U18272 (N_18272,N_14172,N_12674);
xor U18273 (N_18273,N_13288,N_11435);
xor U18274 (N_18274,N_13849,N_13312);
and U18275 (N_18275,N_13935,N_10976);
xor U18276 (N_18276,N_14430,N_13199);
or U18277 (N_18277,N_13573,N_10022);
and U18278 (N_18278,N_11800,N_14945);
xor U18279 (N_18279,N_12047,N_12864);
and U18280 (N_18280,N_11428,N_11261);
or U18281 (N_18281,N_12897,N_10263);
nor U18282 (N_18282,N_11343,N_14914);
nand U18283 (N_18283,N_10600,N_12444);
and U18284 (N_18284,N_10949,N_14043);
nor U18285 (N_18285,N_14453,N_13183);
xor U18286 (N_18286,N_13476,N_12583);
nand U18287 (N_18287,N_12740,N_13571);
or U18288 (N_18288,N_10060,N_10019);
xnor U18289 (N_18289,N_13764,N_14249);
nand U18290 (N_18290,N_13011,N_14863);
and U18291 (N_18291,N_11418,N_14510);
nand U18292 (N_18292,N_13882,N_10587);
and U18293 (N_18293,N_10368,N_10094);
xnor U18294 (N_18294,N_10399,N_11844);
xnor U18295 (N_18295,N_10240,N_13930);
xnor U18296 (N_18296,N_14503,N_14955);
and U18297 (N_18297,N_12295,N_13219);
or U18298 (N_18298,N_13393,N_14120);
nand U18299 (N_18299,N_14742,N_10995);
xor U18300 (N_18300,N_10168,N_10851);
nor U18301 (N_18301,N_10333,N_10984);
and U18302 (N_18302,N_10601,N_10188);
nor U18303 (N_18303,N_12493,N_11943);
and U18304 (N_18304,N_10948,N_14084);
nand U18305 (N_18305,N_10120,N_10773);
xor U18306 (N_18306,N_13184,N_11600);
xnor U18307 (N_18307,N_11013,N_12592);
nand U18308 (N_18308,N_12129,N_13383);
nand U18309 (N_18309,N_12298,N_10127);
nand U18310 (N_18310,N_13833,N_12278);
xor U18311 (N_18311,N_14393,N_11562);
nor U18312 (N_18312,N_13886,N_13720);
or U18313 (N_18313,N_11107,N_12595);
or U18314 (N_18314,N_13685,N_13682);
and U18315 (N_18315,N_11492,N_13836);
nor U18316 (N_18316,N_13768,N_10018);
xnor U18317 (N_18317,N_14974,N_14657);
and U18318 (N_18318,N_10796,N_11542);
or U18319 (N_18319,N_13852,N_12613);
nor U18320 (N_18320,N_11996,N_11094);
xor U18321 (N_18321,N_14972,N_12243);
nand U18322 (N_18322,N_14486,N_10176);
or U18323 (N_18323,N_14701,N_11337);
or U18324 (N_18324,N_12154,N_10469);
xor U18325 (N_18325,N_12503,N_12689);
nand U18326 (N_18326,N_14943,N_13884);
nand U18327 (N_18327,N_10954,N_12624);
xor U18328 (N_18328,N_10276,N_12096);
or U18329 (N_18329,N_10838,N_14922);
and U18330 (N_18330,N_10888,N_11105);
xnor U18331 (N_18331,N_12235,N_13846);
nor U18332 (N_18332,N_10811,N_13299);
nor U18333 (N_18333,N_10358,N_10781);
or U18334 (N_18334,N_10234,N_11564);
nor U18335 (N_18335,N_12185,N_14292);
xor U18336 (N_18336,N_14021,N_10825);
nand U18337 (N_18337,N_13577,N_14716);
and U18338 (N_18338,N_13831,N_13828);
or U18339 (N_18339,N_11043,N_11822);
and U18340 (N_18340,N_11435,N_13947);
nor U18341 (N_18341,N_12150,N_12310);
and U18342 (N_18342,N_12488,N_13752);
and U18343 (N_18343,N_14710,N_14694);
nor U18344 (N_18344,N_11600,N_11491);
nand U18345 (N_18345,N_13402,N_13804);
xor U18346 (N_18346,N_10348,N_10155);
xor U18347 (N_18347,N_14137,N_14792);
nand U18348 (N_18348,N_11307,N_10298);
or U18349 (N_18349,N_13291,N_13713);
nor U18350 (N_18350,N_12429,N_11722);
xor U18351 (N_18351,N_12253,N_12623);
nand U18352 (N_18352,N_14292,N_10317);
and U18353 (N_18353,N_10260,N_13435);
nor U18354 (N_18354,N_14993,N_10645);
and U18355 (N_18355,N_14954,N_14187);
xor U18356 (N_18356,N_10679,N_14321);
or U18357 (N_18357,N_10865,N_11379);
or U18358 (N_18358,N_11350,N_10754);
nor U18359 (N_18359,N_13588,N_10333);
and U18360 (N_18360,N_12234,N_13051);
or U18361 (N_18361,N_13824,N_10650);
nand U18362 (N_18362,N_14511,N_11070);
nand U18363 (N_18363,N_11495,N_10518);
or U18364 (N_18364,N_10413,N_13628);
and U18365 (N_18365,N_12675,N_10943);
or U18366 (N_18366,N_14808,N_10869);
nor U18367 (N_18367,N_14673,N_13104);
or U18368 (N_18368,N_10535,N_13392);
xor U18369 (N_18369,N_10698,N_14302);
nand U18370 (N_18370,N_13130,N_12029);
xor U18371 (N_18371,N_14587,N_14517);
or U18372 (N_18372,N_13912,N_14211);
or U18373 (N_18373,N_10964,N_13432);
nor U18374 (N_18374,N_12964,N_10220);
xnor U18375 (N_18375,N_11668,N_12802);
nand U18376 (N_18376,N_11588,N_11004);
nor U18377 (N_18377,N_14610,N_14040);
xnor U18378 (N_18378,N_11848,N_13905);
nor U18379 (N_18379,N_13917,N_13528);
and U18380 (N_18380,N_10716,N_14726);
xor U18381 (N_18381,N_12512,N_13287);
nand U18382 (N_18382,N_12668,N_10149);
nand U18383 (N_18383,N_11174,N_14049);
nor U18384 (N_18384,N_10984,N_12701);
xor U18385 (N_18385,N_10611,N_14568);
xor U18386 (N_18386,N_10273,N_13869);
or U18387 (N_18387,N_14751,N_13071);
and U18388 (N_18388,N_14775,N_10567);
xnor U18389 (N_18389,N_12583,N_13696);
and U18390 (N_18390,N_13358,N_10417);
or U18391 (N_18391,N_13690,N_14840);
xnor U18392 (N_18392,N_11592,N_11157);
xor U18393 (N_18393,N_12538,N_12497);
and U18394 (N_18394,N_10477,N_13295);
nor U18395 (N_18395,N_13459,N_10003);
and U18396 (N_18396,N_11752,N_13868);
or U18397 (N_18397,N_14391,N_14303);
and U18398 (N_18398,N_10402,N_11417);
nor U18399 (N_18399,N_11496,N_10890);
nor U18400 (N_18400,N_13078,N_14617);
xnor U18401 (N_18401,N_14457,N_13828);
nand U18402 (N_18402,N_13077,N_11887);
or U18403 (N_18403,N_12652,N_13229);
or U18404 (N_18404,N_11158,N_13271);
xor U18405 (N_18405,N_11516,N_10436);
xor U18406 (N_18406,N_11130,N_14582);
and U18407 (N_18407,N_13044,N_11841);
xor U18408 (N_18408,N_12451,N_13686);
or U18409 (N_18409,N_13930,N_11348);
nand U18410 (N_18410,N_10813,N_10630);
nor U18411 (N_18411,N_11999,N_11274);
or U18412 (N_18412,N_13344,N_12171);
nand U18413 (N_18413,N_14027,N_14341);
nand U18414 (N_18414,N_12011,N_11685);
nor U18415 (N_18415,N_12591,N_12108);
and U18416 (N_18416,N_10938,N_13167);
nor U18417 (N_18417,N_11008,N_11330);
xor U18418 (N_18418,N_14715,N_11343);
and U18419 (N_18419,N_10156,N_12352);
or U18420 (N_18420,N_13818,N_14412);
or U18421 (N_18421,N_13489,N_13595);
xnor U18422 (N_18422,N_11094,N_13546);
and U18423 (N_18423,N_10594,N_10336);
nand U18424 (N_18424,N_11946,N_12152);
and U18425 (N_18425,N_11090,N_11794);
or U18426 (N_18426,N_10369,N_12966);
nand U18427 (N_18427,N_10988,N_14360);
xor U18428 (N_18428,N_13359,N_10214);
and U18429 (N_18429,N_12042,N_11358);
nor U18430 (N_18430,N_13902,N_11343);
xor U18431 (N_18431,N_11947,N_13163);
and U18432 (N_18432,N_11739,N_14304);
nor U18433 (N_18433,N_10831,N_13709);
xor U18434 (N_18434,N_13952,N_14044);
xor U18435 (N_18435,N_12699,N_11377);
nand U18436 (N_18436,N_13629,N_10877);
nor U18437 (N_18437,N_12395,N_13987);
nand U18438 (N_18438,N_11838,N_11426);
and U18439 (N_18439,N_11000,N_10768);
xnor U18440 (N_18440,N_13346,N_12687);
nand U18441 (N_18441,N_13946,N_12342);
and U18442 (N_18442,N_12173,N_10576);
xnor U18443 (N_18443,N_12832,N_13847);
or U18444 (N_18444,N_13284,N_11530);
or U18445 (N_18445,N_12886,N_10240);
or U18446 (N_18446,N_10368,N_14830);
nor U18447 (N_18447,N_10014,N_13924);
or U18448 (N_18448,N_10519,N_11807);
nor U18449 (N_18449,N_12198,N_12985);
xor U18450 (N_18450,N_11203,N_12907);
or U18451 (N_18451,N_11924,N_10158);
nand U18452 (N_18452,N_12071,N_12040);
xnor U18453 (N_18453,N_10169,N_10306);
nand U18454 (N_18454,N_13462,N_12608);
nand U18455 (N_18455,N_13563,N_13142);
nand U18456 (N_18456,N_14734,N_14794);
nand U18457 (N_18457,N_14769,N_12932);
nor U18458 (N_18458,N_14469,N_10493);
and U18459 (N_18459,N_13510,N_10364);
and U18460 (N_18460,N_13311,N_12377);
nand U18461 (N_18461,N_10094,N_10633);
xor U18462 (N_18462,N_14714,N_10045);
and U18463 (N_18463,N_12694,N_11623);
or U18464 (N_18464,N_12296,N_12303);
or U18465 (N_18465,N_12138,N_14073);
or U18466 (N_18466,N_10752,N_11302);
xnor U18467 (N_18467,N_13108,N_11615);
nand U18468 (N_18468,N_12109,N_14039);
and U18469 (N_18469,N_11230,N_12452);
nand U18470 (N_18470,N_10282,N_14019);
and U18471 (N_18471,N_11277,N_13645);
xnor U18472 (N_18472,N_13778,N_11290);
nand U18473 (N_18473,N_10375,N_10242);
and U18474 (N_18474,N_14322,N_14059);
nand U18475 (N_18475,N_10882,N_14870);
xor U18476 (N_18476,N_12907,N_11008);
nor U18477 (N_18477,N_12187,N_12270);
or U18478 (N_18478,N_13475,N_11205);
nand U18479 (N_18479,N_13117,N_11890);
or U18480 (N_18480,N_12677,N_14896);
xnor U18481 (N_18481,N_14752,N_12756);
and U18482 (N_18482,N_10869,N_11799);
or U18483 (N_18483,N_11784,N_12658);
or U18484 (N_18484,N_14448,N_13235);
nor U18485 (N_18485,N_11968,N_11911);
nor U18486 (N_18486,N_12205,N_13165);
and U18487 (N_18487,N_11966,N_10521);
nor U18488 (N_18488,N_12739,N_13950);
nand U18489 (N_18489,N_11566,N_12528);
nand U18490 (N_18490,N_14232,N_11145);
and U18491 (N_18491,N_11813,N_12380);
and U18492 (N_18492,N_12001,N_12437);
nand U18493 (N_18493,N_11296,N_13371);
or U18494 (N_18494,N_12552,N_12296);
nand U18495 (N_18495,N_13987,N_11951);
nor U18496 (N_18496,N_14076,N_12604);
or U18497 (N_18497,N_10474,N_12263);
and U18498 (N_18498,N_12373,N_13613);
and U18499 (N_18499,N_10755,N_13870);
nor U18500 (N_18500,N_13600,N_14478);
nand U18501 (N_18501,N_11856,N_10434);
or U18502 (N_18502,N_10065,N_14972);
xor U18503 (N_18503,N_13833,N_10810);
nor U18504 (N_18504,N_14118,N_11422);
or U18505 (N_18505,N_14875,N_11088);
or U18506 (N_18506,N_13460,N_12668);
xor U18507 (N_18507,N_13537,N_12379);
nand U18508 (N_18508,N_13188,N_11789);
xor U18509 (N_18509,N_14052,N_14744);
or U18510 (N_18510,N_13551,N_12813);
nand U18511 (N_18511,N_10747,N_10245);
and U18512 (N_18512,N_10643,N_13769);
nor U18513 (N_18513,N_10746,N_12871);
or U18514 (N_18514,N_12315,N_11460);
xnor U18515 (N_18515,N_13822,N_10249);
nand U18516 (N_18516,N_14638,N_14381);
and U18517 (N_18517,N_11903,N_12230);
nand U18518 (N_18518,N_12004,N_12450);
or U18519 (N_18519,N_11286,N_12882);
xor U18520 (N_18520,N_14937,N_13188);
nor U18521 (N_18521,N_10464,N_13131);
or U18522 (N_18522,N_10085,N_10690);
nand U18523 (N_18523,N_14384,N_11589);
and U18524 (N_18524,N_14159,N_13501);
xor U18525 (N_18525,N_12999,N_11809);
and U18526 (N_18526,N_10972,N_11087);
nand U18527 (N_18527,N_13086,N_10045);
or U18528 (N_18528,N_14238,N_12688);
nand U18529 (N_18529,N_13162,N_14096);
xor U18530 (N_18530,N_10366,N_14354);
and U18531 (N_18531,N_13138,N_12500);
nand U18532 (N_18532,N_14201,N_14271);
nor U18533 (N_18533,N_13261,N_11207);
and U18534 (N_18534,N_14594,N_10673);
nand U18535 (N_18535,N_14487,N_13696);
nor U18536 (N_18536,N_12053,N_12937);
nor U18537 (N_18537,N_10866,N_10445);
or U18538 (N_18538,N_11745,N_13091);
nor U18539 (N_18539,N_11165,N_13664);
and U18540 (N_18540,N_12415,N_10250);
and U18541 (N_18541,N_11198,N_12879);
or U18542 (N_18542,N_13234,N_13342);
xor U18543 (N_18543,N_12881,N_13731);
or U18544 (N_18544,N_12315,N_10826);
xnor U18545 (N_18545,N_13787,N_13986);
nor U18546 (N_18546,N_10767,N_13971);
or U18547 (N_18547,N_11749,N_12959);
or U18548 (N_18548,N_11036,N_14874);
nor U18549 (N_18549,N_11622,N_13666);
nand U18550 (N_18550,N_13760,N_10870);
nor U18551 (N_18551,N_11603,N_14591);
nand U18552 (N_18552,N_13638,N_10688);
and U18553 (N_18553,N_12825,N_12018);
or U18554 (N_18554,N_10342,N_11305);
nand U18555 (N_18555,N_12478,N_12356);
nand U18556 (N_18556,N_14415,N_13144);
nand U18557 (N_18557,N_11606,N_12673);
or U18558 (N_18558,N_12989,N_13779);
nor U18559 (N_18559,N_11702,N_12832);
and U18560 (N_18560,N_13249,N_14961);
nor U18561 (N_18561,N_14250,N_10658);
and U18562 (N_18562,N_10095,N_10345);
or U18563 (N_18563,N_11367,N_10187);
nand U18564 (N_18564,N_13149,N_13026);
xnor U18565 (N_18565,N_11907,N_13505);
nand U18566 (N_18566,N_11659,N_14686);
and U18567 (N_18567,N_11022,N_10181);
nand U18568 (N_18568,N_11939,N_13410);
xor U18569 (N_18569,N_13054,N_13192);
nor U18570 (N_18570,N_12407,N_13634);
and U18571 (N_18571,N_10785,N_13003);
xor U18572 (N_18572,N_10549,N_12563);
or U18573 (N_18573,N_10390,N_10919);
and U18574 (N_18574,N_12619,N_11583);
and U18575 (N_18575,N_14628,N_13560);
or U18576 (N_18576,N_12541,N_10204);
xor U18577 (N_18577,N_13240,N_14473);
and U18578 (N_18578,N_13875,N_11236);
and U18579 (N_18579,N_12013,N_12161);
or U18580 (N_18580,N_12787,N_12332);
nor U18581 (N_18581,N_11650,N_11977);
or U18582 (N_18582,N_13343,N_14547);
or U18583 (N_18583,N_12792,N_13311);
or U18584 (N_18584,N_13818,N_13999);
nor U18585 (N_18585,N_11639,N_14226);
and U18586 (N_18586,N_12839,N_14466);
nor U18587 (N_18587,N_14082,N_12743);
xnor U18588 (N_18588,N_10170,N_14480);
nor U18589 (N_18589,N_13319,N_14338);
xor U18590 (N_18590,N_13136,N_10245);
xor U18591 (N_18591,N_10771,N_13997);
nand U18592 (N_18592,N_13252,N_13346);
and U18593 (N_18593,N_14062,N_10489);
nor U18594 (N_18594,N_13566,N_13862);
and U18595 (N_18595,N_11147,N_12977);
nand U18596 (N_18596,N_14537,N_10761);
and U18597 (N_18597,N_14847,N_14486);
and U18598 (N_18598,N_14807,N_14471);
xnor U18599 (N_18599,N_12794,N_12350);
and U18600 (N_18600,N_10066,N_12760);
and U18601 (N_18601,N_11417,N_14656);
and U18602 (N_18602,N_13571,N_12661);
xnor U18603 (N_18603,N_14756,N_13402);
nor U18604 (N_18604,N_12294,N_14143);
nor U18605 (N_18605,N_11261,N_14696);
or U18606 (N_18606,N_13427,N_11991);
nand U18607 (N_18607,N_14178,N_12667);
or U18608 (N_18608,N_11745,N_14480);
nand U18609 (N_18609,N_13263,N_12815);
nand U18610 (N_18610,N_12749,N_13658);
nor U18611 (N_18611,N_12134,N_14590);
and U18612 (N_18612,N_10111,N_13816);
or U18613 (N_18613,N_10394,N_12155);
xnor U18614 (N_18614,N_13579,N_12600);
nand U18615 (N_18615,N_11641,N_14005);
or U18616 (N_18616,N_12845,N_14283);
xor U18617 (N_18617,N_11787,N_10467);
or U18618 (N_18618,N_10250,N_10783);
and U18619 (N_18619,N_11457,N_13544);
and U18620 (N_18620,N_13652,N_14860);
or U18621 (N_18621,N_10018,N_11288);
xnor U18622 (N_18622,N_11259,N_14948);
nor U18623 (N_18623,N_13610,N_10770);
and U18624 (N_18624,N_11022,N_10822);
and U18625 (N_18625,N_11840,N_14384);
nor U18626 (N_18626,N_11577,N_11755);
xor U18627 (N_18627,N_14691,N_10909);
nor U18628 (N_18628,N_11571,N_13544);
nand U18629 (N_18629,N_10442,N_11908);
and U18630 (N_18630,N_10144,N_10062);
and U18631 (N_18631,N_14224,N_11380);
nor U18632 (N_18632,N_14611,N_12792);
nor U18633 (N_18633,N_14377,N_12377);
or U18634 (N_18634,N_11607,N_14765);
or U18635 (N_18635,N_13180,N_10519);
nand U18636 (N_18636,N_11241,N_14565);
xnor U18637 (N_18637,N_13599,N_14382);
nor U18638 (N_18638,N_11844,N_12412);
and U18639 (N_18639,N_14517,N_14732);
or U18640 (N_18640,N_10050,N_10301);
nand U18641 (N_18641,N_11947,N_11174);
and U18642 (N_18642,N_12027,N_10835);
xor U18643 (N_18643,N_10193,N_13975);
xnor U18644 (N_18644,N_11359,N_13791);
or U18645 (N_18645,N_10343,N_10648);
xor U18646 (N_18646,N_13100,N_14458);
xnor U18647 (N_18647,N_13827,N_14124);
xor U18648 (N_18648,N_14380,N_14926);
and U18649 (N_18649,N_14244,N_12378);
xor U18650 (N_18650,N_10922,N_14670);
and U18651 (N_18651,N_12070,N_10351);
and U18652 (N_18652,N_12950,N_14432);
xor U18653 (N_18653,N_14855,N_10005);
nand U18654 (N_18654,N_12091,N_13096);
nand U18655 (N_18655,N_10917,N_13328);
or U18656 (N_18656,N_11759,N_10756);
or U18657 (N_18657,N_10875,N_13264);
xnor U18658 (N_18658,N_13766,N_12094);
or U18659 (N_18659,N_10497,N_14306);
nand U18660 (N_18660,N_10655,N_13868);
nand U18661 (N_18661,N_12664,N_10078);
or U18662 (N_18662,N_11516,N_14980);
xor U18663 (N_18663,N_10795,N_13511);
and U18664 (N_18664,N_13080,N_10401);
or U18665 (N_18665,N_13873,N_11527);
nor U18666 (N_18666,N_10281,N_14590);
nor U18667 (N_18667,N_11398,N_12388);
or U18668 (N_18668,N_11501,N_12874);
xnor U18669 (N_18669,N_12070,N_11718);
xnor U18670 (N_18670,N_14256,N_12541);
nand U18671 (N_18671,N_10535,N_10233);
or U18672 (N_18672,N_12915,N_10017);
nor U18673 (N_18673,N_11310,N_11492);
xnor U18674 (N_18674,N_14980,N_11518);
and U18675 (N_18675,N_12194,N_10117);
xnor U18676 (N_18676,N_12228,N_14666);
nor U18677 (N_18677,N_10615,N_12657);
and U18678 (N_18678,N_10913,N_10862);
nand U18679 (N_18679,N_13192,N_12340);
nand U18680 (N_18680,N_14351,N_11245);
and U18681 (N_18681,N_12298,N_11524);
or U18682 (N_18682,N_14760,N_14682);
xor U18683 (N_18683,N_10017,N_12280);
xor U18684 (N_18684,N_11120,N_13493);
nor U18685 (N_18685,N_10374,N_11689);
xnor U18686 (N_18686,N_14622,N_12642);
or U18687 (N_18687,N_12199,N_14685);
or U18688 (N_18688,N_10095,N_11637);
or U18689 (N_18689,N_10306,N_11380);
and U18690 (N_18690,N_11076,N_10130);
nor U18691 (N_18691,N_13393,N_14785);
and U18692 (N_18692,N_14067,N_10306);
xor U18693 (N_18693,N_11757,N_10563);
xnor U18694 (N_18694,N_11491,N_13829);
nand U18695 (N_18695,N_13562,N_10919);
xnor U18696 (N_18696,N_14654,N_12411);
nand U18697 (N_18697,N_14708,N_10578);
or U18698 (N_18698,N_13176,N_13314);
nor U18699 (N_18699,N_13381,N_13268);
nand U18700 (N_18700,N_14837,N_13128);
nor U18701 (N_18701,N_12555,N_11239);
or U18702 (N_18702,N_10877,N_10174);
nor U18703 (N_18703,N_11055,N_12749);
and U18704 (N_18704,N_10733,N_13232);
nand U18705 (N_18705,N_10039,N_12341);
nand U18706 (N_18706,N_11285,N_10813);
nand U18707 (N_18707,N_11549,N_14019);
xnor U18708 (N_18708,N_13059,N_13543);
nand U18709 (N_18709,N_13448,N_10509);
or U18710 (N_18710,N_11050,N_13940);
xnor U18711 (N_18711,N_12970,N_11835);
xor U18712 (N_18712,N_14530,N_14858);
and U18713 (N_18713,N_11313,N_10558);
and U18714 (N_18714,N_13185,N_10088);
xnor U18715 (N_18715,N_13247,N_11377);
or U18716 (N_18716,N_11309,N_13742);
xor U18717 (N_18717,N_12512,N_11091);
xnor U18718 (N_18718,N_12616,N_14410);
nand U18719 (N_18719,N_14274,N_14719);
nand U18720 (N_18720,N_12807,N_14029);
nand U18721 (N_18721,N_13402,N_10284);
nor U18722 (N_18722,N_11051,N_12929);
or U18723 (N_18723,N_11821,N_11447);
nand U18724 (N_18724,N_14222,N_11564);
and U18725 (N_18725,N_10390,N_11855);
xnor U18726 (N_18726,N_11963,N_11913);
xor U18727 (N_18727,N_10753,N_11418);
nor U18728 (N_18728,N_12921,N_11075);
and U18729 (N_18729,N_11714,N_10568);
or U18730 (N_18730,N_11668,N_14129);
and U18731 (N_18731,N_10335,N_14323);
or U18732 (N_18732,N_11163,N_10638);
and U18733 (N_18733,N_10661,N_11023);
xor U18734 (N_18734,N_14639,N_10283);
xor U18735 (N_18735,N_10362,N_11870);
or U18736 (N_18736,N_11140,N_13251);
nor U18737 (N_18737,N_12666,N_14501);
or U18738 (N_18738,N_10765,N_13399);
xnor U18739 (N_18739,N_12833,N_10811);
xnor U18740 (N_18740,N_12152,N_14713);
nor U18741 (N_18741,N_14892,N_10761);
or U18742 (N_18742,N_10219,N_11000);
nor U18743 (N_18743,N_12397,N_14900);
nand U18744 (N_18744,N_11106,N_10943);
xnor U18745 (N_18745,N_14772,N_14537);
xnor U18746 (N_18746,N_14692,N_11648);
and U18747 (N_18747,N_14824,N_11046);
nand U18748 (N_18748,N_10568,N_13353);
or U18749 (N_18749,N_11874,N_10154);
nand U18750 (N_18750,N_10101,N_14563);
nand U18751 (N_18751,N_10724,N_10840);
nor U18752 (N_18752,N_12493,N_10695);
or U18753 (N_18753,N_10596,N_10339);
xnor U18754 (N_18754,N_13511,N_10084);
nand U18755 (N_18755,N_12325,N_10186);
nand U18756 (N_18756,N_13643,N_11286);
nor U18757 (N_18757,N_14004,N_13517);
nor U18758 (N_18758,N_13542,N_13270);
and U18759 (N_18759,N_11371,N_11001);
nand U18760 (N_18760,N_12440,N_13073);
nand U18761 (N_18761,N_14772,N_10746);
nand U18762 (N_18762,N_12836,N_12507);
nor U18763 (N_18763,N_14134,N_13999);
nand U18764 (N_18764,N_14540,N_11133);
nand U18765 (N_18765,N_14841,N_10464);
xnor U18766 (N_18766,N_12601,N_12720);
nor U18767 (N_18767,N_13848,N_12687);
nand U18768 (N_18768,N_14743,N_11487);
nor U18769 (N_18769,N_12149,N_14253);
and U18770 (N_18770,N_10724,N_12652);
or U18771 (N_18771,N_10021,N_11816);
or U18772 (N_18772,N_11484,N_10299);
or U18773 (N_18773,N_13232,N_10564);
or U18774 (N_18774,N_14498,N_13055);
nand U18775 (N_18775,N_11845,N_10197);
xnor U18776 (N_18776,N_14581,N_11876);
nand U18777 (N_18777,N_12906,N_10908);
nand U18778 (N_18778,N_13648,N_12712);
and U18779 (N_18779,N_11587,N_14201);
nor U18780 (N_18780,N_13613,N_12474);
nand U18781 (N_18781,N_10866,N_11323);
nand U18782 (N_18782,N_12795,N_11900);
or U18783 (N_18783,N_14432,N_11416);
nand U18784 (N_18784,N_13203,N_10766);
nor U18785 (N_18785,N_11840,N_13824);
xnor U18786 (N_18786,N_10539,N_14756);
xnor U18787 (N_18787,N_13979,N_10996);
nor U18788 (N_18788,N_12284,N_10792);
nand U18789 (N_18789,N_13345,N_10880);
or U18790 (N_18790,N_11160,N_12641);
or U18791 (N_18791,N_11845,N_13585);
or U18792 (N_18792,N_12339,N_13530);
xnor U18793 (N_18793,N_12129,N_14506);
xor U18794 (N_18794,N_13852,N_14018);
or U18795 (N_18795,N_10279,N_10196);
or U18796 (N_18796,N_11828,N_14748);
nor U18797 (N_18797,N_11796,N_13906);
xor U18798 (N_18798,N_13513,N_13035);
nand U18799 (N_18799,N_11638,N_10813);
or U18800 (N_18800,N_13131,N_10504);
nor U18801 (N_18801,N_12115,N_12470);
nand U18802 (N_18802,N_13317,N_11250);
nor U18803 (N_18803,N_10336,N_12333);
nand U18804 (N_18804,N_12228,N_12511);
or U18805 (N_18805,N_14462,N_13092);
nand U18806 (N_18806,N_11219,N_12038);
nor U18807 (N_18807,N_12533,N_10494);
nand U18808 (N_18808,N_10279,N_13117);
nor U18809 (N_18809,N_10012,N_13471);
xor U18810 (N_18810,N_13726,N_14182);
nor U18811 (N_18811,N_11676,N_11530);
and U18812 (N_18812,N_11862,N_10534);
and U18813 (N_18813,N_10944,N_14531);
and U18814 (N_18814,N_11110,N_14851);
and U18815 (N_18815,N_13342,N_13835);
or U18816 (N_18816,N_10063,N_11698);
xnor U18817 (N_18817,N_11491,N_11162);
nor U18818 (N_18818,N_13360,N_14826);
or U18819 (N_18819,N_10700,N_11940);
nand U18820 (N_18820,N_14026,N_12625);
or U18821 (N_18821,N_13968,N_13184);
nor U18822 (N_18822,N_14479,N_13256);
nor U18823 (N_18823,N_14156,N_14263);
nor U18824 (N_18824,N_11187,N_12487);
nor U18825 (N_18825,N_14153,N_12334);
nor U18826 (N_18826,N_13803,N_14095);
and U18827 (N_18827,N_13782,N_14628);
xor U18828 (N_18828,N_13038,N_13207);
or U18829 (N_18829,N_12117,N_12635);
nor U18830 (N_18830,N_10903,N_11862);
xor U18831 (N_18831,N_11697,N_11075);
nand U18832 (N_18832,N_13093,N_11421);
and U18833 (N_18833,N_12275,N_12566);
or U18834 (N_18834,N_10644,N_12151);
nand U18835 (N_18835,N_14213,N_13376);
and U18836 (N_18836,N_11870,N_11134);
or U18837 (N_18837,N_14663,N_14350);
or U18838 (N_18838,N_11456,N_10776);
nand U18839 (N_18839,N_11164,N_10124);
or U18840 (N_18840,N_14414,N_12326);
nand U18841 (N_18841,N_11216,N_14789);
xor U18842 (N_18842,N_12364,N_12767);
or U18843 (N_18843,N_12688,N_14347);
and U18844 (N_18844,N_14677,N_14590);
or U18845 (N_18845,N_12078,N_12356);
and U18846 (N_18846,N_14971,N_11172);
nor U18847 (N_18847,N_13306,N_13166);
nand U18848 (N_18848,N_11285,N_12247);
or U18849 (N_18849,N_12422,N_11705);
or U18850 (N_18850,N_10484,N_12549);
nor U18851 (N_18851,N_13437,N_11542);
nor U18852 (N_18852,N_11267,N_14657);
or U18853 (N_18853,N_12240,N_10887);
and U18854 (N_18854,N_13412,N_11197);
nand U18855 (N_18855,N_11825,N_14324);
and U18856 (N_18856,N_10654,N_10333);
and U18857 (N_18857,N_11710,N_10322);
and U18858 (N_18858,N_14524,N_12648);
or U18859 (N_18859,N_12056,N_14346);
nor U18860 (N_18860,N_13844,N_10776);
or U18861 (N_18861,N_13307,N_12347);
xnor U18862 (N_18862,N_13606,N_14722);
nand U18863 (N_18863,N_12454,N_13431);
or U18864 (N_18864,N_11340,N_14587);
or U18865 (N_18865,N_11227,N_12343);
nor U18866 (N_18866,N_10818,N_13145);
nand U18867 (N_18867,N_14036,N_11351);
and U18868 (N_18868,N_11562,N_10676);
nor U18869 (N_18869,N_12822,N_13283);
nor U18870 (N_18870,N_11700,N_12124);
and U18871 (N_18871,N_13529,N_14674);
and U18872 (N_18872,N_12617,N_10510);
xnor U18873 (N_18873,N_11775,N_13410);
nor U18874 (N_18874,N_12918,N_13217);
and U18875 (N_18875,N_11025,N_13144);
and U18876 (N_18876,N_10353,N_13710);
xnor U18877 (N_18877,N_10832,N_13034);
and U18878 (N_18878,N_13710,N_12223);
nor U18879 (N_18879,N_12123,N_10888);
or U18880 (N_18880,N_12408,N_12868);
and U18881 (N_18881,N_10855,N_14064);
or U18882 (N_18882,N_11219,N_11387);
nor U18883 (N_18883,N_13686,N_13381);
and U18884 (N_18884,N_13759,N_11423);
xnor U18885 (N_18885,N_10670,N_12856);
nand U18886 (N_18886,N_13414,N_11232);
xor U18887 (N_18887,N_13880,N_11672);
nor U18888 (N_18888,N_11269,N_13940);
nor U18889 (N_18889,N_11925,N_14299);
nor U18890 (N_18890,N_11877,N_11552);
and U18891 (N_18891,N_10732,N_13286);
nor U18892 (N_18892,N_14909,N_11089);
xor U18893 (N_18893,N_12319,N_13695);
nor U18894 (N_18894,N_10460,N_11314);
nand U18895 (N_18895,N_12556,N_11247);
and U18896 (N_18896,N_11836,N_14596);
and U18897 (N_18897,N_10075,N_10651);
nand U18898 (N_18898,N_11624,N_11390);
and U18899 (N_18899,N_12854,N_12300);
or U18900 (N_18900,N_10400,N_10062);
or U18901 (N_18901,N_10614,N_13118);
and U18902 (N_18902,N_12623,N_14296);
or U18903 (N_18903,N_14655,N_10108);
nand U18904 (N_18904,N_14074,N_13195);
and U18905 (N_18905,N_11148,N_13066);
xnor U18906 (N_18906,N_11154,N_12130);
nand U18907 (N_18907,N_14032,N_11533);
xnor U18908 (N_18908,N_14700,N_13203);
or U18909 (N_18909,N_10555,N_10713);
nand U18910 (N_18910,N_14862,N_12072);
nor U18911 (N_18911,N_14894,N_10890);
or U18912 (N_18912,N_11603,N_10836);
nand U18913 (N_18913,N_10905,N_12665);
or U18914 (N_18914,N_10378,N_11023);
nand U18915 (N_18915,N_11182,N_10867);
or U18916 (N_18916,N_11297,N_14057);
and U18917 (N_18917,N_11008,N_10802);
xor U18918 (N_18918,N_11484,N_12734);
and U18919 (N_18919,N_13628,N_14829);
and U18920 (N_18920,N_13501,N_14137);
xnor U18921 (N_18921,N_13414,N_11591);
xor U18922 (N_18922,N_10110,N_11974);
or U18923 (N_18923,N_10597,N_12248);
and U18924 (N_18924,N_14341,N_12908);
xor U18925 (N_18925,N_14152,N_14445);
nor U18926 (N_18926,N_10305,N_10140);
nor U18927 (N_18927,N_14966,N_13996);
xor U18928 (N_18928,N_10049,N_13316);
or U18929 (N_18929,N_10934,N_13312);
and U18930 (N_18930,N_13156,N_14147);
xor U18931 (N_18931,N_10435,N_13558);
and U18932 (N_18932,N_10008,N_14636);
nand U18933 (N_18933,N_12219,N_10373);
nand U18934 (N_18934,N_13003,N_13189);
nor U18935 (N_18935,N_10942,N_13897);
or U18936 (N_18936,N_14476,N_11524);
nor U18937 (N_18937,N_14149,N_14360);
nor U18938 (N_18938,N_11715,N_10068);
or U18939 (N_18939,N_10671,N_10999);
nor U18940 (N_18940,N_12584,N_13653);
or U18941 (N_18941,N_12351,N_12413);
or U18942 (N_18942,N_10889,N_10674);
xnor U18943 (N_18943,N_11982,N_13284);
nor U18944 (N_18944,N_11529,N_13674);
nor U18945 (N_18945,N_12802,N_10688);
nand U18946 (N_18946,N_14608,N_12616);
and U18947 (N_18947,N_10541,N_13016);
or U18948 (N_18948,N_13757,N_12843);
nand U18949 (N_18949,N_10382,N_13370);
or U18950 (N_18950,N_12568,N_11520);
and U18951 (N_18951,N_12461,N_11748);
nor U18952 (N_18952,N_10271,N_11727);
and U18953 (N_18953,N_10466,N_11782);
nor U18954 (N_18954,N_14720,N_12380);
and U18955 (N_18955,N_10951,N_12080);
xnor U18956 (N_18956,N_11817,N_10727);
nand U18957 (N_18957,N_10752,N_12890);
nand U18958 (N_18958,N_12919,N_10459);
and U18959 (N_18959,N_10726,N_12548);
xnor U18960 (N_18960,N_12419,N_14540);
nand U18961 (N_18961,N_12333,N_11139);
and U18962 (N_18962,N_11613,N_12297);
and U18963 (N_18963,N_11746,N_14115);
nand U18964 (N_18964,N_14751,N_10248);
or U18965 (N_18965,N_10975,N_13019);
nand U18966 (N_18966,N_12041,N_11122);
nand U18967 (N_18967,N_10055,N_11886);
xor U18968 (N_18968,N_14756,N_14831);
nand U18969 (N_18969,N_11843,N_12439);
nor U18970 (N_18970,N_12598,N_14983);
nor U18971 (N_18971,N_13522,N_10544);
or U18972 (N_18972,N_12156,N_13555);
or U18973 (N_18973,N_10328,N_10171);
or U18974 (N_18974,N_14806,N_14731);
or U18975 (N_18975,N_12023,N_12890);
nor U18976 (N_18976,N_14989,N_11944);
nor U18977 (N_18977,N_13592,N_13661);
nand U18978 (N_18978,N_14986,N_11652);
nand U18979 (N_18979,N_14929,N_13196);
and U18980 (N_18980,N_14145,N_13570);
or U18981 (N_18981,N_10814,N_13113);
and U18982 (N_18982,N_12986,N_14270);
nand U18983 (N_18983,N_12090,N_13728);
nand U18984 (N_18984,N_10272,N_13399);
nor U18985 (N_18985,N_14716,N_13799);
or U18986 (N_18986,N_11665,N_12213);
nor U18987 (N_18987,N_11122,N_11243);
and U18988 (N_18988,N_12660,N_10342);
and U18989 (N_18989,N_10206,N_14566);
nor U18990 (N_18990,N_11270,N_12207);
and U18991 (N_18991,N_10056,N_13258);
nand U18992 (N_18992,N_12049,N_12102);
or U18993 (N_18993,N_13809,N_12279);
and U18994 (N_18994,N_14118,N_13692);
or U18995 (N_18995,N_12201,N_12020);
xor U18996 (N_18996,N_11529,N_12015);
xor U18997 (N_18997,N_12154,N_11631);
nor U18998 (N_18998,N_11722,N_11401);
nor U18999 (N_18999,N_10575,N_12283);
xor U19000 (N_19000,N_11922,N_12522);
or U19001 (N_19001,N_14796,N_12045);
or U19002 (N_19002,N_13557,N_10349);
and U19003 (N_19003,N_13635,N_14066);
xor U19004 (N_19004,N_14400,N_14614);
or U19005 (N_19005,N_12280,N_11307);
nor U19006 (N_19006,N_13018,N_10829);
nand U19007 (N_19007,N_13393,N_12981);
nand U19008 (N_19008,N_13826,N_13297);
and U19009 (N_19009,N_14587,N_14156);
nand U19010 (N_19010,N_11962,N_10559);
or U19011 (N_19011,N_13110,N_12399);
nor U19012 (N_19012,N_13219,N_13913);
nor U19013 (N_19013,N_13551,N_12616);
xor U19014 (N_19014,N_10340,N_14333);
xor U19015 (N_19015,N_10993,N_14869);
and U19016 (N_19016,N_14550,N_12665);
and U19017 (N_19017,N_12217,N_10230);
nor U19018 (N_19018,N_13868,N_14032);
nor U19019 (N_19019,N_11167,N_13662);
nand U19020 (N_19020,N_13126,N_13529);
or U19021 (N_19021,N_14952,N_13949);
nor U19022 (N_19022,N_14849,N_11502);
xor U19023 (N_19023,N_10143,N_14778);
xor U19024 (N_19024,N_13913,N_13587);
nor U19025 (N_19025,N_12239,N_13037);
or U19026 (N_19026,N_14804,N_14778);
xor U19027 (N_19027,N_12855,N_14406);
xnor U19028 (N_19028,N_14124,N_10511);
and U19029 (N_19029,N_13752,N_12684);
xnor U19030 (N_19030,N_12855,N_12142);
and U19031 (N_19031,N_12077,N_14854);
and U19032 (N_19032,N_13956,N_10908);
and U19033 (N_19033,N_12920,N_13198);
xor U19034 (N_19034,N_10467,N_12972);
and U19035 (N_19035,N_14527,N_11341);
xnor U19036 (N_19036,N_13249,N_13110);
or U19037 (N_19037,N_14981,N_10730);
and U19038 (N_19038,N_14734,N_12889);
xnor U19039 (N_19039,N_12385,N_12011);
and U19040 (N_19040,N_13422,N_10344);
nor U19041 (N_19041,N_14721,N_14847);
nand U19042 (N_19042,N_11029,N_14794);
nand U19043 (N_19043,N_13435,N_13844);
and U19044 (N_19044,N_14891,N_12008);
or U19045 (N_19045,N_13815,N_11982);
xnor U19046 (N_19046,N_12006,N_11601);
or U19047 (N_19047,N_13877,N_11861);
xnor U19048 (N_19048,N_14901,N_12894);
nor U19049 (N_19049,N_13837,N_10735);
nor U19050 (N_19050,N_10659,N_13400);
xnor U19051 (N_19051,N_13319,N_13257);
nor U19052 (N_19052,N_10074,N_13972);
nor U19053 (N_19053,N_14304,N_12455);
nand U19054 (N_19054,N_12527,N_10981);
xnor U19055 (N_19055,N_14952,N_12704);
nor U19056 (N_19056,N_11293,N_10751);
or U19057 (N_19057,N_12836,N_11712);
or U19058 (N_19058,N_11065,N_12269);
and U19059 (N_19059,N_11362,N_11077);
and U19060 (N_19060,N_11659,N_13189);
nand U19061 (N_19061,N_14653,N_13703);
and U19062 (N_19062,N_12750,N_13496);
nor U19063 (N_19063,N_12642,N_12337);
or U19064 (N_19064,N_14690,N_12588);
nand U19065 (N_19065,N_13519,N_13302);
nor U19066 (N_19066,N_11958,N_13932);
and U19067 (N_19067,N_12417,N_12137);
xor U19068 (N_19068,N_13932,N_14046);
xnor U19069 (N_19069,N_13935,N_10451);
and U19070 (N_19070,N_11892,N_12934);
nand U19071 (N_19071,N_14784,N_13870);
or U19072 (N_19072,N_12817,N_13712);
or U19073 (N_19073,N_13267,N_12380);
nor U19074 (N_19074,N_13072,N_14715);
or U19075 (N_19075,N_11138,N_10917);
nand U19076 (N_19076,N_10458,N_10891);
nor U19077 (N_19077,N_12759,N_12017);
and U19078 (N_19078,N_13617,N_12589);
xnor U19079 (N_19079,N_10142,N_12675);
and U19080 (N_19080,N_11092,N_11716);
nand U19081 (N_19081,N_14200,N_10716);
or U19082 (N_19082,N_14507,N_14026);
and U19083 (N_19083,N_10028,N_14370);
nand U19084 (N_19084,N_10766,N_13963);
or U19085 (N_19085,N_10250,N_10424);
nand U19086 (N_19086,N_13410,N_14050);
nor U19087 (N_19087,N_12416,N_13592);
xnor U19088 (N_19088,N_10452,N_10416);
or U19089 (N_19089,N_12909,N_13932);
nor U19090 (N_19090,N_14116,N_12085);
nor U19091 (N_19091,N_12968,N_11603);
nor U19092 (N_19092,N_12995,N_11089);
or U19093 (N_19093,N_12536,N_13247);
nor U19094 (N_19094,N_12787,N_12933);
nand U19095 (N_19095,N_10522,N_14040);
xnor U19096 (N_19096,N_13347,N_10045);
nand U19097 (N_19097,N_13523,N_13874);
or U19098 (N_19098,N_10713,N_12319);
and U19099 (N_19099,N_10643,N_10208);
or U19100 (N_19100,N_11533,N_12038);
xor U19101 (N_19101,N_14653,N_10877);
nand U19102 (N_19102,N_11436,N_10565);
nand U19103 (N_19103,N_10921,N_11237);
nor U19104 (N_19104,N_11295,N_11634);
and U19105 (N_19105,N_14106,N_11686);
or U19106 (N_19106,N_10334,N_14015);
nor U19107 (N_19107,N_11045,N_11650);
and U19108 (N_19108,N_10242,N_11786);
xor U19109 (N_19109,N_12449,N_14108);
nand U19110 (N_19110,N_10486,N_14807);
xnor U19111 (N_19111,N_10873,N_10382);
nand U19112 (N_19112,N_10508,N_10513);
nand U19113 (N_19113,N_12526,N_12284);
and U19114 (N_19114,N_10259,N_10160);
or U19115 (N_19115,N_11092,N_11578);
nand U19116 (N_19116,N_10421,N_11079);
nor U19117 (N_19117,N_13343,N_13948);
or U19118 (N_19118,N_12579,N_12103);
nor U19119 (N_19119,N_12331,N_13289);
nand U19120 (N_19120,N_14203,N_13894);
and U19121 (N_19121,N_13446,N_11956);
xor U19122 (N_19122,N_11639,N_13116);
nor U19123 (N_19123,N_11335,N_12068);
nand U19124 (N_19124,N_13198,N_11997);
and U19125 (N_19125,N_11163,N_13735);
and U19126 (N_19126,N_11215,N_14287);
xnor U19127 (N_19127,N_10387,N_12350);
xor U19128 (N_19128,N_12738,N_11479);
nor U19129 (N_19129,N_11539,N_12188);
or U19130 (N_19130,N_10471,N_10238);
nor U19131 (N_19131,N_10789,N_10813);
and U19132 (N_19132,N_11817,N_14097);
nand U19133 (N_19133,N_13443,N_14389);
and U19134 (N_19134,N_14863,N_13444);
xor U19135 (N_19135,N_11302,N_14200);
nor U19136 (N_19136,N_14769,N_10899);
nand U19137 (N_19137,N_13121,N_13494);
nor U19138 (N_19138,N_11305,N_14289);
xor U19139 (N_19139,N_10202,N_11403);
xor U19140 (N_19140,N_11146,N_13344);
nor U19141 (N_19141,N_12441,N_13499);
nand U19142 (N_19142,N_10992,N_11319);
or U19143 (N_19143,N_10886,N_10372);
xor U19144 (N_19144,N_13741,N_13104);
nand U19145 (N_19145,N_10612,N_12469);
nand U19146 (N_19146,N_13759,N_14182);
nand U19147 (N_19147,N_10200,N_11838);
nor U19148 (N_19148,N_10966,N_14010);
nor U19149 (N_19149,N_13224,N_12446);
nand U19150 (N_19150,N_11448,N_12950);
and U19151 (N_19151,N_12958,N_10692);
nor U19152 (N_19152,N_13737,N_11405);
xor U19153 (N_19153,N_12912,N_13298);
nor U19154 (N_19154,N_14312,N_10046);
and U19155 (N_19155,N_13608,N_12079);
or U19156 (N_19156,N_12784,N_10410);
nand U19157 (N_19157,N_14222,N_14738);
and U19158 (N_19158,N_10000,N_14935);
and U19159 (N_19159,N_12579,N_12849);
nand U19160 (N_19160,N_12874,N_12792);
nor U19161 (N_19161,N_11514,N_11284);
nor U19162 (N_19162,N_13716,N_14176);
xor U19163 (N_19163,N_11003,N_10864);
nor U19164 (N_19164,N_13895,N_13582);
xor U19165 (N_19165,N_13355,N_14134);
xnor U19166 (N_19166,N_12218,N_11607);
and U19167 (N_19167,N_14421,N_11175);
and U19168 (N_19168,N_10836,N_13320);
and U19169 (N_19169,N_10966,N_12428);
or U19170 (N_19170,N_13313,N_14256);
and U19171 (N_19171,N_10608,N_11006);
xnor U19172 (N_19172,N_12906,N_13052);
nor U19173 (N_19173,N_13025,N_14507);
or U19174 (N_19174,N_11488,N_10387);
and U19175 (N_19175,N_11253,N_11660);
nand U19176 (N_19176,N_10605,N_12335);
nor U19177 (N_19177,N_11453,N_14989);
nand U19178 (N_19178,N_14589,N_13206);
and U19179 (N_19179,N_14828,N_14025);
or U19180 (N_19180,N_13563,N_10798);
xnor U19181 (N_19181,N_10096,N_11283);
nand U19182 (N_19182,N_11398,N_12530);
xnor U19183 (N_19183,N_13592,N_14397);
or U19184 (N_19184,N_10989,N_13945);
xor U19185 (N_19185,N_12218,N_11092);
and U19186 (N_19186,N_10876,N_11976);
xor U19187 (N_19187,N_11626,N_13471);
nor U19188 (N_19188,N_12520,N_13215);
nand U19189 (N_19189,N_14929,N_12079);
nand U19190 (N_19190,N_10267,N_11084);
and U19191 (N_19191,N_12162,N_11226);
nor U19192 (N_19192,N_11252,N_14631);
nand U19193 (N_19193,N_11769,N_12129);
xor U19194 (N_19194,N_12963,N_13093);
nor U19195 (N_19195,N_14831,N_14356);
nand U19196 (N_19196,N_11768,N_14554);
nand U19197 (N_19197,N_10605,N_10293);
and U19198 (N_19198,N_12714,N_13217);
xor U19199 (N_19199,N_14280,N_11563);
or U19200 (N_19200,N_12310,N_11770);
xor U19201 (N_19201,N_10003,N_13832);
or U19202 (N_19202,N_11239,N_12433);
xor U19203 (N_19203,N_12412,N_13628);
nand U19204 (N_19204,N_14459,N_10768);
xor U19205 (N_19205,N_12028,N_13106);
xor U19206 (N_19206,N_14169,N_13194);
xor U19207 (N_19207,N_11729,N_10790);
or U19208 (N_19208,N_14316,N_13531);
nand U19209 (N_19209,N_12117,N_13081);
nand U19210 (N_19210,N_11370,N_12148);
or U19211 (N_19211,N_13499,N_12164);
or U19212 (N_19212,N_10405,N_13526);
xnor U19213 (N_19213,N_14770,N_10141);
and U19214 (N_19214,N_14750,N_10763);
or U19215 (N_19215,N_14053,N_14450);
and U19216 (N_19216,N_14245,N_12968);
and U19217 (N_19217,N_10538,N_11433);
nand U19218 (N_19218,N_13538,N_14278);
nand U19219 (N_19219,N_12850,N_10252);
xnor U19220 (N_19220,N_10894,N_14786);
nor U19221 (N_19221,N_13864,N_14419);
nand U19222 (N_19222,N_12736,N_12933);
xor U19223 (N_19223,N_12799,N_12982);
nor U19224 (N_19224,N_12460,N_10637);
xor U19225 (N_19225,N_13331,N_14058);
nor U19226 (N_19226,N_10292,N_12864);
nor U19227 (N_19227,N_14513,N_11489);
nand U19228 (N_19228,N_13682,N_13587);
nor U19229 (N_19229,N_14759,N_14802);
and U19230 (N_19230,N_10177,N_12716);
nand U19231 (N_19231,N_10413,N_12656);
and U19232 (N_19232,N_11503,N_11634);
and U19233 (N_19233,N_10092,N_14726);
nand U19234 (N_19234,N_14118,N_14897);
nor U19235 (N_19235,N_13504,N_10178);
xor U19236 (N_19236,N_10527,N_12871);
and U19237 (N_19237,N_12100,N_13093);
xor U19238 (N_19238,N_10379,N_11859);
nor U19239 (N_19239,N_13469,N_11948);
or U19240 (N_19240,N_13137,N_11707);
nand U19241 (N_19241,N_13979,N_13640);
or U19242 (N_19242,N_11976,N_14310);
or U19243 (N_19243,N_11940,N_11241);
xnor U19244 (N_19244,N_12458,N_10566);
nand U19245 (N_19245,N_13980,N_12480);
nand U19246 (N_19246,N_14585,N_12691);
and U19247 (N_19247,N_13029,N_12219);
xnor U19248 (N_19248,N_11307,N_10734);
or U19249 (N_19249,N_12057,N_12167);
xor U19250 (N_19250,N_13888,N_12655);
nor U19251 (N_19251,N_11077,N_13977);
xnor U19252 (N_19252,N_11701,N_11393);
xnor U19253 (N_19253,N_11633,N_10205);
nor U19254 (N_19254,N_13735,N_14359);
or U19255 (N_19255,N_13974,N_12155);
xor U19256 (N_19256,N_10692,N_14485);
nand U19257 (N_19257,N_14811,N_13987);
and U19258 (N_19258,N_12842,N_12184);
or U19259 (N_19259,N_10573,N_13037);
nor U19260 (N_19260,N_11352,N_11268);
and U19261 (N_19261,N_10208,N_13016);
nand U19262 (N_19262,N_12680,N_12127);
xnor U19263 (N_19263,N_14281,N_10887);
or U19264 (N_19264,N_12490,N_13355);
xor U19265 (N_19265,N_11192,N_11977);
and U19266 (N_19266,N_12377,N_13813);
and U19267 (N_19267,N_11525,N_14742);
xor U19268 (N_19268,N_12708,N_13383);
or U19269 (N_19269,N_13641,N_11621);
and U19270 (N_19270,N_10700,N_12611);
and U19271 (N_19271,N_13761,N_12976);
or U19272 (N_19272,N_13457,N_12935);
and U19273 (N_19273,N_12026,N_10061);
nor U19274 (N_19274,N_11020,N_11175);
xor U19275 (N_19275,N_10505,N_12544);
nand U19276 (N_19276,N_11094,N_14913);
nor U19277 (N_19277,N_14464,N_13409);
nor U19278 (N_19278,N_12111,N_11541);
or U19279 (N_19279,N_10556,N_10744);
or U19280 (N_19280,N_11792,N_14170);
nand U19281 (N_19281,N_14351,N_13051);
or U19282 (N_19282,N_12324,N_13103);
or U19283 (N_19283,N_14254,N_11154);
nand U19284 (N_19284,N_14623,N_11378);
or U19285 (N_19285,N_14630,N_10368);
nand U19286 (N_19286,N_14407,N_13049);
nor U19287 (N_19287,N_11897,N_12310);
or U19288 (N_19288,N_14982,N_11106);
nor U19289 (N_19289,N_13062,N_12701);
or U19290 (N_19290,N_12180,N_13866);
nand U19291 (N_19291,N_10302,N_12159);
or U19292 (N_19292,N_14510,N_10602);
nor U19293 (N_19293,N_14729,N_11900);
xor U19294 (N_19294,N_11351,N_12936);
or U19295 (N_19295,N_11131,N_13069);
and U19296 (N_19296,N_13619,N_10551);
or U19297 (N_19297,N_13896,N_10408);
and U19298 (N_19298,N_12455,N_10726);
nor U19299 (N_19299,N_10704,N_11258);
and U19300 (N_19300,N_12090,N_12225);
nand U19301 (N_19301,N_11408,N_11929);
nand U19302 (N_19302,N_12606,N_12664);
nor U19303 (N_19303,N_12724,N_13634);
and U19304 (N_19304,N_14091,N_14369);
or U19305 (N_19305,N_10962,N_14449);
nand U19306 (N_19306,N_12901,N_12785);
and U19307 (N_19307,N_14552,N_10409);
or U19308 (N_19308,N_14795,N_13810);
nand U19309 (N_19309,N_10847,N_11482);
nand U19310 (N_19310,N_14989,N_12691);
or U19311 (N_19311,N_13828,N_11339);
nor U19312 (N_19312,N_12519,N_10180);
nand U19313 (N_19313,N_10593,N_10910);
or U19314 (N_19314,N_13425,N_12024);
nand U19315 (N_19315,N_11574,N_13542);
and U19316 (N_19316,N_14634,N_13624);
and U19317 (N_19317,N_14515,N_12812);
nor U19318 (N_19318,N_14094,N_12869);
or U19319 (N_19319,N_10021,N_14198);
nand U19320 (N_19320,N_11033,N_10341);
or U19321 (N_19321,N_10718,N_14585);
and U19322 (N_19322,N_10812,N_10317);
nor U19323 (N_19323,N_12694,N_10043);
or U19324 (N_19324,N_12133,N_14642);
and U19325 (N_19325,N_11818,N_13176);
and U19326 (N_19326,N_13935,N_13768);
nor U19327 (N_19327,N_13242,N_10540);
nand U19328 (N_19328,N_13630,N_14085);
nor U19329 (N_19329,N_14850,N_13429);
xor U19330 (N_19330,N_14523,N_12556);
or U19331 (N_19331,N_11577,N_14849);
nand U19332 (N_19332,N_14716,N_10775);
nand U19333 (N_19333,N_14907,N_12995);
or U19334 (N_19334,N_14009,N_11281);
and U19335 (N_19335,N_12538,N_13444);
or U19336 (N_19336,N_13132,N_14137);
and U19337 (N_19337,N_14550,N_13629);
nand U19338 (N_19338,N_12226,N_12854);
nand U19339 (N_19339,N_14439,N_12578);
or U19340 (N_19340,N_13189,N_12939);
xor U19341 (N_19341,N_13558,N_10788);
or U19342 (N_19342,N_13025,N_14117);
nand U19343 (N_19343,N_13640,N_14758);
or U19344 (N_19344,N_10918,N_12817);
xnor U19345 (N_19345,N_12105,N_11074);
and U19346 (N_19346,N_13239,N_11517);
nand U19347 (N_19347,N_13819,N_14604);
nor U19348 (N_19348,N_13480,N_12777);
xnor U19349 (N_19349,N_12194,N_10066);
nor U19350 (N_19350,N_12079,N_13120);
nand U19351 (N_19351,N_11526,N_11433);
or U19352 (N_19352,N_14955,N_13183);
nand U19353 (N_19353,N_13564,N_10534);
nor U19354 (N_19354,N_10933,N_13300);
nand U19355 (N_19355,N_12940,N_12504);
nand U19356 (N_19356,N_13375,N_12847);
and U19357 (N_19357,N_10605,N_10730);
xor U19358 (N_19358,N_11616,N_11315);
and U19359 (N_19359,N_14043,N_13029);
xor U19360 (N_19360,N_12318,N_13017);
and U19361 (N_19361,N_11966,N_13584);
nand U19362 (N_19362,N_10669,N_12346);
nand U19363 (N_19363,N_11891,N_13298);
nand U19364 (N_19364,N_10198,N_12586);
nand U19365 (N_19365,N_11279,N_13396);
or U19366 (N_19366,N_10649,N_13648);
xor U19367 (N_19367,N_13155,N_12166);
nand U19368 (N_19368,N_12934,N_11317);
nor U19369 (N_19369,N_11375,N_13351);
or U19370 (N_19370,N_12946,N_14528);
nand U19371 (N_19371,N_11387,N_12708);
or U19372 (N_19372,N_13534,N_14701);
and U19373 (N_19373,N_12765,N_12634);
or U19374 (N_19374,N_14662,N_12104);
nand U19375 (N_19375,N_13167,N_10229);
nor U19376 (N_19376,N_12900,N_11489);
and U19377 (N_19377,N_14712,N_12757);
nor U19378 (N_19378,N_14883,N_12433);
and U19379 (N_19379,N_14149,N_13252);
nand U19380 (N_19380,N_13634,N_14987);
or U19381 (N_19381,N_12650,N_13101);
or U19382 (N_19382,N_13617,N_14138);
nor U19383 (N_19383,N_12365,N_13083);
or U19384 (N_19384,N_11432,N_13279);
xnor U19385 (N_19385,N_13085,N_10311);
xor U19386 (N_19386,N_14873,N_10594);
nor U19387 (N_19387,N_10947,N_12824);
xor U19388 (N_19388,N_10940,N_14566);
and U19389 (N_19389,N_14974,N_12029);
nor U19390 (N_19390,N_14119,N_11075);
and U19391 (N_19391,N_13033,N_14925);
or U19392 (N_19392,N_13047,N_12791);
nand U19393 (N_19393,N_12848,N_11759);
or U19394 (N_19394,N_13700,N_13839);
nand U19395 (N_19395,N_10361,N_13906);
xor U19396 (N_19396,N_13963,N_10180);
nand U19397 (N_19397,N_11119,N_14902);
or U19398 (N_19398,N_10729,N_13638);
xor U19399 (N_19399,N_14351,N_13085);
xor U19400 (N_19400,N_10704,N_11955);
and U19401 (N_19401,N_11447,N_10632);
or U19402 (N_19402,N_12136,N_10769);
and U19403 (N_19403,N_14731,N_11625);
xnor U19404 (N_19404,N_10940,N_13308);
xor U19405 (N_19405,N_10441,N_10570);
or U19406 (N_19406,N_10388,N_14645);
and U19407 (N_19407,N_10564,N_11394);
nand U19408 (N_19408,N_14191,N_14142);
nand U19409 (N_19409,N_11659,N_14223);
or U19410 (N_19410,N_14761,N_12891);
xnor U19411 (N_19411,N_14524,N_11250);
nor U19412 (N_19412,N_11386,N_10799);
nand U19413 (N_19413,N_14941,N_11961);
xor U19414 (N_19414,N_14717,N_10763);
nand U19415 (N_19415,N_10205,N_10663);
nand U19416 (N_19416,N_14255,N_12141);
xor U19417 (N_19417,N_13171,N_11635);
or U19418 (N_19418,N_13252,N_13597);
and U19419 (N_19419,N_14704,N_12000);
nor U19420 (N_19420,N_12511,N_11729);
and U19421 (N_19421,N_13939,N_14301);
and U19422 (N_19422,N_13554,N_13680);
or U19423 (N_19423,N_13783,N_10723);
nand U19424 (N_19424,N_11476,N_10750);
or U19425 (N_19425,N_12035,N_12324);
nor U19426 (N_19426,N_11645,N_13277);
nand U19427 (N_19427,N_11969,N_14184);
nor U19428 (N_19428,N_14838,N_12932);
xor U19429 (N_19429,N_10518,N_13859);
nor U19430 (N_19430,N_11883,N_12872);
nand U19431 (N_19431,N_11961,N_10578);
or U19432 (N_19432,N_13513,N_14037);
nor U19433 (N_19433,N_12837,N_10952);
or U19434 (N_19434,N_11825,N_12581);
or U19435 (N_19435,N_14643,N_10268);
or U19436 (N_19436,N_12770,N_14742);
nor U19437 (N_19437,N_13453,N_11428);
xor U19438 (N_19438,N_12420,N_14256);
nor U19439 (N_19439,N_14139,N_12374);
nor U19440 (N_19440,N_10551,N_14217);
xnor U19441 (N_19441,N_14541,N_11736);
or U19442 (N_19442,N_14344,N_11652);
and U19443 (N_19443,N_13706,N_14922);
xnor U19444 (N_19444,N_10010,N_14130);
or U19445 (N_19445,N_10398,N_11699);
and U19446 (N_19446,N_10192,N_12695);
xor U19447 (N_19447,N_10587,N_11235);
or U19448 (N_19448,N_10860,N_13636);
nor U19449 (N_19449,N_14929,N_14625);
xor U19450 (N_19450,N_13830,N_12900);
and U19451 (N_19451,N_10925,N_13666);
and U19452 (N_19452,N_12946,N_13147);
or U19453 (N_19453,N_13580,N_10030);
nand U19454 (N_19454,N_11928,N_14910);
and U19455 (N_19455,N_11723,N_14084);
or U19456 (N_19456,N_13285,N_14772);
nor U19457 (N_19457,N_10518,N_11546);
xor U19458 (N_19458,N_12596,N_13223);
nand U19459 (N_19459,N_11697,N_14495);
or U19460 (N_19460,N_14395,N_12975);
nor U19461 (N_19461,N_11041,N_14762);
nor U19462 (N_19462,N_12915,N_12196);
nor U19463 (N_19463,N_12969,N_10224);
and U19464 (N_19464,N_14253,N_12657);
nand U19465 (N_19465,N_12876,N_12162);
nor U19466 (N_19466,N_10504,N_14369);
xnor U19467 (N_19467,N_13663,N_14016);
xor U19468 (N_19468,N_11636,N_11678);
xnor U19469 (N_19469,N_11759,N_10248);
and U19470 (N_19470,N_12108,N_13198);
xor U19471 (N_19471,N_11399,N_10757);
and U19472 (N_19472,N_11641,N_13229);
or U19473 (N_19473,N_14860,N_12489);
nand U19474 (N_19474,N_14314,N_10950);
or U19475 (N_19475,N_11603,N_12959);
nand U19476 (N_19476,N_10418,N_10364);
nor U19477 (N_19477,N_12230,N_12757);
xor U19478 (N_19478,N_10460,N_14828);
xor U19479 (N_19479,N_12660,N_13773);
xor U19480 (N_19480,N_14695,N_11187);
xor U19481 (N_19481,N_10860,N_13712);
or U19482 (N_19482,N_10392,N_12371);
and U19483 (N_19483,N_10476,N_12003);
or U19484 (N_19484,N_14445,N_13242);
nor U19485 (N_19485,N_13532,N_13628);
nand U19486 (N_19486,N_13606,N_11822);
and U19487 (N_19487,N_13725,N_13319);
and U19488 (N_19488,N_10255,N_11861);
nand U19489 (N_19489,N_13814,N_13473);
or U19490 (N_19490,N_13829,N_13524);
nor U19491 (N_19491,N_10650,N_12150);
and U19492 (N_19492,N_11625,N_14960);
nor U19493 (N_19493,N_10264,N_13450);
xor U19494 (N_19494,N_11292,N_13518);
or U19495 (N_19495,N_14811,N_11612);
nor U19496 (N_19496,N_13633,N_13148);
nor U19497 (N_19497,N_14998,N_11140);
xnor U19498 (N_19498,N_13044,N_11692);
nor U19499 (N_19499,N_13571,N_11574);
or U19500 (N_19500,N_10550,N_13058);
or U19501 (N_19501,N_10205,N_14470);
nor U19502 (N_19502,N_13730,N_11692);
or U19503 (N_19503,N_12889,N_13102);
and U19504 (N_19504,N_12794,N_11808);
nand U19505 (N_19505,N_13380,N_13033);
nor U19506 (N_19506,N_14202,N_10779);
xnor U19507 (N_19507,N_12804,N_12423);
or U19508 (N_19508,N_11636,N_13499);
and U19509 (N_19509,N_13994,N_10724);
and U19510 (N_19510,N_11731,N_13046);
or U19511 (N_19511,N_13185,N_12017);
xnor U19512 (N_19512,N_11772,N_14760);
nor U19513 (N_19513,N_11059,N_12713);
nor U19514 (N_19514,N_10327,N_14113);
nand U19515 (N_19515,N_14680,N_14356);
nor U19516 (N_19516,N_11836,N_14055);
nand U19517 (N_19517,N_10915,N_14102);
nand U19518 (N_19518,N_14725,N_11003);
nor U19519 (N_19519,N_14481,N_12576);
and U19520 (N_19520,N_10020,N_13041);
or U19521 (N_19521,N_12195,N_13168);
nand U19522 (N_19522,N_14049,N_12760);
nor U19523 (N_19523,N_11453,N_12210);
xnor U19524 (N_19524,N_13803,N_14826);
xor U19525 (N_19525,N_14923,N_14677);
nand U19526 (N_19526,N_10595,N_12790);
or U19527 (N_19527,N_10945,N_10833);
and U19528 (N_19528,N_14319,N_14772);
nor U19529 (N_19529,N_11635,N_14549);
xor U19530 (N_19530,N_13166,N_10035);
nor U19531 (N_19531,N_12027,N_14009);
and U19532 (N_19532,N_14815,N_12260);
xnor U19533 (N_19533,N_13835,N_12097);
and U19534 (N_19534,N_11245,N_10789);
nand U19535 (N_19535,N_12061,N_12245);
or U19536 (N_19536,N_11576,N_10396);
nand U19537 (N_19537,N_12226,N_10779);
nand U19538 (N_19538,N_12637,N_14391);
or U19539 (N_19539,N_11856,N_10986);
nor U19540 (N_19540,N_10412,N_10770);
xnor U19541 (N_19541,N_11769,N_14415);
nor U19542 (N_19542,N_12830,N_11760);
nand U19543 (N_19543,N_11525,N_11322);
and U19544 (N_19544,N_10357,N_12848);
and U19545 (N_19545,N_12236,N_12702);
or U19546 (N_19546,N_13352,N_14376);
nand U19547 (N_19547,N_10804,N_10279);
nand U19548 (N_19548,N_12234,N_11553);
and U19549 (N_19549,N_11123,N_10511);
or U19550 (N_19550,N_13979,N_14713);
nor U19551 (N_19551,N_14333,N_12780);
or U19552 (N_19552,N_11103,N_12848);
and U19553 (N_19553,N_14165,N_11412);
or U19554 (N_19554,N_13119,N_13128);
nor U19555 (N_19555,N_14690,N_11571);
nand U19556 (N_19556,N_10263,N_14658);
and U19557 (N_19557,N_10325,N_12382);
and U19558 (N_19558,N_14770,N_11468);
nor U19559 (N_19559,N_12784,N_13577);
nand U19560 (N_19560,N_11628,N_14880);
nor U19561 (N_19561,N_14491,N_13297);
xor U19562 (N_19562,N_14993,N_11080);
and U19563 (N_19563,N_13634,N_11789);
nand U19564 (N_19564,N_10543,N_11106);
xnor U19565 (N_19565,N_11904,N_11772);
or U19566 (N_19566,N_13964,N_14878);
and U19567 (N_19567,N_10325,N_13438);
nand U19568 (N_19568,N_14347,N_10313);
xnor U19569 (N_19569,N_11766,N_12157);
xnor U19570 (N_19570,N_14930,N_10343);
xnor U19571 (N_19571,N_13380,N_10172);
nand U19572 (N_19572,N_12709,N_14606);
or U19573 (N_19573,N_11328,N_14114);
xor U19574 (N_19574,N_12010,N_11317);
nor U19575 (N_19575,N_12925,N_14844);
or U19576 (N_19576,N_11249,N_11537);
or U19577 (N_19577,N_11905,N_10568);
xor U19578 (N_19578,N_10699,N_10145);
and U19579 (N_19579,N_11236,N_11634);
nor U19580 (N_19580,N_13870,N_10930);
nor U19581 (N_19581,N_13961,N_10138);
nand U19582 (N_19582,N_10130,N_13998);
xnor U19583 (N_19583,N_14313,N_10101);
or U19584 (N_19584,N_13445,N_10267);
nor U19585 (N_19585,N_11468,N_11268);
nand U19586 (N_19586,N_11657,N_10563);
nand U19587 (N_19587,N_11084,N_13225);
nand U19588 (N_19588,N_11638,N_14810);
nor U19589 (N_19589,N_13854,N_14368);
xnor U19590 (N_19590,N_12859,N_11938);
xnor U19591 (N_19591,N_12419,N_11856);
and U19592 (N_19592,N_11214,N_13428);
xnor U19593 (N_19593,N_12786,N_10930);
or U19594 (N_19594,N_13075,N_12435);
nand U19595 (N_19595,N_14147,N_14180);
nor U19596 (N_19596,N_13253,N_12360);
nor U19597 (N_19597,N_10197,N_14998);
or U19598 (N_19598,N_11875,N_14645);
and U19599 (N_19599,N_11437,N_12952);
nand U19600 (N_19600,N_12032,N_11074);
nand U19601 (N_19601,N_10638,N_13812);
and U19602 (N_19602,N_10991,N_13962);
nor U19603 (N_19603,N_13668,N_14386);
or U19604 (N_19604,N_13270,N_11196);
or U19605 (N_19605,N_14202,N_14091);
and U19606 (N_19606,N_14982,N_11516);
and U19607 (N_19607,N_13036,N_13909);
and U19608 (N_19608,N_12561,N_11496);
nor U19609 (N_19609,N_13054,N_11999);
or U19610 (N_19610,N_12212,N_10797);
nor U19611 (N_19611,N_12618,N_14254);
nor U19612 (N_19612,N_12006,N_13596);
nor U19613 (N_19613,N_11200,N_12274);
and U19614 (N_19614,N_10352,N_12859);
xor U19615 (N_19615,N_12335,N_12877);
nand U19616 (N_19616,N_14882,N_14128);
nor U19617 (N_19617,N_14541,N_14165);
and U19618 (N_19618,N_12586,N_13871);
nand U19619 (N_19619,N_12307,N_10299);
nor U19620 (N_19620,N_11474,N_14007);
xor U19621 (N_19621,N_10299,N_12926);
or U19622 (N_19622,N_10674,N_12757);
xor U19623 (N_19623,N_10534,N_12241);
or U19624 (N_19624,N_12424,N_14373);
nand U19625 (N_19625,N_11838,N_13809);
or U19626 (N_19626,N_12726,N_13491);
xnor U19627 (N_19627,N_13853,N_12702);
and U19628 (N_19628,N_10674,N_10142);
or U19629 (N_19629,N_13439,N_13253);
and U19630 (N_19630,N_11211,N_14243);
xnor U19631 (N_19631,N_10846,N_11634);
xor U19632 (N_19632,N_10229,N_14596);
nor U19633 (N_19633,N_12501,N_12756);
or U19634 (N_19634,N_12169,N_12497);
xnor U19635 (N_19635,N_13079,N_12797);
or U19636 (N_19636,N_13719,N_12386);
nor U19637 (N_19637,N_11784,N_10170);
and U19638 (N_19638,N_14914,N_11180);
and U19639 (N_19639,N_14411,N_10621);
or U19640 (N_19640,N_12372,N_12432);
nor U19641 (N_19641,N_13128,N_10532);
nand U19642 (N_19642,N_10606,N_10116);
nor U19643 (N_19643,N_12342,N_14632);
nand U19644 (N_19644,N_10611,N_13065);
xnor U19645 (N_19645,N_11409,N_11972);
nor U19646 (N_19646,N_14627,N_14525);
and U19647 (N_19647,N_11173,N_12530);
nor U19648 (N_19648,N_13294,N_13657);
nor U19649 (N_19649,N_10403,N_14424);
nor U19650 (N_19650,N_12348,N_13793);
xnor U19651 (N_19651,N_14235,N_10435);
xor U19652 (N_19652,N_11167,N_11018);
or U19653 (N_19653,N_11401,N_14093);
xnor U19654 (N_19654,N_11115,N_13624);
nor U19655 (N_19655,N_14930,N_11061);
and U19656 (N_19656,N_13878,N_11875);
nor U19657 (N_19657,N_13998,N_14207);
nand U19658 (N_19658,N_13768,N_10806);
xor U19659 (N_19659,N_13742,N_10320);
nor U19660 (N_19660,N_10351,N_13960);
and U19661 (N_19661,N_13597,N_10826);
nor U19662 (N_19662,N_13834,N_10681);
and U19663 (N_19663,N_11609,N_11220);
and U19664 (N_19664,N_11289,N_11684);
or U19665 (N_19665,N_11229,N_13396);
nor U19666 (N_19666,N_10522,N_13257);
nand U19667 (N_19667,N_13968,N_12901);
or U19668 (N_19668,N_12670,N_12990);
nor U19669 (N_19669,N_13215,N_12223);
xnor U19670 (N_19670,N_12006,N_14013);
nor U19671 (N_19671,N_12153,N_10775);
or U19672 (N_19672,N_10101,N_12413);
or U19673 (N_19673,N_10551,N_10075);
nand U19674 (N_19674,N_11239,N_14264);
nand U19675 (N_19675,N_10770,N_11627);
xnor U19676 (N_19676,N_12747,N_13989);
or U19677 (N_19677,N_14065,N_14653);
and U19678 (N_19678,N_12372,N_12919);
nor U19679 (N_19679,N_13847,N_10192);
or U19680 (N_19680,N_11859,N_12295);
nor U19681 (N_19681,N_12368,N_12268);
nand U19682 (N_19682,N_12860,N_11872);
xnor U19683 (N_19683,N_11884,N_13992);
nor U19684 (N_19684,N_10955,N_12253);
or U19685 (N_19685,N_12482,N_11446);
xor U19686 (N_19686,N_11413,N_13222);
and U19687 (N_19687,N_10492,N_10577);
xor U19688 (N_19688,N_13679,N_12552);
nand U19689 (N_19689,N_13517,N_11547);
xor U19690 (N_19690,N_11669,N_13421);
or U19691 (N_19691,N_13463,N_13392);
xor U19692 (N_19692,N_12321,N_10552);
and U19693 (N_19693,N_13232,N_13016);
nor U19694 (N_19694,N_13510,N_10902);
xor U19695 (N_19695,N_14797,N_11627);
nand U19696 (N_19696,N_13738,N_13223);
nand U19697 (N_19697,N_13505,N_10174);
nand U19698 (N_19698,N_11833,N_12360);
nor U19699 (N_19699,N_10728,N_14064);
and U19700 (N_19700,N_12213,N_12359);
or U19701 (N_19701,N_11268,N_12171);
nand U19702 (N_19702,N_10889,N_11325);
xor U19703 (N_19703,N_10376,N_10754);
xor U19704 (N_19704,N_10034,N_10648);
and U19705 (N_19705,N_11876,N_14751);
xnor U19706 (N_19706,N_14378,N_13745);
or U19707 (N_19707,N_11770,N_14548);
or U19708 (N_19708,N_12812,N_12790);
xor U19709 (N_19709,N_13803,N_12499);
nor U19710 (N_19710,N_11425,N_11705);
nand U19711 (N_19711,N_14168,N_12928);
and U19712 (N_19712,N_10138,N_11692);
nor U19713 (N_19713,N_14910,N_10262);
and U19714 (N_19714,N_12265,N_11283);
or U19715 (N_19715,N_14718,N_11972);
nor U19716 (N_19716,N_11973,N_11610);
nand U19717 (N_19717,N_13654,N_10918);
or U19718 (N_19718,N_14402,N_12698);
nand U19719 (N_19719,N_11858,N_12818);
nand U19720 (N_19720,N_13871,N_10953);
xor U19721 (N_19721,N_12301,N_12698);
and U19722 (N_19722,N_13483,N_11907);
nor U19723 (N_19723,N_11716,N_14519);
and U19724 (N_19724,N_14218,N_14865);
and U19725 (N_19725,N_13852,N_13622);
and U19726 (N_19726,N_14500,N_12283);
xor U19727 (N_19727,N_10772,N_12082);
nand U19728 (N_19728,N_10333,N_10241);
xor U19729 (N_19729,N_11610,N_13740);
nand U19730 (N_19730,N_13698,N_11872);
nor U19731 (N_19731,N_11434,N_13264);
nor U19732 (N_19732,N_12971,N_11807);
and U19733 (N_19733,N_12481,N_14515);
xor U19734 (N_19734,N_13402,N_10312);
nand U19735 (N_19735,N_12546,N_12234);
and U19736 (N_19736,N_11456,N_13722);
nor U19737 (N_19737,N_10152,N_10766);
nand U19738 (N_19738,N_14156,N_11990);
and U19739 (N_19739,N_14302,N_13078);
nand U19740 (N_19740,N_13568,N_11208);
or U19741 (N_19741,N_12442,N_13657);
nand U19742 (N_19742,N_11220,N_10408);
nor U19743 (N_19743,N_13443,N_12992);
or U19744 (N_19744,N_12119,N_14577);
nand U19745 (N_19745,N_10462,N_14061);
xor U19746 (N_19746,N_10866,N_14349);
and U19747 (N_19747,N_12205,N_12202);
nand U19748 (N_19748,N_10702,N_14409);
nand U19749 (N_19749,N_12031,N_10630);
nand U19750 (N_19750,N_14004,N_12772);
or U19751 (N_19751,N_14405,N_14878);
nand U19752 (N_19752,N_14824,N_14401);
nor U19753 (N_19753,N_14163,N_12423);
xor U19754 (N_19754,N_12887,N_12042);
xor U19755 (N_19755,N_10084,N_12082);
and U19756 (N_19756,N_12708,N_11080);
and U19757 (N_19757,N_14104,N_10827);
xnor U19758 (N_19758,N_10103,N_14541);
nand U19759 (N_19759,N_12112,N_12148);
nor U19760 (N_19760,N_14991,N_11443);
or U19761 (N_19761,N_12185,N_14840);
and U19762 (N_19762,N_13313,N_10908);
and U19763 (N_19763,N_14181,N_11660);
and U19764 (N_19764,N_12874,N_10380);
nor U19765 (N_19765,N_12402,N_11867);
nand U19766 (N_19766,N_11528,N_14533);
xor U19767 (N_19767,N_14869,N_12652);
xor U19768 (N_19768,N_10478,N_11102);
nor U19769 (N_19769,N_14494,N_12049);
and U19770 (N_19770,N_11123,N_14178);
nor U19771 (N_19771,N_10863,N_11190);
xnor U19772 (N_19772,N_11729,N_10231);
nor U19773 (N_19773,N_13783,N_13060);
and U19774 (N_19774,N_13991,N_12406);
or U19775 (N_19775,N_14030,N_10505);
and U19776 (N_19776,N_10033,N_11825);
nor U19777 (N_19777,N_12114,N_12254);
nand U19778 (N_19778,N_10926,N_12647);
xor U19779 (N_19779,N_10835,N_14749);
or U19780 (N_19780,N_11934,N_10928);
or U19781 (N_19781,N_14326,N_14378);
or U19782 (N_19782,N_14603,N_10179);
nand U19783 (N_19783,N_12729,N_12636);
xor U19784 (N_19784,N_13931,N_11927);
nor U19785 (N_19785,N_10887,N_12718);
and U19786 (N_19786,N_13675,N_11387);
nor U19787 (N_19787,N_14612,N_12508);
or U19788 (N_19788,N_14180,N_12956);
nand U19789 (N_19789,N_11074,N_13982);
nand U19790 (N_19790,N_13217,N_10307);
nor U19791 (N_19791,N_10736,N_14811);
nor U19792 (N_19792,N_10415,N_13267);
and U19793 (N_19793,N_13483,N_10582);
and U19794 (N_19794,N_14553,N_12560);
nor U19795 (N_19795,N_12956,N_14070);
or U19796 (N_19796,N_13280,N_14078);
nor U19797 (N_19797,N_14121,N_10935);
nand U19798 (N_19798,N_10501,N_12618);
and U19799 (N_19799,N_10284,N_12218);
or U19800 (N_19800,N_14939,N_10742);
and U19801 (N_19801,N_11244,N_12486);
or U19802 (N_19802,N_11875,N_12121);
nor U19803 (N_19803,N_14429,N_13084);
nor U19804 (N_19804,N_12781,N_12722);
nor U19805 (N_19805,N_14195,N_14644);
or U19806 (N_19806,N_13011,N_13346);
nor U19807 (N_19807,N_11561,N_13562);
nor U19808 (N_19808,N_10565,N_11835);
xor U19809 (N_19809,N_13937,N_13267);
xnor U19810 (N_19810,N_13087,N_12086);
nand U19811 (N_19811,N_13318,N_13671);
xor U19812 (N_19812,N_12897,N_10320);
nand U19813 (N_19813,N_12355,N_12901);
and U19814 (N_19814,N_11721,N_12221);
nor U19815 (N_19815,N_10472,N_10043);
xor U19816 (N_19816,N_11238,N_10150);
or U19817 (N_19817,N_10064,N_10203);
nor U19818 (N_19818,N_13920,N_14406);
nor U19819 (N_19819,N_13495,N_11992);
xor U19820 (N_19820,N_12935,N_11553);
and U19821 (N_19821,N_11388,N_14734);
and U19822 (N_19822,N_11244,N_12758);
and U19823 (N_19823,N_12980,N_13082);
xnor U19824 (N_19824,N_13285,N_13401);
nor U19825 (N_19825,N_10881,N_11795);
nor U19826 (N_19826,N_13179,N_11626);
xor U19827 (N_19827,N_12438,N_14154);
nor U19828 (N_19828,N_13015,N_10915);
xnor U19829 (N_19829,N_10855,N_14392);
xor U19830 (N_19830,N_13485,N_14179);
and U19831 (N_19831,N_13803,N_12669);
nand U19832 (N_19832,N_14553,N_12297);
and U19833 (N_19833,N_10321,N_14361);
nor U19834 (N_19834,N_12494,N_11287);
or U19835 (N_19835,N_12099,N_12473);
nor U19836 (N_19836,N_10235,N_13439);
xnor U19837 (N_19837,N_14234,N_14157);
nor U19838 (N_19838,N_11373,N_10908);
or U19839 (N_19839,N_14489,N_10204);
and U19840 (N_19840,N_12877,N_11466);
xnor U19841 (N_19841,N_12055,N_13811);
nor U19842 (N_19842,N_14044,N_14225);
nand U19843 (N_19843,N_14801,N_14955);
xnor U19844 (N_19844,N_11543,N_11080);
xnor U19845 (N_19845,N_13800,N_13835);
and U19846 (N_19846,N_10907,N_12936);
xnor U19847 (N_19847,N_10334,N_13380);
and U19848 (N_19848,N_14918,N_13403);
nor U19849 (N_19849,N_13588,N_13821);
nand U19850 (N_19850,N_14343,N_11786);
nand U19851 (N_19851,N_10778,N_10793);
or U19852 (N_19852,N_10056,N_11767);
nand U19853 (N_19853,N_13794,N_10622);
xnor U19854 (N_19854,N_14049,N_12209);
or U19855 (N_19855,N_13990,N_10447);
nor U19856 (N_19856,N_13792,N_13138);
nor U19857 (N_19857,N_11314,N_13288);
nor U19858 (N_19858,N_10717,N_13674);
or U19859 (N_19859,N_14528,N_14058);
nor U19860 (N_19860,N_10272,N_14036);
and U19861 (N_19861,N_13123,N_14615);
nor U19862 (N_19862,N_13476,N_14120);
nor U19863 (N_19863,N_13143,N_10120);
xor U19864 (N_19864,N_10182,N_10431);
nor U19865 (N_19865,N_14760,N_10963);
xor U19866 (N_19866,N_12925,N_10305);
xor U19867 (N_19867,N_11274,N_10768);
and U19868 (N_19868,N_10667,N_13800);
xnor U19869 (N_19869,N_11747,N_14507);
and U19870 (N_19870,N_10128,N_14421);
or U19871 (N_19871,N_11005,N_12117);
xnor U19872 (N_19872,N_13036,N_12634);
xor U19873 (N_19873,N_12653,N_13965);
nor U19874 (N_19874,N_14151,N_12401);
and U19875 (N_19875,N_13581,N_12405);
and U19876 (N_19876,N_14139,N_11100);
nor U19877 (N_19877,N_11089,N_14013);
or U19878 (N_19878,N_11568,N_11698);
nor U19879 (N_19879,N_10884,N_10314);
nor U19880 (N_19880,N_11260,N_10445);
or U19881 (N_19881,N_10616,N_13694);
nor U19882 (N_19882,N_12418,N_11142);
or U19883 (N_19883,N_12216,N_11313);
nor U19884 (N_19884,N_13403,N_14063);
or U19885 (N_19885,N_11613,N_13993);
and U19886 (N_19886,N_10052,N_10776);
nand U19887 (N_19887,N_14909,N_14430);
nor U19888 (N_19888,N_12944,N_14674);
xor U19889 (N_19889,N_11733,N_10267);
and U19890 (N_19890,N_10831,N_11229);
or U19891 (N_19891,N_14642,N_11560);
and U19892 (N_19892,N_12059,N_10857);
or U19893 (N_19893,N_11486,N_13378);
or U19894 (N_19894,N_14848,N_10978);
nand U19895 (N_19895,N_10073,N_14070);
and U19896 (N_19896,N_13649,N_14077);
xor U19897 (N_19897,N_12950,N_12347);
nand U19898 (N_19898,N_11934,N_10162);
nor U19899 (N_19899,N_12870,N_12922);
xor U19900 (N_19900,N_12930,N_14607);
nand U19901 (N_19901,N_10329,N_13990);
nor U19902 (N_19902,N_14659,N_14662);
or U19903 (N_19903,N_14007,N_14962);
nor U19904 (N_19904,N_12616,N_13601);
nor U19905 (N_19905,N_14417,N_13169);
and U19906 (N_19906,N_13929,N_12807);
nor U19907 (N_19907,N_10840,N_10934);
or U19908 (N_19908,N_12234,N_12183);
and U19909 (N_19909,N_10155,N_14262);
or U19910 (N_19910,N_14948,N_10940);
nand U19911 (N_19911,N_14715,N_14157);
xor U19912 (N_19912,N_13535,N_14128);
nand U19913 (N_19913,N_14381,N_10909);
and U19914 (N_19914,N_13027,N_11893);
or U19915 (N_19915,N_11014,N_12417);
nor U19916 (N_19916,N_12554,N_10637);
or U19917 (N_19917,N_14697,N_12697);
nor U19918 (N_19918,N_12656,N_10613);
and U19919 (N_19919,N_14243,N_10001);
and U19920 (N_19920,N_11660,N_10187);
nand U19921 (N_19921,N_12267,N_11643);
and U19922 (N_19922,N_10884,N_14534);
and U19923 (N_19923,N_11194,N_12744);
nor U19924 (N_19924,N_10031,N_11244);
nand U19925 (N_19925,N_12755,N_14270);
or U19926 (N_19926,N_13732,N_12142);
or U19927 (N_19927,N_12408,N_14761);
nor U19928 (N_19928,N_10727,N_11075);
and U19929 (N_19929,N_14851,N_11639);
or U19930 (N_19930,N_10734,N_10156);
nor U19931 (N_19931,N_12151,N_13075);
or U19932 (N_19932,N_10136,N_10346);
nand U19933 (N_19933,N_14222,N_11414);
xor U19934 (N_19934,N_11007,N_13648);
or U19935 (N_19935,N_10011,N_14044);
xnor U19936 (N_19936,N_12651,N_13494);
xor U19937 (N_19937,N_10717,N_14082);
nand U19938 (N_19938,N_14760,N_12168);
nor U19939 (N_19939,N_14156,N_10350);
xor U19940 (N_19940,N_10425,N_11763);
nand U19941 (N_19941,N_12615,N_10657);
nand U19942 (N_19942,N_13283,N_14927);
or U19943 (N_19943,N_10929,N_10018);
nand U19944 (N_19944,N_14171,N_12850);
xor U19945 (N_19945,N_10647,N_14623);
nor U19946 (N_19946,N_13046,N_11196);
nand U19947 (N_19947,N_14243,N_13822);
xnor U19948 (N_19948,N_14892,N_10386);
and U19949 (N_19949,N_14328,N_13215);
and U19950 (N_19950,N_13572,N_11340);
nor U19951 (N_19951,N_13042,N_13852);
xor U19952 (N_19952,N_11390,N_10101);
or U19953 (N_19953,N_12455,N_11302);
and U19954 (N_19954,N_13979,N_10306);
nand U19955 (N_19955,N_14541,N_12581);
or U19956 (N_19956,N_11173,N_13594);
nor U19957 (N_19957,N_14578,N_10003);
and U19958 (N_19958,N_10713,N_14109);
nand U19959 (N_19959,N_10313,N_14814);
xnor U19960 (N_19960,N_11869,N_14170);
or U19961 (N_19961,N_11556,N_11915);
nor U19962 (N_19962,N_14358,N_12262);
nor U19963 (N_19963,N_10090,N_14129);
xnor U19964 (N_19964,N_13180,N_14829);
and U19965 (N_19965,N_11026,N_14422);
and U19966 (N_19966,N_14064,N_14279);
and U19967 (N_19967,N_12270,N_10517);
nor U19968 (N_19968,N_11913,N_11305);
xnor U19969 (N_19969,N_11456,N_10529);
nand U19970 (N_19970,N_13411,N_11832);
or U19971 (N_19971,N_14941,N_11041);
and U19972 (N_19972,N_14368,N_12271);
nand U19973 (N_19973,N_11442,N_13951);
xnor U19974 (N_19974,N_12254,N_11214);
xnor U19975 (N_19975,N_13922,N_13781);
and U19976 (N_19976,N_12373,N_13426);
or U19977 (N_19977,N_10891,N_14997);
and U19978 (N_19978,N_10384,N_11627);
nand U19979 (N_19979,N_14022,N_13882);
nor U19980 (N_19980,N_14910,N_12451);
nand U19981 (N_19981,N_14989,N_11334);
nor U19982 (N_19982,N_11646,N_14503);
or U19983 (N_19983,N_13672,N_11445);
nand U19984 (N_19984,N_10498,N_13018);
or U19985 (N_19985,N_10019,N_10896);
nand U19986 (N_19986,N_14286,N_11481);
nand U19987 (N_19987,N_14895,N_13298);
xnor U19988 (N_19988,N_13894,N_13585);
and U19989 (N_19989,N_13424,N_11086);
and U19990 (N_19990,N_11772,N_14950);
nor U19991 (N_19991,N_12663,N_14649);
and U19992 (N_19992,N_10279,N_11057);
and U19993 (N_19993,N_11562,N_11462);
and U19994 (N_19994,N_10775,N_13272);
xnor U19995 (N_19995,N_13273,N_13677);
and U19996 (N_19996,N_10046,N_12849);
or U19997 (N_19997,N_12085,N_10490);
nor U19998 (N_19998,N_13689,N_12307);
or U19999 (N_19999,N_12165,N_10833);
nor U20000 (N_20000,N_16455,N_16046);
or U20001 (N_20001,N_15305,N_16875);
xnor U20002 (N_20002,N_15149,N_17715);
or U20003 (N_20003,N_19072,N_17235);
and U20004 (N_20004,N_18038,N_16208);
or U20005 (N_20005,N_19608,N_15201);
nand U20006 (N_20006,N_15555,N_17902);
and U20007 (N_20007,N_19076,N_15457);
nor U20008 (N_20008,N_18718,N_15652);
and U20009 (N_20009,N_18155,N_16191);
nand U20010 (N_20010,N_19572,N_19595);
and U20011 (N_20011,N_15812,N_15725);
and U20012 (N_20012,N_18206,N_19111);
xnor U20013 (N_20013,N_18546,N_15968);
nand U20014 (N_20014,N_16591,N_19253);
xor U20015 (N_20015,N_18180,N_17267);
or U20016 (N_20016,N_17071,N_15281);
xnor U20017 (N_20017,N_18482,N_19776);
xor U20018 (N_20018,N_19600,N_16107);
or U20019 (N_20019,N_17865,N_19470);
or U20020 (N_20020,N_16829,N_15401);
nand U20021 (N_20021,N_16753,N_16346);
nor U20022 (N_20022,N_17953,N_18664);
or U20023 (N_20023,N_15418,N_15164);
nand U20024 (N_20024,N_17882,N_18888);
or U20025 (N_20025,N_15475,N_16968);
and U20026 (N_20026,N_16088,N_18793);
or U20027 (N_20027,N_15801,N_18365);
nor U20028 (N_20028,N_17873,N_15733);
and U20029 (N_20029,N_18489,N_16070);
nand U20030 (N_20030,N_19280,N_19724);
nand U20031 (N_20031,N_18873,N_19794);
nor U20032 (N_20032,N_15240,N_19315);
or U20033 (N_20033,N_19124,N_18896);
xor U20034 (N_20034,N_18390,N_18118);
nand U20035 (N_20035,N_17472,N_17611);
and U20036 (N_20036,N_18802,N_17745);
nand U20037 (N_20037,N_19996,N_19549);
nand U20038 (N_20038,N_15851,N_19486);
and U20039 (N_20039,N_16958,N_16872);
nand U20040 (N_20040,N_18187,N_18071);
nor U20041 (N_20041,N_16659,N_17102);
xor U20042 (N_20042,N_17558,N_15916);
nor U20043 (N_20043,N_19478,N_16501);
nand U20044 (N_20044,N_16527,N_16584);
nand U20045 (N_20045,N_16755,N_19156);
xor U20046 (N_20046,N_18894,N_19363);
or U20047 (N_20047,N_18007,N_19561);
or U20048 (N_20048,N_18198,N_18634);
or U20049 (N_20049,N_15450,N_18490);
nand U20050 (N_20050,N_15207,N_16413);
xnor U20051 (N_20051,N_18231,N_17785);
and U20052 (N_20052,N_18632,N_15501);
and U20053 (N_20053,N_17887,N_19268);
nand U20054 (N_20054,N_19061,N_17288);
and U20055 (N_20055,N_17796,N_16327);
or U20056 (N_20056,N_19224,N_18650);
nand U20057 (N_20057,N_17083,N_19176);
nand U20058 (N_20058,N_16975,N_18004);
xor U20059 (N_20059,N_18125,N_17879);
nand U20060 (N_20060,N_16229,N_18758);
or U20061 (N_20061,N_18767,N_16093);
nand U20062 (N_20062,N_18835,N_17355);
nor U20063 (N_20063,N_17639,N_16378);
xnor U20064 (N_20064,N_17492,N_19093);
nor U20065 (N_20065,N_17268,N_16832);
or U20066 (N_20066,N_16948,N_18436);
and U20067 (N_20067,N_15705,N_18573);
nor U20068 (N_20068,N_18615,N_15712);
nand U20069 (N_20069,N_18417,N_18558);
xor U20070 (N_20070,N_16175,N_17884);
xnor U20071 (N_20071,N_17407,N_15101);
xor U20072 (N_20072,N_18995,N_19181);
xor U20073 (N_20073,N_17219,N_18282);
and U20074 (N_20074,N_16526,N_18566);
nand U20075 (N_20075,N_19946,N_15218);
nor U20076 (N_20076,N_17846,N_15790);
and U20077 (N_20077,N_19381,N_15889);
nor U20078 (N_20078,N_18757,N_19959);
nand U20079 (N_20079,N_17381,N_16538);
nor U20080 (N_20080,N_15408,N_17520);
and U20081 (N_20081,N_19948,N_16807);
nand U20082 (N_20082,N_17425,N_16317);
or U20083 (N_20083,N_19351,N_19547);
xor U20084 (N_20084,N_19443,N_16994);
nand U20085 (N_20085,N_17229,N_19252);
xnor U20086 (N_20086,N_18147,N_19166);
and U20087 (N_20087,N_16903,N_18189);
nand U20088 (N_20088,N_19522,N_16089);
or U20089 (N_20089,N_16788,N_15217);
and U20090 (N_20090,N_15188,N_17194);
nor U20091 (N_20091,N_19021,N_19190);
and U20092 (N_20092,N_17391,N_18322);
nand U20093 (N_20093,N_15148,N_19630);
and U20094 (N_20094,N_16440,N_17678);
or U20095 (N_20095,N_15129,N_19006);
xor U20096 (N_20096,N_17210,N_19922);
or U20097 (N_20097,N_18608,N_15043);
and U20098 (N_20098,N_16113,N_17066);
xor U20099 (N_20099,N_19038,N_15280);
or U20100 (N_20100,N_16028,N_16776);
and U20101 (N_20101,N_17767,N_17203);
nor U20102 (N_20102,N_19282,N_15484);
xnor U20103 (N_20103,N_17113,N_15195);
or U20104 (N_20104,N_18245,N_18841);
or U20105 (N_20105,N_18360,N_17603);
nor U20106 (N_20106,N_15035,N_17868);
nand U20107 (N_20107,N_17711,N_15828);
nor U20108 (N_20108,N_17597,N_15838);
and U20109 (N_20109,N_19047,N_16141);
or U20110 (N_20110,N_16812,N_17314);
nand U20111 (N_20111,N_15206,N_17515);
nand U20112 (N_20112,N_17240,N_19070);
and U20113 (N_20113,N_19951,N_17329);
nand U20114 (N_20114,N_16055,N_15753);
and U20115 (N_20115,N_18585,N_16937);
nor U20116 (N_20116,N_15063,N_15496);
xnor U20117 (N_20117,N_18748,N_19103);
xor U20118 (N_20118,N_16018,N_15593);
and U20119 (N_20119,N_18285,N_16219);
or U20120 (N_20120,N_15056,N_18456);
or U20121 (N_20121,N_17810,N_19267);
nand U20122 (N_20122,N_17260,N_19845);
nor U20123 (N_20123,N_19806,N_16772);
and U20124 (N_20124,N_15514,N_15703);
and U20125 (N_20125,N_17275,N_18715);
or U20126 (N_20126,N_19820,N_17859);
or U20127 (N_20127,N_17590,N_16846);
or U20128 (N_20128,N_17885,N_17814);
xnor U20129 (N_20129,N_19165,N_19403);
xor U20130 (N_20130,N_18750,N_19074);
xor U20131 (N_20131,N_15756,N_18814);
xnor U20132 (N_20132,N_18528,N_19586);
or U20133 (N_20133,N_18240,N_19380);
nor U20134 (N_20134,N_17896,N_18840);
nand U20135 (N_20135,N_18455,N_18296);
and U20136 (N_20136,N_16934,N_18011);
nor U20137 (N_20137,N_17848,N_15465);
or U20138 (N_20138,N_17093,N_18998);
or U20139 (N_20139,N_16890,N_18391);
nor U20140 (N_20140,N_16943,N_15910);
nor U20141 (N_20141,N_15510,N_15880);
nand U20142 (N_20142,N_19968,N_18491);
or U20143 (N_20143,N_19782,N_17759);
xor U20144 (N_20144,N_16740,N_19678);
nor U20145 (N_20145,N_17345,N_19213);
nor U20146 (N_20146,N_15602,N_15476);
xor U20147 (N_20147,N_16822,N_15170);
nand U20148 (N_20148,N_19541,N_19494);
xor U20149 (N_20149,N_17995,N_15692);
nor U20150 (N_20150,N_18570,N_16213);
xor U20151 (N_20151,N_16969,N_15117);
or U20152 (N_20152,N_16759,N_15949);
nand U20153 (N_20153,N_15539,N_19344);
and U20154 (N_20154,N_19923,N_15924);
xor U20155 (N_20155,N_17531,N_16463);
nor U20156 (N_20156,N_17226,N_16879);
nor U20157 (N_20157,N_18920,N_16429);
and U20158 (N_20158,N_15805,N_15367);
and U20159 (N_20159,N_17812,N_17735);
and U20160 (N_20160,N_18041,N_19312);
nand U20161 (N_20161,N_16284,N_19303);
xnor U20162 (N_20162,N_16290,N_19437);
or U20163 (N_20163,N_16108,N_19179);
xnor U20164 (N_20164,N_17933,N_19596);
nand U20165 (N_20165,N_15875,N_15983);
nand U20166 (N_20166,N_17128,N_19565);
nor U20167 (N_20167,N_19877,N_16913);
nor U20168 (N_20168,N_17680,N_16619);
nand U20169 (N_20169,N_18178,N_19276);
nand U20170 (N_20170,N_16823,N_18454);
and U20171 (N_20171,N_17147,N_19854);
or U20172 (N_20172,N_18075,N_18599);
xor U20173 (N_20173,N_16079,N_17955);
nor U20174 (N_20174,N_19762,N_19090);
nand U20175 (N_20175,N_17162,N_17572);
nor U20176 (N_20176,N_18547,N_18830);
or U20177 (N_20177,N_17943,N_15592);
nand U20178 (N_20178,N_17006,N_17914);
or U20179 (N_20179,N_15970,N_19432);
or U20180 (N_20180,N_17251,N_16194);
or U20181 (N_20181,N_16671,N_17893);
or U20182 (N_20182,N_18232,N_16332);
and U20183 (N_20183,N_19399,N_16647);
or U20184 (N_20184,N_19089,N_17794);
nor U20185 (N_20185,N_16187,N_18156);
nand U20186 (N_20186,N_15861,N_19961);
nand U20187 (N_20187,N_17758,N_19429);
xor U20188 (N_20188,N_18336,N_16425);
nor U20189 (N_20189,N_15126,N_19096);
xor U20190 (N_20190,N_18042,N_18527);
nor U20191 (N_20191,N_15553,N_17625);
or U20192 (N_20192,N_18100,N_18465);
and U20193 (N_20193,N_18638,N_17840);
nor U20194 (N_20194,N_19669,N_15283);
and U20195 (N_20195,N_19894,N_19498);
or U20196 (N_20196,N_18500,N_16940);
xnor U20197 (N_20197,N_16092,N_16151);
nand U20198 (N_20198,N_18159,N_19508);
xor U20199 (N_20199,N_19099,N_16736);
or U20200 (N_20200,N_18609,N_15909);
nor U20201 (N_20201,N_15731,N_15893);
or U20202 (N_20202,N_15879,N_15963);
nand U20203 (N_20203,N_15495,N_19775);
nor U20204 (N_20204,N_19689,N_15176);
xor U20205 (N_20205,N_16986,N_15435);
or U20206 (N_20206,N_18225,N_18405);
nand U20207 (N_20207,N_17349,N_16119);
xor U20208 (N_20208,N_16922,N_19200);
xor U20209 (N_20209,N_18483,N_17201);
xor U20210 (N_20210,N_15022,N_16503);
xor U20211 (N_20211,N_19095,N_18526);
or U20212 (N_20212,N_16198,N_17602);
xor U20213 (N_20213,N_17576,N_19605);
nor U20214 (N_20214,N_18452,N_16631);
or U20215 (N_20215,N_15672,N_16997);
nand U20216 (N_20216,N_18622,N_19856);
xor U20217 (N_20217,N_16657,N_18657);
and U20218 (N_20218,N_19926,N_15048);
xnor U20219 (N_20219,N_19274,N_16921);
or U20220 (N_20220,N_16809,N_15862);
xnor U20221 (N_20221,N_18503,N_16827);
and U20222 (N_20222,N_15121,N_16556);
nand U20223 (N_20223,N_19516,N_15980);
nor U20224 (N_20224,N_16794,N_17437);
and U20225 (N_20225,N_16085,N_18906);
nor U20226 (N_20226,N_19874,N_15696);
xor U20227 (N_20227,N_19320,N_17925);
and U20228 (N_20228,N_18374,N_15651);
xnor U20229 (N_20229,N_17718,N_18471);
or U20230 (N_20230,N_17140,N_16916);
nor U20231 (N_20231,N_19699,N_15671);
nand U20232 (N_20232,N_16204,N_15675);
nor U20233 (N_20233,N_18492,N_16318);
xnor U20234 (N_20234,N_18626,N_18843);
xnor U20235 (N_20235,N_15982,N_16241);
xnor U20236 (N_20236,N_18340,N_15603);
nor U20237 (N_20237,N_15444,N_17823);
nand U20238 (N_20238,N_19542,N_15609);
xnor U20239 (N_20239,N_18665,N_16615);
nor U20240 (N_20240,N_19566,N_17648);
xnor U20241 (N_20241,N_15921,N_19206);
nor U20242 (N_20242,N_18025,N_16032);
nand U20243 (N_20243,N_18596,N_18082);
nor U20244 (N_20244,N_19835,N_15704);
and U20245 (N_20245,N_16023,N_17042);
xor U20246 (N_20246,N_16878,N_16133);
or U20247 (N_20247,N_19771,N_18382);
or U20248 (N_20248,N_17212,N_16954);
xor U20249 (N_20249,N_16818,N_15650);
or U20250 (N_20250,N_16730,N_19126);
or U20251 (N_20251,N_15338,N_16163);
nand U20252 (N_20252,N_17408,N_19384);
and U20253 (N_20253,N_15189,N_18164);
or U20254 (N_20254,N_19246,N_17555);
xor U20255 (N_20255,N_19169,N_15220);
xor U20256 (N_20256,N_15831,N_17633);
nand U20257 (N_20257,N_16069,N_16930);
xnor U20258 (N_20258,N_15071,N_18459);
and U20259 (N_20259,N_19515,N_19302);
nor U20260 (N_20260,N_17372,N_18036);
and U20261 (N_20261,N_16140,N_18348);
nor U20262 (N_20262,N_16369,N_19507);
xor U20263 (N_20263,N_15489,N_16273);
nor U20264 (N_20264,N_18811,N_16443);
and U20265 (N_20265,N_17849,N_17365);
and U20266 (N_20266,N_19603,N_15225);
and U20267 (N_20267,N_17522,N_17820);
or U20268 (N_20268,N_17973,N_18263);
nand U20269 (N_20269,N_18303,N_17748);
nor U20270 (N_20270,N_16002,N_18883);
nand U20271 (N_20271,N_17516,N_19199);
nor U20272 (N_20272,N_18555,N_16102);
nor U20273 (N_20273,N_18831,N_15302);
and U20274 (N_20274,N_16644,N_16299);
nand U20275 (N_20275,N_15244,N_19534);
nand U20276 (N_20276,N_17808,N_15318);
nor U20277 (N_20277,N_17374,N_19901);
nand U20278 (N_20278,N_16293,N_17112);
and U20279 (N_20279,N_15449,N_19373);
xnor U20280 (N_20280,N_19598,N_15517);
nor U20281 (N_20281,N_16675,N_17618);
xor U20282 (N_20282,N_18495,N_19532);
xor U20283 (N_20283,N_17709,N_18597);
nand U20284 (N_20284,N_16221,N_15429);
nand U20285 (N_20285,N_17154,N_19406);
xnor U20286 (N_20286,N_15904,N_19488);
xor U20287 (N_20287,N_15908,N_16546);
or U20288 (N_20288,N_15962,N_15422);
nand U20289 (N_20289,N_17048,N_15621);
nor U20290 (N_20290,N_16388,N_15072);
and U20291 (N_20291,N_16248,N_15946);
nand U20292 (N_20292,N_15740,N_17857);
xnor U20293 (N_20293,N_15741,N_19651);
or U20294 (N_20294,N_17111,N_18212);
xnor U20295 (N_20295,N_18955,N_19658);
xnor U20296 (N_20296,N_18305,N_16034);
xnor U20297 (N_20297,N_17412,N_18950);
or U20298 (N_20298,N_17629,N_16166);
nor U20299 (N_20299,N_19855,N_18122);
and U20300 (N_20300,N_18691,N_16033);
nor U20301 (N_20301,N_19864,N_16974);
nand U20302 (N_20302,N_16987,N_17346);
and U20303 (N_20303,N_18891,N_17978);
xor U20304 (N_20304,N_15665,N_18781);
xnor U20305 (N_20305,N_16124,N_19537);
xor U20306 (N_20306,N_15468,N_16328);
nor U20307 (N_20307,N_16439,N_15491);
nor U20308 (N_20308,N_19747,N_18809);
and U20309 (N_20309,N_18525,N_18266);
xnor U20310 (N_20310,N_17155,N_17593);
or U20311 (N_20311,N_18034,N_19029);
and U20312 (N_20312,N_16656,N_19389);
nand U20313 (N_20313,N_15009,N_15549);
xor U20314 (N_20314,N_15407,N_16494);
xnor U20315 (N_20315,N_18307,N_18451);
nor U20316 (N_20316,N_18045,N_16923);
xnor U20317 (N_20317,N_15886,N_15451);
nor U20318 (N_20318,N_18858,N_17187);
nand U20319 (N_20319,N_19256,N_15290);
or U20320 (N_20320,N_17135,N_16300);
or U20321 (N_20321,N_16622,N_16845);
or U20322 (N_20322,N_16808,N_19997);
nor U20323 (N_20323,N_16098,N_18816);
xor U20324 (N_20324,N_16007,N_19628);
nor U20325 (N_20325,N_15850,N_18227);
nand U20326 (N_20326,N_17222,N_17687);
xnor U20327 (N_20327,N_17844,N_17872);
nor U20328 (N_20328,N_15837,N_19388);
nand U20329 (N_20329,N_18580,N_17185);
and U20330 (N_20330,N_16104,N_16607);
nor U20331 (N_20331,N_17538,N_16375);
and U20332 (N_20332,N_15299,N_18229);
nor U20333 (N_20333,N_17689,N_16931);
or U20334 (N_20334,N_17769,N_18397);
nor U20335 (N_20335,N_19920,N_17601);
or U20336 (N_20336,N_15049,N_15682);
xnor U20337 (N_20337,N_19003,N_16022);
or U20338 (N_20338,N_16350,N_17549);
nor U20339 (N_20339,N_15626,N_17526);
nand U20340 (N_20340,N_16574,N_17174);
xnor U20341 (N_20341,N_18532,N_18935);
or U20342 (N_20342,N_16458,N_16478);
and U20343 (N_20343,N_15986,N_16825);
and U20344 (N_20344,N_19697,N_18588);
or U20345 (N_20345,N_19058,N_16233);
and U20346 (N_20346,N_18694,N_15414);
nand U20347 (N_20347,N_16467,N_19191);
or U20348 (N_20348,N_18378,N_18910);
nand U20349 (N_20349,N_17898,N_15421);
nor U20350 (N_20350,N_16596,N_19945);
or U20351 (N_20351,N_15097,N_17254);
nor U20352 (N_20352,N_17191,N_15025);
xor U20353 (N_20353,N_18933,N_16887);
nand U20354 (N_20354,N_19487,N_15782);
or U20355 (N_20355,N_15127,N_15803);
or U20356 (N_20356,N_19196,N_19609);
xnor U20357 (N_20357,N_16760,N_19346);
xnor U20358 (N_20358,N_17904,N_18361);
nand U20359 (N_20359,N_19261,N_15095);
nand U20360 (N_20360,N_16168,N_17188);
and U20361 (N_20361,N_15992,N_17989);
xor U20362 (N_20362,N_17837,N_16843);
xnor U20363 (N_20363,N_15324,N_16705);
nor U20364 (N_20364,N_15300,N_19048);
nor U20365 (N_20365,N_16801,N_16679);
and U20366 (N_20366,N_18496,N_18467);
or U20367 (N_20367,N_18123,N_17511);
nand U20368 (N_20368,N_15387,N_16531);
nor U20369 (N_20369,N_16989,N_16586);
xnor U20370 (N_20370,N_19045,N_15277);
xor U20371 (N_20371,N_18217,N_18044);
xnor U20372 (N_20372,N_19382,N_18519);
nor U20373 (N_20373,N_18362,N_15917);
or U20374 (N_20374,N_19475,N_19777);
xor U20375 (N_20375,N_17471,N_15858);
xnor U20376 (N_20376,N_18683,N_15981);
and U20377 (N_20377,N_17959,N_17836);
or U20378 (N_20378,N_15397,N_16919);
and U20379 (N_20379,N_18902,N_17302);
nor U20380 (N_20380,N_18652,N_16762);
xor U20381 (N_20381,N_15774,N_18511);
or U20382 (N_20382,N_19020,N_19618);
and U20383 (N_20383,N_17273,N_19909);
nor U20384 (N_20384,N_17514,N_16186);
nand U20385 (N_20385,N_18872,N_17775);
nand U20386 (N_20386,N_15957,N_18055);
or U20387 (N_20387,N_16145,N_18333);
and U20388 (N_20388,N_16828,N_17119);
nand U20389 (N_20389,N_19078,N_16949);
xnor U20390 (N_20390,N_19885,N_15051);
and U20391 (N_20391,N_19337,N_15565);
xnor U20392 (N_20392,N_15988,N_17057);
or U20393 (N_20393,N_16642,N_16382);
nand U20394 (N_20394,N_15822,N_19214);
nand U20395 (N_20395,N_17532,N_15003);
or U20396 (N_20396,N_17192,N_16424);
and U20397 (N_20397,N_16540,N_17728);
or U20398 (N_20398,N_16848,N_16988);
xor U20399 (N_20399,N_18523,N_18753);
nor U20400 (N_20400,N_18952,N_17536);
nand U20401 (N_20401,N_17352,N_18969);
or U20402 (N_20402,N_17517,N_19615);
nand U20403 (N_20403,N_18716,N_17905);
nor U20404 (N_20404,N_19913,N_19499);
nand U20405 (N_20405,N_15524,N_16894);
nor U20406 (N_20406,N_18117,N_19573);
or U20407 (N_20407,N_15347,N_17220);
or U20408 (N_20408,N_19583,N_16881);
nor U20409 (N_20409,N_17132,N_15416);
nand U20410 (N_20410,N_16261,N_19435);
nor U20411 (N_20411,N_16539,N_18545);
and U20412 (N_20412,N_16364,N_18326);
nor U20413 (N_20413,N_17109,N_17323);
and U20414 (N_20414,N_17371,N_16851);
and U20415 (N_20415,N_15174,N_18438);
xnor U20416 (N_20416,N_18425,N_15854);
nor U20417 (N_20417,N_16998,N_19447);
and U20418 (N_20418,N_17282,N_15698);
and U20419 (N_20419,N_15033,N_17938);
xnor U20420 (N_20420,N_15105,N_15770);
xnor U20421 (N_20421,N_19819,N_16157);
and U20422 (N_20422,N_19188,N_19841);
and U20423 (N_20423,N_17842,N_16918);
nand U20424 (N_20424,N_18763,N_18332);
and U20425 (N_20425,N_18761,N_17742);
nand U20426 (N_20426,N_19730,N_16372);
nand U20427 (N_20427,N_19980,N_19080);
and U20428 (N_20428,N_17475,N_17403);
or U20429 (N_20429,N_17064,N_17544);
nor U20430 (N_20430,N_18087,N_15202);
nor U20431 (N_20431,N_15469,N_17202);
and U20432 (N_20432,N_19333,N_18542);
or U20433 (N_20433,N_17419,N_18909);
nor U20434 (N_20434,N_18801,N_15474);
nor U20435 (N_20435,N_18138,N_19278);
xnor U20436 (N_20436,N_19789,N_17861);
xor U20437 (N_20437,N_15155,N_17279);
nand U20438 (N_20438,N_19202,N_16123);
xnor U20439 (N_20439,N_15586,N_15527);
and U20440 (N_20440,N_15960,N_16814);
and U20441 (N_20441,N_15434,N_15417);
or U20442 (N_20442,N_18821,N_15800);
and U20443 (N_20443,N_17644,N_16307);
nor U20444 (N_20444,N_19275,N_18863);
xor U20445 (N_20445,N_16353,N_18892);
xor U20446 (N_20446,N_17691,N_15882);
xor U20447 (N_20447,N_16184,N_18593);
nand U20448 (N_20448,N_19121,N_15707);
or U20449 (N_20449,N_19262,N_15848);
nand U20450 (N_20450,N_18053,N_15793);
or U20451 (N_20451,N_19555,N_16831);
xnor U20452 (N_20452,N_15291,N_18137);
or U20453 (N_20453,N_16066,N_15866);
nand U20454 (N_20454,N_18901,N_18017);
and U20455 (N_20455,N_15536,N_16227);
nand U20456 (N_20456,N_16534,N_18331);
nor U20457 (N_20457,N_15409,N_17751);
or U20458 (N_20458,N_18869,N_17473);
and U20459 (N_20459,N_15124,N_16874);
or U20460 (N_20460,N_17491,N_16756);
nor U20461 (N_20461,N_17874,N_19627);
or U20462 (N_20462,N_19787,N_19659);
or U20463 (N_20463,N_17411,N_15273);
and U20464 (N_20464,N_15261,N_19938);
nand U20465 (N_20465,N_19291,N_16286);
xnor U20466 (N_20466,N_15019,N_19013);
nand U20467 (N_20467,N_17047,N_16014);
xor U20468 (N_20468,N_17609,N_17813);
or U20469 (N_20469,N_17432,N_16572);
nor U20470 (N_20470,N_17090,N_19729);
nor U20471 (N_20471,N_19670,N_19872);
and U20472 (N_20472,N_17598,N_17443);
nor U20473 (N_20473,N_16838,N_19438);
nand U20474 (N_20474,N_19958,N_15256);
nand U20475 (N_20475,N_19073,N_19621);
nand U20476 (N_20476,N_17106,N_19813);
nand U20477 (N_20477,N_17004,N_15050);
or U20478 (N_20478,N_18380,N_15406);
or U20479 (N_20479,N_16487,N_18182);
xor U20480 (N_20480,N_16368,N_18766);
nand U20481 (N_20481,N_16763,N_19554);
or U20482 (N_20482,N_18195,N_19408);
xnor U20483 (N_20483,N_15311,N_18899);
nor U20484 (N_20484,N_16668,N_16196);
xnor U20485 (N_20485,N_18795,N_15412);
xor U20486 (N_20486,N_16908,N_15929);
nor U20487 (N_20487,N_19184,N_16739);
nor U20488 (N_20488,N_15065,N_17750);
xor U20489 (N_20489,N_16249,N_16345);
xnor U20490 (N_20490,N_18537,N_16649);
and U20491 (N_20491,N_15702,N_16446);
and U20492 (N_20492,N_16004,N_16427);
or U20493 (N_20493,N_18258,N_18981);
nor U20494 (N_20494,N_17685,N_19891);
and U20495 (N_20495,N_16543,N_19442);
xnor U20496 (N_20496,N_17460,N_15867);
nor U20497 (N_20497,N_16884,N_18329);
xnor U20498 (N_20498,N_18242,N_15445);
and U20499 (N_20499,N_15041,N_16010);
xor U20500 (N_20500,N_16702,N_16689);
or U20501 (N_20501,N_19455,N_15091);
and U20502 (N_20502,N_16161,N_16135);
and U20503 (N_20503,N_18165,N_19803);
nor U20504 (N_20504,N_19809,N_16311);
and U20505 (N_20505,N_19687,N_19154);
or U20506 (N_20506,N_15729,N_15561);
and U20507 (N_20507,N_19266,N_18295);
nor U20508 (N_20508,N_16246,N_19461);
and U20509 (N_20509,N_19342,N_17605);
and U20510 (N_20510,N_16565,N_18889);
and U20511 (N_20511,N_15670,N_16500);
nand U20512 (N_20512,N_15374,N_15958);
nor U20513 (N_20513,N_19263,N_15552);
and U20514 (N_20514,N_16064,N_16337);
nand U20515 (N_20515,N_17054,N_18399);
xnor U20516 (N_20516,N_18563,N_19748);
and U20517 (N_20517,N_18447,N_18518);
and U20518 (N_20518,N_16789,N_18944);
and U20519 (N_20519,N_19796,N_17741);
and U20520 (N_20520,N_19490,N_16871);
and U20521 (N_20521,N_19402,N_17831);
nor U20522 (N_20522,N_18999,N_18866);
nand U20523 (N_20523,N_17667,N_17005);
or U20524 (N_20524,N_17197,N_15947);
nor U20525 (N_20525,N_16235,N_17012);
and U20526 (N_20526,N_15485,N_17638);
nor U20527 (N_20527,N_17918,N_15020);
xnor U20528 (N_20528,N_18008,N_15316);
nor U20529 (N_20529,N_17799,N_15143);
or U20530 (N_20530,N_16059,N_15508);
nor U20531 (N_20531,N_18444,N_19919);
xor U20532 (N_20532,N_15656,N_17175);
nand U20533 (N_20533,N_19599,N_19513);
xnor U20534 (N_20534,N_18068,N_16432);
nor U20535 (N_20535,N_16143,N_16376);
xor U20536 (N_20536,N_16356,N_15221);
nand U20537 (N_20537,N_19299,N_19613);
xor U20538 (N_20538,N_18091,N_15855);
nand U20539 (N_20539,N_18635,N_16225);
nor U20540 (N_20540,N_15312,N_16431);
or U20541 (N_20541,N_18148,N_18112);
and U20542 (N_20542,N_17506,N_18660);
nor U20543 (N_20543,N_16562,N_16274);
nor U20544 (N_20544,N_16258,N_16043);
xnor U20545 (N_20545,N_17650,N_18162);
nand U20546 (N_20546,N_19870,N_15590);
or U20547 (N_20547,N_15781,N_19726);
or U20548 (N_20548,N_15658,N_17205);
nand U20549 (N_20549,N_18111,N_15115);
nand U20550 (N_20550,N_18515,N_18721);
or U20551 (N_20551,N_17830,N_18375);
nor U20552 (N_20552,N_19300,N_16481);
xor U20553 (N_20553,N_18705,N_18880);
xor U20554 (N_20554,N_18719,N_15404);
and U20555 (N_20555,N_19394,N_15039);
xnor U20556 (N_20556,N_16605,N_15697);
and U20557 (N_20557,N_15490,N_16506);
and U20558 (N_20558,N_19497,N_16724);
nor U20559 (N_20559,N_19007,N_19986);
nand U20560 (N_20560,N_16365,N_15606);
nor U20561 (N_20561,N_16402,N_18048);
nand U20562 (N_20562,N_19847,N_19036);
or U20563 (N_20563,N_18449,N_15826);
or U20564 (N_20564,N_15827,N_16497);
or U20565 (N_20565,N_16722,N_17131);
and U20566 (N_20566,N_16484,N_17714);
and U20567 (N_20567,N_19100,N_19718);
nand U20568 (N_20568,N_15266,N_19112);
and U20569 (N_20569,N_16557,N_18393);
or U20570 (N_20570,N_16938,N_18269);
nor U20571 (N_20571,N_18330,N_15876);
xor U20572 (N_20572,N_16054,N_18236);
nor U20573 (N_20573,N_19527,N_15341);
or U20574 (N_20574,N_17947,N_16276);
or U20575 (N_20575,N_19859,N_16090);
nand U20576 (N_20576,N_15177,N_15190);
or U20577 (N_20577,N_17024,N_15940);
xnor U20578 (N_20578,N_16990,N_19136);
or U20579 (N_20579,N_17073,N_16624);
xor U20580 (N_20580,N_17583,N_18559);
nand U20581 (N_20581,N_18176,N_17604);
xnor U20582 (N_20582,N_18643,N_15197);
or U20583 (N_20583,N_17247,N_19876);
nor U20584 (N_20584,N_18640,N_16880);
nor U20585 (N_20585,N_19039,N_16272);
and U20586 (N_20586,N_15974,N_19560);
or U20587 (N_20587,N_18696,N_17353);
or U20588 (N_20588,N_18824,N_17449);
and U20589 (N_20589,N_19964,N_19348);
or U20590 (N_20590,N_17701,N_19028);
and U20591 (N_20591,N_17284,N_18898);
xnor U20592 (N_20592,N_18003,N_18109);
xnor U20593 (N_20593,N_19883,N_15506);
xnor U20594 (N_20594,N_17014,N_17551);
nand U20595 (N_20595,N_16857,N_17541);
nand U20596 (N_20596,N_18141,N_15994);
nand U20597 (N_20597,N_17161,N_19294);
or U20598 (N_20598,N_16169,N_17241);
nor U20599 (N_20599,N_17866,N_15248);
or U20600 (N_20600,N_15157,N_17002);
or U20601 (N_20601,N_15171,N_15928);
or U20602 (N_20602,N_15259,N_17152);
or U20603 (N_20603,N_15955,N_19652);
xnor U20604 (N_20604,N_15158,N_17429);
or U20605 (N_20605,N_16533,N_18557);
xor U20606 (N_20606,N_16991,N_17646);
nor U20607 (N_20607,N_17708,N_19982);
or U20608 (N_20608,N_16254,N_15515);
nand U20609 (N_20609,N_16952,N_18723);
nand U20610 (N_20610,N_15094,N_16853);
xor U20611 (N_20611,N_18280,N_17296);
and U20612 (N_20612,N_15138,N_16426);
or U20613 (N_20613,N_17428,N_16685);
nor U20614 (N_20614,N_17299,N_16452);
nor U20615 (N_20615,N_15328,N_17744);
or U20616 (N_20616,N_18768,N_19395);
and U20617 (N_20617,N_15423,N_19973);
and U20618 (N_20618,N_16688,N_17032);
nand U20619 (N_20619,N_19321,N_18413);
or U20620 (N_20620,N_18062,N_16547);
and U20621 (N_20621,N_15556,N_17682);
or U20622 (N_20622,N_15722,N_15236);
xor U20623 (N_20623,N_17041,N_17945);
and U20624 (N_20624,N_19293,N_15676);
or U20625 (N_20625,N_16966,N_19692);
or U20626 (N_20626,N_18246,N_16640);
and U20627 (N_20627,N_19998,N_17439);
nor U20628 (N_20628,N_18470,N_19145);
or U20629 (N_20629,N_16524,N_19327);
nor U20630 (N_20630,N_16901,N_19479);
nor U20631 (N_20631,N_15926,N_17825);
nor U20632 (N_20632,N_18059,N_19183);
and U20633 (N_20633,N_17231,N_18601);
nor U20634 (N_20634,N_19104,N_19842);
nor U20635 (N_20635,N_18612,N_19120);
and U20636 (N_20636,N_17760,N_17738);
nand U20637 (N_20637,N_18578,N_17712);
xor U20638 (N_20638,N_19535,N_19939);
nand U20639 (N_20639,N_18047,N_17971);
nand U20640 (N_20640,N_15153,N_15905);
or U20641 (N_20641,N_19836,N_17803);
nand U20642 (N_20642,N_17243,N_18679);
and U20643 (N_20643,N_19744,N_15724);
nand U20644 (N_20644,N_16933,N_16103);
and U20645 (N_20645,N_19457,N_17434);
nor U20646 (N_20646,N_15122,N_16433);
or U20647 (N_20647,N_19960,N_18403);
nand U20648 (N_20648,N_16544,N_18056);
nor U20649 (N_20649,N_15734,N_18404);
nand U20650 (N_20650,N_18063,N_19170);
nand U20651 (N_20651,N_19465,N_17436);
nor U20652 (N_20652,N_19323,N_16182);
nand U20653 (N_20653,N_16232,N_19310);
xnor U20654 (N_20654,N_17636,N_17903);
nor U20655 (N_20655,N_18319,N_18868);
nor U20656 (N_20656,N_15991,N_18663);
nand U20657 (N_20657,N_19826,N_17822);
nand U20658 (N_20658,N_18544,N_18905);
xor U20659 (N_20659,N_18215,N_19420);
or U20660 (N_20660,N_16076,N_16520);
and U20661 (N_20661,N_17787,N_15016);
xnor U20662 (N_20662,N_18254,N_17567);
xnor U20663 (N_20663,N_16928,N_15364);
and U20664 (N_20664,N_15522,N_15535);
and U20665 (N_20665,N_15638,N_19059);
nor U20666 (N_20666,N_17060,N_19837);
xor U20667 (N_20667,N_17668,N_17962);
nand U20668 (N_20668,N_15802,N_16891);
nor U20669 (N_20669,N_16780,N_19518);
nor U20670 (N_20670,N_18780,N_18140);
nor U20671 (N_20671,N_19311,N_18325);
or U20672 (N_20672,N_18862,N_18987);
xnor U20673 (N_20673,N_16456,N_15820);
nor U20674 (N_20674,N_19756,N_16821);
xor U20675 (N_20675,N_19064,N_17496);
and U20676 (N_20676,N_16164,N_18341);
nor U20677 (N_20677,N_18357,N_15425);
nand U20678 (N_20678,N_19387,N_19807);
nor U20679 (N_20679,N_16834,N_17963);
and U20680 (N_20680,N_19220,N_19257);
nor U20681 (N_20681,N_17422,N_15642);
nor U20682 (N_20682,N_19705,N_17886);
or U20683 (N_20683,N_16256,N_16582);
xnor U20684 (N_20684,N_15732,N_16265);
xor U20685 (N_20685,N_15894,N_17941);
and U20686 (N_20686,N_16109,N_16121);
xnor U20687 (N_20687,N_15680,N_19460);
or U20688 (N_20688,N_19753,N_19269);
nor U20689 (N_20689,N_15113,N_15006);
nor U20690 (N_20690,N_18787,N_15394);
xnor U20691 (N_20691,N_19580,N_17207);
nand U20692 (N_20692,N_19009,N_17450);
xnor U20693 (N_20693,N_16067,N_15868);
or U20694 (N_20694,N_15282,N_15079);
or U20695 (N_20695,N_19236,N_18418);
nor U20696 (N_20696,N_16844,N_17923);
or U20697 (N_20697,N_16600,N_16550);
or U20698 (N_20698,N_16053,N_18688);
xnor U20699 (N_20699,N_19174,N_19458);
xor U20700 (N_20700,N_15270,N_18172);
or U20701 (N_20701,N_18817,N_19423);
nand U20702 (N_20702,N_18288,N_17483);
and U20703 (N_20703,N_17754,N_15896);
or U20704 (N_20704,N_15687,N_17485);
and U20705 (N_20705,N_19553,N_15996);
nor U20706 (N_20706,N_16960,N_15183);
and U20707 (N_20707,N_16291,N_18453);
and U20708 (N_20708,N_18169,N_16083);
nand U20709 (N_20709,N_18583,N_15613);
nor U20710 (N_20710,N_17277,N_16263);
and U20711 (N_20711,N_17944,N_15550);
nor U20712 (N_20712,N_18370,N_19211);
nand U20713 (N_20713,N_16692,N_17440);
nand U20714 (N_20714,N_15078,N_15276);
and U20715 (N_20715,N_19229,N_15534);
or U20716 (N_20716,N_17620,N_15605);
nand U20717 (N_20717,N_18006,N_19758);
nand U20718 (N_20718,N_16980,N_15380);
xor U20719 (N_20719,N_15577,N_15737);
xnor U20720 (N_20720,N_17635,N_15459);
nor U20721 (N_20721,N_17081,N_16514);
nor U20722 (N_20722,N_19785,N_19892);
and U20723 (N_20723,N_17510,N_19590);
nand U20724 (N_20724,N_19115,N_19993);
nor U20725 (N_20725,N_19407,N_19832);
xnor U20726 (N_20726,N_18256,N_19614);
nand U20727 (N_20727,N_15109,N_19216);
or U20728 (N_20728,N_18692,N_16224);
nand U20729 (N_20729,N_19390,N_17461);
and U20730 (N_20730,N_17564,N_19866);
or U20731 (N_20731,N_19084,N_16522);
and U20732 (N_20732,N_18791,N_16459);
nand U20733 (N_20733,N_17375,N_18207);
or U20734 (N_20734,N_15932,N_15021);
and U20735 (N_20735,N_17170,N_17610);
or U20736 (N_20736,N_17967,N_19693);
nor U20737 (N_20737,N_17557,N_19301);
nand U20738 (N_20738,N_16144,N_16051);
and U20739 (N_20739,N_19101,N_17974);
xor U20740 (N_20740,N_15254,N_16793);
nor U20741 (N_20741,N_18535,N_16435);
xnor U20742 (N_20742,N_15952,N_15611);
nor U20743 (N_20743,N_15814,N_17936);
xnor U20744 (N_20744,N_17166,N_18353);
nand U20745 (N_20745,N_19283,N_19632);
xor U20746 (N_20746,N_18339,N_15106);
nand U20747 (N_20747,N_17988,N_18481);
and U20748 (N_20748,N_17015,N_17493);
xor U20749 (N_20749,N_18666,N_18179);
or U20750 (N_20750,N_15622,N_16334);
nor U20751 (N_20751,N_17530,N_15985);
or U20752 (N_20752,N_16488,N_19338);
nor U20753 (N_20753,N_16742,N_17423);
and U20754 (N_20754,N_15114,N_18363);
or U20755 (N_20755,N_18107,N_18421);
nor U20756 (N_20756,N_16012,N_16939);
or U20757 (N_20757,N_17757,N_19130);
nor U20758 (N_20758,N_19625,N_18359);
and U20759 (N_20759,N_15509,N_19526);
or U20760 (N_20760,N_15120,N_17780);
or U20761 (N_20761,N_16951,N_18110);
or U20762 (N_20762,N_15075,N_17915);
or U20763 (N_20763,N_16301,N_16850);
xor U20764 (N_20764,N_18427,N_19289);
nor U20765 (N_20765,N_19340,N_18653);
nor U20766 (N_20766,N_19077,N_16461);
or U20767 (N_20767,N_15247,N_16895);
nor U20768 (N_20768,N_19336,N_19034);
and U20769 (N_20769,N_16472,N_17599);
or U20770 (N_20770,N_19426,N_18709);
and U20771 (N_20771,N_15245,N_18291);
or U20772 (N_20772,N_19709,N_17743);
or U20773 (N_20773,N_19931,N_15162);
nor U20774 (N_20774,N_17817,N_18671);
nor U20775 (N_20775,N_17634,N_19117);
nor U20776 (N_20776,N_17395,N_15648);
nand U20777 (N_20777,N_18002,N_15654);
or U20778 (N_20778,N_17975,N_19149);
or U20779 (N_20779,N_16528,N_16183);
nor U20780 (N_20780,N_15199,N_19393);
xor U20781 (N_20781,N_18230,N_17070);
nand U20782 (N_20782,N_15745,N_19242);
nand U20783 (N_20783,N_16197,N_16324);
or U20784 (N_20784,N_17591,N_15209);
xnor U20785 (N_20785,N_15255,N_17125);
or U20786 (N_20786,N_19633,N_17547);
nor U20787 (N_20787,N_17357,N_18571);
and U20788 (N_20788,N_17930,N_19306);
and U20789 (N_20789,N_17637,N_17911);
nand U20790 (N_20790,N_19671,N_15856);
and U20791 (N_20791,N_18556,N_18297);
nand U20792 (N_20792,N_16149,N_15521);
nand U20793 (N_20793,N_19057,N_19831);
or U20794 (N_20794,N_15865,N_19168);
nor U20795 (N_20795,N_15797,N_19052);
nor U20796 (N_20796,N_15070,N_16660);
and U20797 (N_20797,N_15965,N_15739);
nand U20798 (N_20798,N_15333,N_15187);
xor U20799 (N_20799,N_19933,N_16267);
and U20800 (N_20800,N_18922,N_17939);
nor U20801 (N_20801,N_16945,N_15872);
xor U20802 (N_20802,N_16451,N_16779);
and U20803 (N_20803,N_15242,N_18347);
nor U20804 (N_20804,N_16535,N_19251);
xnor U20805 (N_20805,N_15604,N_17431);
nor U20806 (N_20806,N_15504,N_17778);
and U20807 (N_20807,N_16266,N_17901);
xor U20808 (N_20808,N_15751,N_15877);
xnor U20809 (N_20809,N_18493,N_19701);
nor U20810 (N_20810,N_19489,N_15104);
nand U20811 (N_20811,N_17335,N_15554);
and U20812 (N_20812,N_19231,N_17038);
and U20813 (N_20813,N_15036,N_16097);
nor U20814 (N_20814,N_18783,N_19025);
and U20815 (N_20815,N_17786,N_19287);
nor U20816 (N_20816,N_15579,N_16518);
and U20817 (N_20817,N_16806,N_17578);
or U20818 (N_20818,N_18916,N_17149);
or U20819 (N_20819,N_16302,N_18774);
xnor U20820 (N_20820,N_19882,N_18770);
xnor U20821 (N_20821,N_18560,N_17684);
or U20822 (N_20822,N_17232,N_19896);
nor U20823 (N_20823,N_17151,N_18312);
and U20824 (N_20824,N_17924,N_19715);
nor U20825 (N_20825,N_17107,N_19296);
and U20826 (N_20826,N_18521,N_18050);
or U20827 (N_20827,N_17631,N_19362);
nand U20828 (N_20828,N_18818,N_16729);
xnor U20829 (N_20829,N_19349,N_15040);
or U20830 (N_20830,N_17972,N_16925);
nand U20831 (N_20831,N_17942,N_19792);
nor U20832 (N_20832,N_17360,N_17392);
nor U20833 (N_20833,N_16700,N_17080);
nand U20834 (N_20834,N_15499,N_15863);
nand U20835 (N_20835,N_19440,N_18376);
xnor U20836 (N_20836,N_17791,N_15337);
xor U20837 (N_20837,N_17084,N_18116);
or U20838 (N_20838,N_19132,N_15513);
nor U20839 (N_20839,N_16652,N_16005);
and U20840 (N_20840,N_16201,N_15296);
and U20841 (N_20841,N_15062,N_18913);
or U20842 (N_20842,N_18623,N_19122);
xor U20843 (N_20843,N_15540,N_16096);
xnor U20844 (N_20844,N_17693,N_17069);
and U20845 (N_20845,N_19163,N_15287);
and U20846 (N_20846,N_18021,N_15743);
and U20847 (N_20847,N_18619,N_18414);
nor U20848 (N_20848,N_17292,N_15666);
xnor U20849 (N_20849,N_19880,N_17761);
and U20850 (N_20850,N_15026,N_15156);
nand U20851 (N_20851,N_16728,N_17688);
xor U20852 (N_20852,N_16548,N_16062);
or U20853 (N_20853,N_19906,N_15585);
and U20854 (N_20854,N_17805,N_17897);
or U20855 (N_20855,N_15146,N_18985);
nand U20856 (N_20856,N_15525,N_15567);
xor U20857 (N_20857,N_18589,N_19279);
and U20858 (N_20858,N_17580,N_17354);
nand U20859 (N_20859,N_18161,N_18067);
or U20860 (N_20860,N_16165,N_18392);
nor U20861 (N_20861,N_19019,N_17659);
or U20862 (N_20862,N_19375,N_18158);
nand U20863 (N_20863,N_16329,N_18243);
xor U20864 (N_20864,N_16902,N_18014);
nor U20865 (N_20865,N_17263,N_16638);
xnor U20866 (N_20866,N_16347,N_17417);
and U20867 (N_20867,N_19405,N_15230);
nor U20868 (N_20868,N_15596,N_16465);
xor U20869 (N_20869,N_17076,N_19811);
nand U20870 (N_20870,N_18054,N_15204);
nor U20871 (N_20871,N_18967,N_17075);
nand U20872 (N_20872,N_18914,N_15978);
or U20873 (N_20873,N_18079,N_16594);
nor U20874 (N_20874,N_15785,N_18426);
and U20875 (N_20875,N_15251,N_15288);
or U20876 (N_20876,N_18674,N_19514);
and U20877 (N_20877,N_17363,N_19162);
xnor U20878 (N_20878,N_18113,N_18900);
and U20879 (N_20879,N_17074,N_16352);
nand U20880 (N_20880,N_15799,N_19483);
nand U20881 (N_20881,N_16953,N_19482);
xnor U20882 (N_20882,N_16490,N_17906);
xor U20883 (N_20883,N_15128,N_17912);
nand U20884 (N_20884,N_19650,N_19784);
or U20885 (N_20885,N_16519,N_16703);
or U20886 (N_20886,N_18857,N_15630);
nand U20887 (N_20887,N_16861,N_17716);
or U20888 (N_20888,N_17478,N_18209);
nor U20889 (N_20889,N_15180,N_16752);
nor U20890 (N_20890,N_19656,N_19409);
nor U20891 (N_20891,N_17426,N_15472);
nor U20892 (N_20892,N_17008,N_18832);
or U20893 (N_20893,N_19317,N_16120);
nand U20894 (N_20894,N_17847,N_18611);
xor U20895 (N_20895,N_15085,N_15100);
and U20896 (N_20896,N_19557,N_16618);
xor U20897 (N_20897,N_16577,N_19197);
or U20898 (N_20898,N_18090,N_16826);
and U20899 (N_20899,N_15231,N_18203);
xnor U20900 (N_20900,N_18746,N_19054);
and U20901 (N_20901,N_16731,N_18685);
or U20902 (N_20902,N_17983,N_16489);
xnor U20903 (N_20903,N_17828,N_17482);
xnor U20904 (N_20904,N_19148,N_18501);
nand U20905 (N_20905,N_16840,N_16602);
and U20906 (N_20906,N_17325,N_18092);
nor U20907 (N_20907,N_19904,N_19681);
nor U20908 (N_20908,N_16129,N_15331);
and U20909 (N_20909,N_15766,N_19619);
and U20910 (N_20910,N_15643,N_15263);
xnor U20911 (N_20911,N_18304,N_15322);
and U20912 (N_20912,N_18487,N_16824);
xnor U20913 (N_20913,N_19441,N_19193);
or U20914 (N_20914,N_15662,N_16218);
xnor U20915 (N_20915,N_17179,N_18401);
and U20916 (N_20916,N_19694,N_17733);
and U20917 (N_20917,N_17890,N_18072);
and U20918 (N_20918,N_16892,N_19577);
nor U20919 (N_20919,N_17169,N_18929);
nand U20920 (N_20920,N_19075,N_18514);
or U20921 (N_20921,N_18874,N_17533);
or U20922 (N_20922,N_18810,N_18435);
and U20923 (N_20923,N_17158,N_15336);
xor U20924 (N_20924,N_19365,N_16160);
nand U20925 (N_20925,N_19999,N_15047);
or U20926 (N_20926,N_17052,N_16377);
nand U20927 (N_20927,N_17479,N_15589);
and U20928 (N_20928,N_18937,N_15292);
and U20929 (N_20929,N_16750,N_19816);
xnor U20930 (N_20930,N_18534,N_15279);
nand U20931 (N_20931,N_18554,N_16178);
or U20932 (N_20932,N_17013,N_19824);
and U20933 (N_20933,N_18251,N_17776);
and U20934 (N_20934,N_15477,N_18625);
nor U20935 (N_20935,N_15998,N_19319);
and U20936 (N_20936,N_17274,N_16418);
or U20937 (N_20937,N_19281,N_16162);
xor U20938 (N_20938,N_19592,N_18081);
nand U20939 (N_20939,N_17876,N_17237);
nand U20940 (N_20940,N_16349,N_18020);
or U20941 (N_20941,N_15748,N_19721);
nand U20942 (N_20942,N_15152,N_16015);
xnor U20943 (N_20943,N_16228,N_17922);
nand U20944 (N_20944,N_19239,N_16511);
xnor U20945 (N_20945,N_19746,N_19046);
xnor U20946 (N_20946,N_18108,N_16150);
or U20947 (N_20947,N_19593,N_18784);
nor U20948 (N_20948,N_15081,N_15843);
and U20949 (N_20949,N_16052,N_17762);
nor U20950 (N_20950,N_18605,N_16084);
nor U20951 (N_20951,N_18096,N_15262);
nor U20952 (N_20952,N_18292,N_18755);
nand U20953 (N_20953,N_17387,N_18029);
nand U20954 (N_20954,N_19629,N_18335);
or U20955 (N_20955,N_18350,N_18499);
nand U20956 (N_20956,N_15730,N_19720);
and U20957 (N_20957,N_17937,N_17632);
or U20958 (N_20958,N_16116,N_17512);
or U20959 (N_20959,N_17142,N_17376);
or U20960 (N_20960,N_19934,N_19088);
nand U20961 (N_20961,N_18850,N_15780);
and U20962 (N_20962,N_18538,N_17783);
nand U20963 (N_20963,N_15726,N_17195);
or U20964 (N_20964,N_18764,N_18727);
nor U20965 (N_20965,N_18129,N_17921);
nand U20966 (N_20966,N_17710,N_16226);
or U20967 (N_20967,N_17852,N_16549);
or U20968 (N_20968,N_17262,N_18439);
and U20969 (N_20969,N_16217,N_18529);
nand U20970 (N_20970,N_15005,N_19195);
nor U20971 (N_20971,N_17441,N_17199);
nand U20972 (N_20972,N_17178,N_15096);
or U20973 (N_20973,N_15467,N_16616);
xor U20974 (N_20974,N_16889,N_15925);
nand U20975 (N_20975,N_16710,N_18224);
nand U20976 (N_20976,N_16910,N_18576);
nor U20977 (N_20977,N_15795,N_16674);
nand U20978 (N_20978,N_16499,N_16171);
nand U20979 (N_20979,N_18502,N_15610);
and U20980 (N_20980,N_19427,N_16781);
xnor U20981 (N_20981,N_17448,N_17990);
nand U20982 (N_20982,N_19918,N_19524);
xnor U20983 (N_20983,N_19750,N_19649);
xor U20984 (N_20984,N_18702,N_19233);
nor U20985 (N_20985,N_15452,N_17337);
nor U20986 (N_20986,N_16906,N_19002);
and U20987 (N_20987,N_18946,N_16156);
nor U20988 (N_20988,N_15392,N_18822);
xor U20989 (N_20989,N_18364,N_15644);
nor U20990 (N_20990,N_16498,N_19893);
nor U20991 (N_20991,N_17869,N_15816);
nor U20992 (N_20992,N_19448,N_18651);
and U20993 (N_20993,N_15987,N_17065);
and U20994 (N_20994,N_15356,N_16045);
or U20995 (N_20995,N_15927,N_16508);
nor U20996 (N_20996,N_19308,N_18932);
or U20997 (N_20997,N_15386,N_18722);
or U20998 (N_20998,N_17756,N_17246);
nor U20999 (N_20999,N_16259,N_18815);
xor U21000 (N_21000,N_15243,N_17926);
nor U21001 (N_21001,N_15182,N_19313);
nand U21002 (N_21002,N_19916,N_15844);
or U21003 (N_21003,N_17739,N_17058);
or U21004 (N_21004,N_15623,N_19474);
and U21005 (N_21005,N_17800,N_18260);
xnor U21006 (N_21006,N_16996,N_17839);
nand U21007 (N_21007,N_18799,N_16065);
and U21008 (N_21008,N_19808,N_18772);
or U21009 (N_21009,N_17347,N_17768);
nand U21010 (N_21010,N_18979,N_17304);
nand U21011 (N_21011,N_18098,N_18028);
or U21012 (N_21012,N_19543,N_19662);
or U21013 (N_21013,N_19157,N_16992);
and U21014 (N_21014,N_17996,N_19079);
and U21015 (N_21015,N_18468,N_15498);
nand U21016 (N_21016,N_17480,N_17293);
nor U21017 (N_21017,N_16741,N_16442);
nand U21018 (N_21018,N_18473,N_16118);
or U21019 (N_21019,N_16590,N_19728);
nand U21020 (N_21020,N_18777,N_17171);
and U21021 (N_21021,N_18211,N_18549);
or U21022 (N_21022,N_19624,N_16950);
xnor U21023 (N_21023,N_15326,N_16253);
or U21024 (N_21024,N_15829,N_19125);
xnor U21025 (N_21025,N_19504,N_17527);
nand U21026 (N_21026,N_17094,N_15934);
xor U21027 (N_21027,N_17562,N_16532);
nor U21028 (N_21028,N_17675,N_15754);
or U21029 (N_21029,N_18504,N_17225);
or U21030 (N_21030,N_16641,N_19738);
or U21031 (N_21031,N_18150,N_19827);
or U21032 (N_21032,N_16320,N_16698);
or U21033 (N_21033,N_16799,N_18250);
and U21034 (N_21034,N_17851,N_17655);
nand U21035 (N_21035,N_16308,N_19035);
and U21036 (N_21036,N_16112,N_16130);
and U21037 (N_21037,N_15215,N_18982);
and U21038 (N_21038,N_16190,N_16009);
or U21039 (N_21039,N_16155,N_19223);
xnor U21040 (N_21040,N_16836,N_17806);
xnor U21041 (N_21041,N_19462,N_17729);
nand U21042 (N_21042,N_17888,N_19155);
nor U21043 (N_21043,N_18420,N_15391);
nand U21044 (N_21044,N_17404,N_19601);
nor U21045 (N_21045,N_17798,N_19367);
xnor U21046 (N_21046,N_19778,N_16684);
or U21047 (N_21047,N_15437,N_17464);
and U21048 (N_21048,N_18592,N_19660);
or U21049 (N_21049,N_15358,N_19767);
and U21050 (N_21050,N_18876,N_16786);
nor U21051 (N_21051,N_19235,N_15314);
or U21052 (N_21052,N_19345,N_18713);
or U21053 (N_21053,N_19745,N_15482);
and U21054 (N_21054,N_18334,N_19840);
xor U21055 (N_21055,N_16325,N_17498);
nand U21056 (N_21056,N_16575,N_19454);
nor U21057 (N_21057,N_17186,N_19118);
or U21058 (N_21058,N_19967,N_15439);
xor U21059 (N_21059,N_17088,N_16732);
nor U21060 (N_21060,N_17505,N_18200);
or U21061 (N_21061,N_17916,N_17850);
nor U21062 (N_21062,N_17871,N_15454);
nand U21063 (N_21063,N_19667,N_18486);
or U21064 (N_21064,N_16645,N_17969);
xor U21065 (N_21065,N_16000,N_17317);
nand U21066 (N_21066,N_18591,N_18119);
xor U21067 (N_21067,N_15546,N_18976);
nand U21068 (N_21068,N_15232,N_17245);
nand U21069 (N_21069,N_19341,N_15557);
nand U21070 (N_21070,N_18971,N_18167);
nand U21071 (N_21071,N_16738,N_16632);
and U21072 (N_21072,N_19696,N_18698);
nand U21073 (N_21073,N_17287,N_17730);
nand U21074 (N_21074,N_15649,N_17695);
and U21075 (N_21075,N_18235,N_19378);
nor U21076 (N_21076,N_16185,N_15599);
nand U21077 (N_21077,N_19050,N_17003);
and U21078 (N_21078,N_16495,N_18302);
nand U21079 (N_21079,N_19116,N_19331);
nand U21080 (N_21080,N_19530,N_18498);
nand U21081 (N_21081,N_18834,N_16691);
xnor U21082 (N_21082,N_15984,N_17312);
nor U21083 (N_21083,N_18294,N_17534);
nand U21084 (N_21084,N_19546,N_18497);
or U21085 (N_21085,N_19468,N_19941);
nor U21086 (N_21086,N_15890,N_15131);
xnor U21087 (N_21087,N_16654,N_18077);
xor U21088 (N_21088,N_19292,N_15308);
or U21089 (N_21089,N_17315,N_15950);
nor U21090 (N_21090,N_17265,N_18102);
and U21091 (N_21091,N_19793,N_18262);
nor U21092 (N_21092,N_17253,N_19937);
or U21093 (N_21093,N_16315,N_15237);
nand U21094 (N_21094,N_15637,N_19971);
and U21095 (N_21095,N_16341,N_17011);
xor U21096 (N_21096,N_15769,N_15529);
xor U21097 (N_21097,N_19594,N_19329);
or U21098 (N_21098,N_16078,N_15912);
or U21099 (N_21099,N_19929,N_17280);
nor U21100 (N_21100,N_17255,N_15286);
nand U21101 (N_21101,N_16585,N_19905);
nor U21102 (N_21102,N_18984,N_16896);
or U21103 (N_21103,N_15870,N_15685);
xor U21104 (N_21104,N_18928,N_19881);
or U21105 (N_21105,N_17982,N_17559);
nand U21106 (N_21106,N_16566,N_16278);
nor U21107 (N_21107,N_19568,N_19114);
nand U21108 (N_21108,N_17579,N_19602);
nor U21109 (N_21109,N_16110,N_17184);
nand U21110 (N_21110,N_16236,N_16798);
and U21111 (N_21111,N_17326,N_16658);
xor U21112 (N_21112,N_15951,N_18153);
xor U21113 (N_21113,N_18567,N_17016);
and U21114 (N_21114,N_16957,N_16146);
or U21115 (N_21115,N_19930,N_18895);
xnor U21116 (N_21116,N_18349,N_16653);
nand U21117 (N_21117,N_16509,N_17156);
nand U21118 (N_21118,N_15086,N_16961);
nor U21119 (N_21119,N_19977,N_17454);
xnor U21120 (N_21120,N_17824,N_17486);
and U21121 (N_21121,N_18463,N_18676);
or U21122 (N_21122,N_16245,N_15575);
nand U21123 (N_21123,N_15185,N_18144);
nor U21124 (N_21124,N_15269,N_16437);
nor U21125 (N_21125,N_19903,N_19812);
nor U21126 (N_21126,N_15294,N_16541);
and U21127 (N_21127,N_19898,N_17833);
or U21128 (N_21128,N_18949,N_18124);
nor U21129 (N_21129,N_15573,N_15371);
xor U21130 (N_21130,N_15786,N_15563);
and U21131 (N_21131,N_19158,N_18099);
nand U21132 (N_21132,N_18697,N_17405);
nand U21133 (N_21133,N_15845,N_18046);
xnor U21134 (N_21134,N_18170,N_17266);
nor U21135 (N_21135,N_17476,N_17368);
xnor U21136 (N_21136,N_15953,N_19326);
and U21137 (N_21137,N_18136,N_19853);
or U21138 (N_21138,N_16551,N_17991);
nor U21139 (N_21139,N_16436,N_15931);
nor U21140 (N_21140,N_18616,N_19422);
and U21141 (N_21141,N_15438,N_18145);
nor U21142 (N_21142,N_15767,N_17818);
nor U21143 (N_21143,N_19640,N_19722);
nor U21144 (N_21144,N_16154,N_15092);
nor U21145 (N_21145,N_19172,N_18742);
xnor U21146 (N_21146,N_16833,N_15399);
nand U21147 (N_21147,N_16977,N_17819);
nand U21148 (N_21148,N_16941,N_19500);
xnor U21149 (N_21149,N_18273,N_15321);
nor U21150 (N_21150,N_15757,N_15388);
nor U21151 (N_21151,N_18631,N_18083);
or U21152 (N_21152,N_16414,N_19071);
nor U21153 (N_21153,N_15902,N_16460);
and U21154 (N_21154,N_16784,N_16373);
or U21155 (N_21155,N_18373,N_17010);
and U21156 (N_21156,N_16967,N_15518);
nor U21157 (N_21157,N_17121,N_19983);
and U21158 (N_21158,N_17489,N_16180);
and U21159 (N_21159,N_17832,N_18479);
nand U21160 (N_21160,N_19673,N_18396);
nor U21161 (N_21161,N_17153,N_15873);
nor U21162 (N_21162,N_18846,N_15233);
xor U21163 (N_21163,N_19821,N_17122);
and U21164 (N_21164,N_17616,N_18219);
or U21165 (N_21165,N_18289,N_17019);
and U21166 (N_21166,N_17215,N_18628);
xnor U21167 (N_21167,N_17777,N_15393);
and U21168 (N_21168,N_16008,N_15601);
nand U21169 (N_21169,N_17881,N_18974);
xor U21170 (N_21170,N_19956,N_19943);
or U21171 (N_21171,N_15058,N_19867);
xnor U21172 (N_21172,N_19851,N_19900);
xnor U21173 (N_21173,N_18562,N_18415);
nand U21174 (N_21174,N_18893,N_15683);
or U21175 (N_21175,N_19452,N_16726);
nor U21176 (N_21176,N_15357,N_17160);
xor U21177 (N_21177,N_19421,N_19886);
or U21178 (N_21178,N_19255,N_17595);
and U21179 (N_21179,N_17797,N_18564);
nand U21180 (N_21180,N_15028,N_19675);
and U21181 (N_21181,N_18572,N_17272);
or U21182 (N_21182,N_19570,N_16393);
xnor U21183 (N_21183,N_16247,N_16363);
nand U21184 (N_21184,N_16068,N_15349);
and U21185 (N_21185,N_19418,N_16912);
nand U21186 (N_21186,N_16105,N_19719);
xnor U21187 (N_21187,N_16222,N_18642);
and U21188 (N_21188,N_17950,N_16039);
and U21189 (N_21189,N_16725,N_16981);
or U21190 (N_21190,N_17053,N_17218);
and U21191 (N_21191,N_19875,N_15268);
nor U21192 (N_21192,N_17853,N_15663);
and U21193 (N_21193,N_15813,N_17660);
and U21194 (N_21194,N_16737,N_18677);
or U21195 (N_21195,N_17727,N_15226);
or U21196 (N_21196,N_16361,N_16920);
or U21197 (N_21197,N_19307,N_16797);
nor U21198 (N_21198,N_16017,N_16697);
xnor U21199 (N_21199,N_15718,N_18166);
and U21200 (N_21200,N_18708,N_18813);
and U21201 (N_21201,N_15210,N_18268);
xnor U21202 (N_21202,N_18785,N_17462);
and U21203 (N_21203,N_18536,N_17018);
or U21204 (N_21204,N_19450,N_17176);
nor U21205 (N_21205,N_17344,N_17841);
nand U21206 (N_21206,N_19022,N_18253);
nor U21207 (N_21207,N_19412,N_17196);
or U21208 (N_21208,N_15993,N_18060);
and U21209 (N_21209,N_18151,N_19297);
xnor U21210 (N_21210,N_18115,N_18394);
xor U21211 (N_21211,N_18086,N_15181);
and U21212 (N_21212,N_17110,N_16769);
nand U21213 (N_21213,N_19607,N_15749);
xor U21214 (N_21214,N_15853,N_16595);
nand U21215 (N_21215,N_16686,N_16959);
or U21216 (N_21216,N_17764,N_19911);
and U21217 (N_21217,N_15690,N_16058);
xnor U21218 (N_21218,N_15833,N_15411);
nor U21219 (N_21219,N_16074,N_19218);
or U21220 (N_21220,N_15548,N_19225);
xor U21221 (N_21221,N_18135,N_17789);
or U21222 (N_21222,N_15372,N_15798);
xnor U21223 (N_21223,N_15922,N_17717);
xor U21224 (N_21224,N_19716,N_17781);
and U21225 (N_21225,N_19953,N_18733);
or U21226 (N_21226,N_16630,N_18171);
xnor U21227 (N_21227,N_16087,N_17976);
nor U21228 (N_21228,N_17792,N_19464);
xor U21229 (N_21229,N_17651,N_16646);
nor U21230 (N_21230,N_16792,N_19343);
nor U21231 (N_21231,N_16517,N_18695);
or U21232 (N_21232,N_18838,N_16136);
and U21233 (N_21233,N_15384,N_18234);
xnor U21234 (N_21234,N_16626,N_18133);
nor U21235 (N_21235,N_15376,N_18267);
nand U21236 (N_21236,N_15307,N_16946);
nor U21237 (N_21237,N_16877,N_15789);
and U21238 (N_21238,N_18973,N_15583);
xor U21239 (N_21239,N_19539,N_16864);
or U21240 (N_21240,N_16275,N_18104);
or U21241 (N_21241,N_15493,N_19760);
nand U21242 (N_21242,N_17043,N_17295);
or U21243 (N_21243,N_19786,N_16768);
xor U21244 (N_21244,N_18191,N_18948);
and U21245 (N_21245,N_15888,N_17617);
nor U21246 (N_21246,N_18699,N_17148);
and U21247 (N_21247,N_18327,N_18693);
or U21248 (N_21248,N_16745,N_18281);
or U21249 (N_21249,N_16537,N_15898);
xor U21250 (N_21250,N_18126,N_18745);
nor U21251 (N_21251,N_15907,N_16706);
and U21252 (N_21252,N_19372,N_19779);
nand U21253 (N_21253,N_17607,N_16359);
nor U21254 (N_21254,N_17935,N_16735);
or U21255 (N_21255,N_16239,N_19700);
nand U21256 (N_21256,N_18033,N_17809);
nand U21257 (N_21257,N_16927,N_15304);
xor U21258 (N_21258,N_17746,N_18606);
and U21259 (N_21259,N_19356,N_18759);
nand U21260 (N_21260,N_16554,N_15107);
and U21261 (N_21261,N_16419,N_19083);
and U21262 (N_21262,N_19410,N_19243);
nand U21263 (N_21263,N_18851,N_16709);
xor U21264 (N_21264,N_19032,N_19755);
xor U21265 (N_21265,N_17957,N_15999);
or U21266 (N_21266,N_18747,N_16552);
or U21267 (N_21267,N_19141,N_18019);
xor U21268 (N_21268,N_16173,N_19734);
and U21269 (N_21269,N_18798,N_18154);
nor U21270 (N_21270,N_17669,N_15582);
nor U21271 (N_21271,N_15420,N_17394);
nand U21272 (N_21272,N_17700,N_19682);
xnor U21273 (N_21273,N_19932,N_16979);
xor U21274 (N_21274,N_16962,N_17692);
nor U21275 (N_21275,N_17997,N_15560);
nor U21276 (N_21276,N_15859,N_17600);
and U21277 (N_21277,N_18550,N_17586);
nand U21278 (N_21278,N_17722,N_19339);
nor U21279 (N_21279,N_16885,N_16553);
nor U21280 (N_21280,N_18735,N_17321);
nand U21281 (N_21281,N_15486,N_19033);
xnor U21282 (N_21282,N_17679,N_19846);
and U21283 (N_21283,N_16858,N_17749);
and U21284 (N_21284,N_18645,N_15990);
nor U21285 (N_21285,N_18197,N_16723);
xnor U21286 (N_21286,N_16386,N_18614);
nor U21287 (N_21287,N_16839,N_16099);
nand U21288 (N_21288,N_16900,N_19612);
or U21289 (N_21289,N_17883,N_15787);
nand U21290 (N_21290,N_17430,N_15923);
or U21291 (N_21291,N_15382,N_15580);
xor U21292 (N_21292,N_15046,N_19466);
nor U21293 (N_21293,N_15335,N_18704);
xor U21294 (N_21294,N_16082,N_16678);
xnor U21295 (N_21295,N_17524,N_16771);
and U21296 (N_21296,N_18321,N_16583);
xor U21297 (N_21297,N_19723,N_18954);
nand U21298 (N_21298,N_19376,N_15436);
or U21299 (N_21299,N_18249,N_16970);
or U21300 (N_21300,N_16223,N_15044);
xnor U21301 (N_21301,N_17168,N_18076);
nor U21302 (N_21302,N_18842,N_18032);
nand U21303 (N_21303,N_18477,N_16813);
nor U21304 (N_21304,N_17463,N_15246);
xnor U21305 (N_21305,N_17802,N_19473);
and U21306 (N_21306,N_15746,N_15334);
nor U21307 (N_21307,N_19416,N_18419);
nand U21308 (N_21308,N_17986,N_16179);
xor U21309 (N_21309,N_19445,N_16181);
or U21310 (N_21310,N_19000,N_19081);
or U21311 (N_21311,N_17341,N_16568);
nor U21312 (N_21312,N_16765,N_19097);
or U21313 (N_21313,N_17670,N_19509);
nor U21314 (N_21314,N_19091,N_16716);
nor U21315 (N_21315,N_18856,N_17980);
nand U21316 (N_21316,N_18970,N_18717);
and U21317 (N_21317,N_19708,N_19023);
nor U21318 (N_21318,N_15234,N_16561);
and U21319 (N_21319,N_16573,N_16255);
xor U21320 (N_21320,N_17621,N_17987);
or U21321 (N_21321,N_17252,N_17642);
nor U21322 (N_21322,N_19496,N_17307);
nor U21323 (N_21323,N_19417,N_17752);
nor U21324 (N_21324,N_15693,N_18085);
nand U21325 (N_21325,N_15140,N_19717);
nand U21326 (N_21326,N_16269,N_15574);
or U21327 (N_21327,N_16306,N_19463);
and U21328 (N_21328,N_16862,N_18073);
and U21329 (N_21329,N_18271,N_15860);
nor U21330 (N_21330,N_17089,N_18885);
xnor U21331 (N_21331,N_18966,N_18997);
xor U21332 (N_21332,N_15470,N_15060);
nand U21333 (N_21333,N_16720,N_16421);
or U21334 (N_21334,N_17189,N_15110);
or U21335 (N_21335,N_18744,N_19506);
and U21336 (N_21336,N_16803,N_18345);
nor U21337 (N_21337,N_15572,N_16633);
or U21338 (N_21338,N_18907,N_18897);
nor U21339 (N_21339,N_18193,N_19288);
or U21340 (N_21340,N_16397,N_16733);
xor U21341 (N_21341,N_17338,N_19529);
or U21342 (N_21342,N_15395,N_19759);
and U21343 (N_21343,N_19131,N_17726);
nand U21344 (N_21344,N_19984,N_19978);
nor U21345 (N_21345,N_16578,N_15284);
nand U21346 (N_21346,N_17612,N_18743);
nor U21347 (N_21347,N_17519,N_16295);
nor U21348 (N_21348,N_18105,N_17348);
and U21349 (N_21349,N_19123,N_15531);
nand U21350 (N_21350,N_19749,N_15791);
or U21351 (N_21351,N_19995,N_18223);
nand U21352 (N_21352,N_19519,N_17095);
or U21353 (N_21353,N_17641,N_19208);
nand U21354 (N_21354,N_19902,N_19954);
nand U21355 (N_21355,N_19334,N_15061);
nand U21356 (N_21356,N_17686,N_19804);
nor U21357 (N_21357,N_19051,N_15616);
or U21358 (N_21358,N_15150,N_15133);
xor U21359 (N_21359,N_16338,N_18338);
nor U21360 (N_21360,N_17545,N_18261);
or U21361 (N_21361,N_19829,N_17308);
xnor U21362 (N_21362,N_19105,N_16153);
or U21363 (N_21363,N_19451,N_17137);
or U21364 (N_21364,N_19766,N_19545);
nand U21365 (N_21365,N_17029,N_16749);
nor U21366 (N_21366,N_17870,N_16748);
nor U21367 (N_21367,N_17537,N_17082);
nand U21368 (N_21368,N_15806,N_17662);
xor U21369 (N_21369,N_16708,N_18598);
or U21370 (N_21370,N_16898,N_15645);
or U21371 (N_21371,N_15507,N_16973);
nand U21372 (N_21372,N_15976,N_18797);
or U21373 (N_21373,N_19142,N_17130);
and U21374 (N_21374,N_17497,N_17367);
and U21375 (N_21375,N_19010,N_18385);
xnor U21376 (N_21376,N_15030,N_15608);
xnor U21377 (N_21377,N_15238,N_17676);
or U21378 (N_21378,N_17009,N_15173);
or U21379 (N_21379,N_15512,N_16870);
and U21380 (N_21380,N_17770,N_18429);
nor U21381 (N_21381,N_17970,N_18058);
nand U21382 (N_21382,N_15008,N_18962);
or U21383 (N_21383,N_19016,N_15297);
or U21384 (N_21384,N_18272,N_17674);
nand U21385 (N_21385,N_17290,N_15455);
xor U21386 (N_21386,N_15640,N_17213);
or U21387 (N_21387,N_18942,N_15775);
and U21388 (N_21388,N_16075,N_16392);
and U21389 (N_21389,N_18016,N_17305);
and U21390 (N_21390,N_19167,N_17568);
nand U21391 (N_21391,N_19533,N_19360);
and U21392 (N_21392,N_19147,N_15010);
and U21393 (N_21393,N_15456,N_19247);
nor U21394 (N_21394,N_18431,N_15659);
and U21395 (N_21395,N_17427,N_17096);
or U21396 (N_21396,N_16746,N_17230);
and U21397 (N_21397,N_19005,N_16563);
nor U21398 (N_21398,N_18094,N_17172);
nor U21399 (N_21399,N_16071,N_19503);
and U21400 (N_21400,N_17459,N_18201);
xor U21401 (N_21401,N_17723,N_16680);
xor U21402 (N_21402,N_19110,N_17037);
nand U21403 (N_21403,N_18024,N_16719);
or U21404 (N_21404,N_17320,N_18958);
xnor U21405 (N_21405,N_17827,N_17596);
nand U21406 (N_21406,N_17892,N_16214);
and U21407 (N_21407,N_15306,N_15037);
and U21408 (N_21408,N_19538,N_18286);
and U21409 (N_21409,N_18656,N_18707);
nor U21410 (N_21410,N_16072,N_16496);
nand U21411 (N_21411,N_15569,N_18700);
nor U21412 (N_21412,N_16873,N_18714);
or U21413 (N_21413,N_18134,N_18213);
nand U21414 (N_21414,N_18630,N_18386);
xnor U21415 (N_21415,N_19564,N_19135);
or U21416 (N_21416,N_17129,N_15351);
nand U21417 (N_21417,N_17481,N_16220);
or U21418 (N_21418,N_16917,N_18963);
nor U21419 (N_21419,N_19053,N_18649);
or U21420 (N_21420,N_15701,N_18194);
and U21421 (N_21421,N_15842,N_16985);
or U21422 (N_21422,N_16766,N_15918);
xor U21423 (N_21423,N_15839,N_19563);
xnor U21424 (N_21424,N_18577,N_16690);
nor U21425 (N_21425,N_15660,N_18884);
or U21426 (N_21426,N_15172,N_18210);
nand U21427 (N_21427,N_15973,N_16485);
or U21428 (N_21428,N_17309,N_19511);
and U21429 (N_21429,N_17396,N_16091);
nor U21430 (N_21430,N_17445,N_19727);
nand U21431 (N_21431,N_16343,N_16391);
or U21432 (N_21432,N_15497,N_18729);
nor U21433 (N_21433,N_15344,N_16856);
nand U21434 (N_21434,N_17118,N_19970);
nor U21435 (N_21435,N_15768,N_15141);
nor U21436 (N_21436,N_18819,N_16935);
and U21437 (N_21437,N_17269,N_18446);
nor U21438 (N_21438,N_17433,N_18977);
nand U21439 (N_21439,N_17713,N_16027);
nand U21440 (N_21440,N_16965,N_19887);
xor U21441 (N_21441,N_15668,N_15528);
nor U21442 (N_21442,N_16268,N_17062);
and U21443 (N_21443,N_18505,N_19833);
or U21444 (N_21444,N_18912,N_18216);
nand U21445 (N_21445,N_15543,N_18760);
nand U21446 (N_21446,N_15566,N_15742);
xnor U21447 (N_21447,N_19805,N_16867);
xor U21448 (N_21448,N_15310,N_18887);
and U21449 (N_21449,N_19137,N_17574);
nor U21450 (N_21450,N_15112,N_15462);
nor U21451 (N_21451,N_15530,N_17451);
xnor U21452 (N_21452,N_16681,N_15519);
or U21453 (N_21453,N_15631,N_15398);
or U21454 (N_21454,N_19467,N_17801);
nand U21455 (N_21455,N_15943,N_18627);
nor U21456 (N_21456,N_17453,N_19198);
and U21457 (N_21457,N_17420,N_15721);
nor U21458 (N_21458,N_17899,N_17223);
or U21459 (N_21459,N_19354,N_15419);
and U21460 (N_21460,N_15505,N_18992);
nand U21461 (N_21461,N_15494,N_15989);
and U21462 (N_21462,N_19668,N_15361);
and U21463 (N_21463,N_18488,N_18513);
nand U21464 (N_21464,N_16422,N_17501);
nor U21465 (N_21465,N_17456,N_18485);
xor U21466 (N_21466,N_18823,N_19258);
and U21467 (N_21467,N_19521,N_17114);
and U21468 (N_21468,N_17928,N_17704);
nor U21469 (N_21469,N_17233,N_15379);
nor U21470 (N_21470,N_15479,N_15516);
or U21471 (N_21471,N_18779,N_18849);
nor U21472 (N_21472,N_19620,N_18829);
or U21473 (N_21473,N_19173,N_16492);
or U21474 (N_21474,N_15967,N_15607);
nor U21475 (N_21475,N_18241,N_18313);
nor U21476 (N_21476,N_16137,N_18106);
nor U21477 (N_21477,N_18655,N_18035);
xnor U21478 (N_21478,N_17061,N_16448);
nor U21479 (N_21479,N_16466,N_18568);
xor U21480 (N_21480,N_16234,N_17416);
nand U21481 (N_21481,N_15674,N_18517);
or U21482 (N_21482,N_15964,N_15151);
and U21483 (N_21483,N_15480,N_18725);
nand U21484 (N_21484,N_19591,N_17182);
nand U21485 (N_21485,N_18416,N_19817);
or U21486 (N_21486,N_18595,N_16370);
nand U21487 (N_21487,N_15614,N_17180);
nand U21488 (N_21488,N_18366,N_15448);
or U21489 (N_21489,N_18867,N_17438);
nor U21490 (N_21490,N_16412,N_16430);
or U21491 (N_21491,N_19732,N_17400);
or U21492 (N_21492,N_19014,N_16240);
and U21493 (N_21493,N_16115,N_17115);
and U21494 (N_21494,N_18730,N_15169);
nor U21495 (N_21495,N_16608,N_17816);
and U21496 (N_21496,N_17264,N_18190);
and U21497 (N_21497,N_17619,N_18177);
xor U21498 (N_21498,N_18808,N_17965);
or U21499 (N_21499,N_15588,N_16001);
nor U21500 (N_21500,N_17452,N_17257);
and U21501 (N_21501,N_17350,N_19138);
xor U21502 (N_21502,N_18026,N_19780);
nor U21503 (N_21503,N_19680,N_16170);
xor U21504 (N_21504,N_17242,N_19801);
and U21505 (N_21505,N_17956,N_19436);
nor U21506 (N_21506,N_18320,N_16206);
and U21507 (N_21507,N_19587,N_15653);
xnor U21508 (N_21508,N_16795,N_17649);
and U21509 (N_21509,N_17864,N_18734);
xor U21510 (N_21510,N_16077,N_17030);
nand U21511 (N_21511,N_19698,N_18972);
or U21512 (N_21512,N_15424,N_17049);
or U21513 (N_21513,N_18163,N_18771);
nand U21514 (N_21514,N_18915,N_15551);
xor U21515 (N_21515,N_19040,N_16513);
xor U21516 (N_21516,N_18644,N_19260);
xor U21517 (N_21517,N_19860,N_19921);
nor U21518 (N_21518,N_19209,N_19702);
nand U21519 (N_21519,N_19068,N_17377);
nand U21520 (N_21520,N_19161,N_18015);
nor U21521 (N_21521,N_18712,N_19674);
nor U21522 (N_21522,N_17656,N_19431);
and U21523 (N_21523,N_15432,N_16013);
nor U21524 (N_21524,N_17763,N_16635);
or U21525 (N_21525,N_17877,N_15165);
xnor U21526 (N_21526,N_18097,N_19037);
xnor U21527 (N_21527,N_18687,N_15103);
nand U21528 (N_21528,N_18461,N_19810);
xor U21529 (N_21529,N_19379,N_19314);
nand U21530 (N_21530,N_16314,N_18080);
nor U21531 (N_21531,N_17141,N_19910);
xnor U21532 (N_21532,N_19392,N_15995);
nand U21533 (N_21533,N_18012,N_16037);
and U21534 (N_21534,N_15857,N_15542);
nand U21535 (N_21535,N_18581,N_15309);
nor U21536 (N_21536,N_17402,N_15116);
nor U21537 (N_21537,N_17815,N_17333);
or U21538 (N_21538,N_15168,N_18607);
nand U21539 (N_21539,N_17063,N_15639);
xor U21540 (N_21540,N_16417,N_19571);
nor U21541 (N_21541,N_16601,N_15034);
and U21542 (N_21542,N_19030,N_15661);
nand U21543 (N_21543,N_18728,N_18854);
xor U21544 (N_21544,N_15031,N_17098);
nor U21545 (N_21545,N_18101,N_17913);
nor U21546 (N_21546,N_19012,N_15134);
xor U21547 (N_21547,N_17289,N_15166);
or U21548 (N_21548,N_17022,N_16125);
xnor U21549 (N_21549,N_18629,N_15979);
or U21550 (N_21550,N_19972,N_15178);
or U21551 (N_21551,N_19994,N_15350);
xnor U21552 (N_21552,N_16614,N_16199);
nand U21553 (N_21553,N_16172,N_19711);
nor U21554 (N_21554,N_17699,N_19735);
xor U21555 (N_21555,N_15684,N_15823);
nand U21556 (N_21556,N_16038,N_19215);
and U21557 (N_21557,N_19230,N_17258);
nand U21558 (N_21558,N_19781,N_16423);
nor U21559 (N_21559,N_18855,N_19385);
nor U21560 (N_21560,N_15997,N_15711);
xor U21561 (N_21561,N_16100,N_15186);
or U21562 (N_21562,N_16305,N_15241);
xor U21563 (N_21563,N_17384,N_16693);
and U21564 (N_21564,N_16664,N_19371);
nor U21565 (N_21565,N_18658,N_18114);
and U21566 (N_21566,N_15773,N_16288);
xor U21567 (N_21567,N_16405,N_15192);
nand U21568 (N_21568,N_17285,N_17127);
or U21569 (N_21569,N_19952,N_19858);
nor U21570 (N_21570,N_16303,N_17144);
or U21571 (N_21571,N_15390,N_17056);
and U21572 (N_21572,N_16474,N_19585);
or U21573 (N_21573,N_19574,N_16778);
or U21574 (N_21574,N_15956,N_17665);
or U21575 (N_21575,N_16073,N_15198);
xnor U21576 (N_21576,N_19396,N_17653);
or U21577 (N_21577,N_18617,N_17343);
nand U21578 (N_21578,N_16049,N_18244);
and U21579 (N_21579,N_19129,N_15834);
nor U21580 (N_21580,N_19834,N_15353);
and U21581 (N_21581,N_15271,N_19815);
nor U21582 (N_21582,N_16159,N_15067);
nand U21583 (N_21583,N_16243,N_18924);
xnor U21584 (N_21584,N_18300,N_19062);
nand U21585 (N_21585,N_17683,N_15914);
nor U21586 (N_21586,N_17389,N_18988);
nand U21587 (N_21587,N_15396,N_16515);
or U21588 (N_21588,N_16505,N_15811);
and U21589 (N_21589,N_15345,N_16476);
nand U21590 (N_21590,N_15135,N_17190);
or U21591 (N_21591,N_19528,N_18437);
or U21592 (N_21592,N_16580,N_15808);
nor U21593 (N_21593,N_17563,N_17103);
xnor U21594 (N_21594,N_19383,N_19604);
nor U21595 (N_21595,N_19617,N_19055);
xor U21596 (N_21596,N_18377,N_16855);
and U21597 (N_21597,N_19976,N_15772);
nand U21598 (N_21598,N_16040,N_16031);
nor U21599 (N_21599,N_18684,N_19686);
nand U21600 (N_21600,N_16139,N_15045);
or U21601 (N_21601,N_16639,N_15634);
and U21602 (N_21602,N_17694,N_19638);
nand U21603 (N_21603,N_17772,N_16404);
nand U21604 (N_21604,N_15403,N_19189);
nand U21605 (N_21605,N_18953,N_17736);
and U21606 (N_21606,N_16387,N_15002);
or U21607 (N_21607,N_15317,N_19328);
or U21608 (N_21608,N_17504,N_17588);
nor U21609 (N_21609,N_19477,N_16416);
or U21610 (N_21610,N_17677,N_19066);
or U21611 (N_21611,N_16056,N_15430);
or U21612 (N_21612,N_19042,N_15278);
and U21613 (N_21613,N_18061,N_17523);
or U21614 (N_21614,N_19770,N_17804);
and U21615 (N_21615,N_17286,N_16238);
nor U21616 (N_21616,N_15119,N_19802);
xor U21617 (N_21617,N_18283,N_19425);
nor U21618 (N_21618,N_17927,N_17278);
nand U21619 (N_21619,N_17863,N_19370);
or U21620 (N_21620,N_15179,N_18199);
nand U21621 (N_21621,N_17829,N_18095);
xor U21622 (N_21622,N_16982,N_18740);
nand U21623 (N_21623,N_17334,N_16696);
and U21624 (N_21624,N_17542,N_17979);
nand U21625 (N_21625,N_16428,N_19108);
nor U21626 (N_21626,N_16473,N_19523);
nand U21627 (N_21627,N_19004,N_17092);
xor U21628 (N_21628,N_17031,N_18214);
and U21629 (N_21629,N_15267,N_16335);
xor U21630 (N_21630,N_16231,N_17369);
nand U21631 (N_21631,N_16924,N_15600);
nor U21632 (N_21632,N_17875,N_16995);
nor U21633 (N_21633,N_19309,N_16025);
nor U21634 (N_21634,N_16721,N_19127);
or U21635 (N_21635,N_18812,N_15883);
nand U21636 (N_21636,N_19707,N_15713);
or U21637 (N_21637,N_17961,N_17193);
xor U21638 (N_21638,N_15219,N_19113);
or U21639 (N_21639,N_16292,N_19476);
xor U21640 (N_21640,N_17838,N_16734);
and U21641 (N_21641,N_19159,N_15728);
xnor U21642 (N_21642,N_18480,N_17681);
nor U21643 (N_21643,N_16371,N_19950);
and U21644 (N_21644,N_16457,N_16167);
and U21645 (N_21645,N_15118,N_19201);
nand U21646 (N_21646,N_17410,N_19690);
xnor U21647 (N_21647,N_17647,N_18422);
nand U21648 (N_21648,N_16095,N_15108);
nor U21649 (N_21649,N_19160,N_18247);
nand U21650 (N_21650,N_19219,N_16449);
nand U21651 (N_21651,N_15975,N_19133);
or U21652 (N_21652,N_17585,N_17488);
and U21653 (N_21653,N_18252,N_16888);
and U21654 (N_21654,N_16883,N_17078);
nand U21655 (N_21655,N_18603,N_18993);
xor U21656 (N_21656,N_18579,N_16604);
and U21657 (N_21657,N_16321,N_15595);
or U21658 (N_21658,N_16462,N_19634);
and U21659 (N_21659,N_19942,N_17067);
xor U21660 (N_21660,N_17867,N_18400);
nand U21661 (N_21661,N_16830,N_19676);
and U21662 (N_21662,N_19647,N_16665);
and U21663 (N_21663,N_17383,N_16628);
and U21664 (N_21664,N_19731,N_15881);
nor U21665 (N_21665,N_18800,N_15736);
nand U21666 (N_21666,N_15442,N_15488);
and U21667 (N_21667,N_19204,N_17587);
xnor U21668 (N_21668,N_16344,N_18881);
xor U21669 (N_21669,N_18921,N_15779);
nor U21670 (N_21670,N_17719,N_19661);
or U21671 (N_21671,N_15874,N_18142);
and U21672 (N_21672,N_16999,N_17550);
nand U21673 (N_21673,N_17105,N_19207);
xor U21674 (N_21674,N_17958,N_19576);
xnor U21675 (N_21675,N_17657,N_19914);
and U21676 (N_21676,N_15054,N_19752);
xnor U21677 (N_21677,N_17920,N_17779);
or U21678 (N_21678,N_17068,N_17211);
xnor U21679 (N_21679,N_18139,N_19015);
and U21680 (N_21680,N_17023,N_15915);
nor U21681 (N_21681,N_19411,N_17931);
nand U21682 (N_21682,N_15368,N_15836);
and U21683 (N_21683,N_18265,N_19927);
and U21684 (N_21684,N_19830,N_19552);
and U21685 (N_21685,N_18903,N_18548);
xor U21686 (N_21686,N_17424,N_18184);
or U21687 (N_21687,N_19569,N_18931);
nor U21688 (N_21688,N_15846,N_16453);
and U21689 (N_21689,N_18408,N_18847);
xor U21690 (N_21690,N_17359,N_19456);
and U21691 (N_21691,N_19086,N_17993);
xor U21692 (N_21692,N_19525,N_18183);
or U21693 (N_21693,N_19825,N_17104);
and U21694 (N_21694,N_15145,N_16567);
nand U21695 (N_21695,N_16192,N_19666);
nand U21696 (N_21696,N_19579,N_16570);
or U21697 (N_21697,N_18904,N_17546);
xor U21698 (N_21698,N_16131,N_16663);
nand U21699 (N_21699,N_15213,N_15913);
or U21700 (N_21700,N_16510,N_18052);
and U21701 (N_21701,N_19400,N_17702);
nand U21702 (N_21702,N_17159,N_18442);
nor U21703 (N_21703,N_19791,N_19501);
or U21704 (N_21704,N_18939,N_18188);
and U21705 (N_21705,N_16122,N_17087);
or U21706 (N_21706,N_18315,N_18264);
nor U21707 (N_21707,N_18553,N_18736);
xnor U21708 (N_21708,N_18860,N_18531);
or U21709 (N_21709,N_15453,N_15017);
and U21710 (N_21710,N_15700,N_19398);
and U21711 (N_21711,N_19575,N_17654);
xnor U21712 (N_21712,N_18344,N_18270);
nor U21713 (N_21713,N_16312,N_15571);
xnor U21714 (N_21714,N_18923,N_18318);
nand U21715 (N_21715,N_19094,N_15260);
nand U21716 (N_21716,N_17985,N_15089);
xnor U21717 (N_21717,N_17281,N_19862);
nor U21718 (N_21718,N_17484,N_15686);
nor U21719 (N_21719,N_16914,N_15066);
and U21720 (N_21720,N_16773,N_17124);
or U21721 (N_21721,N_16904,N_16029);
nor U21722 (N_21722,N_16174,N_15618);
nand U21723 (N_21723,N_17720,N_17784);
xnor U21724 (N_21724,N_15694,N_19861);
xnor U21725 (N_21725,N_18069,N_19899);
nand U21726 (N_21726,N_18120,N_19008);
or U21727 (N_21727,N_16277,N_18886);
xnor U21728 (N_21728,N_18541,N_19623);
xor U21729 (N_21729,N_15632,N_16687);
nor U21730 (N_21730,N_17330,N_15617);
nand U21731 (N_21731,N_16360,N_18371);
nand U21732 (N_21732,N_18221,N_15765);
xnor U21733 (N_21733,N_15849,N_19472);
and U21734 (N_21734,N_18383,N_16035);
and U21735 (N_21735,N_15776,N_17303);
nor U21736 (N_21736,N_19512,N_19178);
xnor U21737 (N_21737,N_18845,N_16718);
nor U21738 (N_21738,N_18673,N_17608);
nor U21739 (N_21739,N_15212,N_15446);
nor U21740 (N_21740,N_16947,N_16905);
nand U21741 (N_21741,N_18574,N_17518);
xor U21742 (N_21742,N_16929,N_17581);
xnor U21743 (N_21743,N_19657,N_17774);
and U21744 (N_21744,N_15503,N_17575);
nand U21745 (N_21745,N_15184,N_17415);
nand U21746 (N_21746,N_16390,N_16336);
nor U21747 (N_21747,N_17771,N_17356);
nor U21748 (N_21748,N_19245,N_15007);
or U21749 (N_21749,N_17934,N_19277);
and U21750 (N_21750,N_16610,N_17138);
xnor U21751 (N_21751,N_19639,N_19646);
and U21752 (N_21752,N_19818,N_15945);
nor U21753 (N_21753,N_18983,N_17626);
nand U21754 (N_21754,N_18132,N_17821);
nor U21755 (N_21755,N_17556,N_19397);
or U21756 (N_21756,N_19857,N_19248);
nand U21757 (N_21757,N_16620,N_19558);
xnor U21758 (N_21758,N_16354,N_19352);
xor U21759 (N_21759,N_16926,N_15966);
or U21760 (N_21760,N_18828,N_16651);
nor U21761 (N_21761,N_17000,N_18522);
nand U21762 (N_21762,N_16876,N_19773);
nand U21763 (N_21763,N_18407,N_15541);
nor U21764 (N_21764,N_18690,N_17994);
and U21765 (N_21765,N_19092,N_16623);
or U21766 (N_21766,N_19873,N_17525);
nor U21767 (N_21767,N_16559,N_17500);
xor U21768 (N_21768,N_19648,N_15715);
nor U21769 (N_21769,N_17447,N_19056);
and U21770 (N_21770,N_18794,N_15744);
and U21771 (N_21771,N_17157,N_19844);
xor U21772 (N_21772,N_15369,N_17217);
or U21773 (N_21773,N_18543,N_16670);
or U21774 (N_21774,N_19098,N_18594);
xnor U21775 (N_21775,N_17385,N_17077);
and U21776 (N_21776,N_18918,N_18587);
nand U21777 (N_21777,N_16403,N_16835);
xnor U21778 (N_21778,N_16847,N_18826);
nand U21779 (N_21779,N_18472,N_19374);
xor U21780 (N_21780,N_16581,N_18441);
and U21781 (N_21781,N_18039,N_19871);
xor U21782 (N_21782,N_16627,N_15389);
nand U21783 (N_21783,N_17907,N_15352);
nor U21784 (N_21784,N_19060,N_16331);
xor U21785 (N_21785,N_19979,N_17055);
nor U21786 (N_21786,N_19936,N_15074);
nand U21787 (N_21787,N_16701,N_18356);
and U21788 (N_21788,N_17206,N_17300);
or U21789 (N_21789,N_18879,N_15961);
xor U21790 (N_21790,N_19889,N_15664);
nand U21791 (N_21791,N_19510,N_19540);
and U21792 (N_21792,N_16200,N_15920);
and U21793 (N_21793,N_16790,N_18352);
nand U21794 (N_21794,N_19863,N_15971);
or U21795 (N_21795,N_19226,N_17690);
and U21796 (N_21796,N_17910,N_18384);
or U21797 (N_21797,N_16396,N_16800);
nand U21798 (N_21798,N_16893,N_19548);
and U21799 (N_21799,N_16355,N_17238);
xnor U21800 (N_21800,N_18255,N_18806);
and U21801 (N_21801,N_17724,N_19228);
or U21802 (N_21802,N_16011,N_15760);
xor U21803 (N_21803,N_16956,N_16932);
nor U21804 (N_21804,N_15059,N_16057);
nand U21805 (N_21805,N_15919,N_16447);
or U21806 (N_21806,N_15629,N_18430);
nand U21807 (N_21807,N_18610,N_19895);
and U21808 (N_21808,N_17143,N_15224);
and U21809 (N_21809,N_15014,N_15948);
or U21810 (N_21810,N_19763,N_17455);
or U21811 (N_21811,N_19655,N_15794);
xor U21812 (N_21812,N_16915,N_19065);
or U21813 (N_21813,N_16019,N_19171);
xnor U21814 (N_21814,N_16666,N_18354);
or U21815 (N_21815,N_17319,N_15142);
nor U21816 (N_21816,N_16406,N_16955);
or U21817 (N_21817,N_18160,N_19761);
or U21818 (N_21818,N_16542,N_17418);
nand U21819 (N_21819,N_16148,N_17540);
or U21820 (N_21820,N_18130,N_17548);
and U21821 (N_21821,N_17856,N_18870);
and U21822 (N_21822,N_19241,N_18031);
xor U21823 (N_21823,N_15084,N_19757);
xnor U21824 (N_21824,N_18458,N_16106);
or U21825 (N_21825,N_17033,N_18293);
nor U21826 (N_21826,N_18936,N_17740);
nand U21827 (N_21827,N_16132,N_17782);
or U21828 (N_21828,N_16081,N_15159);
xnor U21829 (N_21829,N_17079,N_17561);
nor U21830 (N_21830,N_17707,N_16791);
xor U21831 (N_21831,N_17697,N_19449);
xor U21832 (N_21832,N_19679,N_15747);
xor U21833 (N_21833,N_19069,N_19663);
xor U21834 (N_21834,N_15473,N_16003);
nor U21835 (N_21835,N_15930,N_15487);
nor U21836 (N_21836,N_17878,N_17571);
nor U21837 (N_21837,N_16279,N_17091);
nor U21838 (N_21838,N_18358,N_18228);
nand U21839 (N_21839,N_19358,N_15239);
or U21840 (N_21840,N_18956,N_15385);
nand U21841 (N_21841,N_19139,N_19912);
or U21842 (N_21842,N_16598,N_15378);
xnor U21843 (N_21843,N_15810,N_15080);
xor U21844 (N_21844,N_15111,N_18074);
nand U21845 (N_21845,N_18959,N_19710);
nor U21846 (N_21846,N_15228,N_15492);
xor U21847 (N_21847,N_19469,N_18290);
nor U21848 (N_21848,N_18070,N_19290);
and U21849 (N_21849,N_16747,N_19264);
and U21850 (N_21850,N_16707,N_16576);
nor U21851 (N_21851,N_19322,N_19581);
and U21852 (N_21852,N_19907,N_18181);
xor U21853 (N_21853,N_15323,N_18309);
and U21854 (N_21854,N_16297,N_19185);
xor U21855 (N_21855,N_15764,N_15483);
and U21856 (N_21856,N_19366,N_17535);
nor U21857 (N_21857,N_19324,N_19082);
nand U21858 (N_21858,N_15360,N_15906);
or U21859 (N_21859,N_16477,N_17146);
and U21860 (N_21860,N_19259,N_16971);
and U21861 (N_21861,N_15481,N_17592);
xnor U21862 (N_21862,N_15203,N_17658);
or U21863 (N_21863,N_16637,N_17929);
nand U21864 (N_21864,N_16260,N_15564);
or U21865 (N_21865,N_17378,N_18732);
or U21866 (N_21866,N_19672,N_18208);
nor U21867 (N_21867,N_15677,N_18741);
xnor U21868 (N_21868,N_15627,N_18367);
or U21869 (N_21869,N_19879,N_17773);
and U21870 (N_21870,N_19799,N_16262);
or U21871 (N_21871,N_18805,N_19865);
or U21872 (N_21872,N_18968,N_16264);
xnor U21873 (N_21873,N_19491,N_16787);
nand U21874 (N_21874,N_17311,N_17204);
or U21875 (N_21875,N_16491,N_19869);
or U21876 (N_21876,N_15878,N_16128);
and U21877 (N_21877,N_16480,N_15578);
nand U21878 (N_21878,N_18796,N_16796);
xnor U21879 (N_21879,N_18788,N_16783);
nor U21880 (N_21880,N_16655,N_18661);
or U21881 (N_21881,N_19347,N_16617);
nor U21882 (N_21882,N_16865,N_19194);
nand U21883 (N_21883,N_16469,N_19210);
nand U21884 (N_21884,N_17457,N_19270);
nor U21885 (N_21885,N_19713,N_19850);
nand U21886 (N_21886,N_15972,N_19359);
xor U21887 (N_21887,N_16358,N_19227);
nand U21888 (N_21888,N_18836,N_15410);
xor U21889 (N_21889,N_17732,N_16504);
nand U21890 (N_21890,N_17380,N_16804);
nand U21891 (N_21891,N_15426,N_17507);
xnor U21892 (N_21892,N_17007,N_18689);
xnor U21893 (N_21893,N_18103,N_19774);
xor U21894 (N_21894,N_19353,N_19908);
and U21895 (N_21895,N_15264,N_18964);
and U21896 (N_21896,N_17627,N_19325);
nand U21897 (N_21897,N_18328,N_16525);
xor U21898 (N_21898,N_17393,N_15274);
xor U21899 (N_21899,N_18220,N_16271);
or U21900 (N_21900,N_18395,N_15847);
or U21901 (N_21901,N_16754,N_15227);
nand U21902 (N_21902,N_17613,N_15348);
and U21903 (N_21903,N_19852,N_18355);
nand U21904 (N_21904,N_19611,N_19364);
nor U21905 (N_21905,N_16613,N_15933);
nand U21906 (N_21906,N_16978,N_19556);
and U21907 (N_21907,N_15763,N_18343);
or U21908 (N_21908,N_18751,N_17566);
xor U21909 (N_21909,N_15762,N_19271);
nor U21910 (N_21910,N_19485,N_18089);
xnor U21911 (N_21911,N_15655,N_16316);
or U21912 (N_21912,N_15864,N_17891);
and U21913 (N_21913,N_18590,N_18509);
nor U21914 (N_21914,N_19401,N_16529);
nor U21915 (N_21915,N_17584,N_16389);
and U21916 (N_21916,N_19249,N_16379);
and U21917 (N_21917,N_19635,N_18996);
nand U21918 (N_21918,N_17766,N_17040);
nand U21919 (N_21919,N_19684,N_18428);
and U21920 (N_21920,N_19153,N_18440);
and U21921 (N_21921,N_16044,N_17340);
xor U21922 (N_21922,N_18484,N_17552);
nor U21923 (N_21923,N_15678,N_17606);
xor U21924 (N_21924,N_17502,N_18088);
nand U21925 (N_21925,N_18943,N_18882);
or U21926 (N_21926,N_16047,N_16661);
or U21927 (N_21927,N_18865,N_19550);
nand U21928 (N_21928,N_17503,N_18668);
and U21929 (N_21929,N_18317,N_17020);
nand U21930 (N_21930,N_15533,N_17133);
and U21931 (N_21931,N_16536,N_18978);
or U21932 (N_21932,N_19304,N_17366);
nor U21933 (N_21933,N_16767,N_15431);
xnor U21934 (N_21934,N_16339,N_17442);
nand U21935 (N_21935,N_17569,N_19203);
and U21936 (N_21936,N_18277,N_19305);
xnor U21937 (N_21937,N_15405,N_15383);
xnor U21938 (N_21938,N_17964,N_19828);
or U21939 (N_21939,N_17216,N_16493);
nand U21940 (N_21940,N_17214,N_16777);
and U21941 (N_21941,N_16193,N_16061);
xor U21942 (N_21942,N_15778,N_19049);
nor U21943 (N_21943,N_19597,N_16441);
nor U21944 (N_21944,N_16643,N_16215);
xnor U21945 (N_21945,N_15029,N_15636);
and U21946 (N_21946,N_17468,N_16351);
and U21947 (N_21947,N_15076,N_18618);
nand U21948 (N_21948,N_19152,N_15160);
nand U21949 (N_21949,N_18369,N_15620);
nand U21950 (N_21950,N_15818,N_18450);
nor U21951 (N_21951,N_16048,N_16111);
xor U21952 (N_21952,N_19642,N_16603);
nand U21953 (N_21953,N_19878,N_18790);
or U21954 (N_21954,N_18703,N_19404);
nand U21955 (N_21955,N_15558,N_19567);
or U21956 (N_21956,N_19369,N_15591);
xor U21957 (N_21957,N_15869,N_15123);
or U21958 (N_21958,N_15625,N_15175);
xor U21959 (N_21959,N_16408,N_18613);
and U21960 (N_21960,N_16571,N_19645);
xor U21961 (N_21961,N_19027,N_16593);
xor U21962 (N_21962,N_16606,N_19102);
or U21963 (N_21963,N_15313,N_18278);
or U21964 (N_21964,N_15807,N_15130);
nand U21965 (N_21965,N_17554,N_17001);
nor U21966 (N_21966,N_16711,N_16415);
or U21967 (N_21967,N_16289,N_15235);
nor U21968 (N_21968,N_18871,N_15400);
nand U21969 (N_21969,N_15941,N_19286);
nor U21970 (N_21970,N_18582,N_18930);
nand U21971 (N_21971,N_15461,N_19544);
nor U21972 (N_21972,N_19244,N_17940);
or U21973 (N_21973,N_15777,N_16398);
or U21974 (N_21974,N_17444,N_18051);
and U21975 (N_21975,N_15568,N_17652);
nand U21976 (N_21976,N_17908,N_17615);
and U21977 (N_21977,N_15415,N_19164);
nor U21978 (N_21978,N_18476,N_15265);
nand U21979 (N_21979,N_16859,N_17406);
xnor U21980 (N_21980,N_15633,N_15093);
nor U21981 (N_21981,N_18754,N_16545);
nand U21982 (N_21982,N_18411,N_18776);
or U21983 (N_21983,N_15216,N_16560);
or U21984 (N_21984,N_16101,N_16041);
xnor U21985 (N_21985,N_18049,N_19962);
or U21986 (N_21986,N_19589,N_19063);
nand U21987 (N_21987,N_17035,N_19664);
nand U21988 (N_21988,N_15788,N_15954);
nand U21989 (N_21989,N_18157,N_16209);
xor U21990 (N_21990,N_19087,N_15099);
nand U21991 (N_21991,N_17072,N_16381);
and U21992 (N_21992,N_15735,N_15673);
nor U21993 (N_21993,N_18237,N_15832);
or U21994 (N_21994,N_17854,N_15433);
and U21995 (N_21995,N_16281,N_16134);
nand U21996 (N_21996,N_16394,N_19783);
nand U21997 (N_21997,N_15939,N_17465);
nor U21998 (N_21998,N_17528,N_17508);
nor U21999 (N_21999,N_18018,N_17099);
nand U22000 (N_22000,N_19481,N_16770);
nor U22001 (N_22001,N_16126,N_17399);
or U22002 (N_22002,N_18670,N_19205);
or U22003 (N_22003,N_18443,N_18648);
nand U22004 (N_22004,N_15325,N_18752);
or U22005 (N_22005,N_15825,N_17421);
or U22006 (N_22006,N_16842,N_18308);
nand U22007 (N_22007,N_15624,N_17283);
nor U22008 (N_22008,N_16016,N_18388);
or U22009 (N_22009,N_19536,N_15471);
nor U22010 (N_22010,N_18146,N_17458);
or U22011 (N_22011,N_18324,N_18084);
or U22012 (N_22012,N_16963,N_17181);
nor U22013 (N_22013,N_18827,N_15013);
nor U22014 (N_22014,N_19582,N_19616);
or U22015 (N_22015,N_18287,N_15706);
nand U22016 (N_22016,N_17318,N_16964);
nand U22017 (N_22017,N_16471,N_16410);
nand U22018 (N_22018,N_16802,N_16717);
and U22019 (N_22019,N_15088,N_16907);
nor U22020 (N_22020,N_18859,N_17362);
nor U22021 (N_22021,N_16897,N_18346);
nand U22022 (N_22022,N_17577,N_16211);
xnor U22023 (N_22023,N_15257,N_15375);
nor U22024 (N_22024,N_18934,N_18680);
nor U22025 (N_22025,N_16374,N_18947);
and U22026 (N_22026,N_18001,N_18510);
xnor U22027 (N_22027,N_19691,N_19187);
and U22028 (N_22028,N_18222,N_18233);
xnor U22029 (N_22029,N_17734,N_15891);
or U22030 (N_22030,N_15942,N_15402);
or U22031 (N_22031,N_18927,N_16757);
xor U22032 (N_22032,N_17117,N_16287);
nand U22033 (N_22033,N_17336,N_19742);
xor U22034 (N_22034,N_17358,N_19495);
or U22035 (N_22035,N_17034,N_18646);
and U22036 (N_22036,N_18778,N_18941);
xor U22037 (N_22037,N_18769,N_18848);
nand U22038 (N_22038,N_17788,N_18624);
xnor U22039 (N_22039,N_19517,N_17952);
or U22040 (N_22040,N_17086,N_16761);
or U22041 (N_22041,N_18000,N_19924);
nor U22042 (N_22042,N_18551,N_18878);
nor U22043 (N_22043,N_19641,N_17666);
xnor U22044 (N_22044,N_16810,N_15587);
nor U22045 (N_22045,N_18602,N_18877);
or U22046 (N_22046,N_17097,N_16819);
nor U22047 (N_22047,N_18030,N_15669);
xor U22048 (N_22048,N_19966,N_19800);
or U22049 (N_22049,N_18561,N_15042);
nand U22050 (N_22050,N_17951,N_17145);
or U22051 (N_22051,N_17966,N_18765);
xnor U22052 (N_22052,N_19428,N_19041);
nand U22053 (N_22053,N_16257,N_17858);
or U22054 (N_22054,N_18351,N_18792);
and U22055 (N_22055,N_16868,N_19143);
xor U22056 (N_22056,N_15796,N_17332);
xor U22057 (N_22057,N_15154,N_18462);
nor U22058 (N_22058,N_19285,N_18078);
and U22059 (N_22059,N_19150,N_19330);
xnor U22060 (N_22060,N_18311,N_18584);
xor U22061 (N_22061,N_16516,N_15597);
and U22062 (N_22062,N_15750,N_15901);
and U22063 (N_22063,N_16380,N_16142);
nor U22064 (N_22064,N_15841,N_15038);
or U22065 (N_22065,N_16811,N_19221);
xor U22066 (N_22066,N_19318,N_15783);
nor U22067 (N_22067,N_18013,N_18423);
or U22068 (N_22068,N_18507,N_16483);
or U22069 (N_22069,N_19192,N_16673);
or U22070 (N_22070,N_15211,N_17565);
xnor U22071 (N_22071,N_19520,N_15460);
nand U22072 (N_22072,N_15285,N_19843);
or U22073 (N_22073,N_16911,N_18040);
nor U22074 (N_22074,N_15657,N_18945);
xnor U22075 (N_22075,N_17467,N_16650);
nand U22076 (N_22076,N_17474,N_18316);
and U22077 (N_22077,N_16695,N_18986);
and U22078 (N_22078,N_18520,N_15969);
nor U22079 (N_22079,N_16176,N_19295);
xnor U22080 (N_22080,N_18911,N_15792);
or U22081 (N_22081,N_17294,N_16609);
and U22082 (N_22082,N_15911,N_17855);
xor U22083 (N_22083,N_19928,N_16330);
xor U22084 (N_22084,N_17860,N_15272);
and U22085 (N_22085,N_17671,N_17490);
nand U22086 (N_22086,N_15719,N_17765);
and U22087 (N_22087,N_15193,N_16094);
or U22088 (N_22088,N_19665,N_18409);
nand U22089 (N_22089,N_17834,N_16588);
or U22090 (N_22090,N_15937,N_15087);
or U22091 (N_22091,N_16634,N_18786);
and U22092 (N_22092,N_18875,N_15229);
or U22093 (N_22093,N_17529,N_17276);
and U22094 (N_22094,N_19350,N_15214);
nor U22095 (N_22095,N_15381,N_19128);
or U22096 (N_22096,N_18990,N_16507);
nand U22097 (N_22097,N_18009,N_16348);
xnor U22098 (N_22098,N_16775,N_16636);
xor U22099 (N_22099,N_16774,N_18669);
nor U22100 (N_22100,N_18731,N_17589);
or U22101 (N_22101,N_17116,N_19988);
or U22102 (N_22102,N_15635,N_16589);
or U22103 (N_22103,N_19890,N_15502);
or U22104 (N_22104,N_15011,N_17900);
nand U22105 (N_22105,N_17968,N_15069);
nor U22106 (N_22106,N_15887,N_15208);
xor U22107 (N_22107,N_19011,N_19622);
and U22108 (N_22108,N_15441,N_15817);
nor U22109 (N_22109,N_18284,N_15250);
xnor U22110 (N_22110,N_18782,N_17521);
xnor U22111 (N_22111,N_19754,N_15944);
or U22112 (N_22112,N_18720,N_15716);
xor U22113 (N_22113,N_15903,N_15647);
xor U22114 (N_22114,N_15205,N_16837);
nor U22115 (N_22115,N_15136,N_18323);
nor U22116 (N_22116,N_19712,N_17050);
and U22117 (N_22117,N_19332,N_15723);
and U22118 (N_22118,N_19768,N_19839);
and U22119 (N_22119,N_18833,N_19386);
nor U22120 (N_22120,N_15339,N_16323);
and U22121 (N_22121,N_17198,N_17306);
xnor U22122 (N_22122,N_19985,N_17123);
and U22123 (N_22123,N_18389,N_18057);
nand U22124 (N_22124,N_19947,N_19272);
xor U22125 (N_22125,N_19685,N_16230);
nor U22126 (N_22126,N_18276,N_17271);
nor U22127 (N_22127,N_19814,N_19957);
nand U22128 (N_22128,N_19186,N_15359);
and U22129 (N_22129,N_18238,N_18460);
and U22130 (N_22130,N_17361,N_18965);
or U22131 (N_22131,N_15576,N_18516);
and U22132 (N_22132,N_15373,N_15303);
nand U22133 (N_22133,N_15073,N_15526);
nand U22134 (N_22134,N_18474,N_16782);
nor U22135 (N_22135,N_15194,N_18494);
and U22136 (N_22136,N_16751,N_18569);
nor U22137 (N_22137,N_18093,N_19637);
nor U22138 (N_22138,N_19067,N_16383);
nor U22139 (N_22139,N_17021,N_18186);
nor U22140 (N_22140,N_15370,N_19897);
nor U22141 (N_22141,N_18604,N_15223);
nor U22142 (N_22142,N_19018,N_18530);
and U22143 (N_22143,N_17322,N_18565);
and U22144 (N_22144,N_19085,N_15330);
xnor U22145 (N_22145,N_16854,N_19222);
nor U22146 (N_22146,N_19654,N_19298);
nor U22147 (N_22147,N_16662,N_17919);
nor U22148 (N_22148,N_17477,N_17150);
xnor U22149 (N_22149,N_15646,N_17382);
nand U22150 (N_22150,N_19433,N_18275);
nand U22151 (N_22151,N_16621,N_17351);
nand U22152 (N_22152,N_15000,N_17028);
or U22153 (N_22153,N_16444,N_19265);
nand U22154 (N_22154,N_15559,N_17932);
and U22155 (N_22155,N_19849,N_16202);
nand U22156 (N_22156,N_18724,N_16409);
xnor U22157 (N_22157,N_19175,N_15824);
nor U22158 (N_22158,N_17236,N_17977);
nor U22159 (N_22159,N_16704,N_19180);
xnor U22160 (N_22160,N_16207,N_17364);
and U22161 (N_22161,N_18773,N_18205);
and U22162 (N_22162,N_18121,N_19703);
nor U22163 (N_22163,N_17324,N_18681);
and U22164 (N_22164,N_19884,N_19415);
nand U22165 (N_22165,N_15301,N_18925);
nor U22166 (N_22166,N_16210,N_16454);
and U22167 (N_22167,N_15840,N_18710);
and U22168 (N_22168,N_17981,N_17807);
nor U22169 (N_22169,N_15689,N_17388);
and U22170 (N_22170,N_15709,N_19026);
or U22171 (N_22171,N_16313,N_18466);
xor U22172 (N_22172,N_15167,N_15819);
or U22173 (N_22173,N_18820,N_17200);
xnor U22174 (N_22174,N_19653,N_15520);
nor U22175 (N_22175,N_15082,N_17446);
nor U22176 (N_22176,N_15362,N_18372);
nand U22177 (N_22177,N_16667,N_19109);
or U22178 (N_22178,N_18196,N_19991);
xor U22179 (N_22179,N_15936,N_16984);
or U22180 (N_22180,N_18804,N_17316);
nor U22181 (N_22181,N_17039,N_17249);
nand U22182 (N_22182,N_18128,N_18410);
or U22183 (N_22183,N_16625,N_18738);
or U22184 (N_22184,N_18398,N_19357);
nor U22185 (N_22185,N_18027,N_19316);
nor U22186 (N_22186,N_19584,N_16715);
nor U22187 (N_22187,N_18739,N_17640);
xor U22188 (N_22188,N_15667,N_16936);
nor U22189 (N_22189,N_16189,N_15977);
xnor U22190 (N_22190,N_18552,N_18994);
nor U22191 (N_22191,N_16629,N_15427);
xnor U22192 (N_22192,N_16205,N_17999);
nor U22193 (N_22193,N_19610,N_15784);
xor U22194 (N_22194,N_15253,N_19531);
nand U22195 (N_22195,N_19502,N_18310);
nor U22196 (N_22196,N_15804,N_18991);
xor U22197 (N_22197,N_18762,N_15052);
nand U22198 (N_22198,N_17895,N_16569);
xor U22199 (N_22199,N_16450,N_18938);
and U22200 (N_22200,N_18803,N_15545);
or U22201 (N_22201,N_17946,N_18839);
nand U22202 (N_22202,N_15090,N_16237);
xnor U22203 (N_22203,N_15852,N_15897);
and U22204 (N_22204,N_19981,N_16310);
and U22205 (N_22205,N_17643,N_16006);
nand U22206 (N_22206,N_19644,N_19217);
nand U22207 (N_22207,N_18218,N_18448);
or U22208 (N_22208,N_15594,N_18636);
xnor U22209 (N_22209,N_19043,N_16758);
and U22210 (N_22210,N_19238,N_16699);
nor U22211 (N_22211,N_18701,N_15562);
or U22212 (N_22212,N_18951,N_18917);
or U22213 (N_22213,N_17227,N_19434);
nand U22214 (N_22214,N_15363,N_15717);
or U22215 (N_22215,N_16860,N_17409);
xor U22216 (N_22216,N_17862,N_19471);
xor U22217 (N_22217,N_16805,N_16558);
and U22218 (N_22218,N_19377,N_17164);
or U22219 (N_22219,N_15710,N_16333);
nor U22220 (N_22220,N_19492,N_15761);
and U22221 (N_22221,N_16502,N_18127);
and U22222 (N_22222,N_15163,N_15463);
or U22223 (N_22223,N_16177,N_16244);
nand U22224 (N_22224,N_16555,N_17499);
nor U22225 (N_22225,N_19480,N_18406);
nor U22226 (N_22226,N_18686,N_16587);
nand U22227 (N_22227,N_16294,N_17044);
nand U22228 (N_22228,N_15752,N_19888);
or U22229 (N_22229,N_19562,N_17661);
xor U22230 (N_22230,N_16147,N_17880);
nor U22231 (N_22231,N_16366,N_17582);
nor U22232 (N_22232,N_16117,N_17835);
and U22233 (N_22233,N_15720,N_16309);
nand U22234 (N_22234,N_18433,N_18852);
or U22235 (N_22235,N_18066,N_19588);
nand U22236 (N_22236,N_18539,N_19182);
or U22237 (N_22237,N_19969,N_19940);
and U22238 (N_22238,N_17126,N_18457);
nand U22239 (N_22239,N_16866,N_15004);
nor U22240 (N_22240,N_16682,N_17183);
nor U22241 (N_22241,N_17397,N_17894);
nor U22242 (N_22242,N_17539,N_15053);
nand U22243 (N_22243,N_15755,N_17414);
nand U22244 (N_22244,N_18475,N_18853);
and U22245 (N_22245,N_19797,N_19974);
nand U22246 (N_22246,N_19146,N_15619);
nor U22247 (N_22247,N_19631,N_18524);
nor U22248 (N_22248,N_15057,N_18837);
nand U22249 (N_22249,N_15679,N_18957);
nand U22250 (N_22250,N_16579,N_18174);
nor U22251 (N_22251,N_19739,N_18807);
or U22252 (N_22252,N_18647,N_15598);
xor U22253 (N_22253,N_19737,N_19024);
or U22254 (N_22254,N_15295,N_17339);
nand U22255 (N_22255,N_19413,N_18975);
xor U22256 (N_22256,N_19391,N_15612);
nor U22257 (N_22257,N_19733,N_18445);
or U22258 (N_22258,N_15714,N_15681);
nor U22259 (N_22259,N_15275,N_15320);
nand U22260 (N_22260,N_15935,N_16319);
or U22261 (N_22261,N_18023,N_17698);
xor U22262 (N_22262,N_16712,N_19414);
xnor U22263 (N_22263,N_18131,N_16817);
xor U22264 (N_22264,N_15532,N_17721);
nand U22265 (N_22265,N_15068,N_19559);
nand U22266 (N_22266,N_19704,N_17301);
or U22267 (N_22267,N_17889,N_17553);
and U22268 (N_22268,N_19736,N_15892);
and U22269 (N_22269,N_18298,N_19444);
nand U22270 (N_22270,N_16714,N_15147);
nand U22271 (N_22271,N_17045,N_16983);
or U22272 (N_22272,N_16407,N_16599);
nand U22273 (N_22273,N_15628,N_18512);
nor U22274 (N_22274,N_18424,N_18204);
xnor U22275 (N_22275,N_17327,N_17960);
nand U22276 (N_22276,N_15083,N_19459);
or U22277 (N_22277,N_18633,N_17755);
xor U22278 (N_22278,N_17747,N_15885);
and U22279 (N_22279,N_18726,N_19935);
nand U22280 (N_22280,N_16899,N_19484);
and U22281 (N_22281,N_19134,N_17663);
nor U22282 (N_22282,N_19453,N_16322);
nand U22283 (N_22283,N_16024,N_16713);
nor U22284 (N_22284,N_17228,N_19606);
or U22285 (N_22285,N_18202,N_18508);
or U22286 (N_22286,N_15830,N_18756);
xnor U22287 (N_22287,N_15413,N_19424);
nand U22288 (N_22288,N_17046,N_15161);
nand U22289 (N_22289,N_16869,N_16021);
and U22290 (N_22290,N_16114,N_19254);
and U22291 (N_22291,N_15191,N_17573);
nand U22292 (N_22292,N_19990,N_18152);
and U22293 (N_22293,N_17398,N_17753);
nor U22294 (N_22294,N_15144,N_17173);
nand U22295 (N_22295,N_19355,N_16270);
and U22296 (N_22296,N_17386,N_17494);
nor U22297 (N_22297,N_18043,N_16340);
xnor U22298 (N_22298,N_19868,N_15001);
and U22299 (N_22299,N_16475,N_19965);
xor U22300 (N_22300,N_19683,N_17313);
xnor U22301 (N_22301,N_16367,N_19772);
xnor U22302 (N_22302,N_17948,N_15258);
or U22303 (N_22303,N_18175,N_18412);
nand U22304 (N_22304,N_17466,N_17177);
and U22305 (N_22305,N_17731,N_18314);
nor U22306 (N_22306,N_16530,N_15547);
nand U22307 (N_22307,N_16849,N_17614);
xnor U22308 (N_22308,N_15366,N_19031);
xnor U22309 (N_22309,N_15252,N_15293);
and U22310 (N_22310,N_15343,N_16479);
or U22311 (N_22311,N_15511,N_18540);
nand U22312 (N_22312,N_17630,N_16882);
nand U22313 (N_22313,N_19106,N_17101);
nor U22314 (N_22314,N_17085,N_16283);
and U22315 (N_22315,N_16063,N_17139);
nor U22316 (N_22316,N_16399,N_18506);
nor U22317 (N_22317,N_19107,N_17239);
xnor U22318 (N_22318,N_17624,N_17672);
xor U22319 (N_22319,N_19419,N_18381);
nand U22320 (N_22320,N_18908,N_18306);
nor U22321 (N_22321,N_19284,N_16342);
or U22322 (N_22322,N_17209,N_15137);
and U22323 (N_22323,N_18149,N_15544);
nand U22324 (N_22324,N_17390,N_16785);
or U22325 (N_22325,N_15959,N_18387);
nor U22326 (N_22326,N_18533,N_18434);
xnor U22327 (N_22327,N_16127,N_16676);
nand U22328 (N_22328,N_17998,N_16611);
nor U22329 (N_22329,N_16384,N_17790);
or U22330 (N_22330,N_19975,N_15428);
nor U22331 (N_22331,N_16886,N_19001);
xnor U22332 (N_22332,N_15377,N_19949);
nand U22333 (N_22333,N_15222,N_15018);
nand U22334 (N_22334,N_17261,N_15464);
nor U22335 (N_22335,N_16976,N_19044);
xnor U22336 (N_22336,N_17793,N_18861);
and U22337 (N_22337,N_18586,N_17594);
nor U22338 (N_22338,N_15023,N_15346);
xnor U22339 (N_22339,N_16036,N_16060);
or U22340 (N_22340,N_18678,N_15688);
xnor U22341 (N_22341,N_19237,N_18010);
nor U22342 (N_22342,N_17025,N_15443);
or U22343 (N_22343,N_17017,N_16648);
xor U22344 (N_22344,N_17811,N_16152);
and U22345 (N_22345,N_16242,N_15708);
nor U22346 (N_22346,N_15500,N_19250);
or U22347 (N_22347,N_17560,N_18337);
xor U22348 (N_22348,N_18637,N_17845);
xor U22349 (N_22349,N_17435,N_15329);
or U22350 (N_22350,N_19788,N_18368);
or U22351 (N_22351,N_16030,N_19140);
and U22352 (N_22352,N_17664,N_19955);
xor U22353 (N_22353,N_17909,N_18248);
xor U22354 (N_22354,N_16841,N_19764);
xor U22355 (N_22355,N_17413,N_16216);
nand U22356 (N_22356,N_17543,N_19335);
xnor U22357 (N_22357,N_18600,N_17270);
and U22358 (N_22358,N_16464,N_16592);
nand U22359 (N_22359,N_16385,N_19240);
nor U22360 (N_22360,N_19795,N_16138);
and U22361 (N_22361,N_17992,N_16612);
or U22362 (N_22362,N_15570,N_19769);
nor U22363 (N_22363,N_19578,N_16086);
nor U22364 (N_22364,N_17165,N_16972);
nor U22365 (N_22365,N_15478,N_16251);
and U22366 (N_22366,N_18168,N_16438);
and U22367 (N_22367,N_15691,N_18620);
xnor U22368 (N_22368,N_18662,N_17259);
nor U22369 (N_22369,N_19151,N_15538);
or U22370 (N_22370,N_16026,N_18844);
nand U22371 (N_22371,N_19636,N_16909);
nor U22372 (N_22372,N_16820,N_18432);
or U22373 (N_22373,N_17622,N_16298);
or U22374 (N_22374,N_15581,N_18621);
xnor U22375 (N_22375,N_18469,N_15938);
nand U22376 (N_22376,N_17051,N_18737);
nand U22377 (N_22377,N_19232,N_17250);
or U22378 (N_22378,N_19798,N_17100);
and U22379 (N_22379,N_18022,N_19177);
nor U22380 (N_22380,N_16401,N_15015);
nor U22381 (N_22381,N_18940,N_19505);
xor U22382 (N_22382,N_17843,N_15727);
nand U22383 (N_22383,N_15615,N_19987);
xor U22384 (N_22384,N_16815,N_17725);
and U22385 (N_22385,N_16942,N_19493);
xnor U22386 (N_22386,N_15871,N_18259);
nor U22387 (N_22387,N_18749,N_18064);
and U22388 (N_22388,N_17108,N_19989);
nand U22389 (N_22389,N_18065,N_18143);
xnor U22390 (N_22390,N_17136,N_18890);
or U22391 (N_22391,N_16203,N_16250);
or U22392 (N_22392,N_19944,N_16944);
and U22393 (N_22393,N_18654,N_19838);
or U22394 (N_22394,N_18789,N_16252);
xor U22395 (N_22395,N_16357,N_15024);
xor U22396 (N_22396,N_18706,N_18342);
and U22397 (N_22397,N_15064,N_17469);
nor U22398 (N_22398,N_16486,N_17949);
or U22399 (N_22399,N_17645,N_19925);
nand U22400 (N_22400,N_15332,N_18960);
or U22401 (N_22401,N_15249,N_19626);
or U22402 (N_22402,N_17513,N_18037);
xor U22403 (N_22403,N_16158,N_15809);
or U22404 (N_22404,N_17120,N_19643);
xnor U22405 (N_22405,N_16434,N_16050);
nor U22406 (N_22406,N_15340,N_19740);
or U22407 (N_22407,N_16764,N_16445);
nand U22408 (N_22408,N_17370,N_19822);
xor U22409 (N_22409,N_17401,N_19234);
nor U22410 (N_22410,N_18299,N_17224);
and U22411 (N_22411,N_18192,N_18402);
nand U22412 (N_22412,N_15298,N_16564);
or U22413 (N_22413,N_16743,N_17256);
nor U22414 (N_22414,N_16282,N_18005);
xor U22415 (N_22415,N_17208,N_18464);
xnor U22416 (N_22416,N_19361,N_19823);
nor U22417 (N_22417,N_19695,N_19917);
nand U22418 (N_22418,N_18641,N_15466);
nand U22419 (N_22419,N_17673,N_17826);
nor U22420 (N_22420,N_17342,N_17026);
or U22421 (N_22421,N_18667,N_15327);
nand U22422 (N_22422,N_16195,N_16512);
and U22423 (N_22423,N_16280,N_19741);
or U22424 (N_22424,N_17570,N_15900);
nand U22425 (N_22425,N_18961,N_15196);
xnor U22426 (N_22426,N_18864,N_16672);
and U22427 (N_22427,N_15012,N_17628);
nand U22428 (N_22428,N_16304,N_17509);
nor U22429 (N_22429,N_15342,N_18478);
and U22430 (N_22430,N_17705,N_18575);
xor U22431 (N_22431,N_17036,N_15077);
nor U22432 (N_22432,N_16470,N_15537);
nor U22433 (N_22433,N_16020,N_19677);
xor U22434 (N_22434,N_18980,N_16993);
xnor U22435 (N_22435,N_18226,N_18775);
and U22436 (N_22436,N_16863,N_16669);
and U22437 (N_22437,N_18379,N_17487);
or U22438 (N_22438,N_15098,N_17291);
xnor U22439 (N_22439,N_18279,N_16468);
nand U22440 (N_22440,N_15319,N_17244);
xnor U22441 (N_22441,N_15365,N_18926);
nand U22442 (N_22442,N_17373,N_17495);
nand U22443 (N_22443,N_15759,N_17706);
xor U22444 (N_22444,N_15355,N_16188);
xnor U22445 (N_22445,N_15354,N_15027);
nand U22446 (N_22446,N_15032,N_15289);
nor U22447 (N_22447,N_19551,N_15315);
or U22448 (N_22448,N_15132,N_15699);
nor U22449 (N_22449,N_17703,N_18185);
nor U22450 (N_22450,N_15102,N_17954);
xor U22451 (N_22451,N_15200,N_17696);
or U22452 (N_22452,N_15447,N_19212);
and U22453 (N_22453,N_18675,N_15758);
or U22454 (N_22454,N_18989,N_18711);
and U22455 (N_22455,N_18274,N_19714);
nand U22456 (N_22456,N_19017,N_19743);
or U22457 (N_22457,N_17331,N_17737);
nand U22458 (N_22458,N_18659,N_15458);
xor U22459 (N_22459,N_17167,N_16285);
xnor U22460 (N_22460,N_17310,N_19273);
or U22461 (N_22461,N_18173,N_18919);
nor U22462 (N_22462,N_15139,N_16212);
nor U22463 (N_22463,N_15815,N_19706);
and U22464 (N_22464,N_19790,N_17623);
and U22465 (N_22465,N_15641,N_19119);
xor U22466 (N_22466,N_15895,N_19848);
or U22467 (N_22467,N_19915,N_15055);
xnor U22468 (N_22468,N_17027,N_18239);
nor U22469 (N_22469,N_19963,N_16683);
or U22470 (N_22470,N_15771,N_19439);
nor U22471 (N_22471,N_18639,N_16411);
or U22472 (N_22472,N_17059,N_16597);
nor U22473 (N_22473,N_15835,N_16400);
or U22474 (N_22474,N_15125,N_15738);
nand U22475 (N_22475,N_17379,N_16296);
nand U22476 (N_22476,N_19446,N_16395);
or U22477 (N_22477,N_17134,N_17795);
xnor U22478 (N_22478,N_17984,N_18257);
nor U22479 (N_22479,N_18682,N_19430);
xor U22480 (N_22480,N_15523,N_16326);
or U22481 (N_22481,N_16420,N_17328);
nor U22482 (N_22482,N_15695,N_16080);
xnor U22483 (N_22483,N_16677,N_19688);
nor U22484 (N_22484,N_16852,N_17221);
nor U22485 (N_22485,N_18672,N_17298);
and U22486 (N_22486,N_19725,N_15584);
or U22487 (N_22487,N_16362,N_17297);
or U22488 (N_22488,N_16523,N_15821);
or U22489 (N_22489,N_17470,N_19992);
nor U22490 (N_22490,N_16816,N_17248);
nor U22491 (N_22491,N_16521,N_19765);
or U22492 (N_22492,N_18301,N_16727);
nor U22493 (N_22493,N_15884,N_18825);
nand U22494 (N_22494,N_15440,N_19144);
and U22495 (N_22495,N_17163,N_16744);
xnor U22496 (N_22496,N_16482,N_16042);
nand U22497 (N_22497,N_17234,N_19368);
xor U22498 (N_22498,N_15899,N_19751);
and U22499 (N_22499,N_16694,N_17917);
nor U22500 (N_22500,N_17878,N_15804);
xnor U22501 (N_22501,N_17094,N_18402);
nand U22502 (N_22502,N_17407,N_17731);
nor U22503 (N_22503,N_16521,N_15513);
nor U22504 (N_22504,N_19466,N_19584);
and U22505 (N_22505,N_19868,N_16217);
xor U22506 (N_22506,N_17201,N_16088);
or U22507 (N_22507,N_15368,N_18173);
nand U22508 (N_22508,N_15591,N_16201);
and U22509 (N_22509,N_15563,N_17844);
xor U22510 (N_22510,N_19281,N_15078);
or U22511 (N_22511,N_19461,N_15753);
xor U22512 (N_22512,N_18651,N_17041);
xor U22513 (N_22513,N_16519,N_17656);
nor U22514 (N_22514,N_16066,N_15713);
nor U22515 (N_22515,N_18413,N_19135);
xnor U22516 (N_22516,N_17772,N_15841);
and U22517 (N_22517,N_18723,N_17000);
nor U22518 (N_22518,N_17997,N_18106);
nand U22519 (N_22519,N_15340,N_19436);
nand U22520 (N_22520,N_18767,N_16538);
xnor U22521 (N_22521,N_19948,N_18707);
nand U22522 (N_22522,N_18763,N_16676);
nand U22523 (N_22523,N_17746,N_16455);
or U22524 (N_22524,N_17243,N_18881);
nand U22525 (N_22525,N_17173,N_17862);
and U22526 (N_22526,N_15196,N_19148);
or U22527 (N_22527,N_15396,N_16930);
or U22528 (N_22528,N_19872,N_16686);
xnor U22529 (N_22529,N_19291,N_15492);
or U22530 (N_22530,N_19769,N_17742);
or U22531 (N_22531,N_15117,N_19954);
nand U22532 (N_22532,N_17367,N_18906);
nor U22533 (N_22533,N_19222,N_18470);
xnor U22534 (N_22534,N_15072,N_17641);
and U22535 (N_22535,N_18280,N_15732);
nor U22536 (N_22536,N_18305,N_16964);
and U22537 (N_22537,N_19142,N_15833);
nand U22538 (N_22538,N_18127,N_17716);
nor U22539 (N_22539,N_19153,N_18396);
nand U22540 (N_22540,N_18113,N_15461);
nor U22541 (N_22541,N_17301,N_18070);
nor U22542 (N_22542,N_16478,N_17152);
or U22543 (N_22543,N_15270,N_15751);
and U22544 (N_22544,N_17961,N_15948);
or U22545 (N_22545,N_17228,N_15865);
or U22546 (N_22546,N_16146,N_18726);
and U22547 (N_22547,N_15495,N_18035);
nand U22548 (N_22548,N_15238,N_18636);
nand U22549 (N_22549,N_17078,N_19263);
nand U22550 (N_22550,N_15240,N_18608);
nand U22551 (N_22551,N_15079,N_16929);
nand U22552 (N_22552,N_19506,N_16827);
xnor U22553 (N_22553,N_15473,N_19748);
nand U22554 (N_22554,N_19507,N_17447);
xor U22555 (N_22555,N_15039,N_17727);
or U22556 (N_22556,N_16793,N_17914);
nand U22557 (N_22557,N_16023,N_17962);
nor U22558 (N_22558,N_16659,N_19215);
xor U22559 (N_22559,N_18741,N_19816);
or U22560 (N_22560,N_15469,N_17013);
xor U22561 (N_22561,N_17525,N_16585);
or U22562 (N_22562,N_19825,N_18475);
and U22563 (N_22563,N_17483,N_16277);
or U22564 (N_22564,N_17707,N_17099);
and U22565 (N_22565,N_19830,N_16766);
nor U22566 (N_22566,N_18960,N_18879);
or U22567 (N_22567,N_18784,N_18967);
or U22568 (N_22568,N_18049,N_16664);
xor U22569 (N_22569,N_17643,N_18706);
xnor U22570 (N_22570,N_18931,N_18474);
nor U22571 (N_22571,N_19506,N_19090);
and U22572 (N_22572,N_18686,N_17728);
and U22573 (N_22573,N_16738,N_19927);
xor U22574 (N_22574,N_18020,N_18865);
or U22575 (N_22575,N_18902,N_17802);
nand U22576 (N_22576,N_17259,N_16506);
or U22577 (N_22577,N_16892,N_15901);
nor U22578 (N_22578,N_19498,N_18887);
nand U22579 (N_22579,N_18316,N_16122);
or U22580 (N_22580,N_18637,N_19441);
or U22581 (N_22581,N_16931,N_16607);
or U22582 (N_22582,N_16239,N_17413);
or U22583 (N_22583,N_17268,N_15769);
and U22584 (N_22584,N_17139,N_15650);
nand U22585 (N_22585,N_15886,N_15942);
and U22586 (N_22586,N_15243,N_16476);
and U22587 (N_22587,N_16053,N_18257);
nand U22588 (N_22588,N_15295,N_16067);
nor U22589 (N_22589,N_18119,N_16407);
or U22590 (N_22590,N_19716,N_16360);
nand U22591 (N_22591,N_19315,N_19694);
xnor U22592 (N_22592,N_18276,N_15508);
or U22593 (N_22593,N_16082,N_19593);
and U22594 (N_22594,N_18050,N_16744);
and U22595 (N_22595,N_19453,N_17806);
or U22596 (N_22596,N_18776,N_16132);
and U22597 (N_22597,N_18731,N_17045);
nand U22598 (N_22598,N_19931,N_15671);
xor U22599 (N_22599,N_15755,N_15362);
nand U22600 (N_22600,N_19830,N_15400);
nand U22601 (N_22601,N_16963,N_19764);
nand U22602 (N_22602,N_17792,N_19523);
or U22603 (N_22603,N_15024,N_17061);
xnor U22604 (N_22604,N_18925,N_17070);
nor U22605 (N_22605,N_16927,N_18921);
and U22606 (N_22606,N_18905,N_15610);
or U22607 (N_22607,N_17698,N_17702);
xnor U22608 (N_22608,N_19347,N_18529);
xnor U22609 (N_22609,N_19959,N_18212);
xnor U22610 (N_22610,N_16666,N_16133);
or U22611 (N_22611,N_18833,N_15132);
or U22612 (N_22612,N_19969,N_16840);
and U22613 (N_22613,N_15890,N_19331);
or U22614 (N_22614,N_19501,N_19733);
xnor U22615 (N_22615,N_17124,N_18033);
nor U22616 (N_22616,N_17412,N_17769);
or U22617 (N_22617,N_19064,N_18969);
nand U22618 (N_22618,N_18876,N_19233);
xnor U22619 (N_22619,N_19214,N_17556);
nor U22620 (N_22620,N_15055,N_17523);
or U22621 (N_22621,N_16200,N_16491);
nor U22622 (N_22622,N_19611,N_15795);
and U22623 (N_22623,N_19507,N_19072);
xnor U22624 (N_22624,N_19040,N_19933);
nor U22625 (N_22625,N_16351,N_15295);
or U22626 (N_22626,N_19856,N_15441);
or U22627 (N_22627,N_15851,N_15891);
nand U22628 (N_22628,N_18278,N_16427);
or U22629 (N_22629,N_15930,N_19608);
and U22630 (N_22630,N_15800,N_15734);
xnor U22631 (N_22631,N_18048,N_15679);
and U22632 (N_22632,N_18906,N_16125);
and U22633 (N_22633,N_18592,N_15935);
xor U22634 (N_22634,N_19821,N_19915);
xnor U22635 (N_22635,N_16214,N_17846);
and U22636 (N_22636,N_15348,N_18752);
xnor U22637 (N_22637,N_16092,N_16127);
or U22638 (N_22638,N_19872,N_16035);
nand U22639 (N_22639,N_19727,N_16902);
and U22640 (N_22640,N_17261,N_19684);
xnor U22641 (N_22641,N_15374,N_16128);
or U22642 (N_22642,N_16132,N_19396);
nand U22643 (N_22643,N_16117,N_17955);
nand U22644 (N_22644,N_16783,N_17616);
and U22645 (N_22645,N_18263,N_19019);
nor U22646 (N_22646,N_18703,N_19079);
nand U22647 (N_22647,N_18069,N_18623);
or U22648 (N_22648,N_17908,N_16920);
xnor U22649 (N_22649,N_19443,N_17114);
xor U22650 (N_22650,N_17744,N_16027);
or U22651 (N_22651,N_15093,N_18871);
and U22652 (N_22652,N_16517,N_17510);
xnor U22653 (N_22653,N_18808,N_15526);
xnor U22654 (N_22654,N_16602,N_19739);
nor U22655 (N_22655,N_18543,N_17688);
xor U22656 (N_22656,N_16954,N_19565);
nand U22657 (N_22657,N_19244,N_16932);
xnor U22658 (N_22658,N_16184,N_15595);
and U22659 (N_22659,N_18351,N_19068);
or U22660 (N_22660,N_15990,N_17510);
nor U22661 (N_22661,N_19412,N_16295);
nand U22662 (N_22662,N_16045,N_16454);
nand U22663 (N_22663,N_17124,N_18438);
and U22664 (N_22664,N_16446,N_18694);
nor U22665 (N_22665,N_17914,N_17338);
nand U22666 (N_22666,N_18013,N_18813);
xor U22667 (N_22667,N_18800,N_15812);
nor U22668 (N_22668,N_18791,N_16932);
nor U22669 (N_22669,N_18758,N_15143);
nor U22670 (N_22670,N_15683,N_19257);
or U22671 (N_22671,N_16939,N_19950);
nand U22672 (N_22672,N_19177,N_17773);
and U22673 (N_22673,N_16706,N_16442);
xnor U22674 (N_22674,N_16218,N_16117);
and U22675 (N_22675,N_15606,N_16687);
nand U22676 (N_22676,N_16036,N_15898);
nor U22677 (N_22677,N_15115,N_18527);
nand U22678 (N_22678,N_19007,N_15072);
nand U22679 (N_22679,N_16375,N_17257);
nand U22680 (N_22680,N_17760,N_17567);
or U22681 (N_22681,N_17327,N_19970);
nor U22682 (N_22682,N_16574,N_19134);
and U22683 (N_22683,N_15984,N_18693);
and U22684 (N_22684,N_17340,N_16245);
xor U22685 (N_22685,N_19542,N_17752);
nand U22686 (N_22686,N_19794,N_19276);
nand U22687 (N_22687,N_17771,N_18398);
nor U22688 (N_22688,N_16653,N_15214);
nand U22689 (N_22689,N_18666,N_18753);
or U22690 (N_22690,N_15443,N_16076);
and U22691 (N_22691,N_15489,N_17481);
nor U22692 (N_22692,N_15052,N_15257);
nand U22693 (N_22693,N_15872,N_19838);
nor U22694 (N_22694,N_17928,N_18233);
nor U22695 (N_22695,N_17210,N_17309);
xor U22696 (N_22696,N_18442,N_17729);
nand U22697 (N_22697,N_18564,N_16790);
and U22698 (N_22698,N_15283,N_18391);
nand U22699 (N_22699,N_15157,N_18991);
xnor U22700 (N_22700,N_17482,N_15253);
and U22701 (N_22701,N_19787,N_16949);
xor U22702 (N_22702,N_15571,N_18372);
or U22703 (N_22703,N_19948,N_16827);
nor U22704 (N_22704,N_19130,N_15284);
xnor U22705 (N_22705,N_17532,N_18501);
nor U22706 (N_22706,N_16593,N_15199);
or U22707 (N_22707,N_16570,N_15023);
nor U22708 (N_22708,N_19458,N_15408);
nand U22709 (N_22709,N_17907,N_15544);
nor U22710 (N_22710,N_16385,N_15569);
and U22711 (N_22711,N_19561,N_16059);
or U22712 (N_22712,N_16829,N_15111);
and U22713 (N_22713,N_18422,N_17708);
nor U22714 (N_22714,N_19700,N_18337);
or U22715 (N_22715,N_16118,N_17587);
and U22716 (N_22716,N_18216,N_17641);
nor U22717 (N_22717,N_16110,N_16226);
nand U22718 (N_22718,N_15311,N_15728);
and U22719 (N_22719,N_16892,N_15227);
nor U22720 (N_22720,N_16651,N_19142);
or U22721 (N_22721,N_16549,N_17410);
xor U22722 (N_22722,N_18646,N_17033);
nand U22723 (N_22723,N_16085,N_17413);
or U22724 (N_22724,N_18159,N_18815);
xnor U22725 (N_22725,N_19319,N_18957);
nand U22726 (N_22726,N_17963,N_16954);
and U22727 (N_22727,N_15866,N_19583);
or U22728 (N_22728,N_19386,N_15584);
or U22729 (N_22729,N_15314,N_18503);
nand U22730 (N_22730,N_17771,N_16716);
xor U22731 (N_22731,N_16099,N_17004);
xor U22732 (N_22732,N_18218,N_19960);
nor U22733 (N_22733,N_15901,N_17175);
and U22734 (N_22734,N_17423,N_16310);
xor U22735 (N_22735,N_16979,N_19418);
xor U22736 (N_22736,N_19862,N_17233);
nor U22737 (N_22737,N_19511,N_16589);
nor U22738 (N_22738,N_18173,N_19693);
and U22739 (N_22739,N_16125,N_16858);
or U22740 (N_22740,N_15166,N_16342);
and U22741 (N_22741,N_17646,N_18042);
xor U22742 (N_22742,N_15779,N_15851);
nand U22743 (N_22743,N_19408,N_17619);
nand U22744 (N_22744,N_16756,N_17048);
nand U22745 (N_22745,N_18205,N_19088);
nor U22746 (N_22746,N_17839,N_19558);
and U22747 (N_22747,N_16844,N_19594);
and U22748 (N_22748,N_16289,N_19949);
xnor U22749 (N_22749,N_18063,N_16736);
nand U22750 (N_22750,N_15951,N_17514);
nor U22751 (N_22751,N_16552,N_15192);
xor U22752 (N_22752,N_16043,N_15123);
xor U22753 (N_22753,N_16765,N_17837);
and U22754 (N_22754,N_19246,N_15228);
nand U22755 (N_22755,N_16246,N_15201);
xnor U22756 (N_22756,N_17903,N_15802);
nand U22757 (N_22757,N_16047,N_15810);
nor U22758 (N_22758,N_16822,N_19979);
or U22759 (N_22759,N_18757,N_19482);
and U22760 (N_22760,N_19697,N_17494);
or U22761 (N_22761,N_19149,N_15762);
or U22762 (N_22762,N_19290,N_15682);
or U22763 (N_22763,N_17770,N_15727);
nor U22764 (N_22764,N_19992,N_16816);
and U22765 (N_22765,N_15598,N_19097);
xor U22766 (N_22766,N_15467,N_19377);
or U22767 (N_22767,N_16009,N_17370);
and U22768 (N_22768,N_16292,N_19910);
nand U22769 (N_22769,N_17294,N_17022);
xor U22770 (N_22770,N_15931,N_15675);
nor U22771 (N_22771,N_17945,N_16176);
xor U22772 (N_22772,N_17464,N_17764);
nor U22773 (N_22773,N_15996,N_16640);
or U22774 (N_22774,N_15573,N_17974);
or U22775 (N_22775,N_18651,N_16020);
and U22776 (N_22776,N_19274,N_19384);
xnor U22777 (N_22777,N_17119,N_19390);
or U22778 (N_22778,N_18186,N_19967);
or U22779 (N_22779,N_17028,N_18999);
nor U22780 (N_22780,N_15123,N_19431);
or U22781 (N_22781,N_17242,N_19599);
nand U22782 (N_22782,N_19681,N_15355);
nor U22783 (N_22783,N_19791,N_19824);
nor U22784 (N_22784,N_17837,N_17885);
or U22785 (N_22785,N_18308,N_17646);
or U22786 (N_22786,N_19165,N_15999);
or U22787 (N_22787,N_17776,N_15657);
xnor U22788 (N_22788,N_15252,N_17224);
nor U22789 (N_22789,N_19550,N_16788);
and U22790 (N_22790,N_19173,N_16249);
nor U22791 (N_22791,N_15352,N_19382);
nand U22792 (N_22792,N_15925,N_15717);
xnor U22793 (N_22793,N_15336,N_17278);
or U22794 (N_22794,N_16324,N_18297);
nand U22795 (N_22795,N_18783,N_18545);
or U22796 (N_22796,N_19722,N_18286);
nor U22797 (N_22797,N_16568,N_15964);
or U22798 (N_22798,N_15155,N_16821);
nor U22799 (N_22799,N_17853,N_15468);
nand U22800 (N_22800,N_16530,N_16269);
or U22801 (N_22801,N_19221,N_17125);
nand U22802 (N_22802,N_15201,N_18113);
and U22803 (N_22803,N_18872,N_17340);
and U22804 (N_22804,N_18289,N_18413);
or U22805 (N_22805,N_19091,N_17328);
nand U22806 (N_22806,N_15698,N_19434);
nand U22807 (N_22807,N_15007,N_15571);
or U22808 (N_22808,N_17020,N_19711);
and U22809 (N_22809,N_16109,N_15547);
and U22810 (N_22810,N_15278,N_17072);
and U22811 (N_22811,N_16521,N_16193);
nand U22812 (N_22812,N_19031,N_17937);
nand U22813 (N_22813,N_16774,N_18156);
xnor U22814 (N_22814,N_17355,N_16696);
xnor U22815 (N_22815,N_17223,N_15018);
xor U22816 (N_22816,N_15787,N_16896);
xnor U22817 (N_22817,N_16781,N_19153);
and U22818 (N_22818,N_18057,N_18280);
nor U22819 (N_22819,N_17548,N_15595);
nor U22820 (N_22820,N_16578,N_15707);
nor U22821 (N_22821,N_19115,N_18498);
nor U22822 (N_22822,N_19800,N_15086);
nor U22823 (N_22823,N_17785,N_15315);
or U22824 (N_22824,N_19179,N_19308);
nor U22825 (N_22825,N_19405,N_17512);
nor U22826 (N_22826,N_19608,N_18258);
and U22827 (N_22827,N_17499,N_19985);
nand U22828 (N_22828,N_19418,N_17502);
nor U22829 (N_22829,N_15243,N_15981);
nand U22830 (N_22830,N_15250,N_18739);
xnor U22831 (N_22831,N_17238,N_19441);
nor U22832 (N_22832,N_18126,N_19095);
or U22833 (N_22833,N_18890,N_19980);
nor U22834 (N_22834,N_16086,N_16455);
or U22835 (N_22835,N_17127,N_15188);
or U22836 (N_22836,N_16729,N_16635);
nor U22837 (N_22837,N_15577,N_16660);
nor U22838 (N_22838,N_15277,N_18812);
xor U22839 (N_22839,N_19142,N_16689);
nor U22840 (N_22840,N_15507,N_16950);
and U22841 (N_22841,N_19756,N_19035);
xor U22842 (N_22842,N_16249,N_18357);
and U22843 (N_22843,N_18118,N_17456);
nor U22844 (N_22844,N_15827,N_19287);
and U22845 (N_22845,N_15863,N_18712);
nor U22846 (N_22846,N_17736,N_17326);
xnor U22847 (N_22847,N_19173,N_15233);
and U22848 (N_22848,N_15248,N_17763);
or U22849 (N_22849,N_16544,N_19262);
nand U22850 (N_22850,N_16674,N_18634);
and U22851 (N_22851,N_19295,N_16404);
and U22852 (N_22852,N_17634,N_18453);
and U22853 (N_22853,N_17222,N_18390);
and U22854 (N_22854,N_18826,N_19173);
and U22855 (N_22855,N_19878,N_16682);
nor U22856 (N_22856,N_17078,N_15062);
or U22857 (N_22857,N_17757,N_17570);
or U22858 (N_22858,N_17727,N_15782);
and U22859 (N_22859,N_17988,N_16343);
xor U22860 (N_22860,N_16302,N_18464);
nor U22861 (N_22861,N_18963,N_17628);
xnor U22862 (N_22862,N_15348,N_18865);
xor U22863 (N_22863,N_16614,N_18994);
nor U22864 (N_22864,N_18002,N_19242);
nand U22865 (N_22865,N_19758,N_16068);
and U22866 (N_22866,N_19785,N_19463);
or U22867 (N_22867,N_17566,N_15213);
or U22868 (N_22868,N_19964,N_15356);
and U22869 (N_22869,N_18975,N_17942);
nor U22870 (N_22870,N_19371,N_16312);
and U22871 (N_22871,N_15257,N_15193);
nor U22872 (N_22872,N_17336,N_16335);
or U22873 (N_22873,N_19788,N_19793);
or U22874 (N_22874,N_19833,N_19585);
and U22875 (N_22875,N_19152,N_18058);
and U22876 (N_22876,N_19416,N_18816);
nand U22877 (N_22877,N_18120,N_15961);
xnor U22878 (N_22878,N_17207,N_16990);
xor U22879 (N_22879,N_15324,N_18668);
nor U22880 (N_22880,N_16412,N_19256);
nor U22881 (N_22881,N_16713,N_17713);
xnor U22882 (N_22882,N_15321,N_15574);
nand U22883 (N_22883,N_18417,N_19971);
nand U22884 (N_22884,N_15152,N_17449);
nor U22885 (N_22885,N_18428,N_19261);
and U22886 (N_22886,N_19527,N_16290);
nand U22887 (N_22887,N_19810,N_16838);
nor U22888 (N_22888,N_17727,N_19220);
xor U22889 (N_22889,N_19037,N_15396);
and U22890 (N_22890,N_19503,N_19186);
or U22891 (N_22891,N_16826,N_18667);
or U22892 (N_22892,N_19270,N_18692);
nor U22893 (N_22893,N_17058,N_19018);
nand U22894 (N_22894,N_18333,N_18165);
nor U22895 (N_22895,N_19813,N_15703);
nor U22896 (N_22896,N_17898,N_19749);
and U22897 (N_22897,N_15760,N_17063);
xor U22898 (N_22898,N_17694,N_17001);
and U22899 (N_22899,N_19411,N_15069);
nand U22900 (N_22900,N_17113,N_18907);
xor U22901 (N_22901,N_17208,N_18807);
and U22902 (N_22902,N_19802,N_16261);
xor U22903 (N_22903,N_18145,N_19801);
and U22904 (N_22904,N_15881,N_15499);
xnor U22905 (N_22905,N_17304,N_18975);
or U22906 (N_22906,N_16869,N_18836);
or U22907 (N_22907,N_16819,N_16390);
nor U22908 (N_22908,N_15188,N_15504);
xor U22909 (N_22909,N_15941,N_17597);
and U22910 (N_22910,N_19592,N_15814);
or U22911 (N_22911,N_16944,N_18845);
nor U22912 (N_22912,N_16444,N_17156);
nor U22913 (N_22913,N_17082,N_17383);
or U22914 (N_22914,N_17288,N_18792);
nor U22915 (N_22915,N_18579,N_16235);
xnor U22916 (N_22916,N_16484,N_16938);
nor U22917 (N_22917,N_16820,N_16821);
or U22918 (N_22918,N_19256,N_16521);
xor U22919 (N_22919,N_17512,N_18274);
xor U22920 (N_22920,N_19740,N_16594);
nand U22921 (N_22921,N_17607,N_16001);
xor U22922 (N_22922,N_18883,N_16835);
and U22923 (N_22923,N_16827,N_15594);
nand U22924 (N_22924,N_16435,N_19395);
nand U22925 (N_22925,N_16760,N_16701);
and U22926 (N_22926,N_17571,N_18214);
nand U22927 (N_22927,N_17756,N_19650);
nor U22928 (N_22928,N_15086,N_17183);
or U22929 (N_22929,N_18166,N_19619);
nand U22930 (N_22930,N_15654,N_16958);
nor U22931 (N_22931,N_15047,N_19216);
or U22932 (N_22932,N_19699,N_19089);
nor U22933 (N_22933,N_16163,N_19303);
xnor U22934 (N_22934,N_16418,N_15438);
and U22935 (N_22935,N_16446,N_19390);
nor U22936 (N_22936,N_19344,N_15669);
xnor U22937 (N_22937,N_19527,N_17946);
and U22938 (N_22938,N_19892,N_18671);
xnor U22939 (N_22939,N_15032,N_15540);
or U22940 (N_22940,N_19712,N_17521);
nand U22941 (N_22941,N_16292,N_18570);
or U22942 (N_22942,N_19435,N_19604);
nand U22943 (N_22943,N_19530,N_16461);
nor U22944 (N_22944,N_16111,N_15412);
nor U22945 (N_22945,N_19057,N_17065);
nor U22946 (N_22946,N_16950,N_17547);
nor U22947 (N_22947,N_15136,N_17558);
and U22948 (N_22948,N_15725,N_17687);
or U22949 (N_22949,N_15619,N_17464);
xnor U22950 (N_22950,N_16712,N_15629);
nand U22951 (N_22951,N_16069,N_16301);
or U22952 (N_22952,N_19586,N_16956);
or U22953 (N_22953,N_17753,N_15367);
nor U22954 (N_22954,N_15636,N_15327);
or U22955 (N_22955,N_19458,N_18475);
nand U22956 (N_22956,N_19644,N_19070);
nor U22957 (N_22957,N_17921,N_17517);
or U22958 (N_22958,N_18501,N_18808);
xor U22959 (N_22959,N_15748,N_19763);
and U22960 (N_22960,N_17730,N_17674);
nand U22961 (N_22961,N_18061,N_16970);
nand U22962 (N_22962,N_19970,N_18007);
xnor U22963 (N_22963,N_16350,N_15802);
or U22964 (N_22964,N_18555,N_17551);
nor U22965 (N_22965,N_17752,N_16426);
nor U22966 (N_22966,N_18144,N_19796);
nand U22967 (N_22967,N_17707,N_16711);
nor U22968 (N_22968,N_16390,N_19564);
nor U22969 (N_22969,N_18438,N_16782);
or U22970 (N_22970,N_19752,N_17623);
or U22971 (N_22971,N_16428,N_15312);
and U22972 (N_22972,N_15359,N_16827);
nand U22973 (N_22973,N_18591,N_19935);
nor U22974 (N_22974,N_18027,N_19139);
nor U22975 (N_22975,N_17556,N_16583);
and U22976 (N_22976,N_19569,N_15185);
and U22977 (N_22977,N_19764,N_19668);
xor U22978 (N_22978,N_15148,N_19725);
and U22979 (N_22979,N_19504,N_19429);
xor U22980 (N_22980,N_18260,N_18893);
nor U22981 (N_22981,N_18937,N_19454);
nand U22982 (N_22982,N_19773,N_18679);
or U22983 (N_22983,N_19562,N_17863);
and U22984 (N_22984,N_19813,N_15592);
nor U22985 (N_22985,N_15543,N_16936);
xor U22986 (N_22986,N_15493,N_17449);
nor U22987 (N_22987,N_17018,N_18288);
and U22988 (N_22988,N_18787,N_17112);
xnor U22989 (N_22989,N_17384,N_18122);
xor U22990 (N_22990,N_15865,N_17870);
nand U22991 (N_22991,N_19051,N_19951);
or U22992 (N_22992,N_17530,N_19925);
xnor U22993 (N_22993,N_18192,N_17018);
xor U22994 (N_22994,N_18877,N_17020);
nand U22995 (N_22995,N_16524,N_19052);
and U22996 (N_22996,N_19523,N_19333);
and U22997 (N_22997,N_19195,N_19587);
nor U22998 (N_22998,N_16387,N_15695);
nand U22999 (N_22999,N_17011,N_18767);
xnor U23000 (N_23000,N_16487,N_17224);
xor U23001 (N_23001,N_18632,N_19024);
nand U23002 (N_23002,N_17882,N_16144);
xnor U23003 (N_23003,N_15967,N_19073);
xnor U23004 (N_23004,N_16740,N_19952);
or U23005 (N_23005,N_19233,N_19335);
or U23006 (N_23006,N_16787,N_16489);
nor U23007 (N_23007,N_15650,N_18657);
or U23008 (N_23008,N_17536,N_15457);
and U23009 (N_23009,N_19418,N_16239);
xnor U23010 (N_23010,N_15738,N_16356);
nand U23011 (N_23011,N_18494,N_17518);
or U23012 (N_23012,N_19454,N_16208);
and U23013 (N_23013,N_16037,N_17976);
nor U23014 (N_23014,N_19274,N_18028);
nor U23015 (N_23015,N_17412,N_19636);
and U23016 (N_23016,N_19424,N_17445);
or U23017 (N_23017,N_16908,N_19454);
nand U23018 (N_23018,N_16438,N_18579);
and U23019 (N_23019,N_17925,N_17598);
and U23020 (N_23020,N_16329,N_19560);
nand U23021 (N_23021,N_19832,N_17657);
and U23022 (N_23022,N_18524,N_16032);
and U23023 (N_23023,N_19370,N_15482);
xnor U23024 (N_23024,N_19740,N_17765);
or U23025 (N_23025,N_19755,N_18676);
nor U23026 (N_23026,N_16627,N_17935);
and U23027 (N_23027,N_16466,N_19479);
nor U23028 (N_23028,N_16946,N_19239);
xnor U23029 (N_23029,N_16368,N_15163);
xor U23030 (N_23030,N_19859,N_17278);
nand U23031 (N_23031,N_16310,N_16975);
xor U23032 (N_23032,N_19463,N_16148);
nor U23033 (N_23033,N_15530,N_15442);
nor U23034 (N_23034,N_18866,N_18057);
nand U23035 (N_23035,N_16975,N_19620);
nor U23036 (N_23036,N_18732,N_18151);
nand U23037 (N_23037,N_19402,N_19120);
xor U23038 (N_23038,N_19627,N_15585);
and U23039 (N_23039,N_19313,N_15730);
nand U23040 (N_23040,N_17479,N_19840);
or U23041 (N_23041,N_15076,N_18589);
nand U23042 (N_23042,N_17312,N_18930);
xnor U23043 (N_23043,N_16666,N_18865);
nand U23044 (N_23044,N_17994,N_17006);
and U23045 (N_23045,N_16859,N_18119);
nor U23046 (N_23046,N_19715,N_18562);
nor U23047 (N_23047,N_16494,N_15640);
nor U23048 (N_23048,N_15252,N_16022);
nor U23049 (N_23049,N_18800,N_19076);
nand U23050 (N_23050,N_16181,N_18589);
nand U23051 (N_23051,N_17430,N_18483);
nor U23052 (N_23052,N_19114,N_15835);
and U23053 (N_23053,N_18267,N_19351);
nand U23054 (N_23054,N_15213,N_16898);
xor U23055 (N_23055,N_16286,N_19783);
nor U23056 (N_23056,N_15772,N_15660);
nand U23057 (N_23057,N_16676,N_15613);
nand U23058 (N_23058,N_15461,N_18534);
or U23059 (N_23059,N_15134,N_15681);
nor U23060 (N_23060,N_15141,N_16127);
nor U23061 (N_23061,N_19388,N_15984);
nand U23062 (N_23062,N_18729,N_16356);
or U23063 (N_23063,N_16016,N_16894);
and U23064 (N_23064,N_17116,N_19915);
or U23065 (N_23065,N_19409,N_15770);
and U23066 (N_23066,N_18206,N_19948);
nor U23067 (N_23067,N_17028,N_19547);
and U23068 (N_23068,N_15136,N_16737);
nor U23069 (N_23069,N_17827,N_19663);
nor U23070 (N_23070,N_17597,N_18029);
nor U23071 (N_23071,N_15944,N_19537);
nand U23072 (N_23072,N_18536,N_17848);
nand U23073 (N_23073,N_18196,N_15991);
or U23074 (N_23074,N_15026,N_19586);
xor U23075 (N_23075,N_19643,N_16679);
or U23076 (N_23076,N_16537,N_16594);
nand U23077 (N_23077,N_16876,N_17369);
xnor U23078 (N_23078,N_18279,N_19177);
or U23079 (N_23079,N_18498,N_17768);
nand U23080 (N_23080,N_17296,N_16314);
nand U23081 (N_23081,N_15476,N_17324);
or U23082 (N_23082,N_18306,N_18531);
xnor U23083 (N_23083,N_18766,N_17463);
xnor U23084 (N_23084,N_19729,N_19191);
nand U23085 (N_23085,N_18489,N_15910);
nor U23086 (N_23086,N_15496,N_17624);
or U23087 (N_23087,N_17939,N_18791);
and U23088 (N_23088,N_18192,N_15709);
and U23089 (N_23089,N_16003,N_16627);
xnor U23090 (N_23090,N_17052,N_19811);
xor U23091 (N_23091,N_18939,N_15170);
xnor U23092 (N_23092,N_15265,N_16892);
or U23093 (N_23093,N_15927,N_16603);
or U23094 (N_23094,N_18423,N_19201);
nand U23095 (N_23095,N_19830,N_16250);
nand U23096 (N_23096,N_16300,N_16389);
or U23097 (N_23097,N_19838,N_16933);
nand U23098 (N_23098,N_18645,N_17358);
nor U23099 (N_23099,N_16996,N_16199);
nor U23100 (N_23100,N_16532,N_16030);
and U23101 (N_23101,N_17671,N_16418);
nand U23102 (N_23102,N_15095,N_19361);
and U23103 (N_23103,N_19602,N_16990);
nor U23104 (N_23104,N_17851,N_15124);
nand U23105 (N_23105,N_16038,N_18083);
nand U23106 (N_23106,N_17617,N_17553);
and U23107 (N_23107,N_16411,N_17233);
nand U23108 (N_23108,N_19541,N_17800);
nand U23109 (N_23109,N_19530,N_16733);
xnor U23110 (N_23110,N_16529,N_18229);
and U23111 (N_23111,N_19091,N_18164);
nand U23112 (N_23112,N_16896,N_18291);
or U23113 (N_23113,N_17831,N_19813);
and U23114 (N_23114,N_15142,N_16727);
nor U23115 (N_23115,N_18930,N_15306);
nor U23116 (N_23116,N_16472,N_19773);
nor U23117 (N_23117,N_19346,N_18203);
nor U23118 (N_23118,N_16048,N_17401);
nand U23119 (N_23119,N_16467,N_19921);
xnor U23120 (N_23120,N_18067,N_16238);
xor U23121 (N_23121,N_15320,N_18835);
nand U23122 (N_23122,N_15012,N_15590);
xor U23123 (N_23123,N_17031,N_18852);
nand U23124 (N_23124,N_17531,N_16893);
nand U23125 (N_23125,N_16906,N_17564);
xor U23126 (N_23126,N_19635,N_15068);
and U23127 (N_23127,N_18992,N_16116);
nand U23128 (N_23128,N_17989,N_18741);
nand U23129 (N_23129,N_15891,N_17933);
xnor U23130 (N_23130,N_16588,N_17439);
and U23131 (N_23131,N_17395,N_16339);
nand U23132 (N_23132,N_19529,N_15831);
and U23133 (N_23133,N_16790,N_16973);
nand U23134 (N_23134,N_18444,N_15503);
nand U23135 (N_23135,N_17501,N_17741);
and U23136 (N_23136,N_19566,N_15861);
and U23137 (N_23137,N_15239,N_18072);
nand U23138 (N_23138,N_19484,N_16872);
xor U23139 (N_23139,N_15154,N_16883);
nand U23140 (N_23140,N_18650,N_19683);
xnor U23141 (N_23141,N_19986,N_19109);
and U23142 (N_23142,N_19517,N_19784);
nor U23143 (N_23143,N_16564,N_16114);
or U23144 (N_23144,N_17487,N_18542);
nand U23145 (N_23145,N_15165,N_19391);
or U23146 (N_23146,N_15933,N_15250);
and U23147 (N_23147,N_19810,N_15053);
nand U23148 (N_23148,N_15569,N_16570);
and U23149 (N_23149,N_18461,N_17623);
and U23150 (N_23150,N_18254,N_19078);
nand U23151 (N_23151,N_17023,N_19139);
xnor U23152 (N_23152,N_18893,N_16824);
and U23153 (N_23153,N_19468,N_19787);
nand U23154 (N_23154,N_17188,N_19243);
or U23155 (N_23155,N_19713,N_19448);
or U23156 (N_23156,N_15263,N_17991);
or U23157 (N_23157,N_18578,N_18078);
nand U23158 (N_23158,N_16523,N_18925);
and U23159 (N_23159,N_16699,N_16001);
or U23160 (N_23160,N_17724,N_18715);
and U23161 (N_23161,N_18686,N_16142);
nand U23162 (N_23162,N_15223,N_19327);
and U23163 (N_23163,N_18113,N_19274);
or U23164 (N_23164,N_19912,N_19637);
nor U23165 (N_23165,N_19032,N_18349);
or U23166 (N_23166,N_18299,N_16278);
or U23167 (N_23167,N_19193,N_15470);
nand U23168 (N_23168,N_15962,N_18295);
xor U23169 (N_23169,N_15609,N_15619);
nor U23170 (N_23170,N_17756,N_15944);
and U23171 (N_23171,N_17311,N_16177);
xor U23172 (N_23172,N_15302,N_17325);
nand U23173 (N_23173,N_16570,N_15608);
and U23174 (N_23174,N_17413,N_16027);
nor U23175 (N_23175,N_15064,N_15027);
xor U23176 (N_23176,N_19029,N_15118);
nand U23177 (N_23177,N_18791,N_18642);
and U23178 (N_23178,N_15976,N_16857);
nand U23179 (N_23179,N_15418,N_19549);
xnor U23180 (N_23180,N_18233,N_15605);
or U23181 (N_23181,N_18397,N_18328);
nand U23182 (N_23182,N_17542,N_17814);
or U23183 (N_23183,N_15136,N_16402);
xnor U23184 (N_23184,N_17442,N_18565);
and U23185 (N_23185,N_15746,N_15810);
and U23186 (N_23186,N_16473,N_15123);
nand U23187 (N_23187,N_15029,N_17585);
or U23188 (N_23188,N_15255,N_17578);
xor U23189 (N_23189,N_18030,N_18999);
nor U23190 (N_23190,N_15045,N_19797);
xnor U23191 (N_23191,N_19697,N_18186);
xnor U23192 (N_23192,N_18199,N_15570);
and U23193 (N_23193,N_18513,N_17682);
nor U23194 (N_23194,N_18980,N_17270);
nand U23195 (N_23195,N_16942,N_19875);
and U23196 (N_23196,N_17709,N_16297);
xnor U23197 (N_23197,N_18572,N_17360);
nand U23198 (N_23198,N_16797,N_18413);
nand U23199 (N_23199,N_17875,N_19112);
and U23200 (N_23200,N_19257,N_18559);
nor U23201 (N_23201,N_16009,N_17637);
xnor U23202 (N_23202,N_16504,N_15794);
or U23203 (N_23203,N_19807,N_16968);
and U23204 (N_23204,N_16359,N_15603);
xnor U23205 (N_23205,N_19925,N_16773);
or U23206 (N_23206,N_16991,N_18849);
or U23207 (N_23207,N_16077,N_19592);
or U23208 (N_23208,N_17647,N_19950);
nand U23209 (N_23209,N_18263,N_19186);
or U23210 (N_23210,N_17721,N_16739);
xor U23211 (N_23211,N_19966,N_16983);
nor U23212 (N_23212,N_16113,N_16427);
nand U23213 (N_23213,N_15532,N_17868);
nand U23214 (N_23214,N_19443,N_19529);
xor U23215 (N_23215,N_16201,N_19268);
or U23216 (N_23216,N_18707,N_17345);
or U23217 (N_23217,N_16798,N_16030);
nand U23218 (N_23218,N_19363,N_19087);
nand U23219 (N_23219,N_18156,N_19337);
and U23220 (N_23220,N_18438,N_18974);
nand U23221 (N_23221,N_16573,N_17047);
nand U23222 (N_23222,N_17583,N_17761);
xor U23223 (N_23223,N_18730,N_18321);
and U23224 (N_23224,N_18899,N_16344);
or U23225 (N_23225,N_15726,N_19372);
or U23226 (N_23226,N_15618,N_15007);
and U23227 (N_23227,N_18482,N_19148);
nand U23228 (N_23228,N_15075,N_17106);
nor U23229 (N_23229,N_16018,N_19534);
or U23230 (N_23230,N_16418,N_15225);
nand U23231 (N_23231,N_17283,N_19754);
or U23232 (N_23232,N_16505,N_19519);
or U23233 (N_23233,N_15707,N_18384);
xor U23234 (N_23234,N_16753,N_18072);
or U23235 (N_23235,N_16586,N_15390);
xor U23236 (N_23236,N_15837,N_15852);
and U23237 (N_23237,N_15550,N_16615);
and U23238 (N_23238,N_16268,N_17641);
or U23239 (N_23239,N_16009,N_18130);
nor U23240 (N_23240,N_15611,N_19916);
xnor U23241 (N_23241,N_18932,N_16502);
and U23242 (N_23242,N_19165,N_16120);
and U23243 (N_23243,N_17464,N_16880);
nand U23244 (N_23244,N_16253,N_15440);
nor U23245 (N_23245,N_16182,N_19647);
and U23246 (N_23246,N_15022,N_17647);
and U23247 (N_23247,N_15161,N_18660);
xor U23248 (N_23248,N_16934,N_19168);
xor U23249 (N_23249,N_17126,N_19456);
nand U23250 (N_23250,N_18618,N_15199);
nand U23251 (N_23251,N_19398,N_15745);
and U23252 (N_23252,N_16567,N_18117);
and U23253 (N_23253,N_16342,N_15256);
nand U23254 (N_23254,N_18780,N_15065);
xnor U23255 (N_23255,N_17559,N_15713);
nand U23256 (N_23256,N_19314,N_15345);
xnor U23257 (N_23257,N_18983,N_19200);
nand U23258 (N_23258,N_19858,N_18996);
nor U23259 (N_23259,N_19907,N_15294);
and U23260 (N_23260,N_18422,N_15800);
xnor U23261 (N_23261,N_18855,N_17921);
nor U23262 (N_23262,N_16691,N_18961);
nor U23263 (N_23263,N_16137,N_19008);
xnor U23264 (N_23264,N_19614,N_17274);
or U23265 (N_23265,N_19666,N_17125);
nand U23266 (N_23266,N_16777,N_19828);
and U23267 (N_23267,N_18213,N_16191);
nor U23268 (N_23268,N_15464,N_19998);
nor U23269 (N_23269,N_17685,N_17788);
nand U23270 (N_23270,N_19508,N_17544);
xnor U23271 (N_23271,N_18026,N_18627);
and U23272 (N_23272,N_15243,N_18557);
or U23273 (N_23273,N_17872,N_15582);
or U23274 (N_23274,N_17597,N_19925);
or U23275 (N_23275,N_17077,N_15877);
nor U23276 (N_23276,N_18616,N_16564);
xnor U23277 (N_23277,N_15178,N_19999);
and U23278 (N_23278,N_18561,N_19589);
and U23279 (N_23279,N_17399,N_16241);
nand U23280 (N_23280,N_17160,N_17777);
or U23281 (N_23281,N_15311,N_16731);
or U23282 (N_23282,N_16442,N_18276);
and U23283 (N_23283,N_17520,N_16899);
nor U23284 (N_23284,N_19373,N_19545);
nor U23285 (N_23285,N_18460,N_17120);
or U23286 (N_23286,N_16042,N_15041);
nor U23287 (N_23287,N_19324,N_19263);
xnor U23288 (N_23288,N_15254,N_15310);
or U23289 (N_23289,N_18718,N_16999);
and U23290 (N_23290,N_17091,N_15742);
or U23291 (N_23291,N_15188,N_18386);
and U23292 (N_23292,N_18253,N_18303);
nor U23293 (N_23293,N_17035,N_18222);
xnor U23294 (N_23294,N_15927,N_15019);
nand U23295 (N_23295,N_17700,N_19428);
xor U23296 (N_23296,N_18723,N_17498);
xnor U23297 (N_23297,N_17851,N_17952);
or U23298 (N_23298,N_16884,N_15585);
nand U23299 (N_23299,N_16267,N_15437);
or U23300 (N_23300,N_15460,N_15231);
and U23301 (N_23301,N_18835,N_19274);
nand U23302 (N_23302,N_19795,N_18653);
nor U23303 (N_23303,N_18130,N_16145);
or U23304 (N_23304,N_17072,N_18881);
and U23305 (N_23305,N_19060,N_15938);
xnor U23306 (N_23306,N_15431,N_19313);
or U23307 (N_23307,N_19267,N_16385);
nand U23308 (N_23308,N_16584,N_17579);
or U23309 (N_23309,N_15061,N_19992);
nor U23310 (N_23310,N_19152,N_19718);
nand U23311 (N_23311,N_19413,N_17530);
nor U23312 (N_23312,N_17195,N_19979);
nor U23313 (N_23313,N_19382,N_17809);
nor U23314 (N_23314,N_15211,N_19108);
or U23315 (N_23315,N_18951,N_15654);
nor U23316 (N_23316,N_19902,N_16761);
nor U23317 (N_23317,N_17896,N_18075);
xor U23318 (N_23318,N_15380,N_17067);
xnor U23319 (N_23319,N_15211,N_18522);
or U23320 (N_23320,N_17461,N_15618);
nand U23321 (N_23321,N_18230,N_19680);
and U23322 (N_23322,N_15812,N_18597);
or U23323 (N_23323,N_18928,N_15469);
nor U23324 (N_23324,N_16241,N_15797);
or U23325 (N_23325,N_17597,N_18322);
xor U23326 (N_23326,N_15955,N_17871);
xnor U23327 (N_23327,N_15536,N_16891);
xor U23328 (N_23328,N_17788,N_16004);
or U23329 (N_23329,N_17879,N_16117);
xnor U23330 (N_23330,N_17582,N_19128);
xor U23331 (N_23331,N_17893,N_15004);
xor U23332 (N_23332,N_16767,N_19274);
or U23333 (N_23333,N_19561,N_17007);
or U23334 (N_23334,N_16528,N_18170);
and U23335 (N_23335,N_17581,N_17773);
and U23336 (N_23336,N_17871,N_16308);
and U23337 (N_23337,N_18619,N_19052);
and U23338 (N_23338,N_17061,N_17385);
or U23339 (N_23339,N_18409,N_15408);
or U23340 (N_23340,N_17751,N_16842);
xnor U23341 (N_23341,N_18543,N_18646);
nor U23342 (N_23342,N_19944,N_18857);
nor U23343 (N_23343,N_17519,N_19425);
xor U23344 (N_23344,N_16580,N_16079);
or U23345 (N_23345,N_18743,N_19096);
or U23346 (N_23346,N_16372,N_19626);
nor U23347 (N_23347,N_19377,N_18041);
nor U23348 (N_23348,N_17933,N_19206);
or U23349 (N_23349,N_19269,N_16983);
or U23350 (N_23350,N_16920,N_15280);
and U23351 (N_23351,N_18464,N_18421);
xnor U23352 (N_23352,N_19750,N_19540);
and U23353 (N_23353,N_18667,N_17179);
xor U23354 (N_23354,N_17479,N_16565);
xnor U23355 (N_23355,N_18493,N_17672);
and U23356 (N_23356,N_18112,N_17868);
nand U23357 (N_23357,N_15437,N_19458);
xnor U23358 (N_23358,N_19920,N_17257);
nand U23359 (N_23359,N_18189,N_17179);
and U23360 (N_23360,N_19569,N_16098);
xnor U23361 (N_23361,N_18205,N_19986);
and U23362 (N_23362,N_17122,N_18920);
or U23363 (N_23363,N_18685,N_18082);
nand U23364 (N_23364,N_18289,N_17948);
xnor U23365 (N_23365,N_19735,N_15617);
or U23366 (N_23366,N_16342,N_19740);
xor U23367 (N_23367,N_16296,N_16354);
or U23368 (N_23368,N_18877,N_15378);
xnor U23369 (N_23369,N_19422,N_19837);
or U23370 (N_23370,N_17600,N_16208);
nor U23371 (N_23371,N_15846,N_16866);
xor U23372 (N_23372,N_17938,N_18058);
nor U23373 (N_23373,N_15259,N_19211);
and U23374 (N_23374,N_18122,N_19993);
and U23375 (N_23375,N_15216,N_15494);
nand U23376 (N_23376,N_15210,N_16438);
nor U23377 (N_23377,N_18249,N_19266);
nand U23378 (N_23378,N_16476,N_16041);
xnor U23379 (N_23379,N_19696,N_16194);
nand U23380 (N_23380,N_17574,N_17379);
nand U23381 (N_23381,N_19112,N_16118);
nand U23382 (N_23382,N_19577,N_15851);
and U23383 (N_23383,N_18138,N_15027);
nor U23384 (N_23384,N_17414,N_19725);
nor U23385 (N_23385,N_17645,N_17371);
xor U23386 (N_23386,N_16782,N_16728);
nor U23387 (N_23387,N_17653,N_16039);
nand U23388 (N_23388,N_19574,N_16908);
and U23389 (N_23389,N_15800,N_15473);
nor U23390 (N_23390,N_19314,N_16784);
nand U23391 (N_23391,N_17000,N_15342);
xor U23392 (N_23392,N_16779,N_17690);
and U23393 (N_23393,N_18683,N_19261);
xor U23394 (N_23394,N_16536,N_15774);
nor U23395 (N_23395,N_16537,N_17454);
or U23396 (N_23396,N_15049,N_16823);
nand U23397 (N_23397,N_17749,N_16236);
and U23398 (N_23398,N_17002,N_15413);
xor U23399 (N_23399,N_19671,N_19077);
and U23400 (N_23400,N_17938,N_19335);
and U23401 (N_23401,N_15458,N_19635);
xnor U23402 (N_23402,N_19468,N_18876);
xnor U23403 (N_23403,N_19534,N_17174);
and U23404 (N_23404,N_15898,N_18319);
or U23405 (N_23405,N_19053,N_17065);
xor U23406 (N_23406,N_16753,N_17313);
xnor U23407 (N_23407,N_17354,N_15474);
or U23408 (N_23408,N_16460,N_17714);
or U23409 (N_23409,N_15582,N_17483);
and U23410 (N_23410,N_18235,N_15183);
nand U23411 (N_23411,N_18657,N_18273);
nand U23412 (N_23412,N_15729,N_15870);
or U23413 (N_23413,N_16892,N_15726);
xnor U23414 (N_23414,N_15282,N_17497);
and U23415 (N_23415,N_16457,N_16280);
nand U23416 (N_23416,N_16513,N_18694);
xor U23417 (N_23417,N_16303,N_15211);
nand U23418 (N_23418,N_15877,N_17466);
nand U23419 (N_23419,N_17702,N_16511);
or U23420 (N_23420,N_17874,N_19927);
or U23421 (N_23421,N_15591,N_18993);
xnor U23422 (N_23422,N_18966,N_17369);
and U23423 (N_23423,N_15018,N_16907);
or U23424 (N_23424,N_17079,N_19575);
or U23425 (N_23425,N_17571,N_16606);
xor U23426 (N_23426,N_17760,N_19241);
xnor U23427 (N_23427,N_17155,N_17817);
nor U23428 (N_23428,N_15393,N_15211);
nor U23429 (N_23429,N_18781,N_19046);
nand U23430 (N_23430,N_15896,N_18695);
xor U23431 (N_23431,N_19144,N_18439);
and U23432 (N_23432,N_19669,N_18176);
xor U23433 (N_23433,N_18420,N_18039);
or U23434 (N_23434,N_16632,N_16433);
and U23435 (N_23435,N_17026,N_17513);
or U23436 (N_23436,N_19904,N_16524);
nor U23437 (N_23437,N_18195,N_18584);
xnor U23438 (N_23438,N_17246,N_15470);
xor U23439 (N_23439,N_15643,N_19637);
nor U23440 (N_23440,N_18569,N_18857);
nand U23441 (N_23441,N_17342,N_17693);
and U23442 (N_23442,N_16280,N_15639);
or U23443 (N_23443,N_19160,N_16650);
and U23444 (N_23444,N_16367,N_18693);
nand U23445 (N_23445,N_17851,N_17205);
nand U23446 (N_23446,N_18233,N_18460);
xor U23447 (N_23447,N_18908,N_19978);
or U23448 (N_23448,N_16847,N_15388);
and U23449 (N_23449,N_16733,N_18209);
xor U23450 (N_23450,N_15408,N_16144);
or U23451 (N_23451,N_15099,N_19606);
nand U23452 (N_23452,N_18990,N_19921);
and U23453 (N_23453,N_17408,N_18643);
xnor U23454 (N_23454,N_17818,N_18115);
nand U23455 (N_23455,N_16860,N_15381);
or U23456 (N_23456,N_16145,N_17532);
xor U23457 (N_23457,N_17740,N_15724);
nor U23458 (N_23458,N_15456,N_15972);
xor U23459 (N_23459,N_17396,N_15725);
or U23460 (N_23460,N_15042,N_17009);
nand U23461 (N_23461,N_18232,N_15412);
xor U23462 (N_23462,N_19163,N_19565);
xor U23463 (N_23463,N_16686,N_19123);
and U23464 (N_23464,N_15030,N_17248);
nand U23465 (N_23465,N_15647,N_19996);
or U23466 (N_23466,N_16756,N_18033);
nand U23467 (N_23467,N_17960,N_19538);
nand U23468 (N_23468,N_17647,N_17948);
and U23469 (N_23469,N_18993,N_15726);
xnor U23470 (N_23470,N_15216,N_15621);
nor U23471 (N_23471,N_17368,N_16416);
and U23472 (N_23472,N_19241,N_15986);
nor U23473 (N_23473,N_16967,N_17179);
and U23474 (N_23474,N_19107,N_17557);
or U23475 (N_23475,N_19738,N_18342);
nor U23476 (N_23476,N_15259,N_15990);
nor U23477 (N_23477,N_19919,N_19649);
nand U23478 (N_23478,N_18223,N_19062);
or U23479 (N_23479,N_18022,N_17363);
or U23480 (N_23480,N_19272,N_15145);
nor U23481 (N_23481,N_18820,N_15521);
or U23482 (N_23482,N_15908,N_16039);
or U23483 (N_23483,N_17907,N_16289);
nor U23484 (N_23484,N_15480,N_19761);
or U23485 (N_23485,N_15767,N_19642);
nand U23486 (N_23486,N_17183,N_19590);
or U23487 (N_23487,N_18054,N_19739);
nor U23488 (N_23488,N_19793,N_16734);
nor U23489 (N_23489,N_17495,N_15029);
or U23490 (N_23490,N_19711,N_19243);
nand U23491 (N_23491,N_16248,N_16258);
and U23492 (N_23492,N_18724,N_19746);
xnor U23493 (N_23493,N_15410,N_15380);
xor U23494 (N_23494,N_15999,N_15282);
and U23495 (N_23495,N_17137,N_18127);
and U23496 (N_23496,N_16245,N_17833);
nand U23497 (N_23497,N_15655,N_15605);
nand U23498 (N_23498,N_19639,N_17230);
and U23499 (N_23499,N_17150,N_17819);
and U23500 (N_23500,N_18236,N_15855);
xnor U23501 (N_23501,N_16600,N_18509);
or U23502 (N_23502,N_17098,N_15799);
and U23503 (N_23503,N_17880,N_18727);
xnor U23504 (N_23504,N_17376,N_17233);
nand U23505 (N_23505,N_18455,N_16215);
nand U23506 (N_23506,N_17056,N_19946);
or U23507 (N_23507,N_15732,N_18881);
or U23508 (N_23508,N_15031,N_17639);
xor U23509 (N_23509,N_17575,N_19365);
xor U23510 (N_23510,N_18528,N_16708);
xor U23511 (N_23511,N_15879,N_19112);
or U23512 (N_23512,N_18268,N_15496);
and U23513 (N_23513,N_19284,N_17501);
xnor U23514 (N_23514,N_16462,N_15945);
or U23515 (N_23515,N_18869,N_15206);
xor U23516 (N_23516,N_16413,N_16466);
nand U23517 (N_23517,N_16144,N_18344);
nand U23518 (N_23518,N_19394,N_16057);
and U23519 (N_23519,N_17913,N_16942);
xnor U23520 (N_23520,N_17728,N_15149);
or U23521 (N_23521,N_18284,N_17749);
nand U23522 (N_23522,N_16621,N_18219);
nand U23523 (N_23523,N_16813,N_18425);
and U23524 (N_23524,N_18135,N_19270);
nor U23525 (N_23525,N_18227,N_18935);
nor U23526 (N_23526,N_19900,N_18866);
and U23527 (N_23527,N_18047,N_18640);
xor U23528 (N_23528,N_15482,N_18303);
nand U23529 (N_23529,N_18248,N_18350);
nand U23530 (N_23530,N_16996,N_17618);
nor U23531 (N_23531,N_18735,N_19257);
and U23532 (N_23532,N_19111,N_15991);
nand U23533 (N_23533,N_19091,N_19131);
or U23534 (N_23534,N_15451,N_18574);
nor U23535 (N_23535,N_15479,N_18947);
nor U23536 (N_23536,N_17382,N_15811);
nand U23537 (N_23537,N_19791,N_17152);
nand U23538 (N_23538,N_15417,N_15217);
xor U23539 (N_23539,N_16651,N_18395);
xor U23540 (N_23540,N_19625,N_15483);
and U23541 (N_23541,N_19571,N_16687);
nand U23542 (N_23542,N_17305,N_16419);
or U23543 (N_23543,N_18350,N_18532);
nor U23544 (N_23544,N_17382,N_17812);
xnor U23545 (N_23545,N_17024,N_15135);
or U23546 (N_23546,N_16399,N_18751);
xnor U23547 (N_23547,N_17703,N_15546);
and U23548 (N_23548,N_17823,N_15365);
nor U23549 (N_23549,N_18031,N_17366);
xnor U23550 (N_23550,N_17815,N_15017);
and U23551 (N_23551,N_15860,N_15460);
nor U23552 (N_23552,N_16325,N_18552);
nand U23553 (N_23553,N_16833,N_19823);
and U23554 (N_23554,N_18354,N_19301);
nor U23555 (N_23555,N_16833,N_17013);
or U23556 (N_23556,N_15365,N_19273);
nor U23557 (N_23557,N_17363,N_16824);
nand U23558 (N_23558,N_16764,N_16318);
and U23559 (N_23559,N_16881,N_19922);
and U23560 (N_23560,N_15905,N_18296);
nor U23561 (N_23561,N_18167,N_18083);
xor U23562 (N_23562,N_18942,N_18814);
or U23563 (N_23563,N_16759,N_19342);
or U23564 (N_23564,N_18014,N_18620);
nor U23565 (N_23565,N_16614,N_18872);
and U23566 (N_23566,N_19775,N_17027);
or U23567 (N_23567,N_15558,N_15778);
nor U23568 (N_23568,N_15597,N_17235);
nand U23569 (N_23569,N_19545,N_19662);
nor U23570 (N_23570,N_19529,N_17613);
nand U23571 (N_23571,N_15750,N_19097);
nand U23572 (N_23572,N_15453,N_15677);
nor U23573 (N_23573,N_16862,N_16131);
or U23574 (N_23574,N_17360,N_17640);
nor U23575 (N_23575,N_19690,N_18635);
xnor U23576 (N_23576,N_18336,N_17266);
and U23577 (N_23577,N_16575,N_16764);
and U23578 (N_23578,N_16104,N_16961);
nand U23579 (N_23579,N_19544,N_18894);
xnor U23580 (N_23580,N_16591,N_16371);
or U23581 (N_23581,N_18144,N_18291);
xor U23582 (N_23582,N_19241,N_19075);
nor U23583 (N_23583,N_18083,N_18889);
or U23584 (N_23584,N_18173,N_17754);
xnor U23585 (N_23585,N_17282,N_16108);
nand U23586 (N_23586,N_17945,N_19909);
nand U23587 (N_23587,N_19767,N_15194);
and U23588 (N_23588,N_15850,N_17779);
or U23589 (N_23589,N_16804,N_18646);
xnor U23590 (N_23590,N_19727,N_15373);
xor U23591 (N_23591,N_18876,N_17026);
and U23592 (N_23592,N_19908,N_19242);
or U23593 (N_23593,N_17142,N_16408);
nor U23594 (N_23594,N_18285,N_18151);
nand U23595 (N_23595,N_16499,N_17700);
nand U23596 (N_23596,N_17930,N_17703);
nand U23597 (N_23597,N_18771,N_17062);
and U23598 (N_23598,N_16972,N_18228);
and U23599 (N_23599,N_16897,N_19860);
or U23600 (N_23600,N_19035,N_15061);
or U23601 (N_23601,N_16310,N_16919);
xnor U23602 (N_23602,N_17629,N_19802);
and U23603 (N_23603,N_15721,N_19751);
and U23604 (N_23604,N_19417,N_18265);
or U23605 (N_23605,N_19187,N_15586);
xor U23606 (N_23606,N_15415,N_16725);
xnor U23607 (N_23607,N_19727,N_15988);
or U23608 (N_23608,N_15915,N_15496);
or U23609 (N_23609,N_16532,N_16323);
and U23610 (N_23610,N_19607,N_17269);
and U23611 (N_23611,N_15204,N_17219);
xor U23612 (N_23612,N_15623,N_15878);
or U23613 (N_23613,N_17470,N_19304);
xnor U23614 (N_23614,N_18572,N_17327);
nor U23615 (N_23615,N_18195,N_19785);
nor U23616 (N_23616,N_18212,N_16443);
xor U23617 (N_23617,N_18294,N_16615);
xnor U23618 (N_23618,N_19892,N_15764);
nor U23619 (N_23619,N_16427,N_17087);
and U23620 (N_23620,N_16135,N_19399);
nand U23621 (N_23621,N_17290,N_17105);
nand U23622 (N_23622,N_18218,N_19332);
nor U23623 (N_23623,N_19691,N_17038);
xnor U23624 (N_23624,N_17531,N_16077);
xnor U23625 (N_23625,N_19244,N_18618);
or U23626 (N_23626,N_15680,N_17302);
and U23627 (N_23627,N_19664,N_15132);
or U23628 (N_23628,N_15415,N_18851);
nor U23629 (N_23629,N_18262,N_19742);
nor U23630 (N_23630,N_19208,N_16389);
nand U23631 (N_23631,N_16603,N_15513);
nor U23632 (N_23632,N_19492,N_19449);
and U23633 (N_23633,N_16796,N_18182);
and U23634 (N_23634,N_19508,N_15206);
nor U23635 (N_23635,N_16668,N_18980);
or U23636 (N_23636,N_16508,N_19202);
nor U23637 (N_23637,N_17779,N_16123);
or U23638 (N_23638,N_17383,N_19386);
nand U23639 (N_23639,N_18714,N_19103);
xnor U23640 (N_23640,N_15208,N_18463);
nand U23641 (N_23641,N_15418,N_17739);
nand U23642 (N_23642,N_19138,N_18270);
and U23643 (N_23643,N_19280,N_15191);
or U23644 (N_23644,N_17264,N_17676);
and U23645 (N_23645,N_16788,N_17191);
xnor U23646 (N_23646,N_17178,N_19210);
nand U23647 (N_23647,N_18252,N_19014);
and U23648 (N_23648,N_16033,N_17241);
nand U23649 (N_23649,N_17632,N_18439);
or U23650 (N_23650,N_16042,N_15114);
and U23651 (N_23651,N_17377,N_19333);
or U23652 (N_23652,N_17553,N_18677);
nand U23653 (N_23653,N_16154,N_16150);
nor U23654 (N_23654,N_16396,N_18958);
nor U23655 (N_23655,N_17720,N_18602);
xnor U23656 (N_23656,N_19204,N_15568);
nor U23657 (N_23657,N_15892,N_17756);
nor U23658 (N_23658,N_15758,N_18752);
or U23659 (N_23659,N_17967,N_17760);
xnor U23660 (N_23660,N_19045,N_17063);
or U23661 (N_23661,N_16286,N_15404);
or U23662 (N_23662,N_16303,N_19346);
nor U23663 (N_23663,N_16069,N_18155);
nor U23664 (N_23664,N_19452,N_19753);
nand U23665 (N_23665,N_15683,N_19397);
or U23666 (N_23666,N_19504,N_16804);
or U23667 (N_23667,N_17909,N_17845);
or U23668 (N_23668,N_15575,N_18988);
nand U23669 (N_23669,N_19001,N_15076);
xor U23670 (N_23670,N_15731,N_19522);
nand U23671 (N_23671,N_17416,N_19420);
xnor U23672 (N_23672,N_15458,N_17116);
xor U23673 (N_23673,N_15594,N_17141);
nor U23674 (N_23674,N_17011,N_18991);
xnor U23675 (N_23675,N_16238,N_19125);
nor U23676 (N_23676,N_19144,N_16553);
nor U23677 (N_23677,N_15295,N_19449);
xor U23678 (N_23678,N_16587,N_15364);
xnor U23679 (N_23679,N_17551,N_19715);
or U23680 (N_23680,N_18045,N_17838);
nor U23681 (N_23681,N_19220,N_18851);
nand U23682 (N_23682,N_17891,N_17206);
or U23683 (N_23683,N_18944,N_15287);
or U23684 (N_23684,N_15860,N_18643);
or U23685 (N_23685,N_16184,N_16861);
or U23686 (N_23686,N_15286,N_17297);
or U23687 (N_23687,N_19562,N_17178);
or U23688 (N_23688,N_18268,N_16342);
nor U23689 (N_23689,N_17727,N_15041);
or U23690 (N_23690,N_17572,N_15458);
nor U23691 (N_23691,N_17088,N_18380);
nor U23692 (N_23692,N_16048,N_18890);
and U23693 (N_23693,N_16111,N_19061);
or U23694 (N_23694,N_19524,N_16979);
xor U23695 (N_23695,N_18614,N_16239);
and U23696 (N_23696,N_17208,N_18362);
xor U23697 (N_23697,N_18040,N_19886);
and U23698 (N_23698,N_15375,N_16073);
nand U23699 (N_23699,N_16514,N_18724);
or U23700 (N_23700,N_15326,N_15175);
nand U23701 (N_23701,N_16030,N_18753);
xor U23702 (N_23702,N_18532,N_19430);
xnor U23703 (N_23703,N_16609,N_19062);
xor U23704 (N_23704,N_18802,N_16535);
nand U23705 (N_23705,N_16623,N_19606);
xnor U23706 (N_23706,N_18903,N_19284);
xor U23707 (N_23707,N_15352,N_16227);
and U23708 (N_23708,N_16647,N_18740);
and U23709 (N_23709,N_17040,N_16300);
or U23710 (N_23710,N_16879,N_16434);
nor U23711 (N_23711,N_15069,N_15172);
nand U23712 (N_23712,N_18374,N_19488);
and U23713 (N_23713,N_19598,N_17027);
nor U23714 (N_23714,N_15395,N_16515);
xor U23715 (N_23715,N_18342,N_19519);
xor U23716 (N_23716,N_16561,N_17493);
and U23717 (N_23717,N_18394,N_16018);
xnor U23718 (N_23718,N_19711,N_16179);
and U23719 (N_23719,N_16189,N_16803);
or U23720 (N_23720,N_15272,N_17446);
or U23721 (N_23721,N_16804,N_19305);
nor U23722 (N_23722,N_15698,N_18062);
and U23723 (N_23723,N_15867,N_16357);
nor U23724 (N_23724,N_17534,N_16998);
nand U23725 (N_23725,N_18283,N_17790);
or U23726 (N_23726,N_19205,N_17988);
or U23727 (N_23727,N_19454,N_17195);
nand U23728 (N_23728,N_16760,N_16767);
and U23729 (N_23729,N_19002,N_18388);
and U23730 (N_23730,N_16197,N_17543);
xor U23731 (N_23731,N_15124,N_19147);
nor U23732 (N_23732,N_18995,N_17820);
and U23733 (N_23733,N_15366,N_16288);
nor U23734 (N_23734,N_16506,N_16306);
xnor U23735 (N_23735,N_16809,N_19600);
or U23736 (N_23736,N_16809,N_19623);
and U23737 (N_23737,N_16199,N_19369);
nor U23738 (N_23738,N_18481,N_18146);
and U23739 (N_23739,N_19549,N_18084);
and U23740 (N_23740,N_15495,N_15616);
xor U23741 (N_23741,N_16102,N_18160);
nor U23742 (N_23742,N_19977,N_19923);
or U23743 (N_23743,N_18940,N_15088);
nor U23744 (N_23744,N_16110,N_16882);
xor U23745 (N_23745,N_16104,N_17956);
and U23746 (N_23746,N_16332,N_17353);
and U23747 (N_23747,N_19772,N_17045);
nand U23748 (N_23748,N_16978,N_15533);
nand U23749 (N_23749,N_18819,N_15365);
nand U23750 (N_23750,N_16701,N_17557);
and U23751 (N_23751,N_17276,N_16937);
nor U23752 (N_23752,N_16485,N_18068);
and U23753 (N_23753,N_15220,N_16511);
xor U23754 (N_23754,N_16634,N_17541);
nand U23755 (N_23755,N_18011,N_15749);
and U23756 (N_23756,N_18117,N_17746);
nor U23757 (N_23757,N_18973,N_17094);
or U23758 (N_23758,N_17338,N_19934);
or U23759 (N_23759,N_17277,N_17318);
xnor U23760 (N_23760,N_17488,N_15573);
or U23761 (N_23761,N_17494,N_18515);
or U23762 (N_23762,N_15276,N_19107);
xnor U23763 (N_23763,N_17711,N_18793);
or U23764 (N_23764,N_17747,N_19250);
nand U23765 (N_23765,N_17209,N_18357);
nand U23766 (N_23766,N_18495,N_17313);
or U23767 (N_23767,N_19435,N_18940);
nand U23768 (N_23768,N_17051,N_15756);
or U23769 (N_23769,N_16160,N_19687);
nor U23770 (N_23770,N_18278,N_18174);
xor U23771 (N_23771,N_17135,N_18785);
xnor U23772 (N_23772,N_19845,N_18544);
and U23773 (N_23773,N_15282,N_19396);
or U23774 (N_23774,N_19402,N_16751);
and U23775 (N_23775,N_18965,N_18280);
nand U23776 (N_23776,N_18189,N_15135);
xnor U23777 (N_23777,N_17042,N_18223);
xnor U23778 (N_23778,N_18245,N_19742);
nor U23779 (N_23779,N_16295,N_16181);
and U23780 (N_23780,N_16371,N_19701);
nor U23781 (N_23781,N_18537,N_15132);
xor U23782 (N_23782,N_17598,N_17950);
xor U23783 (N_23783,N_16791,N_16326);
nor U23784 (N_23784,N_16996,N_15077);
xor U23785 (N_23785,N_19504,N_19718);
xnor U23786 (N_23786,N_17699,N_17214);
nor U23787 (N_23787,N_16478,N_17437);
xor U23788 (N_23788,N_17057,N_19008);
or U23789 (N_23789,N_16169,N_17028);
xor U23790 (N_23790,N_17732,N_17098);
xnor U23791 (N_23791,N_17284,N_19211);
xnor U23792 (N_23792,N_16234,N_18041);
nand U23793 (N_23793,N_19950,N_19012);
xor U23794 (N_23794,N_19974,N_17177);
nand U23795 (N_23795,N_19033,N_16566);
xor U23796 (N_23796,N_16778,N_17348);
nor U23797 (N_23797,N_19034,N_15457);
and U23798 (N_23798,N_16899,N_16461);
or U23799 (N_23799,N_16328,N_19366);
xor U23800 (N_23800,N_16649,N_16019);
nor U23801 (N_23801,N_19403,N_17213);
xor U23802 (N_23802,N_18449,N_17624);
or U23803 (N_23803,N_18122,N_17510);
nand U23804 (N_23804,N_18304,N_17798);
nor U23805 (N_23805,N_17623,N_17125);
nor U23806 (N_23806,N_16736,N_19791);
nor U23807 (N_23807,N_15887,N_17176);
and U23808 (N_23808,N_19110,N_15225);
or U23809 (N_23809,N_15361,N_15165);
nand U23810 (N_23810,N_18567,N_16670);
xnor U23811 (N_23811,N_15351,N_16227);
nor U23812 (N_23812,N_18191,N_18332);
nand U23813 (N_23813,N_18286,N_15457);
or U23814 (N_23814,N_16486,N_19984);
xor U23815 (N_23815,N_19446,N_15549);
nor U23816 (N_23816,N_16626,N_19297);
or U23817 (N_23817,N_19527,N_16476);
xnor U23818 (N_23818,N_15744,N_17046);
nor U23819 (N_23819,N_17639,N_15101);
and U23820 (N_23820,N_15396,N_15288);
nor U23821 (N_23821,N_18695,N_19392);
and U23822 (N_23822,N_17759,N_15596);
xor U23823 (N_23823,N_18669,N_18890);
or U23824 (N_23824,N_19266,N_17911);
xnor U23825 (N_23825,N_16503,N_17636);
xor U23826 (N_23826,N_19939,N_18010);
nand U23827 (N_23827,N_19328,N_16161);
nor U23828 (N_23828,N_15197,N_17717);
and U23829 (N_23829,N_19071,N_17607);
and U23830 (N_23830,N_17624,N_18596);
or U23831 (N_23831,N_16356,N_15104);
or U23832 (N_23832,N_16020,N_17368);
or U23833 (N_23833,N_17152,N_16404);
nor U23834 (N_23834,N_15569,N_19150);
nand U23835 (N_23835,N_18463,N_18276);
or U23836 (N_23836,N_15935,N_16960);
xnor U23837 (N_23837,N_17172,N_19043);
nand U23838 (N_23838,N_16487,N_17603);
nand U23839 (N_23839,N_15179,N_17796);
nor U23840 (N_23840,N_16549,N_16980);
or U23841 (N_23841,N_18731,N_18470);
or U23842 (N_23842,N_15736,N_18988);
nor U23843 (N_23843,N_16895,N_15568);
nor U23844 (N_23844,N_16602,N_18313);
xor U23845 (N_23845,N_15778,N_18461);
and U23846 (N_23846,N_19124,N_18296);
xor U23847 (N_23847,N_17907,N_18034);
nand U23848 (N_23848,N_15072,N_15151);
nand U23849 (N_23849,N_16920,N_16901);
xor U23850 (N_23850,N_19768,N_17321);
nor U23851 (N_23851,N_18548,N_17948);
and U23852 (N_23852,N_18101,N_15701);
and U23853 (N_23853,N_16160,N_15532);
nand U23854 (N_23854,N_19628,N_17127);
xor U23855 (N_23855,N_15034,N_17611);
or U23856 (N_23856,N_19906,N_19787);
xor U23857 (N_23857,N_16880,N_18239);
xnor U23858 (N_23858,N_19097,N_19449);
or U23859 (N_23859,N_19768,N_19926);
nand U23860 (N_23860,N_17887,N_18608);
or U23861 (N_23861,N_18085,N_16979);
xor U23862 (N_23862,N_19116,N_15306);
and U23863 (N_23863,N_19435,N_18710);
nor U23864 (N_23864,N_17010,N_17881);
xnor U23865 (N_23865,N_15362,N_19909);
nand U23866 (N_23866,N_16331,N_17458);
nand U23867 (N_23867,N_17816,N_18157);
nand U23868 (N_23868,N_16599,N_17888);
nor U23869 (N_23869,N_16712,N_18978);
xor U23870 (N_23870,N_18497,N_17889);
and U23871 (N_23871,N_15715,N_16758);
nand U23872 (N_23872,N_18266,N_16779);
or U23873 (N_23873,N_19076,N_16837);
or U23874 (N_23874,N_15335,N_19419);
nand U23875 (N_23875,N_19687,N_17186);
or U23876 (N_23876,N_17798,N_17406);
nor U23877 (N_23877,N_19445,N_16971);
nor U23878 (N_23878,N_17890,N_17873);
nand U23879 (N_23879,N_15925,N_17337);
or U23880 (N_23880,N_19007,N_19575);
xor U23881 (N_23881,N_15567,N_18946);
or U23882 (N_23882,N_17991,N_17731);
or U23883 (N_23883,N_17408,N_15556);
or U23884 (N_23884,N_16263,N_17593);
or U23885 (N_23885,N_16623,N_18686);
or U23886 (N_23886,N_15613,N_19501);
xor U23887 (N_23887,N_17675,N_16383);
and U23888 (N_23888,N_17292,N_15523);
and U23889 (N_23889,N_18950,N_15189);
or U23890 (N_23890,N_15324,N_19408);
or U23891 (N_23891,N_16634,N_15005);
and U23892 (N_23892,N_16794,N_16100);
nor U23893 (N_23893,N_17174,N_15302);
nor U23894 (N_23894,N_16261,N_16967);
nor U23895 (N_23895,N_18496,N_18626);
xnor U23896 (N_23896,N_17161,N_15850);
and U23897 (N_23897,N_15734,N_15205);
xnor U23898 (N_23898,N_16931,N_19885);
or U23899 (N_23899,N_18369,N_15586);
nand U23900 (N_23900,N_15242,N_15979);
xor U23901 (N_23901,N_19637,N_17046);
and U23902 (N_23902,N_18675,N_16131);
or U23903 (N_23903,N_16690,N_16272);
and U23904 (N_23904,N_15815,N_15502);
nand U23905 (N_23905,N_16013,N_17691);
or U23906 (N_23906,N_16728,N_19400);
or U23907 (N_23907,N_18909,N_18764);
or U23908 (N_23908,N_15079,N_16941);
or U23909 (N_23909,N_15694,N_19137);
or U23910 (N_23910,N_16916,N_17241);
nand U23911 (N_23911,N_19587,N_19842);
nor U23912 (N_23912,N_17070,N_18172);
nor U23913 (N_23913,N_15075,N_19269);
or U23914 (N_23914,N_18152,N_17884);
nor U23915 (N_23915,N_19078,N_18742);
and U23916 (N_23916,N_19528,N_17549);
or U23917 (N_23917,N_17394,N_18676);
nor U23918 (N_23918,N_19621,N_18624);
xor U23919 (N_23919,N_18744,N_16594);
xor U23920 (N_23920,N_18939,N_17451);
and U23921 (N_23921,N_17330,N_15967);
or U23922 (N_23922,N_17817,N_19909);
nand U23923 (N_23923,N_19028,N_15482);
or U23924 (N_23924,N_17860,N_16363);
nor U23925 (N_23925,N_16020,N_18212);
xnor U23926 (N_23926,N_18343,N_15480);
nand U23927 (N_23927,N_19432,N_18607);
xnor U23928 (N_23928,N_18615,N_15879);
xnor U23929 (N_23929,N_19817,N_15208);
or U23930 (N_23930,N_16382,N_19078);
nand U23931 (N_23931,N_16793,N_19677);
xor U23932 (N_23932,N_17913,N_19745);
or U23933 (N_23933,N_18969,N_18602);
nor U23934 (N_23934,N_15321,N_17498);
nor U23935 (N_23935,N_17471,N_18012);
nand U23936 (N_23936,N_18949,N_18349);
nand U23937 (N_23937,N_19813,N_17907);
and U23938 (N_23938,N_16031,N_16066);
nor U23939 (N_23939,N_17538,N_19843);
nand U23940 (N_23940,N_18535,N_17821);
nor U23941 (N_23941,N_17490,N_18179);
nor U23942 (N_23942,N_19221,N_16457);
and U23943 (N_23943,N_15183,N_18377);
nor U23944 (N_23944,N_19948,N_19713);
nor U23945 (N_23945,N_15814,N_17818);
nor U23946 (N_23946,N_15473,N_17283);
xnor U23947 (N_23947,N_16380,N_19951);
nor U23948 (N_23948,N_17324,N_16938);
nor U23949 (N_23949,N_15718,N_15733);
xnor U23950 (N_23950,N_16994,N_18677);
xnor U23951 (N_23951,N_19232,N_16976);
nor U23952 (N_23952,N_19910,N_17125);
nand U23953 (N_23953,N_18219,N_19045);
nand U23954 (N_23954,N_16484,N_17674);
xnor U23955 (N_23955,N_17391,N_18634);
nor U23956 (N_23956,N_16850,N_15144);
nand U23957 (N_23957,N_17481,N_18912);
nor U23958 (N_23958,N_15549,N_19986);
xnor U23959 (N_23959,N_19576,N_18419);
nor U23960 (N_23960,N_15703,N_18120);
or U23961 (N_23961,N_17410,N_15012);
nor U23962 (N_23962,N_18641,N_16010);
nand U23963 (N_23963,N_18350,N_17585);
nor U23964 (N_23964,N_18957,N_17524);
nand U23965 (N_23965,N_16183,N_17221);
or U23966 (N_23966,N_17930,N_16834);
nor U23967 (N_23967,N_18380,N_19303);
nor U23968 (N_23968,N_16473,N_16335);
or U23969 (N_23969,N_16083,N_16403);
or U23970 (N_23970,N_17306,N_15196);
or U23971 (N_23971,N_19806,N_18509);
and U23972 (N_23972,N_18688,N_16754);
xor U23973 (N_23973,N_15549,N_17080);
nor U23974 (N_23974,N_15266,N_16389);
and U23975 (N_23975,N_19367,N_16290);
and U23976 (N_23976,N_15010,N_18550);
nand U23977 (N_23977,N_16153,N_19394);
and U23978 (N_23978,N_16340,N_18435);
or U23979 (N_23979,N_15979,N_17896);
nor U23980 (N_23980,N_18249,N_18769);
or U23981 (N_23981,N_15979,N_16583);
or U23982 (N_23982,N_18949,N_19076);
nor U23983 (N_23983,N_15009,N_17675);
and U23984 (N_23984,N_16284,N_15253);
nand U23985 (N_23985,N_18715,N_18464);
nor U23986 (N_23986,N_18738,N_16368);
nand U23987 (N_23987,N_17666,N_17906);
and U23988 (N_23988,N_18990,N_17627);
or U23989 (N_23989,N_18913,N_17333);
nand U23990 (N_23990,N_18541,N_18194);
nor U23991 (N_23991,N_19063,N_17484);
and U23992 (N_23992,N_18518,N_18048);
nand U23993 (N_23993,N_18803,N_15897);
and U23994 (N_23994,N_18016,N_16458);
nand U23995 (N_23995,N_16944,N_15922);
xor U23996 (N_23996,N_15303,N_15394);
or U23997 (N_23997,N_15477,N_15615);
nand U23998 (N_23998,N_19813,N_18928);
and U23999 (N_23999,N_18639,N_19524);
nand U24000 (N_24000,N_16015,N_18552);
nand U24001 (N_24001,N_19777,N_19412);
or U24002 (N_24002,N_19914,N_15970);
nor U24003 (N_24003,N_18132,N_17778);
or U24004 (N_24004,N_17784,N_15878);
and U24005 (N_24005,N_18961,N_18082);
nand U24006 (N_24006,N_17257,N_17258);
xnor U24007 (N_24007,N_16545,N_16377);
nand U24008 (N_24008,N_17271,N_19417);
and U24009 (N_24009,N_19845,N_19966);
and U24010 (N_24010,N_15575,N_15715);
and U24011 (N_24011,N_19257,N_17800);
xor U24012 (N_24012,N_18596,N_17064);
nor U24013 (N_24013,N_18246,N_17042);
nor U24014 (N_24014,N_17860,N_18592);
xnor U24015 (N_24015,N_15503,N_18581);
xnor U24016 (N_24016,N_19800,N_19852);
or U24017 (N_24017,N_17030,N_16751);
nor U24018 (N_24018,N_16872,N_16136);
nand U24019 (N_24019,N_17989,N_19924);
xnor U24020 (N_24020,N_16047,N_19434);
nand U24021 (N_24021,N_18467,N_19343);
xnor U24022 (N_24022,N_17886,N_15053);
xnor U24023 (N_24023,N_19085,N_19531);
xor U24024 (N_24024,N_19321,N_18078);
nand U24025 (N_24025,N_16253,N_19774);
or U24026 (N_24026,N_17500,N_19344);
nand U24027 (N_24027,N_19118,N_17562);
nor U24028 (N_24028,N_15448,N_19603);
nand U24029 (N_24029,N_16240,N_19616);
xor U24030 (N_24030,N_15107,N_18187);
nand U24031 (N_24031,N_17148,N_16853);
xor U24032 (N_24032,N_15996,N_16723);
nand U24033 (N_24033,N_18174,N_16504);
and U24034 (N_24034,N_19664,N_17411);
nand U24035 (N_24035,N_17389,N_17948);
or U24036 (N_24036,N_19828,N_15630);
nand U24037 (N_24037,N_17251,N_16061);
and U24038 (N_24038,N_17012,N_16354);
nand U24039 (N_24039,N_19793,N_17331);
and U24040 (N_24040,N_15826,N_18788);
xor U24041 (N_24041,N_19895,N_19285);
and U24042 (N_24042,N_15056,N_17966);
nand U24043 (N_24043,N_18471,N_16234);
nor U24044 (N_24044,N_18684,N_18343);
or U24045 (N_24045,N_18796,N_16419);
and U24046 (N_24046,N_17850,N_18802);
nor U24047 (N_24047,N_19827,N_16853);
or U24048 (N_24048,N_19788,N_19015);
and U24049 (N_24049,N_16780,N_17132);
and U24050 (N_24050,N_18516,N_18479);
or U24051 (N_24051,N_16024,N_19338);
and U24052 (N_24052,N_19144,N_19792);
nand U24053 (N_24053,N_17341,N_18596);
and U24054 (N_24054,N_16631,N_15142);
and U24055 (N_24055,N_16793,N_16153);
xor U24056 (N_24056,N_18019,N_19547);
and U24057 (N_24057,N_19486,N_15814);
xor U24058 (N_24058,N_17367,N_15680);
and U24059 (N_24059,N_16056,N_19944);
nand U24060 (N_24060,N_17191,N_15287);
or U24061 (N_24061,N_17466,N_15787);
xor U24062 (N_24062,N_16974,N_19542);
and U24063 (N_24063,N_17427,N_15119);
or U24064 (N_24064,N_17553,N_19041);
or U24065 (N_24065,N_15176,N_19309);
or U24066 (N_24066,N_16789,N_17133);
and U24067 (N_24067,N_19208,N_17259);
xor U24068 (N_24068,N_19956,N_16714);
or U24069 (N_24069,N_17943,N_19186);
and U24070 (N_24070,N_17478,N_18334);
nor U24071 (N_24071,N_15803,N_15881);
nand U24072 (N_24072,N_19060,N_18572);
xnor U24073 (N_24073,N_15338,N_19620);
or U24074 (N_24074,N_16159,N_15095);
or U24075 (N_24075,N_17627,N_17259);
xnor U24076 (N_24076,N_15291,N_19053);
nand U24077 (N_24077,N_16553,N_17789);
nor U24078 (N_24078,N_15193,N_16722);
nor U24079 (N_24079,N_16507,N_17415);
and U24080 (N_24080,N_18073,N_15264);
nand U24081 (N_24081,N_15168,N_15866);
xor U24082 (N_24082,N_19042,N_15644);
nor U24083 (N_24083,N_18072,N_16852);
xnor U24084 (N_24084,N_15310,N_16922);
nor U24085 (N_24085,N_16300,N_15358);
nor U24086 (N_24086,N_18823,N_18741);
and U24087 (N_24087,N_15700,N_15250);
and U24088 (N_24088,N_19867,N_17379);
nand U24089 (N_24089,N_17162,N_18851);
or U24090 (N_24090,N_15133,N_16213);
nor U24091 (N_24091,N_19882,N_18615);
and U24092 (N_24092,N_15670,N_19753);
nor U24093 (N_24093,N_16417,N_15951);
and U24094 (N_24094,N_18711,N_15578);
nor U24095 (N_24095,N_18096,N_18444);
and U24096 (N_24096,N_19745,N_15165);
nor U24097 (N_24097,N_15775,N_17028);
nor U24098 (N_24098,N_15254,N_19749);
xnor U24099 (N_24099,N_18848,N_18287);
and U24100 (N_24100,N_19860,N_16513);
nand U24101 (N_24101,N_17058,N_15767);
nor U24102 (N_24102,N_18856,N_16703);
nand U24103 (N_24103,N_16656,N_17742);
or U24104 (N_24104,N_16293,N_16999);
nor U24105 (N_24105,N_15502,N_17529);
xor U24106 (N_24106,N_17747,N_17093);
and U24107 (N_24107,N_19724,N_17996);
or U24108 (N_24108,N_18525,N_15965);
or U24109 (N_24109,N_16546,N_15942);
xnor U24110 (N_24110,N_18411,N_16305);
or U24111 (N_24111,N_19206,N_18423);
or U24112 (N_24112,N_17696,N_15278);
xor U24113 (N_24113,N_17501,N_17830);
nor U24114 (N_24114,N_19089,N_16238);
xnor U24115 (N_24115,N_16561,N_15241);
or U24116 (N_24116,N_18339,N_18875);
nor U24117 (N_24117,N_19682,N_15419);
or U24118 (N_24118,N_17475,N_15874);
nor U24119 (N_24119,N_17762,N_18362);
xor U24120 (N_24120,N_16896,N_19202);
or U24121 (N_24121,N_15480,N_19900);
and U24122 (N_24122,N_16483,N_16316);
or U24123 (N_24123,N_18518,N_19551);
and U24124 (N_24124,N_16594,N_16836);
or U24125 (N_24125,N_15517,N_18138);
and U24126 (N_24126,N_19076,N_18152);
nand U24127 (N_24127,N_16365,N_15468);
xor U24128 (N_24128,N_15299,N_16866);
nand U24129 (N_24129,N_16036,N_19725);
and U24130 (N_24130,N_16988,N_16479);
xor U24131 (N_24131,N_16112,N_16265);
nor U24132 (N_24132,N_17149,N_15252);
nand U24133 (N_24133,N_16810,N_17371);
xor U24134 (N_24134,N_15919,N_17501);
and U24135 (N_24135,N_19321,N_17460);
and U24136 (N_24136,N_18311,N_17185);
or U24137 (N_24137,N_15136,N_17295);
nand U24138 (N_24138,N_18526,N_18466);
and U24139 (N_24139,N_19268,N_15650);
nand U24140 (N_24140,N_16781,N_18919);
or U24141 (N_24141,N_18823,N_19396);
xnor U24142 (N_24142,N_15174,N_17831);
and U24143 (N_24143,N_17110,N_19591);
or U24144 (N_24144,N_16955,N_19973);
xor U24145 (N_24145,N_15633,N_19849);
nor U24146 (N_24146,N_15834,N_18546);
nand U24147 (N_24147,N_15108,N_18548);
nor U24148 (N_24148,N_16647,N_17127);
nand U24149 (N_24149,N_18504,N_18159);
or U24150 (N_24150,N_19303,N_17486);
nor U24151 (N_24151,N_18507,N_16987);
nand U24152 (N_24152,N_19886,N_18686);
nand U24153 (N_24153,N_15724,N_18524);
and U24154 (N_24154,N_15186,N_15182);
or U24155 (N_24155,N_15245,N_19600);
nor U24156 (N_24156,N_18253,N_17644);
and U24157 (N_24157,N_15709,N_18291);
xnor U24158 (N_24158,N_15164,N_19510);
xnor U24159 (N_24159,N_19724,N_16827);
xor U24160 (N_24160,N_19073,N_17213);
xor U24161 (N_24161,N_15841,N_18229);
xor U24162 (N_24162,N_17693,N_16262);
xnor U24163 (N_24163,N_16231,N_16515);
xnor U24164 (N_24164,N_15727,N_18543);
and U24165 (N_24165,N_18868,N_16976);
nor U24166 (N_24166,N_16083,N_18463);
nor U24167 (N_24167,N_18536,N_17049);
or U24168 (N_24168,N_18547,N_19071);
xnor U24169 (N_24169,N_15814,N_16832);
or U24170 (N_24170,N_17287,N_18009);
xor U24171 (N_24171,N_17387,N_15132);
xor U24172 (N_24172,N_19160,N_17383);
nand U24173 (N_24173,N_16921,N_19296);
nand U24174 (N_24174,N_15117,N_15783);
or U24175 (N_24175,N_17968,N_16549);
xnor U24176 (N_24176,N_17421,N_16497);
and U24177 (N_24177,N_16547,N_17933);
or U24178 (N_24178,N_19306,N_19759);
or U24179 (N_24179,N_19763,N_15881);
nand U24180 (N_24180,N_16969,N_19676);
xor U24181 (N_24181,N_18510,N_16963);
nor U24182 (N_24182,N_16577,N_18244);
xnor U24183 (N_24183,N_18837,N_17534);
or U24184 (N_24184,N_17847,N_17564);
or U24185 (N_24185,N_15602,N_17852);
or U24186 (N_24186,N_19178,N_17098);
or U24187 (N_24187,N_19400,N_17971);
xnor U24188 (N_24188,N_17832,N_17178);
xnor U24189 (N_24189,N_16192,N_19348);
xnor U24190 (N_24190,N_16566,N_15120);
and U24191 (N_24191,N_15167,N_17137);
nor U24192 (N_24192,N_15795,N_19314);
xnor U24193 (N_24193,N_19058,N_18763);
and U24194 (N_24194,N_19523,N_16032);
and U24195 (N_24195,N_15604,N_18109);
and U24196 (N_24196,N_19451,N_17133);
nor U24197 (N_24197,N_17201,N_15775);
and U24198 (N_24198,N_17327,N_19546);
or U24199 (N_24199,N_16881,N_16116);
or U24200 (N_24200,N_17269,N_17889);
or U24201 (N_24201,N_18862,N_15330);
nor U24202 (N_24202,N_15388,N_16941);
nor U24203 (N_24203,N_19055,N_15663);
nor U24204 (N_24204,N_15858,N_15530);
nor U24205 (N_24205,N_19911,N_19855);
or U24206 (N_24206,N_16922,N_15569);
and U24207 (N_24207,N_19687,N_16497);
nor U24208 (N_24208,N_19745,N_18225);
nand U24209 (N_24209,N_18857,N_17736);
xnor U24210 (N_24210,N_15791,N_17352);
nor U24211 (N_24211,N_17330,N_19405);
or U24212 (N_24212,N_16326,N_18133);
xnor U24213 (N_24213,N_15070,N_15074);
and U24214 (N_24214,N_19566,N_16330);
xor U24215 (N_24215,N_17959,N_16121);
xor U24216 (N_24216,N_15124,N_17484);
nand U24217 (N_24217,N_19410,N_17058);
nand U24218 (N_24218,N_17026,N_18897);
xor U24219 (N_24219,N_17941,N_16393);
xor U24220 (N_24220,N_17911,N_18055);
xor U24221 (N_24221,N_16024,N_17690);
and U24222 (N_24222,N_16409,N_15751);
and U24223 (N_24223,N_17926,N_16370);
nor U24224 (N_24224,N_19262,N_19493);
or U24225 (N_24225,N_17196,N_17041);
or U24226 (N_24226,N_19427,N_17896);
nand U24227 (N_24227,N_15737,N_15218);
and U24228 (N_24228,N_18042,N_16765);
xnor U24229 (N_24229,N_17204,N_17137);
and U24230 (N_24230,N_17831,N_17572);
nor U24231 (N_24231,N_16605,N_15456);
or U24232 (N_24232,N_19092,N_18597);
nor U24233 (N_24233,N_15108,N_18435);
or U24234 (N_24234,N_18199,N_19487);
nand U24235 (N_24235,N_17907,N_18708);
nor U24236 (N_24236,N_16948,N_19219);
or U24237 (N_24237,N_15042,N_18740);
nor U24238 (N_24238,N_19341,N_19510);
nand U24239 (N_24239,N_19242,N_19013);
and U24240 (N_24240,N_19627,N_17003);
xor U24241 (N_24241,N_15675,N_16757);
and U24242 (N_24242,N_19664,N_19318);
nor U24243 (N_24243,N_16744,N_17914);
nand U24244 (N_24244,N_15221,N_16970);
and U24245 (N_24245,N_16007,N_15737);
and U24246 (N_24246,N_15142,N_19796);
xnor U24247 (N_24247,N_17635,N_19958);
nand U24248 (N_24248,N_18238,N_19697);
and U24249 (N_24249,N_18962,N_17535);
nand U24250 (N_24250,N_16562,N_19553);
nand U24251 (N_24251,N_19947,N_17139);
and U24252 (N_24252,N_15087,N_17102);
nand U24253 (N_24253,N_15023,N_15633);
or U24254 (N_24254,N_17790,N_18469);
or U24255 (N_24255,N_17607,N_19608);
xnor U24256 (N_24256,N_19485,N_17720);
nor U24257 (N_24257,N_18508,N_18550);
xnor U24258 (N_24258,N_15120,N_18283);
and U24259 (N_24259,N_19803,N_15333);
xnor U24260 (N_24260,N_16660,N_19258);
nor U24261 (N_24261,N_15351,N_16584);
and U24262 (N_24262,N_16415,N_19534);
or U24263 (N_24263,N_17445,N_18095);
xor U24264 (N_24264,N_19653,N_19670);
xnor U24265 (N_24265,N_15197,N_19972);
nand U24266 (N_24266,N_16456,N_18565);
and U24267 (N_24267,N_16827,N_17638);
nor U24268 (N_24268,N_16210,N_17847);
and U24269 (N_24269,N_16181,N_15581);
and U24270 (N_24270,N_15777,N_18508);
or U24271 (N_24271,N_16798,N_18170);
xor U24272 (N_24272,N_17210,N_15903);
xor U24273 (N_24273,N_18946,N_16061);
or U24274 (N_24274,N_17227,N_17798);
and U24275 (N_24275,N_15293,N_18190);
or U24276 (N_24276,N_19776,N_18639);
and U24277 (N_24277,N_16816,N_18490);
nand U24278 (N_24278,N_16742,N_16917);
nand U24279 (N_24279,N_18033,N_16925);
nand U24280 (N_24280,N_19985,N_17539);
nor U24281 (N_24281,N_17643,N_17319);
and U24282 (N_24282,N_15156,N_17434);
or U24283 (N_24283,N_19546,N_19214);
nand U24284 (N_24284,N_15066,N_19324);
nand U24285 (N_24285,N_16967,N_15083);
nor U24286 (N_24286,N_15142,N_16522);
xor U24287 (N_24287,N_15606,N_17997);
xnor U24288 (N_24288,N_17909,N_18109);
nor U24289 (N_24289,N_16433,N_18914);
nand U24290 (N_24290,N_19371,N_15249);
nand U24291 (N_24291,N_16972,N_15844);
nor U24292 (N_24292,N_19088,N_18664);
xnor U24293 (N_24293,N_17551,N_18136);
nor U24294 (N_24294,N_16440,N_18138);
nand U24295 (N_24295,N_15943,N_15039);
xor U24296 (N_24296,N_16132,N_15609);
nor U24297 (N_24297,N_15179,N_15918);
xor U24298 (N_24298,N_18577,N_16309);
nor U24299 (N_24299,N_17854,N_17427);
nor U24300 (N_24300,N_16289,N_16473);
and U24301 (N_24301,N_19361,N_19312);
xor U24302 (N_24302,N_19252,N_16335);
or U24303 (N_24303,N_16110,N_16301);
xor U24304 (N_24304,N_15883,N_18196);
or U24305 (N_24305,N_18395,N_16239);
nand U24306 (N_24306,N_18628,N_17639);
nor U24307 (N_24307,N_17005,N_16071);
nand U24308 (N_24308,N_16432,N_17263);
nand U24309 (N_24309,N_19572,N_19721);
and U24310 (N_24310,N_17968,N_17197);
and U24311 (N_24311,N_19737,N_16029);
nor U24312 (N_24312,N_17614,N_16385);
or U24313 (N_24313,N_18189,N_17352);
and U24314 (N_24314,N_15867,N_17878);
nand U24315 (N_24315,N_15767,N_15068);
or U24316 (N_24316,N_19578,N_17296);
xor U24317 (N_24317,N_19076,N_17683);
nor U24318 (N_24318,N_16316,N_19356);
and U24319 (N_24319,N_18949,N_19696);
nor U24320 (N_24320,N_19729,N_16460);
or U24321 (N_24321,N_19479,N_17178);
xor U24322 (N_24322,N_16881,N_17286);
nand U24323 (N_24323,N_19349,N_18550);
or U24324 (N_24324,N_16390,N_19450);
xor U24325 (N_24325,N_18329,N_18800);
and U24326 (N_24326,N_15174,N_15033);
xnor U24327 (N_24327,N_15678,N_16702);
nor U24328 (N_24328,N_19045,N_18774);
nand U24329 (N_24329,N_18251,N_15220);
or U24330 (N_24330,N_18282,N_18645);
and U24331 (N_24331,N_17057,N_17504);
xor U24332 (N_24332,N_19222,N_16590);
nor U24333 (N_24333,N_19154,N_17386);
or U24334 (N_24334,N_19815,N_18008);
nand U24335 (N_24335,N_17893,N_19033);
nor U24336 (N_24336,N_17231,N_16479);
nor U24337 (N_24337,N_17037,N_15684);
and U24338 (N_24338,N_15756,N_18771);
or U24339 (N_24339,N_16206,N_18093);
xor U24340 (N_24340,N_19512,N_17347);
or U24341 (N_24341,N_16534,N_17270);
and U24342 (N_24342,N_17933,N_15925);
nand U24343 (N_24343,N_17874,N_18162);
and U24344 (N_24344,N_17611,N_18641);
and U24345 (N_24345,N_19779,N_17294);
and U24346 (N_24346,N_18747,N_15848);
or U24347 (N_24347,N_17136,N_18935);
and U24348 (N_24348,N_17735,N_16463);
or U24349 (N_24349,N_15254,N_16879);
xor U24350 (N_24350,N_19699,N_19737);
nand U24351 (N_24351,N_16631,N_18858);
or U24352 (N_24352,N_19740,N_17248);
xor U24353 (N_24353,N_18041,N_18866);
nor U24354 (N_24354,N_16814,N_19383);
nor U24355 (N_24355,N_19501,N_16572);
nand U24356 (N_24356,N_16733,N_17098);
nand U24357 (N_24357,N_15456,N_18545);
or U24358 (N_24358,N_19471,N_16994);
nand U24359 (N_24359,N_16355,N_19846);
nand U24360 (N_24360,N_16301,N_18507);
nand U24361 (N_24361,N_15781,N_18870);
nand U24362 (N_24362,N_19813,N_19749);
nor U24363 (N_24363,N_15396,N_15168);
nand U24364 (N_24364,N_19067,N_18790);
and U24365 (N_24365,N_19719,N_19071);
or U24366 (N_24366,N_18650,N_15771);
xnor U24367 (N_24367,N_15142,N_17385);
or U24368 (N_24368,N_19102,N_18281);
xor U24369 (N_24369,N_16818,N_17284);
xnor U24370 (N_24370,N_19609,N_19447);
nor U24371 (N_24371,N_17624,N_18808);
nor U24372 (N_24372,N_19560,N_19317);
or U24373 (N_24373,N_17677,N_16301);
or U24374 (N_24374,N_16577,N_15381);
xor U24375 (N_24375,N_15654,N_15245);
or U24376 (N_24376,N_17006,N_16280);
or U24377 (N_24377,N_17129,N_17235);
or U24378 (N_24378,N_17986,N_19311);
or U24379 (N_24379,N_15825,N_16658);
xnor U24380 (N_24380,N_19640,N_17399);
and U24381 (N_24381,N_15338,N_18660);
nand U24382 (N_24382,N_15284,N_17467);
or U24383 (N_24383,N_16803,N_15173);
and U24384 (N_24384,N_16482,N_16764);
nor U24385 (N_24385,N_16244,N_17081);
nor U24386 (N_24386,N_19140,N_16475);
nand U24387 (N_24387,N_15524,N_16883);
nor U24388 (N_24388,N_16445,N_18456);
xnor U24389 (N_24389,N_19520,N_17212);
nand U24390 (N_24390,N_15927,N_15501);
and U24391 (N_24391,N_16747,N_18974);
or U24392 (N_24392,N_17662,N_18877);
or U24393 (N_24393,N_16469,N_18739);
or U24394 (N_24394,N_19544,N_18839);
xnor U24395 (N_24395,N_18047,N_16012);
and U24396 (N_24396,N_19490,N_18465);
and U24397 (N_24397,N_19338,N_17591);
nor U24398 (N_24398,N_15054,N_16370);
or U24399 (N_24399,N_15165,N_18934);
and U24400 (N_24400,N_15586,N_15748);
nand U24401 (N_24401,N_17866,N_18994);
or U24402 (N_24402,N_18530,N_17035);
nand U24403 (N_24403,N_16570,N_17801);
and U24404 (N_24404,N_18437,N_17252);
nor U24405 (N_24405,N_19101,N_19316);
nand U24406 (N_24406,N_16576,N_16648);
and U24407 (N_24407,N_18673,N_19133);
nand U24408 (N_24408,N_16106,N_17797);
xor U24409 (N_24409,N_18181,N_15134);
or U24410 (N_24410,N_18421,N_18792);
nor U24411 (N_24411,N_16299,N_17282);
nand U24412 (N_24412,N_15561,N_18146);
and U24413 (N_24413,N_17646,N_17580);
xor U24414 (N_24414,N_19173,N_19923);
and U24415 (N_24415,N_16650,N_18501);
xnor U24416 (N_24416,N_19970,N_15795);
nand U24417 (N_24417,N_15797,N_15236);
nand U24418 (N_24418,N_16731,N_16526);
nand U24419 (N_24419,N_16267,N_17733);
nand U24420 (N_24420,N_15012,N_16710);
xnor U24421 (N_24421,N_18096,N_17043);
xnor U24422 (N_24422,N_17357,N_15899);
xnor U24423 (N_24423,N_19832,N_15237);
nand U24424 (N_24424,N_19313,N_16392);
xor U24425 (N_24425,N_19107,N_15979);
nor U24426 (N_24426,N_16703,N_18865);
xnor U24427 (N_24427,N_16631,N_16468);
and U24428 (N_24428,N_18214,N_16268);
nor U24429 (N_24429,N_17815,N_16984);
and U24430 (N_24430,N_15088,N_17105);
nand U24431 (N_24431,N_18319,N_18005);
or U24432 (N_24432,N_15621,N_18402);
and U24433 (N_24433,N_17229,N_18782);
xnor U24434 (N_24434,N_19479,N_19013);
xor U24435 (N_24435,N_16334,N_18468);
nor U24436 (N_24436,N_16342,N_16907);
nand U24437 (N_24437,N_17614,N_17078);
nand U24438 (N_24438,N_18339,N_16539);
and U24439 (N_24439,N_16925,N_17446);
xnor U24440 (N_24440,N_18905,N_19435);
and U24441 (N_24441,N_17618,N_17127);
nand U24442 (N_24442,N_17306,N_15072);
nor U24443 (N_24443,N_18394,N_16244);
or U24444 (N_24444,N_15399,N_16924);
and U24445 (N_24445,N_16926,N_15492);
xor U24446 (N_24446,N_19220,N_16261);
nor U24447 (N_24447,N_15672,N_15885);
and U24448 (N_24448,N_18181,N_18798);
nor U24449 (N_24449,N_17283,N_16294);
or U24450 (N_24450,N_17868,N_15830);
nor U24451 (N_24451,N_15468,N_18360);
and U24452 (N_24452,N_15271,N_17469);
nor U24453 (N_24453,N_16552,N_19194);
xnor U24454 (N_24454,N_15393,N_17889);
and U24455 (N_24455,N_16588,N_17828);
nand U24456 (N_24456,N_18918,N_15770);
or U24457 (N_24457,N_17320,N_19097);
xnor U24458 (N_24458,N_18498,N_19868);
xor U24459 (N_24459,N_15757,N_19435);
xnor U24460 (N_24460,N_16803,N_16413);
or U24461 (N_24461,N_15481,N_18079);
nand U24462 (N_24462,N_19430,N_18051);
nor U24463 (N_24463,N_16817,N_15413);
xnor U24464 (N_24464,N_19616,N_15112);
nand U24465 (N_24465,N_15612,N_17873);
nor U24466 (N_24466,N_17645,N_18775);
xnor U24467 (N_24467,N_19022,N_19601);
or U24468 (N_24468,N_17338,N_19790);
xor U24469 (N_24469,N_16695,N_17824);
and U24470 (N_24470,N_15184,N_19845);
or U24471 (N_24471,N_18169,N_19338);
or U24472 (N_24472,N_16007,N_16053);
nor U24473 (N_24473,N_15841,N_18333);
xnor U24474 (N_24474,N_18512,N_18284);
or U24475 (N_24475,N_18611,N_15248);
or U24476 (N_24476,N_19432,N_15212);
or U24477 (N_24477,N_19995,N_15508);
xnor U24478 (N_24478,N_17560,N_19946);
nand U24479 (N_24479,N_16517,N_19589);
xnor U24480 (N_24480,N_17723,N_15400);
or U24481 (N_24481,N_16130,N_15688);
nand U24482 (N_24482,N_17653,N_15640);
nand U24483 (N_24483,N_15339,N_15014);
and U24484 (N_24484,N_19647,N_18818);
and U24485 (N_24485,N_15478,N_15755);
and U24486 (N_24486,N_15072,N_18889);
xnor U24487 (N_24487,N_15491,N_19675);
and U24488 (N_24488,N_17800,N_16777);
or U24489 (N_24489,N_19173,N_18941);
nor U24490 (N_24490,N_16194,N_19318);
xor U24491 (N_24491,N_18009,N_19119);
and U24492 (N_24492,N_16317,N_18687);
xor U24493 (N_24493,N_17958,N_16559);
and U24494 (N_24494,N_16611,N_15176);
nand U24495 (N_24495,N_17983,N_17562);
nor U24496 (N_24496,N_15255,N_18137);
nor U24497 (N_24497,N_17359,N_15254);
xor U24498 (N_24498,N_16266,N_15082);
xor U24499 (N_24499,N_17308,N_15450);
and U24500 (N_24500,N_19375,N_16187);
or U24501 (N_24501,N_18213,N_15695);
xnor U24502 (N_24502,N_16775,N_18544);
nor U24503 (N_24503,N_16113,N_17933);
and U24504 (N_24504,N_15162,N_18835);
or U24505 (N_24505,N_15309,N_17703);
and U24506 (N_24506,N_16647,N_16135);
nor U24507 (N_24507,N_17411,N_19732);
nand U24508 (N_24508,N_17341,N_15986);
xnor U24509 (N_24509,N_15239,N_19523);
or U24510 (N_24510,N_17195,N_15029);
nand U24511 (N_24511,N_15816,N_15283);
or U24512 (N_24512,N_17109,N_18770);
xnor U24513 (N_24513,N_16609,N_16698);
and U24514 (N_24514,N_18838,N_17370);
and U24515 (N_24515,N_16983,N_15369);
nand U24516 (N_24516,N_16835,N_18497);
nor U24517 (N_24517,N_15091,N_17241);
xnor U24518 (N_24518,N_19978,N_15079);
nor U24519 (N_24519,N_15687,N_18816);
nand U24520 (N_24520,N_19541,N_18365);
or U24521 (N_24521,N_19623,N_17282);
nor U24522 (N_24522,N_18388,N_19652);
or U24523 (N_24523,N_17442,N_17053);
xnor U24524 (N_24524,N_19764,N_16198);
xor U24525 (N_24525,N_15024,N_19634);
nor U24526 (N_24526,N_18389,N_15228);
and U24527 (N_24527,N_17116,N_15123);
nor U24528 (N_24528,N_17351,N_17016);
and U24529 (N_24529,N_18444,N_17928);
nor U24530 (N_24530,N_18523,N_17135);
nor U24531 (N_24531,N_16258,N_17466);
xor U24532 (N_24532,N_19125,N_15949);
xor U24533 (N_24533,N_19763,N_18236);
nor U24534 (N_24534,N_19812,N_15083);
nor U24535 (N_24535,N_15687,N_17499);
or U24536 (N_24536,N_17422,N_17395);
nor U24537 (N_24537,N_17593,N_18318);
nand U24538 (N_24538,N_15934,N_15149);
xor U24539 (N_24539,N_19422,N_17638);
xnor U24540 (N_24540,N_17642,N_15006);
or U24541 (N_24541,N_15075,N_19450);
nor U24542 (N_24542,N_15542,N_17261);
nand U24543 (N_24543,N_17379,N_16060);
or U24544 (N_24544,N_18889,N_18604);
and U24545 (N_24545,N_18294,N_18076);
nor U24546 (N_24546,N_15412,N_15500);
nand U24547 (N_24547,N_16213,N_19478);
and U24548 (N_24548,N_16227,N_16554);
nand U24549 (N_24549,N_18922,N_19965);
nand U24550 (N_24550,N_19922,N_16700);
or U24551 (N_24551,N_15393,N_16526);
and U24552 (N_24552,N_15294,N_19303);
and U24553 (N_24553,N_19073,N_16503);
xnor U24554 (N_24554,N_18457,N_15845);
xor U24555 (N_24555,N_17262,N_15949);
nor U24556 (N_24556,N_17677,N_17091);
nor U24557 (N_24557,N_17875,N_17230);
and U24558 (N_24558,N_19665,N_16764);
nor U24559 (N_24559,N_17953,N_15264);
xor U24560 (N_24560,N_16057,N_15634);
nand U24561 (N_24561,N_19998,N_18228);
xnor U24562 (N_24562,N_19186,N_18439);
nand U24563 (N_24563,N_17786,N_16943);
nor U24564 (N_24564,N_19540,N_19302);
and U24565 (N_24565,N_16740,N_17582);
or U24566 (N_24566,N_15341,N_18853);
and U24567 (N_24567,N_17939,N_16120);
and U24568 (N_24568,N_18367,N_19452);
nand U24569 (N_24569,N_18479,N_17780);
nor U24570 (N_24570,N_15900,N_18851);
nand U24571 (N_24571,N_15095,N_15241);
nor U24572 (N_24572,N_17559,N_16977);
nand U24573 (N_24573,N_16305,N_15063);
xnor U24574 (N_24574,N_15116,N_19446);
and U24575 (N_24575,N_15089,N_15189);
xor U24576 (N_24576,N_16349,N_17172);
nor U24577 (N_24577,N_15874,N_18569);
nor U24578 (N_24578,N_18460,N_17018);
or U24579 (N_24579,N_16467,N_17036);
xnor U24580 (N_24580,N_19177,N_18699);
nand U24581 (N_24581,N_16340,N_17151);
nand U24582 (N_24582,N_15904,N_18414);
or U24583 (N_24583,N_16859,N_18597);
nor U24584 (N_24584,N_18141,N_15595);
xnor U24585 (N_24585,N_17934,N_16335);
nor U24586 (N_24586,N_15808,N_16883);
and U24587 (N_24587,N_19033,N_19423);
xor U24588 (N_24588,N_18825,N_19181);
nor U24589 (N_24589,N_15390,N_17859);
xor U24590 (N_24590,N_16814,N_18842);
nor U24591 (N_24591,N_19279,N_18784);
xor U24592 (N_24592,N_19074,N_17505);
nand U24593 (N_24593,N_18283,N_15995);
xor U24594 (N_24594,N_18212,N_18713);
nor U24595 (N_24595,N_18846,N_16081);
and U24596 (N_24596,N_19586,N_16166);
nand U24597 (N_24597,N_17873,N_17760);
and U24598 (N_24598,N_16246,N_18015);
nand U24599 (N_24599,N_16135,N_15771);
xor U24600 (N_24600,N_18940,N_19415);
nand U24601 (N_24601,N_17968,N_17077);
nand U24602 (N_24602,N_16917,N_16214);
xor U24603 (N_24603,N_19249,N_19629);
xnor U24604 (N_24604,N_17900,N_19813);
nand U24605 (N_24605,N_16506,N_15862);
xnor U24606 (N_24606,N_18126,N_19097);
and U24607 (N_24607,N_19122,N_17021);
nand U24608 (N_24608,N_15222,N_18040);
and U24609 (N_24609,N_15742,N_15476);
xnor U24610 (N_24610,N_18543,N_17432);
nor U24611 (N_24611,N_19702,N_17242);
nand U24612 (N_24612,N_15208,N_18721);
xnor U24613 (N_24613,N_18239,N_18287);
xor U24614 (N_24614,N_18347,N_18918);
nand U24615 (N_24615,N_15617,N_18974);
or U24616 (N_24616,N_19972,N_17044);
xor U24617 (N_24617,N_19958,N_16069);
nand U24618 (N_24618,N_17571,N_15826);
or U24619 (N_24619,N_18034,N_17705);
and U24620 (N_24620,N_15726,N_17587);
nand U24621 (N_24621,N_17572,N_19820);
nand U24622 (N_24622,N_15801,N_15138);
xor U24623 (N_24623,N_17929,N_15637);
nor U24624 (N_24624,N_16780,N_19023);
or U24625 (N_24625,N_16084,N_16792);
or U24626 (N_24626,N_19473,N_15622);
or U24627 (N_24627,N_19460,N_16845);
and U24628 (N_24628,N_15433,N_15340);
nand U24629 (N_24629,N_18274,N_17802);
nor U24630 (N_24630,N_16576,N_17440);
and U24631 (N_24631,N_16358,N_17374);
and U24632 (N_24632,N_19571,N_18008);
nand U24633 (N_24633,N_16991,N_16279);
or U24634 (N_24634,N_18563,N_19340);
or U24635 (N_24635,N_17066,N_16665);
nor U24636 (N_24636,N_18871,N_16859);
xnor U24637 (N_24637,N_17664,N_15587);
and U24638 (N_24638,N_19672,N_19482);
or U24639 (N_24639,N_15822,N_15820);
or U24640 (N_24640,N_15921,N_17549);
and U24641 (N_24641,N_18229,N_15710);
nand U24642 (N_24642,N_15683,N_15015);
nand U24643 (N_24643,N_15230,N_18902);
or U24644 (N_24644,N_19044,N_16306);
nor U24645 (N_24645,N_17588,N_15826);
xnor U24646 (N_24646,N_15223,N_16643);
xor U24647 (N_24647,N_18423,N_18331);
xnor U24648 (N_24648,N_18055,N_18297);
or U24649 (N_24649,N_19777,N_17925);
and U24650 (N_24650,N_18117,N_17321);
nor U24651 (N_24651,N_19983,N_19913);
nor U24652 (N_24652,N_15696,N_15764);
or U24653 (N_24653,N_15292,N_19479);
or U24654 (N_24654,N_15018,N_17206);
nand U24655 (N_24655,N_15382,N_19314);
nor U24656 (N_24656,N_16526,N_19915);
nor U24657 (N_24657,N_17296,N_17223);
or U24658 (N_24658,N_17688,N_19976);
or U24659 (N_24659,N_15557,N_15523);
or U24660 (N_24660,N_18411,N_19720);
or U24661 (N_24661,N_15773,N_15802);
and U24662 (N_24662,N_19078,N_15139);
and U24663 (N_24663,N_19926,N_18584);
nor U24664 (N_24664,N_17361,N_18812);
or U24665 (N_24665,N_19200,N_17784);
and U24666 (N_24666,N_16882,N_16414);
and U24667 (N_24667,N_18525,N_17604);
xor U24668 (N_24668,N_18048,N_16312);
nand U24669 (N_24669,N_19849,N_18619);
xnor U24670 (N_24670,N_19599,N_19816);
nand U24671 (N_24671,N_19196,N_17057);
xor U24672 (N_24672,N_15788,N_18704);
nor U24673 (N_24673,N_16961,N_16650);
nand U24674 (N_24674,N_17379,N_15353);
nand U24675 (N_24675,N_16058,N_18516);
and U24676 (N_24676,N_17256,N_16829);
xor U24677 (N_24677,N_16011,N_18407);
xor U24678 (N_24678,N_19847,N_17012);
and U24679 (N_24679,N_15060,N_15532);
nor U24680 (N_24680,N_16479,N_16035);
xnor U24681 (N_24681,N_15216,N_18053);
and U24682 (N_24682,N_16051,N_16772);
and U24683 (N_24683,N_15770,N_17165);
and U24684 (N_24684,N_15006,N_18131);
and U24685 (N_24685,N_19088,N_17741);
or U24686 (N_24686,N_15499,N_17619);
xnor U24687 (N_24687,N_18415,N_15177);
nor U24688 (N_24688,N_19653,N_18044);
or U24689 (N_24689,N_17624,N_15863);
xor U24690 (N_24690,N_18152,N_19814);
or U24691 (N_24691,N_15367,N_17303);
xnor U24692 (N_24692,N_18330,N_15234);
nand U24693 (N_24693,N_17222,N_16119);
nor U24694 (N_24694,N_16357,N_17025);
or U24695 (N_24695,N_17519,N_19801);
nor U24696 (N_24696,N_16408,N_15920);
nand U24697 (N_24697,N_17438,N_18132);
and U24698 (N_24698,N_17474,N_15906);
nand U24699 (N_24699,N_18095,N_15684);
or U24700 (N_24700,N_16550,N_15715);
or U24701 (N_24701,N_18714,N_19297);
nor U24702 (N_24702,N_18605,N_19558);
and U24703 (N_24703,N_17133,N_15642);
and U24704 (N_24704,N_16855,N_15573);
or U24705 (N_24705,N_18521,N_15898);
xnor U24706 (N_24706,N_15677,N_18196);
or U24707 (N_24707,N_15631,N_15553);
nor U24708 (N_24708,N_18756,N_15864);
nand U24709 (N_24709,N_19773,N_19770);
nor U24710 (N_24710,N_17770,N_16330);
and U24711 (N_24711,N_18169,N_16566);
xnor U24712 (N_24712,N_17907,N_16005);
nor U24713 (N_24713,N_18294,N_19295);
nand U24714 (N_24714,N_17435,N_19993);
nand U24715 (N_24715,N_15721,N_19484);
nor U24716 (N_24716,N_19386,N_17221);
or U24717 (N_24717,N_19532,N_17784);
and U24718 (N_24718,N_16942,N_18560);
or U24719 (N_24719,N_16561,N_18890);
and U24720 (N_24720,N_16833,N_15572);
xnor U24721 (N_24721,N_18967,N_17225);
or U24722 (N_24722,N_16413,N_16667);
nor U24723 (N_24723,N_17995,N_15993);
nand U24724 (N_24724,N_18481,N_19142);
xor U24725 (N_24725,N_18467,N_18161);
nor U24726 (N_24726,N_16252,N_19725);
nand U24727 (N_24727,N_19909,N_15565);
or U24728 (N_24728,N_16286,N_18796);
xor U24729 (N_24729,N_17327,N_15563);
and U24730 (N_24730,N_18712,N_15837);
nor U24731 (N_24731,N_16711,N_17770);
or U24732 (N_24732,N_16127,N_17994);
and U24733 (N_24733,N_17037,N_18038);
or U24734 (N_24734,N_18966,N_16928);
or U24735 (N_24735,N_18548,N_15745);
and U24736 (N_24736,N_16939,N_19479);
nor U24737 (N_24737,N_18026,N_18609);
and U24738 (N_24738,N_17591,N_16829);
nand U24739 (N_24739,N_18401,N_18714);
nor U24740 (N_24740,N_16689,N_17998);
nor U24741 (N_24741,N_15232,N_17877);
and U24742 (N_24742,N_16331,N_16843);
xor U24743 (N_24743,N_19449,N_19656);
xnor U24744 (N_24744,N_15726,N_19564);
nand U24745 (N_24745,N_19300,N_15596);
nor U24746 (N_24746,N_15703,N_17020);
nand U24747 (N_24747,N_15358,N_19312);
nand U24748 (N_24748,N_16261,N_15509);
or U24749 (N_24749,N_18031,N_16614);
xor U24750 (N_24750,N_17783,N_19059);
nand U24751 (N_24751,N_17643,N_16470);
nor U24752 (N_24752,N_18424,N_19263);
or U24753 (N_24753,N_15927,N_19872);
xor U24754 (N_24754,N_19653,N_19625);
and U24755 (N_24755,N_17225,N_18147);
nor U24756 (N_24756,N_17292,N_17670);
xor U24757 (N_24757,N_19909,N_17781);
and U24758 (N_24758,N_15721,N_19382);
nand U24759 (N_24759,N_18290,N_15605);
xor U24760 (N_24760,N_15402,N_19566);
or U24761 (N_24761,N_19029,N_16743);
xnor U24762 (N_24762,N_18628,N_18534);
nor U24763 (N_24763,N_15400,N_15249);
xnor U24764 (N_24764,N_19801,N_16576);
or U24765 (N_24765,N_19335,N_17324);
xnor U24766 (N_24766,N_19920,N_17188);
nand U24767 (N_24767,N_19375,N_17759);
nand U24768 (N_24768,N_19602,N_19273);
nor U24769 (N_24769,N_17994,N_15066);
and U24770 (N_24770,N_16663,N_15402);
xor U24771 (N_24771,N_19368,N_15911);
nor U24772 (N_24772,N_17439,N_15554);
nor U24773 (N_24773,N_19363,N_17640);
xnor U24774 (N_24774,N_16513,N_19090);
or U24775 (N_24775,N_18415,N_19343);
and U24776 (N_24776,N_16980,N_17334);
nor U24777 (N_24777,N_17997,N_19167);
or U24778 (N_24778,N_16874,N_15177);
xor U24779 (N_24779,N_15102,N_19616);
nor U24780 (N_24780,N_17927,N_15439);
and U24781 (N_24781,N_15406,N_16457);
nor U24782 (N_24782,N_19276,N_17145);
nor U24783 (N_24783,N_18917,N_17816);
and U24784 (N_24784,N_16616,N_16875);
nor U24785 (N_24785,N_15434,N_15575);
and U24786 (N_24786,N_15884,N_17904);
nor U24787 (N_24787,N_15226,N_16733);
nand U24788 (N_24788,N_15280,N_17993);
nand U24789 (N_24789,N_19370,N_15440);
xnor U24790 (N_24790,N_16684,N_19000);
xor U24791 (N_24791,N_15553,N_18170);
nand U24792 (N_24792,N_17519,N_16768);
nor U24793 (N_24793,N_16840,N_16588);
and U24794 (N_24794,N_17152,N_16555);
and U24795 (N_24795,N_18506,N_15136);
and U24796 (N_24796,N_19868,N_16053);
xnor U24797 (N_24797,N_18974,N_19261);
and U24798 (N_24798,N_17307,N_19559);
nand U24799 (N_24799,N_15184,N_19606);
or U24800 (N_24800,N_15544,N_17323);
or U24801 (N_24801,N_19586,N_17514);
nor U24802 (N_24802,N_17139,N_19567);
xnor U24803 (N_24803,N_17519,N_17866);
and U24804 (N_24804,N_17567,N_16427);
xnor U24805 (N_24805,N_16487,N_17215);
nor U24806 (N_24806,N_19332,N_18187);
xnor U24807 (N_24807,N_17385,N_15989);
and U24808 (N_24808,N_15210,N_15396);
nand U24809 (N_24809,N_18604,N_18526);
nor U24810 (N_24810,N_16979,N_17788);
or U24811 (N_24811,N_17182,N_19354);
and U24812 (N_24812,N_18109,N_15355);
nand U24813 (N_24813,N_15916,N_19303);
and U24814 (N_24814,N_16299,N_19250);
and U24815 (N_24815,N_16025,N_17829);
or U24816 (N_24816,N_15316,N_18867);
nand U24817 (N_24817,N_19067,N_17241);
nor U24818 (N_24818,N_16129,N_18204);
xor U24819 (N_24819,N_19180,N_18145);
xnor U24820 (N_24820,N_19208,N_17195);
xor U24821 (N_24821,N_19458,N_17071);
xnor U24822 (N_24822,N_15718,N_16684);
xnor U24823 (N_24823,N_18078,N_17268);
or U24824 (N_24824,N_19190,N_15211);
or U24825 (N_24825,N_17127,N_16196);
nand U24826 (N_24826,N_18888,N_18968);
xnor U24827 (N_24827,N_15689,N_18928);
or U24828 (N_24828,N_19636,N_15210);
or U24829 (N_24829,N_15253,N_19315);
nor U24830 (N_24830,N_16165,N_15244);
nor U24831 (N_24831,N_16569,N_16589);
and U24832 (N_24832,N_18328,N_19411);
or U24833 (N_24833,N_19884,N_18898);
or U24834 (N_24834,N_15522,N_15588);
and U24835 (N_24835,N_19280,N_15282);
or U24836 (N_24836,N_19828,N_18353);
or U24837 (N_24837,N_19788,N_15551);
and U24838 (N_24838,N_16881,N_17674);
nor U24839 (N_24839,N_18395,N_18080);
xnor U24840 (N_24840,N_17789,N_18635);
and U24841 (N_24841,N_17523,N_16129);
and U24842 (N_24842,N_17708,N_19984);
xor U24843 (N_24843,N_19150,N_17321);
nand U24844 (N_24844,N_17249,N_17111);
and U24845 (N_24845,N_18247,N_18259);
xnor U24846 (N_24846,N_19353,N_18008);
and U24847 (N_24847,N_16569,N_19352);
xor U24848 (N_24848,N_15722,N_17451);
and U24849 (N_24849,N_18414,N_16025);
nand U24850 (N_24850,N_17325,N_18555);
nand U24851 (N_24851,N_17113,N_19223);
and U24852 (N_24852,N_19885,N_17034);
nor U24853 (N_24853,N_18087,N_19041);
nor U24854 (N_24854,N_17374,N_17221);
xnor U24855 (N_24855,N_16081,N_19682);
and U24856 (N_24856,N_19299,N_17013);
nor U24857 (N_24857,N_18490,N_16982);
nand U24858 (N_24858,N_15806,N_19994);
and U24859 (N_24859,N_17119,N_15111);
and U24860 (N_24860,N_18265,N_19466);
nor U24861 (N_24861,N_18349,N_17308);
or U24862 (N_24862,N_19628,N_19249);
nor U24863 (N_24863,N_19070,N_18541);
nand U24864 (N_24864,N_19412,N_16260);
nor U24865 (N_24865,N_19133,N_17424);
xor U24866 (N_24866,N_19835,N_17367);
and U24867 (N_24867,N_15523,N_16710);
or U24868 (N_24868,N_18267,N_19869);
xnor U24869 (N_24869,N_19328,N_18149);
or U24870 (N_24870,N_18290,N_15399);
nand U24871 (N_24871,N_19941,N_15015);
nand U24872 (N_24872,N_19411,N_15107);
nand U24873 (N_24873,N_15478,N_16900);
xnor U24874 (N_24874,N_15557,N_17241);
and U24875 (N_24875,N_18878,N_19793);
nand U24876 (N_24876,N_19597,N_15089);
nand U24877 (N_24877,N_16147,N_17625);
xnor U24878 (N_24878,N_16670,N_15808);
nor U24879 (N_24879,N_19481,N_16608);
nor U24880 (N_24880,N_17377,N_16453);
or U24881 (N_24881,N_18357,N_18620);
nand U24882 (N_24882,N_17303,N_17118);
and U24883 (N_24883,N_15886,N_15317);
xor U24884 (N_24884,N_17981,N_19885);
nor U24885 (N_24885,N_16744,N_17034);
nor U24886 (N_24886,N_16836,N_16238);
nor U24887 (N_24887,N_18485,N_19635);
or U24888 (N_24888,N_17771,N_18539);
or U24889 (N_24889,N_15234,N_19364);
xnor U24890 (N_24890,N_18609,N_19514);
xor U24891 (N_24891,N_17131,N_15688);
xor U24892 (N_24892,N_19934,N_16886);
xnor U24893 (N_24893,N_18229,N_15016);
nor U24894 (N_24894,N_17700,N_17895);
nand U24895 (N_24895,N_18726,N_17235);
or U24896 (N_24896,N_19852,N_17452);
nand U24897 (N_24897,N_15854,N_17915);
nor U24898 (N_24898,N_17063,N_18138);
and U24899 (N_24899,N_18100,N_16113);
nand U24900 (N_24900,N_16068,N_15250);
nand U24901 (N_24901,N_18219,N_17922);
nand U24902 (N_24902,N_18997,N_17662);
xnor U24903 (N_24903,N_15788,N_18509);
xor U24904 (N_24904,N_19539,N_16508);
and U24905 (N_24905,N_16899,N_17361);
nor U24906 (N_24906,N_16176,N_19074);
nand U24907 (N_24907,N_17490,N_18100);
nand U24908 (N_24908,N_16673,N_17542);
nand U24909 (N_24909,N_19720,N_17842);
xnor U24910 (N_24910,N_18527,N_19889);
or U24911 (N_24911,N_19070,N_15064);
or U24912 (N_24912,N_17786,N_19127);
nand U24913 (N_24913,N_18490,N_16882);
nor U24914 (N_24914,N_18659,N_16008);
nand U24915 (N_24915,N_17059,N_16700);
nand U24916 (N_24916,N_19627,N_17287);
xnor U24917 (N_24917,N_19679,N_16177);
and U24918 (N_24918,N_19437,N_16886);
xor U24919 (N_24919,N_18921,N_15515);
nor U24920 (N_24920,N_15972,N_16289);
nand U24921 (N_24921,N_18304,N_19121);
nor U24922 (N_24922,N_19664,N_18677);
xor U24923 (N_24923,N_15401,N_16052);
and U24924 (N_24924,N_18201,N_16409);
and U24925 (N_24925,N_15119,N_16001);
nand U24926 (N_24926,N_15116,N_17392);
and U24927 (N_24927,N_16792,N_15291);
xor U24928 (N_24928,N_17297,N_18980);
xor U24929 (N_24929,N_17385,N_18898);
and U24930 (N_24930,N_16438,N_19763);
and U24931 (N_24931,N_15866,N_19449);
nor U24932 (N_24932,N_17854,N_16511);
nand U24933 (N_24933,N_19746,N_15821);
xnor U24934 (N_24934,N_19445,N_18528);
or U24935 (N_24935,N_17300,N_15050);
or U24936 (N_24936,N_18214,N_15240);
or U24937 (N_24937,N_19042,N_18076);
nor U24938 (N_24938,N_18095,N_15543);
or U24939 (N_24939,N_19664,N_17216);
and U24940 (N_24940,N_19599,N_18584);
nor U24941 (N_24941,N_17286,N_19906);
nor U24942 (N_24942,N_16915,N_17827);
and U24943 (N_24943,N_16867,N_17460);
nand U24944 (N_24944,N_19915,N_19552);
or U24945 (N_24945,N_18913,N_17074);
nand U24946 (N_24946,N_17468,N_19977);
xor U24947 (N_24947,N_15193,N_17221);
xor U24948 (N_24948,N_15151,N_18092);
or U24949 (N_24949,N_17948,N_16410);
nand U24950 (N_24950,N_18652,N_16674);
nand U24951 (N_24951,N_18424,N_17928);
nand U24952 (N_24952,N_18552,N_19240);
nand U24953 (N_24953,N_16165,N_18223);
nor U24954 (N_24954,N_17131,N_18483);
xnor U24955 (N_24955,N_19579,N_19892);
or U24956 (N_24956,N_17521,N_17904);
nand U24957 (N_24957,N_19838,N_16534);
xor U24958 (N_24958,N_18118,N_18139);
xnor U24959 (N_24959,N_17236,N_17785);
nand U24960 (N_24960,N_15298,N_17489);
xnor U24961 (N_24961,N_19938,N_19251);
and U24962 (N_24962,N_17927,N_18214);
xor U24963 (N_24963,N_19003,N_18683);
and U24964 (N_24964,N_15777,N_16883);
xnor U24965 (N_24965,N_16882,N_16306);
xor U24966 (N_24966,N_18605,N_16961);
xor U24967 (N_24967,N_16068,N_17644);
and U24968 (N_24968,N_19730,N_15546);
nand U24969 (N_24969,N_18504,N_17377);
and U24970 (N_24970,N_19114,N_15089);
or U24971 (N_24971,N_18566,N_18763);
xor U24972 (N_24972,N_17272,N_18634);
xor U24973 (N_24973,N_19894,N_19251);
xnor U24974 (N_24974,N_15868,N_15701);
nor U24975 (N_24975,N_18644,N_19843);
and U24976 (N_24976,N_19574,N_19482);
xnor U24977 (N_24977,N_17708,N_19345);
nand U24978 (N_24978,N_16622,N_19481);
nand U24979 (N_24979,N_15247,N_15642);
nor U24980 (N_24980,N_15304,N_18664);
nand U24981 (N_24981,N_17049,N_17238);
or U24982 (N_24982,N_17899,N_17849);
xor U24983 (N_24983,N_15589,N_16125);
nor U24984 (N_24984,N_19862,N_19224);
nand U24985 (N_24985,N_19196,N_16579);
or U24986 (N_24986,N_18182,N_19398);
or U24987 (N_24987,N_16212,N_18050);
nor U24988 (N_24988,N_15994,N_19424);
xnor U24989 (N_24989,N_19029,N_15384);
nor U24990 (N_24990,N_18957,N_15225);
nor U24991 (N_24991,N_16533,N_16169);
nor U24992 (N_24992,N_17327,N_15389);
or U24993 (N_24993,N_18055,N_17301);
or U24994 (N_24994,N_16637,N_16636);
nand U24995 (N_24995,N_19153,N_19742);
or U24996 (N_24996,N_15833,N_15051);
xnor U24997 (N_24997,N_19908,N_19336);
nand U24998 (N_24998,N_15082,N_15508);
nor U24999 (N_24999,N_15456,N_18644);
and UO_0 (O_0,N_22568,N_23485);
and UO_1 (O_1,N_24953,N_22191);
nand UO_2 (O_2,N_21545,N_20899);
xnor UO_3 (O_3,N_21664,N_22424);
xor UO_4 (O_4,N_22462,N_24854);
and UO_5 (O_5,N_24926,N_23196);
or UO_6 (O_6,N_21230,N_23654);
and UO_7 (O_7,N_20529,N_24747);
and UO_8 (O_8,N_23110,N_20635);
xor UO_9 (O_9,N_20348,N_21048);
and UO_10 (O_10,N_20335,N_20065);
or UO_11 (O_11,N_20722,N_20841);
nor UO_12 (O_12,N_20552,N_24661);
nor UO_13 (O_13,N_24220,N_23496);
nand UO_14 (O_14,N_22924,N_20262);
nor UO_15 (O_15,N_24278,N_20819);
nand UO_16 (O_16,N_21764,N_20693);
xnor UO_17 (O_17,N_22987,N_20416);
or UO_18 (O_18,N_23600,N_20206);
nand UO_19 (O_19,N_24812,N_24343);
nor UO_20 (O_20,N_23574,N_24636);
xnor UO_21 (O_21,N_22877,N_20209);
nand UO_22 (O_22,N_20404,N_24786);
nand UO_23 (O_23,N_20421,N_22305);
nor UO_24 (O_24,N_20746,N_22100);
or UO_25 (O_25,N_23716,N_24690);
or UO_26 (O_26,N_24888,N_22923);
xor UO_27 (O_27,N_22774,N_22037);
nor UO_28 (O_28,N_24622,N_20756);
or UO_29 (O_29,N_21621,N_23165);
nand UO_30 (O_30,N_21487,N_20796);
and UO_31 (O_31,N_24961,N_23910);
xor UO_32 (O_32,N_21742,N_20266);
nor UO_33 (O_33,N_20627,N_20305);
or UO_34 (O_34,N_24190,N_24114);
xnor UO_35 (O_35,N_22115,N_21956);
nand UO_36 (O_36,N_21707,N_22123);
and UO_37 (O_37,N_24225,N_22434);
xnor UO_38 (O_38,N_21753,N_23514);
and UO_39 (O_39,N_24484,N_24852);
and UO_40 (O_40,N_23314,N_23011);
xor UO_41 (O_41,N_22018,N_23401);
xor UO_42 (O_42,N_20223,N_22512);
xor UO_43 (O_43,N_21242,N_23567);
nor UO_44 (O_44,N_24451,N_20770);
nor UO_45 (O_45,N_21321,N_21296);
xnor UO_46 (O_46,N_22164,N_23224);
nor UO_47 (O_47,N_20153,N_23946);
or UO_48 (O_48,N_21273,N_24535);
or UO_49 (O_49,N_23399,N_20343);
and UO_50 (O_50,N_24033,N_22937);
nand UO_51 (O_51,N_22093,N_23377);
nor UO_52 (O_52,N_23743,N_22428);
nand UO_53 (O_53,N_21421,N_24308);
and UO_54 (O_54,N_21770,N_23923);
nand UO_55 (O_55,N_20053,N_20879);
nand UO_56 (O_56,N_21258,N_22366);
and UO_57 (O_57,N_21805,N_22565);
nor UO_58 (O_58,N_21574,N_20917);
nor UO_59 (O_59,N_21915,N_23342);
nand UO_60 (O_60,N_20498,N_22386);
xnor UO_61 (O_61,N_22096,N_24376);
or UO_62 (O_62,N_23641,N_23777);
nand UO_63 (O_63,N_23788,N_20713);
nor UO_64 (O_64,N_23729,N_21370);
nor UO_65 (O_65,N_20540,N_23676);
and UO_66 (O_66,N_22874,N_23131);
and UO_67 (O_67,N_22084,N_24422);
or UO_68 (O_68,N_21138,N_22119);
xnor UO_69 (O_69,N_21969,N_22703);
xor UO_70 (O_70,N_20977,N_23499);
nor UO_71 (O_71,N_24840,N_22656);
xor UO_72 (O_72,N_24553,N_22620);
xor UO_73 (O_73,N_23215,N_21624);
and UO_74 (O_74,N_20547,N_22596);
or UO_75 (O_75,N_24265,N_20138);
nor UO_76 (O_76,N_24629,N_24122);
and UO_77 (O_77,N_22103,N_23116);
and UO_78 (O_78,N_24464,N_20821);
nand UO_79 (O_79,N_20754,N_21694);
xor UO_80 (O_80,N_20385,N_22251);
and UO_81 (O_81,N_21783,N_20414);
xor UO_82 (O_82,N_23697,N_23542);
or UO_83 (O_83,N_23631,N_21306);
nand UO_84 (O_84,N_23249,N_20439);
nor UO_85 (O_85,N_20594,N_24008);
nor UO_86 (O_86,N_24279,N_24657);
xor UO_87 (O_87,N_24152,N_22657);
xor UO_88 (O_88,N_23076,N_23546);
xor UO_89 (O_89,N_21420,N_24663);
nor UO_90 (O_90,N_23603,N_20884);
or UO_91 (O_91,N_22078,N_21367);
xor UO_92 (O_92,N_24654,N_22735);
nand UO_93 (O_93,N_24761,N_22441);
or UO_94 (O_94,N_22856,N_21374);
xnor UO_95 (O_95,N_21024,N_21814);
nand UO_96 (O_96,N_22531,N_20403);
nand UO_97 (O_97,N_22810,N_23101);
nor UO_98 (O_98,N_20241,N_24387);
or UO_99 (O_99,N_21442,N_23674);
nand UO_100 (O_100,N_20064,N_24179);
nor UO_101 (O_101,N_24277,N_24716);
xor UO_102 (O_102,N_21901,N_21887);
and UO_103 (O_103,N_23884,N_24861);
and UO_104 (O_104,N_23859,N_24669);
or UO_105 (O_105,N_22661,N_23559);
and UO_106 (O_106,N_24894,N_22057);
or UO_107 (O_107,N_22275,N_23509);
nand UO_108 (O_108,N_23338,N_20624);
or UO_109 (O_109,N_21137,N_23786);
or UO_110 (O_110,N_20597,N_21727);
xor UO_111 (O_111,N_24899,N_23558);
nor UO_112 (O_112,N_23779,N_24021);
nor UO_113 (O_113,N_23949,N_22396);
nand UO_114 (O_114,N_23590,N_24704);
nand UO_115 (O_115,N_24619,N_21775);
nor UO_116 (O_116,N_22163,N_22367);
or UO_117 (O_117,N_24738,N_22605);
or UO_118 (O_118,N_24943,N_20658);
or UO_119 (O_119,N_22910,N_24016);
xnor UO_120 (O_120,N_20657,N_22347);
or UO_121 (O_121,N_21762,N_22999);
xnor UO_122 (O_122,N_22371,N_20921);
or UO_123 (O_123,N_20025,N_24407);
xor UO_124 (O_124,N_20446,N_23646);
nor UO_125 (O_125,N_22876,N_21142);
nor UO_126 (O_126,N_21350,N_20397);
nor UO_127 (O_127,N_24583,N_20570);
nand UO_128 (O_128,N_21238,N_22209);
or UO_129 (O_129,N_22612,N_20018);
or UO_130 (O_130,N_20853,N_22246);
and UO_131 (O_131,N_24514,N_24784);
nor UO_132 (O_132,N_20393,N_20847);
and UO_133 (O_133,N_20974,N_21113);
and UO_134 (O_134,N_20950,N_24166);
nand UO_135 (O_135,N_20401,N_21106);
nand UO_136 (O_136,N_21553,N_22299);
nand UO_137 (O_137,N_22771,N_22598);
or UO_138 (O_138,N_20164,N_23041);
xor UO_139 (O_139,N_23166,N_21071);
nand UO_140 (O_140,N_20478,N_20792);
and UO_141 (O_141,N_24173,N_22981);
and UO_142 (O_142,N_21922,N_20830);
nand UO_143 (O_143,N_22268,N_23507);
xnor UO_144 (O_144,N_20508,N_21741);
and UO_145 (O_145,N_24141,N_20261);
and UO_146 (O_146,N_24104,N_23890);
and UO_147 (O_147,N_21865,N_22132);
and UO_148 (O_148,N_20121,N_22388);
or UO_149 (O_149,N_22936,N_21479);
or UO_150 (O_150,N_23421,N_24321);
or UO_151 (O_151,N_23580,N_23912);
xor UO_152 (O_152,N_24577,N_22368);
nor UO_153 (O_153,N_23585,N_21047);
nor UO_154 (O_154,N_20285,N_20060);
xnor UO_155 (O_155,N_22785,N_21074);
or UO_156 (O_156,N_23313,N_20212);
or UO_157 (O_157,N_22318,N_23353);
nor UO_158 (O_158,N_21703,N_22146);
and UO_159 (O_159,N_20844,N_24199);
nor UO_160 (O_160,N_23699,N_21403);
nand UO_161 (O_161,N_21299,N_24720);
xnor UO_162 (O_162,N_20311,N_23565);
or UO_163 (O_163,N_22486,N_21265);
nor UO_164 (O_164,N_22733,N_21755);
nand UO_165 (O_165,N_21037,N_23932);
or UO_166 (O_166,N_23067,N_22747);
nand UO_167 (O_167,N_24954,N_21376);
xor UO_168 (O_168,N_24805,N_24349);
nor UO_169 (O_169,N_23982,N_24102);
xor UO_170 (O_170,N_23023,N_23706);
xor UO_171 (O_171,N_22647,N_24071);
xor UO_172 (O_172,N_23944,N_24986);
nand UO_173 (O_173,N_20978,N_21651);
and UO_174 (O_174,N_24841,N_21267);
or UO_175 (O_175,N_21013,N_22862);
nand UO_176 (O_176,N_21986,N_22646);
nor UO_177 (O_177,N_23241,N_24785);
nor UO_178 (O_178,N_20837,N_23024);
or UO_179 (O_179,N_24453,N_23272);
and UO_180 (O_180,N_21114,N_22239);
xnor UO_181 (O_181,N_22896,N_20876);
nand UO_182 (O_182,N_20217,N_23075);
nand UO_183 (O_183,N_22282,N_21186);
nand UO_184 (O_184,N_23169,N_22286);
nand UO_185 (O_185,N_20278,N_20939);
nand UO_186 (O_186,N_20232,N_21638);
xor UO_187 (O_187,N_24649,N_21164);
xor UO_188 (O_188,N_20265,N_23945);
nor UO_189 (O_189,N_21700,N_21540);
nor UO_190 (O_190,N_20320,N_23667);
and UO_191 (O_191,N_20516,N_23091);
nand UO_192 (O_192,N_20264,N_24600);
nand UO_193 (O_193,N_24333,N_22935);
xor UO_194 (O_194,N_20805,N_22963);
xor UO_195 (O_195,N_22709,N_21518);
nor UO_196 (O_196,N_24616,N_20119);
or UO_197 (O_197,N_20398,N_21184);
xor UO_198 (O_198,N_23973,N_20755);
or UO_199 (O_199,N_24253,N_23818);
nand UO_200 (O_200,N_20992,N_20113);
or UO_201 (O_201,N_21368,N_21968);
nor UO_202 (O_202,N_24646,N_21171);
or UO_203 (O_203,N_22508,N_20733);
and UO_204 (O_204,N_23535,N_21493);
and UO_205 (O_205,N_24072,N_23597);
nor UO_206 (O_206,N_22603,N_24470);
nand UO_207 (O_207,N_23883,N_20681);
nor UO_208 (O_208,N_23275,N_20956);
and UO_209 (O_209,N_23727,N_21917);
xor UO_210 (O_210,N_24380,N_23294);
nor UO_211 (O_211,N_23336,N_24260);
and UO_212 (O_212,N_22839,N_22230);
or UO_213 (O_213,N_23301,N_22357);
or UO_214 (O_214,N_22138,N_20461);
nand UO_215 (O_215,N_22304,N_23791);
or UO_216 (O_216,N_24110,N_24196);
and UO_217 (O_217,N_20067,N_23714);
xnor UO_218 (O_218,N_24490,N_22331);
nor UO_219 (O_219,N_24215,N_24069);
xor UO_220 (O_220,N_22290,N_21528);
nor UO_221 (O_221,N_22002,N_22684);
nand UO_222 (O_222,N_23424,N_23137);
nor UO_223 (O_223,N_20730,N_24662);
nor UO_224 (O_224,N_22036,N_21226);
nand UO_225 (O_225,N_24753,N_22801);
and UO_226 (O_226,N_20344,N_21693);
xor UO_227 (O_227,N_21942,N_21434);
and UO_228 (O_228,N_20156,N_21837);
nor UO_229 (O_229,N_20833,N_23135);
and UO_230 (O_230,N_21369,N_22311);
and UO_231 (O_231,N_24755,N_20623);
or UO_232 (O_232,N_24117,N_22705);
xnor UO_233 (O_233,N_22653,N_24419);
nand UO_234 (O_234,N_20584,N_23445);
nand UO_235 (O_235,N_24549,N_21696);
nand UO_236 (O_236,N_23161,N_23007);
nand UO_237 (O_237,N_23010,N_23824);
and UO_238 (O_238,N_24214,N_22086);
nand UO_239 (O_239,N_22830,N_20774);
and UO_240 (O_240,N_21965,N_21132);
and UO_241 (O_241,N_23566,N_20790);
nand UO_242 (O_242,N_20500,N_20134);
and UO_243 (O_243,N_23680,N_24679);
and UO_244 (O_244,N_20896,N_23775);
nand UO_245 (O_245,N_23435,N_23709);
xor UO_246 (O_246,N_21169,N_22613);
nor UO_247 (O_247,N_20184,N_21061);
nand UO_248 (O_248,N_23873,N_24691);
or UO_249 (O_249,N_23929,N_21980);
nor UO_250 (O_250,N_24644,N_22624);
xnor UO_251 (O_251,N_21121,N_23891);
xnor UO_252 (O_252,N_21055,N_24133);
xor UO_253 (O_253,N_21890,N_24287);
nor UO_254 (O_254,N_23254,N_24829);
nand UO_255 (O_255,N_21235,N_20097);
nand UO_256 (O_256,N_22233,N_21019);
or UO_257 (O_257,N_22414,N_24517);
nand UO_258 (O_258,N_23947,N_23164);
and UO_259 (O_259,N_20129,N_24444);
and UO_260 (O_260,N_24292,N_21846);
xnor UO_261 (O_261,N_23831,N_23098);
xor UO_262 (O_262,N_23832,N_21615);
xor UO_263 (O_263,N_24269,N_20709);
nor UO_264 (O_264,N_21556,N_24031);
and UO_265 (O_265,N_21410,N_20870);
and UO_266 (O_266,N_23800,N_21692);
or UO_267 (O_267,N_24729,N_24226);
nor UO_268 (O_268,N_23466,N_22202);
and UO_269 (O_269,N_22600,N_20072);
xnor UO_270 (O_270,N_23820,N_24063);
nand UO_271 (O_271,N_20862,N_22675);
nor UO_272 (O_272,N_23853,N_22677);
nand UO_273 (O_273,N_21852,N_23815);
or UO_274 (O_274,N_22193,N_23359);
or UO_275 (O_275,N_22382,N_22947);
and UO_276 (O_276,N_21924,N_21850);
nand UO_277 (O_277,N_22384,N_23557);
xor UO_278 (O_278,N_21225,N_22676);
and UO_279 (O_279,N_20490,N_22836);
xor UO_280 (O_280,N_22194,N_20910);
nor UO_281 (O_281,N_21402,N_23373);
nor UO_282 (O_282,N_22756,N_24448);
nand UO_283 (O_283,N_20685,N_22348);
nor UO_284 (O_284,N_20903,N_23930);
nand UO_285 (O_285,N_20659,N_20761);
or UO_286 (O_286,N_23615,N_24150);
and UO_287 (O_287,N_21196,N_21888);
xor UO_288 (O_288,N_20962,N_20520);
xnor UO_289 (O_289,N_21529,N_23132);
or UO_290 (O_290,N_24309,N_23413);
nand UO_291 (O_291,N_24138,N_22763);
and UO_292 (O_292,N_23823,N_21052);
or UO_293 (O_293,N_24485,N_20572);
xnor UO_294 (O_294,N_20745,N_24874);
nand UO_295 (O_295,N_20188,N_24780);
and UO_296 (O_296,N_24898,N_22016);
and UO_297 (O_297,N_24182,N_22417);
or UO_298 (O_298,N_23814,N_24251);
xor UO_299 (O_299,N_23194,N_23795);
nor UO_300 (O_300,N_24564,N_21305);
or UO_301 (O_301,N_22764,N_23575);
or UO_302 (O_302,N_23243,N_23372);
nand UO_303 (O_303,N_22732,N_21194);
or UO_304 (O_304,N_23126,N_22315);
nand UO_305 (O_305,N_22853,N_20099);
nor UO_306 (O_306,N_22047,N_21637);
and UO_307 (O_307,N_20583,N_24140);
or UO_308 (O_308,N_24410,N_24394);
or UO_309 (O_309,N_22145,N_21027);
xnor UO_310 (O_310,N_20515,N_24803);
nand UO_311 (O_311,N_23529,N_23971);
nand UO_312 (O_312,N_20866,N_23551);
and UO_313 (O_313,N_23970,N_23203);
xor UO_314 (O_314,N_22476,N_20506);
or UO_315 (O_315,N_20652,N_22931);
xor UO_316 (O_316,N_23809,N_20845);
nand UO_317 (O_317,N_20673,N_24530);
or UO_318 (O_318,N_23456,N_20469);
and UO_319 (O_319,N_22871,N_21801);
or UO_320 (O_320,N_21962,N_21338);
or UO_321 (O_321,N_21578,N_23827);
nand UO_322 (O_322,N_20019,N_24642);
and UO_323 (O_323,N_23368,N_21119);
nand UO_324 (O_324,N_23573,N_20125);
xor UO_325 (O_325,N_21758,N_23283);
nor UO_326 (O_326,N_22177,N_22723);
nand UO_327 (O_327,N_21262,N_22322);
and UO_328 (O_328,N_24159,N_23593);
nand UO_329 (O_329,N_22962,N_22772);
or UO_330 (O_330,N_21398,N_24879);
xnor UO_331 (O_331,N_23304,N_21979);
and UO_332 (O_332,N_23108,N_20943);
and UO_333 (O_333,N_23352,N_22444);
nor UO_334 (O_334,N_24590,N_20486);
xnor UO_335 (O_335,N_23055,N_24536);
xnor UO_336 (O_336,N_20811,N_21339);
or UO_337 (O_337,N_20231,N_24606);
nor UO_338 (O_338,N_21058,N_23491);
xnor UO_339 (O_339,N_24802,N_21038);
or UO_340 (O_340,N_24609,N_21094);
xnor UO_341 (O_341,N_21820,N_23670);
nor UO_342 (O_342,N_22721,N_22008);
nor UO_343 (O_343,N_21345,N_23948);
nor UO_344 (O_344,N_23478,N_22983);
nor UO_345 (O_345,N_20095,N_23479);
nand UO_346 (O_346,N_24067,N_23746);
nor UO_347 (O_347,N_23453,N_22448);
nor UO_348 (O_348,N_24782,N_20519);
nor UO_349 (O_349,N_24696,N_23897);
xor UO_350 (O_350,N_24243,N_22049);
nor UO_351 (O_351,N_21777,N_22574);
xnor UO_352 (O_352,N_21760,N_21355);
nor UO_353 (O_353,N_20985,N_20782);
and UO_354 (O_354,N_23639,N_23668);
xnor UO_355 (O_355,N_23969,N_21531);
xnor UO_356 (O_356,N_24818,N_22160);
nor UO_357 (O_357,N_21630,N_20828);
or UO_358 (O_358,N_21213,N_22150);
xnor UO_359 (O_359,N_20062,N_22590);
and UO_360 (O_360,N_22545,N_22440);
and UO_361 (O_361,N_24825,N_20077);
nor UO_362 (O_362,N_20251,N_21148);
and UO_363 (O_363,N_24043,N_23310);
xnor UO_364 (O_364,N_23036,N_23031);
nor UO_365 (O_365,N_20131,N_23356);
or UO_366 (O_366,N_23351,N_24768);
xnor UO_367 (O_367,N_23903,N_24241);
xnor UO_368 (O_368,N_22288,N_24951);
and UO_369 (O_369,N_21414,N_22429);
nor UO_370 (O_370,N_22475,N_24262);
and UO_371 (O_371,N_20965,N_20400);
or UO_372 (O_372,N_22790,N_22457);
nand UO_373 (O_373,N_20878,N_22988);
nor UO_374 (O_374,N_22083,N_22058);
xor UO_375 (O_375,N_20827,N_22155);
nand UO_376 (O_376,N_22497,N_22564);
or UO_377 (O_377,N_22467,N_23976);
nor UO_378 (O_378,N_23299,N_24762);
and UO_379 (O_379,N_20319,N_21991);
and UO_380 (O_380,N_24326,N_23916);
and UO_381 (O_381,N_24285,N_20700);
xnor UO_382 (O_382,N_24848,N_23703);
and UO_383 (O_383,N_24881,N_20532);
xnor UO_384 (O_384,N_23062,N_20954);
xnor UO_385 (O_385,N_22553,N_21492);
xor UO_386 (O_386,N_21608,N_23140);
and UO_387 (O_387,N_20883,N_21134);
nand UO_388 (O_388,N_23705,N_23695);
or UO_389 (O_389,N_21557,N_24373);
xor UO_390 (O_390,N_24809,N_21733);
nor UO_391 (O_391,N_23657,N_24124);
nand UO_392 (O_392,N_23601,N_22468);
and UO_393 (O_393,N_22865,N_22426);
nand UO_394 (O_394,N_21383,N_23042);
xor UO_395 (O_395,N_22971,N_22761);
nor UO_396 (O_396,N_22128,N_22986);
or UO_397 (O_397,N_21248,N_22217);
or UO_398 (O_398,N_23629,N_20183);
nor UO_399 (O_399,N_23048,N_20438);
or UO_400 (O_400,N_21035,N_23644);
and UO_401 (O_401,N_22717,N_23996);
xnor UO_402 (O_402,N_24900,N_22463);
and UO_403 (O_403,N_24767,N_22823);
and UO_404 (O_404,N_21112,N_20068);
nand UO_405 (O_405,N_21384,N_24358);
nor UO_406 (O_406,N_23189,N_23388);
xor UO_407 (O_407,N_23192,N_20023);
xor UO_408 (O_408,N_20724,N_21261);
nand UO_409 (O_409,N_20885,N_23961);
xor UO_410 (O_410,N_23177,N_23488);
nand UO_411 (O_411,N_22766,N_24950);
nand UO_412 (O_412,N_23588,N_24025);
xnor UO_413 (O_413,N_20863,N_20250);
xor UO_414 (O_414,N_21829,N_20476);
nand UO_415 (O_415,N_23571,N_22715);
or UO_416 (O_416,N_20735,N_24789);
and UO_417 (O_417,N_22206,N_22597);
and UO_418 (O_418,N_22787,N_24781);
and UO_419 (O_419,N_21836,N_23070);
nand UO_420 (O_420,N_22231,N_23157);
nand UO_421 (O_421,N_23874,N_22267);
xnor UO_422 (O_422,N_23017,N_21958);
and UO_423 (O_423,N_23329,N_21159);
nand UO_424 (O_424,N_20058,N_24697);
or UO_425 (O_425,N_20151,N_24458);
xnor UO_426 (O_426,N_22312,N_24955);
nor UO_427 (O_427,N_23684,N_20314);
nor UO_428 (O_428,N_22978,N_24584);
nor UO_429 (O_429,N_21278,N_24779);
xnor UO_430 (O_430,N_20441,N_23669);
nor UO_431 (O_431,N_21092,N_23475);
nand UO_432 (O_432,N_20838,N_23090);
xnor UO_433 (O_433,N_20021,N_20482);
nor UO_434 (O_434,N_23530,N_23708);
and UO_435 (O_435,N_20130,N_21300);
nor UO_436 (O_436,N_22127,N_22355);
or UO_437 (O_437,N_21010,N_21932);
nand UO_438 (O_438,N_21103,N_22688);
and UO_439 (O_439,N_23198,N_20093);
xnor UO_440 (O_440,N_22616,N_23265);
xnor UO_441 (O_441,N_23483,N_22687);
nand UO_442 (O_442,N_21324,N_20558);
and UO_443 (O_443,N_23893,N_23778);
and UO_444 (O_444,N_20366,N_24703);
xnor UO_445 (O_445,N_22994,N_23665);
nand UO_446 (O_446,N_22953,N_23395);
and UO_447 (O_447,N_21373,N_22742);
nand UO_448 (O_448,N_22064,N_21022);
nor UO_449 (O_449,N_24837,N_23502);
nor UO_450 (O_450,N_20925,N_24096);
xnor UO_451 (O_451,N_20229,N_23141);
and UO_452 (O_452,N_22556,N_22767);
nor UO_453 (O_453,N_22437,N_21950);
nor UO_454 (O_454,N_22854,N_21100);
or UO_455 (O_455,N_23562,N_22548);
and UO_456 (O_456,N_23921,N_20383);
nand UO_457 (O_457,N_24819,N_24540);
and UO_458 (O_458,N_23414,N_22234);
or UO_459 (O_459,N_20003,N_21804);
nor UO_460 (O_460,N_20048,N_22136);
xor UO_461 (O_461,N_21964,N_21896);
xor UO_462 (O_462,N_24995,N_21788);
nor UO_463 (O_463,N_24992,N_20424);
nand UO_464 (O_464,N_21216,N_24930);
nor UO_465 (O_465,N_20785,N_22925);
nor UO_466 (O_466,N_22863,N_22375);
nand UO_467 (O_467,N_21600,N_23065);
and UO_468 (O_468,N_22406,N_21007);
nor UO_469 (O_469,N_23187,N_22850);
nor UO_470 (O_470,N_23438,N_20405);
nand UO_471 (O_471,N_22970,N_23980);
or UO_472 (O_472,N_21416,N_21200);
xnor UO_473 (O_473,N_20101,N_24601);
xnor UO_474 (O_474,N_24304,N_22284);
xnor UO_475 (O_475,N_20897,N_21215);
and UO_476 (O_476,N_21743,N_22812);
xor UO_477 (O_477,N_21246,N_20258);
or UO_478 (O_478,N_22249,N_23998);
xor UO_479 (O_479,N_20990,N_23273);
nand UO_480 (O_480,N_22634,N_21625);
or UO_481 (O_481,N_20475,N_24734);
xnor UO_482 (O_482,N_24597,N_21811);
and UO_483 (O_483,N_22706,N_21222);
xnor UO_484 (O_484,N_22210,N_23268);
nand UO_485 (O_485,N_22039,N_24602);
nor UO_486 (O_486,N_20270,N_24252);
xor UO_487 (O_487,N_21417,N_24817);
xor UO_488 (O_488,N_20387,N_21555);
nor UO_489 (O_489,N_23344,N_20290);
nor UO_490 (O_490,N_22835,N_21821);
or UO_491 (O_491,N_20220,N_20810);
nor UO_492 (O_492,N_24533,N_20886);
xor UO_493 (O_493,N_23607,N_20268);
nor UO_494 (O_494,N_21097,N_22946);
nand UO_495 (O_495,N_20808,N_24632);
nand UO_496 (O_496,N_23570,N_20703);
nand UO_497 (O_497,N_20609,N_20315);
nand UO_498 (O_498,N_22180,N_21565);
or UO_499 (O_499,N_21538,N_20781);
nand UO_500 (O_500,N_22498,N_24297);
or UO_501 (O_501,N_23899,N_20322);
and UO_502 (O_502,N_21372,N_20676);
nand UO_503 (O_503,N_22829,N_23333);
or UO_504 (O_504,N_21426,N_21746);
and UO_505 (O_505,N_23812,N_20171);
and UO_506 (O_506,N_20514,N_21672);
and UO_507 (O_507,N_24403,N_22998);
nand UO_508 (O_508,N_21435,N_23472);
or UO_509 (O_509,N_24445,N_24468);
xnor UO_510 (O_510,N_22811,N_22474);
xor UO_511 (O_511,N_24655,N_23555);
nor UO_512 (O_512,N_24798,N_22198);
or UO_513 (O_513,N_20566,N_24421);
nor UO_514 (O_514,N_22555,N_24232);
or UO_515 (O_515,N_20739,N_21361);
nor UO_516 (O_516,N_22402,N_20877);
or UO_517 (O_517,N_22505,N_22930);
or UO_518 (O_518,N_20667,N_22066);
xor UO_519 (O_519,N_23086,N_22737);
and UO_520 (O_520,N_21951,N_23663);
xnor UO_521 (O_521,N_22985,N_20859);
or UO_522 (O_522,N_22557,N_24587);
nor UO_523 (O_523,N_23064,N_22539);
and UO_524 (O_524,N_22302,N_23366);
nor UO_525 (O_525,N_22815,N_22649);
and UO_526 (O_526,N_20959,N_24511);
nand UO_527 (O_527,N_20677,N_24996);
nor UO_528 (O_528,N_24611,N_24933);
and UO_529 (O_529,N_22456,N_23526);
nor UO_530 (O_530,N_20411,N_20347);
nor UO_531 (O_531,N_21747,N_20004);
nand UO_532 (O_532,N_23525,N_21678);
and UO_533 (O_533,N_21893,N_21930);
or UO_534 (O_534,N_24718,N_23410);
xor UO_535 (O_535,N_20436,N_24545);
nor UO_536 (O_536,N_20927,N_20035);
or UO_537 (O_537,N_23463,N_20005);
xor UO_538 (O_538,N_21726,N_20479);
or UO_539 (O_539,N_21342,N_24688);
nor UO_540 (O_540,N_22226,N_21729);
or UO_541 (O_541,N_21876,N_20307);
and UO_542 (O_542,N_23280,N_21670);
xor UO_543 (O_543,N_23470,N_21532);
nor UO_544 (O_544,N_20850,N_24156);
or UO_545 (O_545,N_20891,N_21385);
or UO_546 (O_546,N_24727,N_23707);
or UO_547 (O_547,N_21150,N_20712);
and UO_548 (O_548,N_20435,N_21655);
nor UO_549 (O_549,N_21784,N_20936);
nor UO_550 (O_550,N_21168,N_20671);
or UO_551 (O_551,N_22446,N_21303);
nand UO_552 (O_552,N_23267,N_21899);
nor UO_553 (O_553,N_22798,N_23246);
xor UO_554 (O_554,N_22496,N_24671);
nand UO_555 (O_555,N_23768,N_21304);
or UO_556 (O_556,N_24901,N_20976);
nand UO_557 (O_557,N_24200,N_24694);
xor UO_558 (O_558,N_23690,N_23420);
and UO_559 (O_559,N_21560,N_23087);
or UO_560 (O_560,N_21673,N_23425);
nor UO_561 (O_561,N_24491,N_23860);
and UO_562 (O_562,N_20008,N_23868);
nand UO_563 (O_563,N_24432,N_22845);
nand UO_564 (O_564,N_20273,N_23335);
and UO_565 (O_565,N_23650,N_20626);
nor UO_566 (O_566,N_21067,N_22753);
nor UO_567 (O_567,N_22576,N_24896);
nand UO_568 (O_568,N_21685,N_20971);
nand UO_569 (O_569,N_20094,N_24375);
xnor UO_570 (O_570,N_21697,N_22795);
nand UO_571 (O_571,N_24083,N_24656);
nand UO_572 (O_572,N_24801,N_23852);
nand UO_573 (O_573,N_22011,N_21043);
nor UO_574 (O_574,N_20037,N_23061);
xnor UO_575 (O_575,N_22967,N_22793);
nand UO_576 (O_576,N_22154,N_21274);
nor UO_577 (O_577,N_22698,N_23749);
and UO_578 (O_578,N_23726,N_23094);
xnor UO_579 (O_579,N_20177,N_20534);
nand UO_580 (O_580,N_24137,N_21705);
or UO_581 (O_581,N_22816,N_23568);
nand UO_582 (O_582,N_24902,N_20854);
nand UO_583 (O_583,N_24331,N_22004);
and UO_584 (O_584,N_22625,N_23229);
nor UO_585 (O_585,N_24006,N_23480);
xor UO_586 (O_586,N_22886,N_21552);
xor UO_587 (O_587,N_23465,N_24161);
nand UO_588 (O_588,N_22524,N_21773);
nand UO_589 (O_589,N_24750,N_22328);
nand UO_590 (O_590,N_24229,N_22952);
and UO_591 (O_591,N_20447,N_21605);
or UO_592 (O_592,N_24005,N_21898);
and UO_593 (O_593,N_22861,N_23710);
nand UO_594 (O_594,N_21015,N_21264);
nor UO_595 (O_595,N_24876,N_21290);
nor UO_596 (O_596,N_24686,N_23924);
xor UO_597 (O_597,N_24164,N_23349);
or UO_598 (O_598,N_21090,N_24360);
nand UO_599 (O_599,N_23848,N_22293);
nand UO_600 (O_600,N_22602,N_22566);
xor UO_601 (O_601,N_20339,N_21617);
nor UO_602 (O_602,N_22511,N_22776);
nand UO_603 (O_603,N_24162,N_21704);
xnor UO_604 (O_604,N_20849,N_23581);
nor UO_605 (O_605,N_24344,N_20083);
and UO_606 (O_606,N_20873,N_24764);
xor UO_607 (O_607,N_23125,N_22350);
or UO_608 (O_608,N_20502,N_22063);
nand UO_609 (O_609,N_23564,N_23608);
nand UO_610 (O_610,N_23963,N_21756);
nand UO_611 (O_611,N_20611,N_24054);
nor UO_612 (O_612,N_20535,N_23817);
xor UO_613 (O_613,N_20210,N_22099);
xnor UO_614 (O_614,N_21307,N_22300);
nor UO_615 (O_615,N_23341,N_21268);
or UO_616 (O_616,N_24532,N_20297);
and UO_617 (O_617,N_20768,N_20788);
xor UO_618 (O_618,N_21436,N_23442);
and UO_619 (O_619,N_24744,N_20323);
nor UO_620 (O_620,N_21620,N_23789);
and UO_621 (O_621,N_24291,N_20618);
xnor UO_622 (O_622,N_24512,N_24266);
and UO_623 (O_623,N_21457,N_21044);
nand UO_624 (O_624,N_23941,N_22026);
or UO_625 (O_625,N_22255,N_23621);
nand UO_626 (O_626,N_23220,N_20991);
xnor UO_627 (O_627,N_21653,N_23599);
or UO_628 (O_628,N_21281,N_23328);
nand UO_629 (O_629,N_24446,N_24157);
or UO_630 (O_630,N_20716,N_24171);
and UO_631 (O_631,N_20857,N_20656);
and UO_632 (O_632,N_22218,N_21330);
and UO_633 (O_633,N_22584,N_21875);
nand UO_634 (O_634,N_21149,N_21567);
or UO_635 (O_635,N_22415,N_24498);
or UO_636 (O_636,N_20324,N_22465);
nand UO_637 (O_637,N_22297,N_20395);
or UO_638 (O_638,N_21093,N_24790);
nor UO_639 (O_639,N_24684,N_22730);
nor UO_640 (O_640,N_20726,N_24770);
xor UO_641 (O_641,N_24061,N_20462);
nand UO_642 (O_642,N_21279,N_22250);
xnor UO_643 (O_643,N_24244,N_22518);
xor UO_644 (O_644,N_21412,N_24795);
and UO_645 (O_645,N_23647,N_24233);
nor UO_646 (O_646,N_20536,N_22059);
nand UO_647 (O_647,N_24228,N_20528);
nand UO_648 (O_648,N_20381,N_22101);
or UO_649 (O_649,N_20028,N_21357);
or UO_650 (O_650,N_23544,N_23208);
and UO_651 (O_651,N_23306,N_23870);
nand UO_652 (O_652,N_21155,N_21810);
and UO_653 (O_653,N_21634,N_24289);
nor UO_654 (O_654,N_20608,N_21135);
nand UO_655 (O_655,N_21364,N_24717);
nor UO_656 (O_656,N_24505,N_22540);
nand UO_657 (O_657,N_20425,N_21291);
nor UO_658 (O_658,N_20373,N_22907);
or UO_659 (O_659,N_22822,N_20918);
and UO_660 (O_660,N_23774,N_21452);
nand UO_661 (O_661,N_21586,N_23127);
xor UO_662 (O_662,N_23974,N_24982);
xnor UO_663 (O_663,N_22725,N_24100);
and UO_664 (O_664,N_21245,N_23999);
nor UO_665 (O_665,N_24965,N_20997);
xor UO_666 (O_666,N_24227,N_24793);
nand UO_667 (O_667,N_24293,N_21737);
and UO_668 (O_668,N_23128,N_22151);
and UO_669 (O_669,N_22014,N_21444);
nor UO_670 (O_670,N_22027,N_21014);
nor UO_671 (O_671,N_23252,N_20822);
or UO_672 (O_672,N_20634,N_22919);
nand UO_673 (O_673,N_23350,N_22718);
xor UO_674 (O_674,N_24763,N_24724);
nor UO_675 (O_675,N_21161,N_20731);
and UO_676 (O_676,N_22991,N_23728);
nand UO_677 (O_677,N_22362,N_24135);
xnor UO_678 (O_678,N_24807,N_20283);
nand UO_679 (O_679,N_21381,N_20252);
xnor UO_680 (O_680,N_22133,N_24612);
or UO_681 (O_681,N_20214,N_20617);
and UO_682 (O_682,N_20970,N_23983);
nand UO_683 (O_683,N_22298,N_22633);
nor UO_684 (O_684,N_21719,N_23592);
nand UO_685 (O_685,N_24404,N_21809);
and UO_686 (O_686,N_23416,N_20630);
nor UO_687 (O_687,N_20417,N_24917);
or UO_688 (O_688,N_23846,N_24757);
nor UO_689 (O_689,N_21853,N_21419);
nor UO_690 (O_690,N_23748,N_22961);
and UO_691 (O_691,N_22401,N_22510);
and UO_692 (O_692,N_23956,N_20504);
nor UO_693 (O_693,N_22281,N_23182);
or UO_694 (O_694,N_20079,N_20813);
or UO_695 (O_695,N_24211,N_21576);
and UO_696 (O_696,N_20527,N_20146);
xnor UO_697 (O_697,N_24496,N_24558);
xnor UO_698 (O_698,N_21360,N_21794);
or UO_699 (O_699,N_21791,N_21325);
and UO_700 (O_700,N_20362,N_21877);
nand UO_701 (O_701,N_22431,N_24944);
or UO_702 (O_702,N_22671,N_20686);
nor UO_703 (O_703,N_23582,N_20957);
and UO_704 (O_704,N_24897,N_24402);
xnor UO_705 (O_705,N_23392,N_20279);
nor UO_706 (O_706,N_22944,N_21669);
nor UO_707 (O_707,N_21478,N_24295);
nor UO_708 (O_708,N_20593,N_21250);
or UO_709 (O_709,N_24507,N_20227);
xor UO_710 (O_710,N_23018,N_20795);
and UO_711 (O_711,N_20073,N_23231);
or UO_712 (O_712,N_22263,N_20075);
nor UO_713 (O_713,N_21842,N_22879);
nand UO_714 (O_714,N_24019,N_23911);
and UO_715 (O_715,N_21008,N_23739);
and UO_716 (O_716,N_21827,N_24659);
and UO_717 (O_717,N_22541,N_23053);
or UO_718 (O_718,N_24346,N_20915);
or UO_719 (O_719,N_20987,N_24388);
nor UO_720 (O_720,N_20596,N_24573);
or UO_721 (O_721,N_23020,N_20926);
or UO_722 (O_722,N_21054,N_20642);
or UO_723 (O_723,N_21387,N_21284);
xor UO_724 (O_724,N_22323,N_23207);
xor UO_725 (O_725,N_22044,N_20158);
or UO_726 (O_726,N_24218,N_23422);
or UO_727 (O_727,N_20114,N_24797);
xnor UO_728 (O_728,N_24500,N_20969);
nor UO_729 (O_729,N_23060,N_23158);
nor UO_730 (O_730,N_21450,N_20861);
nand UO_731 (O_731,N_21182,N_24450);
nor UO_732 (O_732,N_20675,N_24339);
nor UO_733 (O_733,N_22549,N_23330);
xor UO_734 (O_734,N_20803,N_23136);
nor UO_735 (O_735,N_24437,N_22820);
nand UO_736 (O_736,N_24390,N_21752);
xnor UO_737 (O_737,N_21590,N_22642);
and UO_738 (O_738,N_20964,N_20371);
nor UO_739 (O_739,N_21490,N_23382);
xor UO_740 (O_740,N_22205,N_21612);
nor UO_741 (O_741,N_24000,N_23513);
and UO_742 (O_742,N_22022,N_20751);
and UO_743 (O_743,N_22980,N_24756);
nor UO_744 (O_744,N_20107,N_23174);
and UO_745 (O_745,N_21496,N_24365);
or UO_746 (O_746,N_24743,N_20407);
xnor UO_747 (O_747,N_21486,N_20033);
or UO_748 (O_748,N_22001,N_24416);
and UO_749 (O_749,N_23212,N_21587);
and UO_750 (O_750,N_22754,N_23990);
nor UO_751 (O_751,N_20329,N_21517);
xor UO_752 (O_752,N_22079,N_24882);
nand UO_753 (O_753,N_22073,N_22933);
and UO_754 (O_754,N_20563,N_21401);
or UO_755 (O_755,N_20382,N_21833);
xor UO_756 (O_756,N_23439,N_23673);
or UO_757 (O_757,N_21331,N_24090);
nor UO_758 (O_758,N_22242,N_23193);
nand UO_759 (O_759,N_20598,N_21346);
nand UO_760 (O_760,N_20380,N_23927);
xor UO_761 (O_761,N_23239,N_21781);
or UO_762 (O_762,N_21807,N_23522);
nand UO_763 (O_763,N_24323,N_20050);
nand UO_764 (O_764,N_21754,N_20355);
nor UO_765 (O_765,N_24497,N_20820);
and UO_766 (O_766,N_24106,N_23078);
nand UO_767 (O_767,N_20239,N_24181);
or UO_768 (O_768,N_20194,N_22489);
or UO_769 (O_769,N_20951,N_20046);
and UO_770 (O_770,N_20249,N_23200);
or UO_771 (O_771,N_22447,N_22430);
nor UO_772 (O_772,N_24101,N_24351);
or UO_773 (O_773,N_24264,N_21389);
nand UO_774 (O_774,N_22021,N_24548);
xor UO_775 (O_775,N_20662,N_21867);
nor UO_776 (O_776,N_20829,N_20544);
and UO_777 (O_777,N_22170,N_23950);
xor UO_778 (O_778,N_21241,N_22680);
and UO_779 (O_779,N_21386,N_24538);
xnor UO_780 (O_780,N_21539,N_21849);
and UO_781 (O_781,N_23842,N_24325);
nor UO_782 (O_782,N_21371,N_22888);
nor UO_783 (O_783,N_21471,N_22172);
xor UO_784 (O_784,N_21218,N_20378);
and UO_785 (O_785,N_23622,N_22724);
nand UO_786 (O_786,N_21166,N_24192);
and UO_787 (O_787,N_22959,N_20872);
nor UO_788 (O_788,N_21614,N_24525);
and UO_789 (O_789,N_22261,N_20496);
nor UO_790 (O_790,N_23181,N_20133);
nor UO_791 (O_791,N_23348,N_24681);
xor UO_792 (O_792,N_20826,N_24041);
and UO_793 (O_793,N_24516,N_21648);
nand UO_794 (O_794,N_21516,N_21739);
or UO_795 (O_795,N_21929,N_21317);
xnor UO_796 (O_796,N_23218,N_24431);
or UO_797 (O_797,N_20484,N_22351);
or UO_798 (O_798,N_21716,N_22762);
and UO_799 (O_799,N_20771,N_23213);
nor UO_800 (O_800,N_20196,N_21584);
xnor UO_801 (O_801,N_23054,N_23679);
and UO_802 (O_802,N_22592,N_21179);
nand UO_803 (O_803,N_22618,N_24283);
nor UO_804 (O_804,N_20763,N_22982);
nor UO_805 (O_805,N_22965,N_23454);
nand UO_806 (O_806,N_21881,N_21356);
xor UO_807 (O_807,N_23202,N_24604);
and UO_808 (O_808,N_24751,N_22975);
or UO_809 (O_809,N_20000,N_23548);
nor UO_810 (O_810,N_23933,N_20904);
nand UO_811 (O_811,N_21713,N_22948);
or UO_812 (O_812,N_24337,N_24306);
xor UO_813 (O_813,N_20390,N_22308);
nand UO_814 (O_814,N_21332,N_21017);
nand UO_815 (O_815,N_24175,N_20326);
and UO_816 (O_816,N_22466,N_22361);
and UO_817 (O_817,N_22700,N_21397);
xnor UO_818 (O_818,N_22069,N_22353);
and UO_819 (O_819,N_21959,N_21140);
xnor UO_820 (O_820,N_22626,N_20198);
nor UO_821 (O_821,N_21506,N_20426);
nand UO_822 (O_822,N_24363,N_23408);
and UO_823 (O_823,N_24769,N_23736);
nor UO_824 (O_824,N_20346,N_20472);
nand UO_825 (O_825,N_22654,N_23426);
nor UO_826 (O_826,N_24993,N_24143);
and UO_827 (O_827,N_22538,N_20391);
or UO_828 (O_828,N_24599,N_22273);
or UO_829 (O_829,N_23833,N_22520);
nor UO_830 (O_830,N_20856,N_23804);
nand UO_831 (O_831,N_24256,N_24465);
xnor UO_832 (O_832,N_24370,N_24664);
xnor UO_833 (O_833,N_24760,N_22523);
nand UO_834 (O_834,N_21728,N_22089);
and UO_835 (O_835,N_21585,N_24438);
and UO_836 (O_836,N_20167,N_23985);
nand UO_837 (O_837,N_24931,N_24909);
nand UO_838 (O_838,N_21458,N_21065);
xnor UO_839 (O_839,N_22235,N_20575);
nand UO_840 (O_840,N_20621,N_21234);
nand UO_841 (O_841,N_23626,N_21089);
or UO_842 (O_842,N_24044,N_20692);
nand UO_843 (O_843,N_22873,N_22818);
and UO_844 (O_844,N_23583,N_22072);
or UO_845 (O_845,N_20350,N_20452);
xnor UO_846 (O_846,N_20152,N_23702);
nand UO_847 (O_847,N_24372,N_22107);
and UO_848 (O_848,N_23074,N_24315);
xnor UO_849 (O_849,N_22528,N_23688);
or UO_850 (O_850,N_20738,N_21025);
xnor UO_851 (O_851,N_20137,N_24541);
or UO_852 (O_852,N_24842,N_20843);
xor UO_853 (O_853,N_21353,N_24434);
nand UO_854 (O_854,N_22964,N_24473);
nand UO_855 (O_855,N_24420,N_20999);
and UO_856 (O_856,N_23534,N_21961);
or UO_857 (O_857,N_20465,N_20942);
nand UO_858 (O_858,N_23045,N_24254);
nor UO_859 (O_859,N_22477,N_20545);
and UO_860 (O_860,N_20967,N_23940);
nand UO_861 (O_861,N_24634,N_20715);
nand UO_862 (O_862,N_24475,N_24060);
nand UO_863 (O_863,N_21575,N_23233);
and UO_864 (O_864,N_22106,N_24307);
and UO_865 (O_865,N_20332,N_23430);
xor UO_866 (O_866,N_24336,N_20234);
nor UO_867 (O_867,N_24223,N_22569);
and UO_868 (O_868,N_24575,N_23097);
and UO_869 (O_869,N_23450,N_23151);
xor UO_870 (O_870,N_21524,N_20481);
and UO_871 (O_871,N_20793,N_24868);
and UO_872 (O_872,N_21911,N_24924);
nor UO_873 (O_873,N_21736,N_22543);
xnor UO_874 (O_874,N_23360,N_22111);
xor UO_875 (O_875,N_21533,N_20587);
or UO_876 (O_876,N_23953,N_24991);
nand UO_877 (O_877,N_20736,N_22552);
nor UO_878 (O_878,N_21118,N_24593);
nand UO_879 (O_879,N_21993,N_21453);
and UO_880 (O_880,N_20636,N_21862);
or UO_881 (O_881,N_20492,N_24971);
or UO_882 (O_882,N_20995,N_21690);
and UO_883 (O_883,N_23757,N_24816);
xnor UO_884 (O_884,N_24570,N_23550);
or UO_885 (O_885,N_24562,N_22751);
xnor UO_886 (O_886,N_22387,N_24730);
or UO_887 (O_887,N_22410,N_24890);
nand UO_888 (O_888,N_22439,N_23498);
and UO_889 (O_889,N_23038,N_22579);
nor UO_890 (O_890,N_23991,N_20695);
and UO_891 (O_891,N_24249,N_21658);
nor UO_892 (O_892,N_20236,N_24341);
nor UO_893 (O_893,N_20613,N_20743);
or UO_894 (O_894,N_20674,N_20045);
nand UO_895 (O_895,N_23609,N_23909);
or UO_896 (O_896,N_24385,N_20902);
and UO_897 (O_897,N_22438,N_20086);
xnor UO_898 (O_898,N_21086,N_23967);
and UO_899 (O_899,N_24721,N_23816);
or UO_900 (O_900,N_22697,N_21593);
nand UO_901 (O_901,N_20010,N_22159);
nand UO_902 (O_902,N_21042,N_20143);
xnor UO_903 (O_903,N_21983,N_21068);
nand UO_904 (O_904,N_21706,N_21424);
nand UO_905 (O_905,N_24011,N_23545);
xor UO_906 (O_906,N_24494,N_23190);
and UO_907 (O_907,N_20780,N_24221);
or UO_908 (O_908,N_23375,N_23843);
or UO_909 (O_909,N_24338,N_20092);
xnor UO_910 (O_910,N_22222,N_21597);
nor UO_911 (O_911,N_21313,N_23877);
nor UO_912 (O_912,N_22773,N_21466);
or UO_913 (O_913,N_23913,N_24911);
nor UO_914 (O_914,N_23602,N_22635);
nand UO_915 (O_915,N_20218,N_22615);
and UO_916 (O_916,N_24371,N_22755);
nor UO_917 (O_917,N_21079,N_24270);
or UO_918 (O_918,N_20599,N_22313);
and UO_919 (O_919,N_21839,N_20334);
xnor UO_920 (O_920,N_20518,N_24074);
xor UO_921 (O_921,N_22416,N_20832);
or UO_922 (O_922,N_24735,N_22973);
and UO_923 (O_923,N_20672,N_22020);
or UO_924 (O_924,N_20263,N_23659);
or UO_925 (O_925,N_24334,N_21271);
xnor UO_926 (O_926,N_24518,N_21859);
nand UO_927 (O_927,N_24578,N_24905);
or UO_928 (O_928,N_21680,N_20860);
or UO_929 (O_929,N_20154,N_22241);
or UO_930 (O_930,N_21914,N_24832);
and UO_931 (O_931,N_24231,N_21500);
nor UO_932 (O_932,N_22636,N_24423);
and UO_933 (O_933,N_22420,N_22922);
and UO_934 (O_934,N_21460,N_21178);
nor UO_935 (O_935,N_20888,N_22452);
xnor UO_936 (O_936,N_20280,N_23835);
or UO_937 (O_937,N_20982,N_22503);
and UO_938 (O_938,N_23027,N_22117);
nor UO_939 (O_939,N_23093,N_23701);
nor UO_940 (O_940,N_23397,N_24369);
and UO_941 (O_941,N_23784,N_20591);
or UO_942 (O_942,N_22645,N_23964);
and UO_943 (O_943,N_23156,N_24176);
or UO_944 (O_944,N_24726,N_20653);
xnor UO_945 (O_945,N_24045,N_22674);
nand UO_946 (O_946,N_20645,N_24170);
xor UO_947 (O_947,N_21341,N_22280);
nand UO_948 (O_948,N_24426,N_21519);
or UO_949 (O_949,N_23481,N_21799);
or UO_950 (O_950,N_24566,N_22662);
or UO_951 (O_951,N_20203,N_20631);
xor UO_952 (O_952,N_23885,N_21938);
or UO_953 (O_953,N_22619,N_22168);
xor UO_954 (O_954,N_23616,N_23878);
nand UO_955 (O_955,N_22148,N_24186);
xor UO_956 (O_956,N_22071,N_21798);
nand UO_957 (O_957,N_24455,N_20647);
nand UO_958 (O_958,N_22734,N_21639);
or UO_959 (O_959,N_21974,N_23477);
or UO_960 (O_960,N_24567,N_23217);
or UO_961 (O_961,N_22669,N_21512);
or UO_962 (O_962,N_24672,N_24313);
nor UO_963 (O_963,N_21660,N_22051);
and UO_964 (O_964,N_24537,N_20980);
nand UO_965 (O_965,N_21484,N_23300);
xor UO_966 (O_966,N_22391,N_20372);
and UO_967 (O_967,N_20670,N_21104);
nor UO_968 (O_968,N_21668,N_21223);
xor UO_969 (O_969,N_23296,N_23718);
or UO_970 (O_970,N_24749,N_22803);
and UO_971 (O_971,N_23751,N_20389);
or UO_972 (O_972,N_20116,N_20026);
or UO_973 (O_973,N_22495,N_23486);
xor UO_974 (O_974,N_22274,N_24887);
nand UO_975 (O_975,N_21208,N_21488);
or UO_976 (O_976,N_20477,N_21408);
nor UO_977 (O_977,N_23618,N_22702);
nor UO_978 (O_978,N_24099,N_22893);
nor UO_979 (O_979,N_24638,N_23787);
and UO_980 (O_980,N_23109,N_23433);
nor UO_981 (O_981,N_21076,N_22957);
nor UO_982 (O_982,N_23464,N_23317);
nand UO_983 (O_983,N_22679,N_24520);
and UO_984 (O_984,N_22190,N_23289);
nand UO_985 (O_985,N_23858,N_22536);
xnor UO_986 (O_986,N_24430,N_20039);
or UO_987 (O_987,N_23807,N_21308);
nor UO_988 (O_988,N_21254,N_22668);
nand UO_989 (O_989,N_21891,N_21869);
or UO_990 (O_990,N_23423,N_21767);
nor UO_991 (O_991,N_20691,N_21431);
or UO_992 (O_992,N_24618,N_21283);
nand UO_993 (O_993,N_23693,N_23291);
or UO_994 (O_994,N_23404,N_20247);
and UO_995 (O_995,N_21206,N_24319);
or UO_996 (O_996,N_22195,N_24920);
xnor UO_997 (O_997,N_21311,N_23347);
nand UO_998 (O_998,N_20704,N_21465);
nand UO_999 (O_999,N_21095,N_21618);
xor UO_1000 (O_1000,N_23648,N_21497);
xnor UO_1001 (O_1001,N_24869,N_24937);
xor UO_1002 (O_1002,N_22121,N_22450);
nor UO_1003 (O_1003,N_22997,N_20409);
and UO_1004 (O_1004,N_24737,N_23678);
xnor UO_1005 (O_1005,N_23642,N_23484);
nor UO_1006 (O_1006,N_22740,N_22769);
nor UO_1007 (O_1007,N_20551,N_24652);
xnor UO_1008 (O_1008,N_22757,N_22364);
nand UO_1009 (O_1009,N_23037,N_20560);
xnor UO_1010 (O_1010,N_21731,N_20088);
or UO_1011 (O_1011,N_23362,N_21288);
xnor UO_1012 (O_1012,N_21769,N_24079);
nor UO_1013 (O_1013,N_21320,N_20846);
or UO_1014 (O_1014,N_21778,N_24858);
and UO_1015 (O_1015,N_24872,N_21201);
xor UO_1016 (O_1016,N_23994,N_22157);
xnor UO_1017 (O_1017,N_22872,N_22587);
and UO_1018 (O_1018,N_23251,N_24502);
xnor UO_1019 (O_1019,N_24258,N_20934);
nand UO_1020 (O_1020,N_22214,N_22714);
and UO_1021 (O_1021,N_20192,N_23596);
xnor UO_1022 (O_1022,N_23142,N_23387);
nand UO_1023 (O_1023,N_20109,N_20179);
nand UO_1024 (O_1024,N_23449,N_23361);
xnor UO_1025 (O_1025,N_24049,N_23606);
or UO_1026 (O_1026,N_20538,N_21430);
or UO_1027 (O_1027,N_23441,N_20620);
nand UO_1028 (O_1028,N_24773,N_22533);
and UO_1029 (O_1029,N_21032,N_24683);
xnor UO_1030 (O_1030,N_22048,N_20396);
nor UO_1031 (O_1031,N_24383,N_22085);
or UO_1032 (O_1032,N_24739,N_24867);
and UO_1033 (O_1033,N_20302,N_21677);
and UO_1034 (O_1034,N_21391,N_22943);
and UO_1035 (O_1035,N_22183,N_23888);
or UO_1036 (O_1036,N_23400,N_23013);
or UO_1037 (O_1037,N_20984,N_21789);
or UO_1038 (O_1038,N_24693,N_24002);
nor UO_1039 (O_1039,N_22356,N_21354);
nand UO_1040 (O_1040,N_20090,N_20629);
and UO_1041 (O_1041,N_24418,N_20036);
and UO_1042 (O_1042,N_24921,N_23129);
and UO_1043 (O_1043,N_21459,N_20531);
nand UO_1044 (O_1044,N_20014,N_21667);
xor UO_1045 (O_1045,N_21404,N_20267);
xnor UO_1046 (O_1046,N_24489,N_22729);
or UO_1047 (O_1047,N_23741,N_20365);
nor UO_1048 (O_1048,N_22254,N_22403);
nor UO_1049 (O_1049,N_22229,N_24526);
xnor UO_1050 (O_1050,N_24424,N_20466);
or UO_1051 (O_1051,N_23894,N_21536);
and UO_1052 (O_1052,N_22377,N_20293);
or UO_1053 (O_1053,N_20649,N_20084);
and UO_1054 (O_1054,N_22149,N_20392);
and UO_1055 (O_1055,N_24082,N_20660);
and UO_1056 (O_1056,N_21170,N_22651);
nor UO_1057 (O_1057,N_22208,N_23543);
and UO_1058 (O_1058,N_20895,N_20972);
xor UO_1059 (O_1059,N_24442,N_23210);
nand UO_1060 (O_1060,N_21772,N_20986);
nor UO_1061 (O_1061,N_20162,N_20698);
xnor UO_1062 (O_1062,N_20728,N_21561);
nand UO_1063 (O_1063,N_22023,N_22213);
nand UO_1064 (O_1064,N_21905,N_24406);
xor UO_1065 (O_1065,N_24778,N_23049);
nor UO_1066 (O_1066,N_21476,N_23307);
nor UO_1067 (O_1067,N_23563,N_20687);
nand UO_1068 (O_1068,N_21569,N_21378);
xor UO_1069 (O_1069,N_23069,N_21405);
or UO_1070 (O_1070,N_24427,N_23516);
nand UO_1071 (O_1071,N_23989,N_24127);
and UO_1072 (O_1072,N_22535,N_21870);
and UO_1073 (O_1073,N_21513,N_22781);
nor UO_1074 (O_1074,N_23469,N_22207);
xor UO_1075 (O_1075,N_24715,N_24748);
and UO_1076 (O_1076,N_24310,N_22252);
nor UO_1077 (O_1077,N_21563,N_21233);
nor UO_1078 (O_1078,N_23691,N_23238);
xor UO_1079 (O_1079,N_22846,N_22722);
nor UO_1080 (O_1080,N_21868,N_21826);
xnor UO_1081 (O_1081,N_21358,N_24701);
nor UO_1082 (O_1082,N_20953,N_23390);
xor UO_1083 (O_1083,N_20556,N_23171);
or UO_1084 (O_1084,N_20442,N_20690);
nand UO_1085 (O_1085,N_24980,N_22102);
or UO_1086 (O_1086,N_20057,N_21708);
or UO_1087 (O_1087,N_24412,N_21635);
and UO_1088 (O_1088,N_21129,N_21334);
and UO_1089 (O_1089,N_23753,N_23685);
xor UO_1090 (O_1090,N_24919,N_21400);
or UO_1091 (O_1091,N_21001,N_24003);
and UO_1092 (O_1092,N_21702,N_20817);
or UO_1093 (O_1093,N_21551,N_24853);
and UO_1094 (O_1094,N_22650,N_21193);
xnor UO_1095 (O_1095,N_24048,N_23118);
or UO_1096 (O_1096,N_23837,N_20301);
nand UO_1097 (O_1097,N_21146,N_21966);
xnor UO_1098 (O_1098,N_22824,N_21858);
or UO_1099 (O_1099,N_22259,N_24217);
nand UO_1100 (O_1100,N_24187,N_22777);
nor UO_1101 (O_1101,N_20721,N_24959);
nand UO_1102 (O_1102,N_20110,N_20081);
nand UO_1103 (O_1103,N_23415,N_21101);
nor UO_1104 (O_1104,N_22792,N_20729);
nand UO_1105 (O_1105,N_24443,N_23286);
and UO_1106 (O_1106,N_24990,N_20549);
nand UO_1107 (O_1107,N_20922,N_22581);
nor UO_1108 (O_1108,N_21831,N_23747);
nor UO_1109 (O_1109,N_24409,N_23088);
nor UO_1110 (O_1110,N_24472,N_23455);
nor UO_1111 (O_1111,N_21892,N_20607);
and UO_1112 (O_1112,N_22563,N_20443);
and UO_1113 (O_1113,N_23199,N_20106);
nand UO_1114 (O_1114,N_24707,N_22211);
and UO_1115 (O_1115,N_21120,N_20144);
xor UO_1116 (O_1116,N_23358,N_20388);
nor UO_1117 (O_1117,N_21380,N_21815);
nor UO_1118 (O_1118,N_22577,N_22345);
xnor UO_1119 (O_1119,N_22749,N_24752);
or UO_1120 (O_1120,N_22042,N_24772);
or UO_1121 (O_1121,N_20663,N_20932);
or UO_1122 (O_1122,N_22665,N_23292);
nand UO_1123 (O_1123,N_22464,N_22483);
nor UO_1124 (O_1124,N_20148,N_22041);
nand UO_1125 (O_1125,N_22197,N_23613);
and UO_1126 (O_1126,N_21636,N_23612);
nor UO_1127 (O_1127,N_22478,N_22909);
nor UO_1128 (O_1128,N_20744,N_24877);
nand UO_1129 (O_1129,N_21683,N_23245);
and UO_1130 (O_1130,N_23857,N_21272);
nand UO_1131 (O_1131,N_24399,N_23440);
nor UO_1132 (O_1132,N_21641,N_23111);
xnor UO_1133 (O_1133,N_21472,N_23476);
or UO_1134 (O_1134,N_23898,N_20567);
nor UO_1135 (O_1135,N_20440,N_24184);
nand UO_1136 (O_1136,N_22945,N_21319);
or UO_1137 (O_1137,N_24969,N_20748);
and UO_1138 (O_1138,N_23248,N_22419);
nor UO_1139 (O_1139,N_22726,N_20328);
xor UO_1140 (O_1140,N_24845,N_22404);
and UO_1141 (O_1141,N_23431,N_22385);
nor UO_1142 (O_1142,N_21040,N_23738);
nor UO_1143 (O_1143,N_22258,N_21425);
nand UO_1144 (O_1144,N_23704,N_24174);
nor UO_1145 (O_1145,N_21577,N_20778);
or UO_1146 (O_1146,N_20030,N_23821);
or UO_1147 (O_1147,N_23914,N_22958);
nor UO_1148 (O_1148,N_23240,N_22024);
nand UO_1149 (O_1149,N_20219,N_21083);
nand UO_1150 (O_1150,N_23619,N_20224);
and UO_1151 (O_1151,N_23719,N_21818);
and UO_1152 (O_1152,N_24092,N_22216);
and UO_1153 (O_1153,N_22310,N_24168);
nand UO_1154 (O_1154,N_20509,N_21069);
or UO_1155 (O_1155,N_21328,N_23123);
and UO_1156 (O_1156,N_21480,N_21790);
nand UO_1157 (O_1157,N_24859,N_24189);
nor UO_1158 (O_1158,N_20711,N_22359);
nand UO_1159 (O_1159,N_23432,N_21423);
or UO_1160 (O_1160,N_23737,N_20104);
nand UO_1161 (O_1161,N_22485,N_20360);
and UO_1162 (O_1162,N_23538,N_24630);
xnor UO_1163 (O_1163,N_23474,N_20303);
or UO_1164 (O_1164,N_24457,N_21158);
xnor UO_1165 (O_1165,N_24364,N_22759);
or UO_1166 (O_1166,N_22232,N_21018);
xor UO_1167 (O_1167,N_20300,N_20289);
xor UO_1168 (O_1168,N_24799,N_24037);
or UO_1169 (O_1169,N_21131,N_24238);
nor UO_1170 (O_1170,N_22256,N_23624);
nand UO_1171 (O_1171,N_22445,N_21469);
nor UO_1172 (O_1172,N_20824,N_20628);
nand UO_1173 (O_1173,N_22112,N_22459);
nor UO_1174 (O_1174,N_20410,N_24105);
xnor UO_1175 (O_1175,N_21502,N_22560);
and UO_1176 (O_1176,N_22052,N_21510);
xnor UO_1177 (O_1177,N_20230,N_22606);
xor UO_1178 (O_1178,N_22908,N_21080);
nor UO_1179 (O_1179,N_20253,N_21970);
and UO_1180 (O_1180,N_20961,N_24719);
and UO_1181 (O_1181,N_22707,N_20683);
nand UO_1182 (O_1182,N_22842,N_22283);
nand UO_1183 (O_1183,N_24705,N_24936);
nor UO_1184 (O_1184,N_24185,N_22828);
and UO_1185 (O_1185,N_22968,N_24462);
and UO_1186 (O_1186,N_24699,N_22247);
nor UO_1187 (O_1187,N_23319,N_21280);
or UO_1188 (O_1188,N_22125,N_21975);
and UO_1189 (O_1189,N_21127,N_20639);
xnor UO_1190 (O_1190,N_22778,N_21990);
nand UO_1191 (O_1191,N_22009,N_20197);
nor UO_1192 (O_1192,N_23533,N_24392);
nand UO_1193 (O_1193,N_22333,N_20043);
nor UO_1194 (O_1194,N_22203,N_24913);
nor UO_1195 (O_1195,N_22561,N_22515);
and UO_1196 (O_1196,N_21269,N_21413);
nor UO_1197 (O_1197,N_23228,N_22484);
and UO_1198 (O_1198,N_24126,N_24172);
nor UO_1199 (O_1199,N_24939,N_20221);
or UO_1200 (O_1200,N_23322,N_23002);
and UO_1201 (O_1201,N_23955,N_24851);
xnor UO_1202 (O_1202,N_23635,N_24395);
and UO_1203 (O_1203,N_23261,N_24335);
or UO_1204 (O_1204,N_23153,N_22814);
xor UO_1205 (O_1205,N_24414,N_22470);
or UO_1206 (O_1206,N_21468,N_24032);
xor UO_1207 (O_1207,N_24856,N_21312);
nor UO_1208 (O_1208,N_21301,N_21774);
nand UO_1209 (O_1209,N_20869,N_21751);
nand UO_1210 (O_1210,N_20423,N_23901);
nor UO_1211 (O_1211,N_20708,N_20379);
nand UO_1212 (O_1212,N_21623,N_24907);
xor UO_1213 (O_1213,N_24281,N_24449);
xor UO_1214 (O_1214,N_20666,N_21796);
and UO_1215 (O_1215,N_24594,N_20701);
xnor UO_1216 (O_1216,N_23781,N_20940);
nand UO_1217 (O_1217,N_21343,N_21503);
xnor UO_1218 (O_1218,N_23332,N_23298);
nand UO_1219 (O_1219,N_23872,N_21765);
nor UO_1220 (O_1220,N_21543,N_22711);
and UO_1221 (O_1221,N_22573,N_20747);
xor UO_1222 (O_1222,N_24271,N_23461);
or UO_1223 (O_1223,N_22142,N_23733);
nor UO_1224 (O_1224,N_24833,N_21963);
nand UO_1225 (O_1225,N_20464,N_24052);
nand UO_1226 (O_1226,N_22327,N_21474);
xor UO_1227 (O_1227,N_21063,N_22223);
and UO_1228 (O_1228,N_24674,N_24940);
nor UO_1229 (O_1229,N_24916,N_20499);
xnor UO_1230 (O_1230,N_22379,N_23936);
nand UO_1231 (O_1231,N_23649,N_21411);
or UO_1232 (O_1232,N_20737,N_23026);
or UO_1233 (O_1233,N_22969,N_21592);
nand UO_1234 (O_1234,N_24588,N_23407);
and UO_1235 (O_1235,N_23500,N_24009);
nand UO_1236 (O_1236,N_21945,N_20237);
or UO_1237 (O_1237,N_22897,N_21583);
nand UO_1238 (O_1238,N_21263,N_21390);
nor UO_1239 (O_1239,N_23770,N_20494);
or UO_1240 (O_1240,N_22849,N_21359);
nand UO_1241 (O_1241,N_20432,N_21187);
or UO_1242 (O_1242,N_23915,N_24850);
and UO_1243 (O_1243,N_20259,N_20887);
nand UO_1244 (O_1244,N_21195,N_24576);
nand UO_1245 (O_1245,N_21210,N_21581);
nand UO_1246 (O_1246,N_22775,N_24963);
and UO_1247 (O_1247,N_24884,N_23008);
and UO_1248 (O_1248,N_21734,N_20699);
xnor UO_1249 (O_1249,N_23549,N_21293);
or UO_1250 (O_1250,N_21318,N_20352);
nand UO_1251 (O_1251,N_23068,N_20076);
and UO_1252 (O_1252,N_20458,N_21606);
nand UO_1253 (O_1253,N_20020,N_23150);
nor UO_1254 (O_1254,N_24527,N_20016);
xnor UO_1255 (O_1255,N_20553,N_20336);
nand UO_1256 (O_1256,N_24653,N_21920);
and UO_1257 (O_1257,N_20459,N_20759);
and UO_1258 (O_1258,N_20806,N_23468);
nand UO_1259 (O_1259,N_23119,N_24481);
or UO_1260 (O_1260,N_21482,N_21295);
and UO_1261 (O_1261,N_20187,N_20605);
or UO_1262 (O_1262,N_23279,N_22339);
xor UO_1263 (O_1263,N_20696,N_24758);
nor UO_1264 (O_1264,N_24510,N_24058);
or UO_1265 (O_1265,N_24878,N_22449);
xor UO_1266 (O_1266,N_20313,N_22369);
and UO_1267 (O_1267,N_22593,N_24627);
or UO_1268 (O_1268,N_22373,N_22604);
and UO_1269 (O_1269,N_24775,N_23255);
and UO_1270 (O_1270,N_22869,N_24393);
xor UO_1271 (O_1271,N_24941,N_21698);
nand UO_1272 (O_1272,N_22889,N_23532);
nor UO_1273 (O_1273,N_23309,N_21123);
xnor UO_1274 (O_1274,N_21546,N_22806);
and UO_1275 (O_1275,N_20979,N_23917);
nand UO_1276 (O_1276,N_20602,N_22060);
or UO_1277 (O_1277,N_23270,N_22493);
nand UO_1278 (O_1278,N_20758,N_23095);
nand UO_1279 (O_1279,N_20564,N_21236);
and UO_1280 (O_1280,N_23205,N_22397);
and UO_1281 (O_1281,N_24984,N_20460);
nand UO_1282 (O_1282,N_20622,N_24246);
or UO_1283 (O_1283,N_22454,N_21927);
nor UO_1284 (O_1284,N_23871,N_20118);
nor UO_1285 (O_1285,N_24378,N_23756);
nand UO_1286 (O_1286,N_20989,N_21462);
nand UO_1287 (O_1287,N_20993,N_23029);
xnor UO_1288 (O_1288,N_21840,N_21939);
and UO_1289 (O_1289,N_22314,N_22501);
xnor UO_1290 (O_1290,N_21594,N_23371);
or UO_1291 (O_1291,N_20199,N_21910);
nand UO_1292 (O_1292,N_22135,N_23661);
and UO_1293 (O_1293,N_23211,N_20889);
nor UO_1294 (O_1294,N_22571,N_21759);
nor UO_1295 (O_1295,N_20202,N_21294);
nand UO_1296 (O_1296,N_23160,N_23721);
xor UO_1297 (O_1297,N_20644,N_24125);
or UO_1298 (O_1298,N_23900,N_20190);
or UO_1299 (O_1299,N_20742,N_22436);
nor UO_1300 (O_1300,N_24250,N_23051);
and UO_1301 (O_1301,N_20988,N_24906);
nand UO_1302 (O_1302,N_20929,N_21550);
nand UO_1303 (O_1303,N_22227,N_21723);
nor UO_1304 (O_1304,N_23856,N_22514);
or UO_1305 (O_1305,N_22622,N_21967);
and UO_1306 (O_1306,N_24725,N_22976);
and UO_1307 (O_1307,N_22547,N_22826);
or UO_1308 (O_1308,N_21116,N_21874);
and UO_1309 (O_1309,N_21530,N_22878);
nand UO_1310 (O_1310,N_20356,N_21779);
xor UO_1311 (O_1311,N_23713,N_22546);
nand UO_1312 (O_1312,N_24284,N_21340);
and UO_1313 (O_1313,N_21851,N_21562);
nand UO_1314 (O_1314,N_21701,N_20565);
xor UO_1315 (O_1315,N_22834,N_24207);
or UO_1316 (O_1316,N_21243,N_24923);
or UO_1317 (O_1317,N_23274,N_22291);
nor UO_1318 (O_1318,N_23755,N_24843);
nand UO_1319 (O_1319,N_21287,N_22088);
and UO_1320 (O_1320,N_24433,N_20679);
nand UO_1321 (O_1321,N_21724,N_20044);
xnor UO_1322 (O_1322,N_20180,N_24483);
xnor UO_1323 (O_1323,N_20061,N_22081);
xnor UO_1324 (O_1324,N_22461,N_22015);
and UO_1325 (O_1325,N_20632,N_22827);
and UO_1326 (O_1326,N_22113,N_22301);
nand UO_1327 (O_1327,N_21023,N_20463);
and UO_1328 (O_1328,N_20937,N_21604);
xnor UO_1329 (O_1329,N_23089,N_21725);
xor UO_1330 (O_1330,N_20981,N_23134);
nor UO_1331 (O_1331,N_22940,N_20055);
nor UO_1332 (O_1332,N_21298,N_23016);
xnor UO_1333 (O_1333,N_23230,N_21352);
nor UO_1334 (O_1334,N_23889,N_24139);
xor UO_1335 (O_1335,N_23505,N_23907);
or UO_1336 (O_1336,N_24055,N_22082);
nor UO_1337 (O_1337,N_21282,N_20448);
nand UO_1338 (O_1338,N_22090,N_24447);
nand UO_1339 (O_1339,N_21163,N_23052);
nand UO_1340 (O_1340,N_20718,N_20952);
nand UO_1341 (O_1341,N_23552,N_20340);
nor UO_1342 (O_1342,N_22899,N_21712);
and UO_1343 (O_1343,N_24469,N_23577);
xnor UO_1344 (O_1344,N_24771,N_21527);
or UO_1345 (O_1345,N_22875,N_24666);
nand UO_1346 (O_1346,N_24787,N_23443);
nor UO_1347 (O_1347,N_23578,N_24550);
nor UO_1348 (O_1348,N_21715,N_24811);
nor UO_1349 (O_1349,N_23834,N_20394);
or UO_1350 (O_1350,N_23005,N_22995);
nand UO_1351 (O_1351,N_23012,N_23085);
and UO_1352 (O_1352,N_23717,N_23206);
and UO_1353 (O_1353,N_22453,N_24633);
or UO_1354 (O_1354,N_24976,N_21177);
xnor UO_1355 (O_1355,N_23115,N_24039);
or UO_1356 (O_1356,N_23343,N_22389);
or UO_1357 (O_1357,N_21717,N_24860);
nor UO_1358 (O_1358,N_22739,N_24613);
or UO_1359 (O_1359,N_23696,N_24036);
or UO_1360 (O_1360,N_20312,N_24213);
xor UO_1361 (O_1361,N_21976,N_22713);
and UO_1362 (O_1362,N_21960,N_23004);
and UO_1363 (O_1363,N_23586,N_24286);
nand UO_1364 (O_1364,N_24628,N_24864);
or UO_1365 (O_1365,N_21447,N_23895);
or UO_1366 (O_1366,N_23030,N_23223);
nand UO_1367 (O_1367,N_20646,N_21663);
nor UO_1368 (O_1368,N_23875,N_24013);
xor UO_1369 (O_1369,N_22794,N_21622);
nand UO_1370 (O_1370,N_20892,N_23235);
nand UO_1371 (O_1371,N_21053,N_24377);
nor UO_1372 (O_1372,N_22716,N_21139);
or UO_1373 (O_1373,N_23237,N_20345);
xor UO_1374 (O_1374,N_20102,N_21688);
or UO_1375 (O_1375,N_22294,N_22562);
and UO_1376 (O_1376,N_21822,N_24345);
or UO_1377 (O_1377,N_20913,N_24320);
and UO_1378 (O_1378,N_24240,N_20581);
or UO_1379 (O_1379,N_20867,N_22610);
xnor UO_1380 (O_1380,N_21081,N_23138);
and UO_1381 (O_1381,N_23102,N_22139);
xor UO_1382 (O_1382,N_22045,N_20580);
and UO_1383 (O_1383,N_20880,N_23124);
and UO_1384 (O_1384,N_23222,N_23656);
xnor UO_1385 (O_1385,N_20308,N_22408);
or UO_1386 (O_1386,N_23627,N_24212);
xor UO_1387 (O_1387,N_21895,N_24210);
and UO_1388 (O_1388,N_22399,N_21363);
nand UO_1389 (O_1389,N_20548,N_20233);
or UO_1390 (O_1390,N_23106,N_20920);
xor UO_1391 (O_1391,N_22621,N_23059);
nor UO_1392 (O_1392,N_21144,N_21889);
and UO_1393 (O_1393,N_23394,N_21337);
or UO_1394 (O_1394,N_23412,N_23799);
nor UO_1395 (O_1395,N_23840,N_20546);
or UO_1396 (O_1396,N_21348,N_23473);
nor UO_1397 (O_1397,N_21695,N_23290);
or UO_1398 (O_1398,N_24188,N_22097);
nor UO_1399 (O_1399,N_22623,N_21157);
and UO_1400 (O_1400,N_24471,N_22296);
xnor UO_1401 (O_1401,N_20571,N_23459);
nor UO_1402 (O_1402,N_24129,N_24682);
nor UO_1403 (O_1403,N_24947,N_24382);
nand UO_1404 (O_1404,N_20122,N_20117);
xnor UO_1405 (O_1405,N_22199,N_21523);
or UO_1406 (O_1406,N_22421,N_23867);
and UO_1407 (O_1407,N_24645,N_23725);
nand UO_1408 (O_1408,N_24746,N_21860);
nor UO_1409 (O_1409,N_23881,N_21031);
nor UO_1410 (O_1410,N_24524,N_22344);
or UO_1411 (O_1411,N_21072,N_21133);
and UO_1412 (O_1412,N_21897,N_22704);
and UO_1413 (O_1413,N_24062,N_20601);
nand UO_1414 (O_1414,N_20787,N_23047);
xor UO_1415 (O_1415,N_21075,N_21073);
and UO_1416 (O_1416,N_22883,N_24732);
nor UO_1417 (O_1417,N_22451,N_20769);
and UO_1418 (O_1418,N_24065,N_24677);
nor UO_1419 (O_1419,N_20433,N_20168);
and UO_1420 (O_1420,N_22819,N_22260);
and UO_1421 (O_1421,N_24544,N_24180);
nand UO_1422 (O_1422,N_20858,N_24714);
and UO_1423 (O_1423,N_20765,N_20525);
and UO_1424 (O_1424,N_20815,N_24968);
and UO_1425 (O_1425,N_23393,N_24838);
nand UO_1426 (O_1426,N_20333,N_21102);
and UO_1427 (O_1427,N_24844,N_20654);
nand UO_1428 (O_1428,N_20485,N_20386);
nand UO_1429 (O_1429,N_20606,N_23698);
and UO_1430 (O_1430,N_21309,N_21776);
and UO_1431 (O_1431,N_23752,N_23735);
or UO_1432 (O_1432,N_21441,N_22005);
nor UO_1433 (O_1433,N_23242,N_24700);
or UO_1434 (O_1434,N_24121,N_23518);
nor UO_1435 (O_1435,N_22966,N_23402);
and UO_1436 (O_1436,N_20797,N_23645);
or UO_1437 (O_1437,N_20059,N_21335);
xor UO_1438 (O_1438,N_24015,N_21882);
nor UO_1439 (O_1439,N_23378,N_24985);
xor UO_1440 (O_1440,N_21676,N_24318);
nand UO_1441 (O_1441,N_21407,N_22825);
nand UO_1442 (O_1442,N_21992,N_24648);
and UO_1443 (O_1443,N_23653,N_20216);
nor UO_1444 (O_1444,N_21643,N_23508);
xnor UO_1445 (O_1445,N_20633,N_21253);
xor UO_1446 (O_1446,N_22689,N_22637);
nand UO_1447 (O_1447,N_21603,N_23880);
or UO_1448 (O_1448,N_20235,N_24579);
nor UO_1449 (O_1449,N_20011,N_20002);
xor UO_1450 (O_1450,N_20160,N_21925);
and UO_1451 (O_1451,N_20257,N_22244);
nor UO_1452 (O_1452,N_21628,N_23829);
or UO_1453 (O_1453,N_24722,N_24311);
nand UO_1454 (O_1454,N_22594,N_23396);
nor UO_1455 (O_1455,N_22960,N_24357);
nor UO_1456 (O_1456,N_22381,N_22509);
nand UO_1457 (O_1457,N_23987,N_23188);
nand UO_1458 (O_1458,N_21588,N_24324);
and UO_1459 (O_1459,N_23978,N_24353);
nand UO_1460 (O_1460,N_21699,N_20376);
or UO_1461 (O_1461,N_20612,N_24639);
or UO_1462 (O_1462,N_23682,N_21088);
and UO_1463 (O_1463,N_21681,N_24792);
nor UO_1464 (O_1464,N_23308,N_21231);
or UO_1465 (O_1465,N_24620,N_21091);
xnor UO_1466 (O_1466,N_23419,N_24608);
and UO_1467 (O_1467,N_24155,N_24131);
and UO_1468 (O_1468,N_20542,N_22507);
nor UO_1469 (O_1469,N_23643,N_24912);
nor UO_1470 (O_1470,N_23227,N_24667);
or UO_1471 (O_1471,N_23324,N_23519);
xor UO_1472 (O_1472,N_21785,N_23072);
and UO_1473 (O_1473,N_22480,N_21750);
nor UO_1474 (O_1474,N_24459,N_20422);
nor UO_1475 (O_1475,N_21998,N_24581);
and UO_1476 (O_1476,N_21203,N_24109);
nor UO_1477 (O_1477,N_23321,N_21940);
xnor UO_1478 (O_1478,N_20933,N_24263);
and UO_1479 (O_1479,N_21847,N_20437);
or UO_1480 (O_1480,N_24400,N_23391);
xor UO_1481 (O_1481,N_20483,N_24925);
nor UO_1482 (O_1482,N_23159,N_21314);
or UO_1483 (O_1483,N_21988,N_21004);
and UO_1484 (O_1484,N_22303,N_23506);
nand UO_1485 (O_1485,N_21147,N_24056);
nor UO_1486 (O_1486,N_23692,N_23745);
nor UO_1487 (O_1487,N_24711,N_22035);
xor UO_1488 (O_1488,N_20963,N_24379);
and UO_1489 (O_1489,N_20912,N_23446);
nor UO_1490 (O_1490,N_23152,N_21598);
nand UO_1491 (O_1491,N_22796,N_23826);
nand UO_1492 (O_1492,N_24572,N_22174);
nor UO_1493 (O_1493,N_24942,N_20052);
nor UO_1494 (O_1494,N_21907,N_22880);
and UO_1495 (O_1495,N_22891,N_24791);
xnor UO_1496 (O_1496,N_24274,N_24477);
nand UO_1497 (O_1497,N_23662,N_21522);
nor UO_1498 (O_1498,N_20001,N_22050);
xor UO_1499 (O_1499,N_24312,N_23960);
and UO_1500 (O_1500,N_20839,N_23633);
xnor UO_1501 (O_1501,N_24408,N_24235);
and UO_1502 (O_1502,N_21626,N_21547);
or UO_1503 (O_1503,N_21036,N_20124);
nand UO_1504 (O_1504,N_24506,N_23772);
nor UO_1505 (O_1505,N_22837,N_20136);
or UO_1506 (O_1506,N_20006,N_20185);
and UO_1507 (O_1507,N_24935,N_23179);
or UO_1508 (O_1508,N_22276,N_20178);
xor UO_1509 (O_1509,N_22182,N_23271);
or UO_1510 (O_1510,N_23302,N_21377);
or UO_1511 (O_1511,N_23981,N_21572);
nor UO_1512 (O_1512,N_21098,N_23436);
nor UO_1513 (O_1513,N_22804,N_23732);
or UO_1514 (O_1514,N_22727,N_23494);
nand UO_1515 (O_1515,N_20286,N_21289);
xor UO_1516 (O_1516,N_24413,N_24479);
or UO_1517 (O_1517,N_24503,N_21251);
and UO_1518 (O_1518,N_22422,N_24515);
nor UO_1519 (O_1519,N_23369,N_20809);
and UO_1520 (O_1520,N_20132,N_20510);
nand UO_1521 (O_1521,N_23379,N_20749);
nand UO_1522 (O_1522,N_23796,N_21440);
xnor UO_1523 (O_1523,N_20031,N_20614);
nand UO_1524 (O_1524,N_24804,N_24892);
or UO_1525 (O_1525,N_23381,N_22640);
nor UO_1526 (O_1526,N_24098,N_24695);
and UO_1527 (O_1527,N_24839,N_20784);
nand UO_1528 (O_1528,N_24820,N_23844);
nor UO_1529 (O_1529,N_20182,N_21130);
nor UO_1530 (O_1530,N_21456,N_24314);
xnor UO_1531 (O_1531,N_20798,N_24086);
and UO_1532 (O_1532,N_24018,N_22712);
and UO_1533 (O_1533,N_24073,N_20941);
nand UO_1534 (O_1534,N_21485,N_21817);
nand UO_1535 (O_1535,N_23214,N_20641);
nand UO_1536 (O_1536,N_20271,N_22595);
and UO_1537 (O_1537,N_23830,N_24650);
nor UO_1538 (O_1538,N_24866,N_24219);
xor UO_1539 (O_1539,N_22608,N_23389);
xnor UO_1540 (O_1540,N_22098,N_22488);
nand UO_1541 (O_1541,N_20725,N_22398);
or UO_1542 (O_1542,N_21467,N_23569);
and UO_1543 (O_1543,N_24332,N_24193);
and UO_1544 (O_1544,N_23028,N_23531);
nor UO_1545 (O_1545,N_21640,N_22162);
and UO_1546 (O_1546,N_24621,N_23882);
nor UO_1547 (O_1547,N_23780,N_22786);
xnor UO_1548 (O_1548,N_21165,N_20893);
nor UO_1549 (O_1549,N_24542,N_22768);
xor UO_1550 (O_1550,N_22409,N_24023);
nor UO_1551 (O_1551,N_24456,N_21982);
nor UO_1552 (O_1552,N_24871,N_21470);
nand UO_1553 (O_1553,N_21662,N_22075);
nor UO_1554 (O_1554,N_24928,N_24531);
nor UO_1555 (O_1555,N_24267,N_20775);
nor UO_1556 (O_1556,N_22309,N_22171);
xnor UO_1557 (O_1557,N_22760,N_23080);
or UO_1558 (O_1558,N_21382,N_20015);
or UO_1559 (O_1559,N_24234,N_23427);
xor UO_1560 (O_1560,N_22161,N_21909);
or UO_1561 (O_1561,N_23185,N_21793);
xor UO_1562 (O_1562,N_20517,N_23367);
xnor UO_1563 (O_1563,N_23576,N_20554);
xor UO_1564 (O_1564,N_22808,N_22692);
nand UO_1565 (O_1565,N_23793,N_21761);
or UO_1566 (O_1566,N_23720,N_21771);
or UO_1567 (O_1567,N_21926,N_24467);
nand UO_1568 (O_1568,N_22655,N_20242);
nor UO_1569 (O_1569,N_21921,N_22394);
or UO_1570 (O_1570,N_22166,N_22236);
and UO_1571 (O_1571,N_22196,N_21152);
or UO_1572 (O_1572,N_23681,N_23954);
nor UO_1573 (O_1573,N_23919,N_20619);
nor UO_1574 (O_1574,N_23965,N_22094);
xnor UO_1575 (O_1575,N_24280,N_23962);
and UO_1576 (O_1576,N_22341,N_24698);
and UO_1577 (O_1577,N_20702,N_23447);
nor UO_1578 (O_1578,N_21489,N_22270);
nand UO_1579 (O_1579,N_23334,N_23482);
or UO_1580 (O_1580,N_23340,N_24501);
or UO_1581 (O_1581,N_20473,N_22374);
and UO_1582 (O_1582,N_22941,N_23452);
nand UO_1583 (O_1583,N_20246,N_24081);
or UO_1584 (O_1584,N_24960,N_24569);
nand UO_1585 (O_1585,N_24115,N_23176);
and UO_1586 (O_1586,N_23797,N_21020);
nor UO_1587 (O_1587,N_23287,N_23262);
nor UO_1588 (O_1588,N_22500,N_22109);
nand UO_1589 (O_1589,N_24028,N_20968);
xor UO_1590 (O_1590,N_24014,N_24004);
xnor UO_1591 (O_1591,N_21229,N_23019);
nand UO_1592 (O_1592,N_24759,N_21463);
or UO_1593 (O_1593,N_23828,N_23117);
or UO_1594 (O_1594,N_23014,N_23839);
or UO_1595 (O_1595,N_24047,N_23277);
and UO_1596 (O_1596,N_23808,N_22627);
and UO_1597 (O_1597,N_21894,N_24130);
xnor UO_1598 (O_1598,N_24012,N_23180);
and UO_1599 (O_1599,N_24846,N_24046);
nor UO_1600 (O_1600,N_21566,N_20804);
or UO_1601 (O_1601,N_24823,N_21439);
xor UO_1602 (O_1602,N_22074,N_20960);
or UO_1603 (O_1603,N_20603,N_22881);
and UO_1604 (O_1604,N_22427,N_23295);
nor UO_1605 (O_1605,N_22220,N_20149);
or UO_1606 (O_1606,N_20142,N_20282);
and UO_1607 (O_1607,N_21564,N_21005);
nor UO_1608 (O_1608,N_24202,N_24386);
or UO_1609 (O_1609,N_22519,N_23758);
xor UO_1610 (O_1610,N_22840,N_23547);
nand UO_1611 (O_1611,N_22215,N_22744);
or UO_1612 (O_1612,N_24617,N_23244);
nor UO_1613 (O_1613,N_24543,N_23232);
and UO_1614 (O_1614,N_22585,N_21832);
nand UO_1615 (O_1615,N_22204,N_22411);
nor UO_1616 (O_1616,N_20415,N_23209);
nand UO_1617 (O_1617,N_23782,N_21240);
nand UO_1618 (O_1618,N_20330,N_23039);
xnor UO_1619 (O_1619,N_24794,N_21631);
nor UO_1620 (O_1620,N_20786,N_24568);
and UO_1621 (O_1621,N_20281,N_20707);
xnor UO_1622 (O_1622,N_24440,N_21333);
or UO_1623 (O_1623,N_20420,N_21078);
nand UO_1624 (O_1624,N_21432,N_24482);
nor UO_1625 (O_1625,N_21952,N_20983);
and UO_1626 (O_1626,N_20875,N_23363);
nand UO_1627 (O_1627,N_20588,N_23957);
nand UO_1628 (O_1628,N_21740,N_20753);
xor UO_1629 (O_1629,N_20812,N_22272);
or UO_1630 (O_1630,N_22124,N_21266);
nand UO_1631 (O_1631,N_21515,N_21947);
or UO_1632 (O_1632,N_23979,N_22129);
xnor UO_1633 (O_1633,N_24706,N_20834);
xnor UO_1634 (O_1634,N_22077,N_22926);
xnor UO_1635 (O_1635,N_23997,N_23966);
nand UO_1636 (O_1636,N_23318,N_23614);
nand UO_1637 (O_1637,N_20740,N_21375);
xor UO_1638 (O_1638,N_21613,N_22504);
nor UO_1639 (O_1639,N_23183,N_22212);
nor UO_1640 (O_1640,N_21228,N_24591);
xor UO_1641 (O_1641,N_20600,N_22289);
xor UO_1642 (O_1642,N_24580,N_20453);
or UO_1643 (O_1643,N_22056,N_22455);
or UO_1644 (O_1644,N_21878,N_22567);
and UO_1645 (O_1645,N_24610,N_22342);
xnor UO_1646 (O_1646,N_22390,N_22525);
or UO_1647 (O_1647,N_20470,N_22187);
and UO_1648 (O_1648,N_21277,N_20358);
nor UO_1649 (O_1649,N_22663,N_24603);
nor UO_1650 (O_1650,N_21122,N_21520);
and UO_1651 (O_1651,N_24673,N_24870);
or UO_1652 (O_1652,N_20900,N_21684);
nand UO_1653 (O_1653,N_24631,N_20562);
nor UO_1654 (O_1654,N_22354,N_21501);
nand UO_1655 (O_1655,N_21629,N_22335);
and UO_1656 (O_1656,N_22365,N_24519);
nand UO_1657 (O_1657,N_23144,N_22200);
and UO_1658 (O_1658,N_24547,N_24222);
nor UO_1659 (O_1659,N_20616,N_21050);
nor UO_1660 (O_1660,N_24398,N_24702);
xor UO_1661 (O_1661,N_24994,N_23236);
and UO_1662 (O_1662,N_22782,N_22307);
nand UO_1663 (O_1663,N_23219,N_20096);
nand UO_1664 (O_1664,N_23595,N_24236);
and UO_1665 (O_1665,N_20276,N_22979);
xor UO_1666 (O_1666,N_23723,N_23798);
nor UO_1667 (O_1667,N_20082,N_21016);
and UO_1668 (O_1668,N_24116,N_24132);
or UO_1669 (O_1669,N_24596,N_20543);
and UO_1670 (O_1670,N_21714,N_23540);
and UO_1671 (O_1671,N_24452,N_23604);
nand UO_1672 (O_1672,N_24094,N_20491);
xnor UO_1673 (O_1673,N_22502,N_20467);
or UO_1674 (O_1674,N_24554,N_24134);
xnor UO_1675 (O_1675,N_22578,N_24972);
nand UO_1676 (O_1676,N_22321,N_21473);
or UO_1677 (O_1677,N_23139,N_24374);
nor UO_1678 (O_1678,N_21428,N_21049);
or UO_1679 (O_1679,N_22638,N_23972);
xor UO_1680 (O_1680,N_20882,N_23617);
and UO_1681 (O_1681,N_21916,N_21711);
and UO_1682 (O_1682,N_21446,N_22809);
xor UO_1683 (O_1683,N_21188,N_21220);
xnor UO_1684 (O_1684,N_22240,N_20836);
or UO_1685 (O_1685,N_20555,N_23762);
or UO_1686 (O_1686,N_21156,N_23374);
or UO_1687 (O_1687,N_22857,N_20041);
nor UO_1688 (O_1688,N_20272,N_22116);
nand UO_1689 (O_1689,N_23822,N_23579);
nor UO_1690 (O_1690,N_24559,N_21199);
and UO_1691 (O_1691,N_21197,N_22110);
xnor UO_1692 (O_1692,N_22831,N_20091);
and UO_1693 (O_1693,N_23553,N_23145);
xnor UO_1694 (O_1694,N_21730,N_20938);
xor UO_1695 (O_1695,N_21507,N_22169);
and UO_1696 (O_1696,N_24391,N_24123);
nand UO_1697 (O_1697,N_22317,N_24488);
nor UO_1698 (O_1698,N_22765,N_24731);
nand UO_1699 (O_1699,N_20316,N_22954);
nand UO_1700 (O_1700,N_24355,N_24294);
nor UO_1701 (O_1701,N_23263,N_24112);
nand UO_1702 (O_1702,N_22728,N_20169);
nor UO_1703 (O_1703,N_21627,N_22678);
xnor UO_1704 (O_1704,N_20243,N_20924);
and UO_1705 (O_1705,N_23168,N_24889);
nand UO_1706 (O_1706,N_20801,N_24436);
xnor UO_1707 (O_1707,N_20100,N_23742);
xor UO_1708 (O_1708,N_24301,N_21949);
and UO_1709 (O_1709,N_24216,N_24886);
or UO_1710 (O_1710,N_20222,N_21931);
nand UO_1711 (O_1711,N_24359,N_20071);
xor UO_1712 (O_1712,N_22010,N_24316);
nand UO_1713 (O_1713,N_23365,N_20568);
xor UO_1714 (O_1714,N_20559,N_22336);
nand UO_1715 (O_1715,N_20098,N_22902);
nand UO_1716 (O_1716,N_21559,N_23297);
and UO_1717 (O_1717,N_21409,N_23406);
or UO_1718 (O_1718,N_22904,N_22152);
and UO_1719 (O_1719,N_21834,N_20684);
xnor UO_1720 (O_1720,N_20495,N_23694);
nand UO_1721 (O_1721,N_21190,N_20277);
xnor UO_1722 (O_1722,N_21205,N_21154);
nand UO_1723 (O_1723,N_24077,N_22884);
nor UO_1724 (O_1724,N_20480,N_20533);
xnor UO_1725 (O_1725,N_21722,N_22262);
or UO_1726 (O_1726,N_20038,N_22900);
or UO_1727 (O_1727,N_22352,N_22046);
or UO_1728 (O_1728,N_22165,N_23628);
or UO_1729 (O_1729,N_24149,N_24108);
and UO_1730 (O_1730,N_22176,N_21838);
nor UO_1731 (O_1731,N_21259,N_24147);
nor UO_1732 (O_1732,N_22095,N_22791);
and UO_1733 (O_1733,N_20406,N_22949);
xor UO_1734 (O_1734,N_23803,N_20342);
nor UO_1735 (O_1735,N_24555,N_20928);
nand UO_1736 (O_1736,N_20361,N_24146);
and UO_1737 (O_1737,N_23315,N_23605);
xor UO_1738 (O_1738,N_23040,N_24136);
and UO_1739 (O_1739,N_24435,N_24676);
xnor UO_1740 (O_1740,N_22188,N_21544);
xnor UO_1741 (O_1741,N_24022,N_20577);
xor UO_1742 (O_1742,N_24298,N_22522);
nand UO_1743 (O_1743,N_24051,N_24945);
xnor UO_1744 (O_1744,N_23316,N_24641);
and UO_1745 (O_1745,N_23640,N_20948);
and UO_1746 (O_1746,N_24191,N_24534);
or UO_1747 (O_1747,N_20191,N_23201);
xnor UO_1748 (O_1748,N_22091,N_21033);
xnor UO_1749 (O_1749,N_21508,N_22458);
nand UO_1750 (O_1750,N_20741,N_22104);
nand UO_1751 (O_1751,N_23493,N_21548);
nor UO_1752 (O_1752,N_22487,N_23370);
nand UO_1753 (O_1753,N_24883,N_22358);
or UO_1754 (O_1754,N_22855,N_21175);
nand UO_1755 (O_1755,N_22783,N_22570);
and UO_1756 (O_1756,N_22559,N_23594);
nand UO_1757 (O_1757,N_22882,N_24026);
nand UO_1758 (O_1758,N_23383,N_22599);
nor UO_1759 (O_1759,N_21498,N_22929);
and UO_1760 (O_1760,N_24988,N_23864);
nor UO_1761 (O_1761,N_21879,N_20024);
nor UO_1762 (O_1762,N_20147,N_24687);
nor UO_1763 (O_1763,N_20287,N_24713);
xnor UO_1764 (O_1764,N_22413,N_20200);
xnor UO_1765 (O_1765,N_24384,N_20569);
or UO_1766 (O_1766,N_20145,N_23066);
or UO_1767 (O_1767,N_21981,N_20186);
or UO_1768 (O_1768,N_21816,N_21445);
and UO_1769 (O_1769,N_21813,N_24460);
and UO_1770 (O_1770,N_22588,N_24822);
nor UO_1771 (O_1771,N_20474,N_24361);
nand UO_1772 (O_1772,N_22720,N_21589);
nand UO_1773 (O_1773,N_22338,N_20363);
nand UO_1774 (O_1774,N_24814,N_23216);
xnor UO_1775 (O_1775,N_22316,N_20069);
nor UO_1776 (O_1776,N_20471,N_23975);
nand UO_1777 (O_1777,N_21933,N_23077);
or UO_1778 (O_1778,N_24340,N_22691);
and UO_1779 (O_1779,N_24728,N_21395);
xnor UO_1780 (O_1780,N_22068,N_21394);
nand UO_1781 (O_1781,N_22122,N_22265);
xor UO_1782 (O_1782,N_23225,N_20505);
and UO_1783 (O_1783,N_24658,N_24007);
or UO_1784 (O_1784,N_20150,N_23988);
nor UO_1785 (O_1785,N_23790,N_24201);
xnor UO_1786 (O_1786,N_23922,N_20842);
nor UO_1787 (O_1787,N_21066,N_23331);
xor UO_1788 (O_1788,N_24571,N_24605);
xor UO_1789 (O_1789,N_21176,N_22156);
and UO_1790 (O_1790,N_20923,N_21845);
xor UO_1791 (O_1791,N_20526,N_24978);
nand UO_1792 (O_1792,N_23147,N_24177);
nand UO_1793 (O_1793,N_22942,N_20640);
xnor UO_1794 (O_1794,N_23836,N_22800);
nor UO_1795 (O_1795,N_22860,N_24615);
and UO_1796 (O_1796,N_24195,N_23591);
xor UO_1797 (O_1797,N_23355,N_22030);
or UO_1798 (O_1798,N_22295,N_24948);
xor UO_1799 (O_1799,N_24974,N_22257);
or UO_1800 (O_1800,N_22143,N_24927);
or UO_1801 (O_1801,N_20906,N_21534);
xnor UO_1802 (O_1802,N_20108,N_20444);
nor UO_1803 (O_1803,N_21214,N_21903);
or UO_1804 (O_1804,N_22334,N_20120);
and UO_1805 (O_1805,N_22780,N_23664);
nor UO_1806 (O_1806,N_24643,N_24463);
and UO_1807 (O_1807,N_24504,N_22412);
or UO_1808 (O_1808,N_20512,N_21944);
xnor UO_1809 (O_1809,N_20450,N_20354);
or UO_1810 (O_1810,N_22802,N_24733);
nor UO_1811 (O_1811,N_24551,N_22092);
xor UO_1812 (O_1812,N_22696,N_21573);
nand UO_1813 (O_1813,N_22617,N_21009);
nand UO_1814 (O_1814,N_23092,N_24053);
and UO_1815 (O_1815,N_21595,N_22225);
or UO_1816 (O_1816,N_23879,N_23554);
nor UO_1817 (O_1817,N_21084,N_23652);
xor UO_1818 (O_1818,N_22013,N_21415);
nand UO_1819 (O_1819,N_24660,N_20274);
or UO_1820 (O_1820,N_24330,N_23234);
xor UO_1821 (O_1821,N_24085,N_20375);
and UO_1822 (O_1822,N_23655,N_21012);
or UO_1823 (O_1823,N_23258,N_20503);
xor UO_1824 (O_1824,N_20225,N_20680);
and UO_1825 (O_1825,N_20240,N_21162);
or UO_1826 (O_1826,N_24997,N_20029);
nand UO_1827 (O_1827,N_20434,N_21351);
and UO_1828 (O_1828,N_23056,N_24949);
and UO_1829 (O_1829,N_24806,N_22558);
nor UO_1830 (O_1830,N_20864,N_22405);
or UO_1831 (O_1831,N_20835,N_21948);
and UO_1832 (O_1832,N_21302,N_24962);
xor UO_1833 (O_1833,N_24508,N_23610);
and UO_1834 (O_1834,N_24557,N_20309);
nor UO_1835 (O_1835,N_24093,N_24849);
or UO_1836 (O_1836,N_21666,N_23683);
xnor UO_1837 (O_1837,N_20349,N_20244);
xnor UO_1838 (O_1838,N_21946,N_21721);
or UO_1839 (O_1839,N_23730,N_22266);
xor UO_1840 (O_1840,N_20174,N_21787);
and UO_1841 (O_1841,N_24461,N_23204);
nor UO_1842 (O_1842,N_22609,N_23100);
and UO_1843 (O_1843,N_20331,N_21686);
nor UO_1844 (O_1844,N_21056,N_24486);
and UO_1845 (O_1845,N_23847,N_20245);
and UO_1846 (O_1846,N_22630,N_22731);
nor UO_1847 (O_1847,N_21227,N_21011);
xor UO_1848 (O_1848,N_22517,N_23813);
or UO_1849 (O_1849,N_24513,N_22491);
or UO_1850 (O_1850,N_21749,N_21570);
and UO_1851 (O_1851,N_21689,N_20374);
and UO_1852 (O_1852,N_20248,N_20455);
xor UO_1853 (O_1853,N_21198,N_22076);
or UO_1854 (O_1854,N_20310,N_20163);
xor UO_1855 (O_1855,N_20682,N_23253);
xor UO_1856 (O_1856,N_20321,N_20557);
and UO_1857 (O_1857,N_21579,N_24290);
or UO_1858 (O_1858,N_24255,N_22144);
nor UO_1859 (O_1859,N_24362,N_24885);
or UO_1860 (O_1860,N_23556,N_24118);
and UO_1861 (O_1861,N_20161,N_24144);
nor UO_1862 (O_1862,N_21365,N_23032);
and UO_1863 (O_1863,N_21735,N_21219);
or UO_1864 (O_1864,N_20907,N_21379);
and UO_1865 (O_1865,N_24381,N_21511);
and UO_1866 (O_1866,N_22695,N_21591);
or UO_1867 (O_1867,N_24091,N_24529);
nor UO_1868 (O_1868,N_22019,N_23354);
nor UO_1869 (O_1869,N_22472,N_21388);
and UO_1870 (O_1870,N_21286,N_22285);
and UO_1871 (O_1871,N_24766,N_22053);
or UO_1872 (O_1872,N_23312,N_24348);
or UO_1873 (O_1873,N_21999,N_21744);
nor UO_1874 (O_1874,N_23107,N_23104);
nor UO_1875 (O_1875,N_20643,N_24487);
or UO_1876 (O_1876,N_21323,N_20288);
nor UO_1877 (O_1877,N_21582,N_24401);
nand UO_1878 (O_1878,N_20157,N_20128);
xnor UO_1879 (O_1879,N_20717,N_20054);
nor UO_1880 (O_1880,N_21064,N_20589);
nand UO_1881 (O_1881,N_24084,N_24640);
or UO_1882 (O_1882,N_21481,N_21464);
or UO_1883 (O_1883,N_24493,N_21738);
and UO_1884 (O_1884,N_20848,N_23276);
xor UO_1885 (O_1885,N_20269,N_20103);
or UO_1886 (O_1886,N_21871,N_23284);
and UO_1887 (O_1887,N_21571,N_20868);
nor UO_1888 (O_1888,N_23939,N_23986);
and UO_1889 (O_1889,N_23952,N_23935);
xor UO_1890 (O_1890,N_24709,N_24855);
nand UO_1891 (O_1891,N_22607,N_22271);
nand UO_1892 (O_1892,N_24910,N_23792);
nor UO_1893 (O_1893,N_24999,N_21718);
nand UO_1894 (O_1894,N_22325,N_23849);
nor UO_1895 (O_1895,N_24828,N_21128);
nor UO_1896 (O_1896,N_21835,N_23278);
nor UO_1897 (O_1897,N_24670,N_21873);
or UO_1898 (O_1898,N_20760,N_20773);
or UO_1899 (O_1899,N_23178,N_23715);
nor UO_1900 (O_1900,N_22867,N_23636);
or UO_1901 (O_1901,N_23926,N_23345);
or UO_1902 (O_1902,N_20032,N_23942);
xor UO_1903 (O_1903,N_22847,N_22178);
and UO_1904 (O_1904,N_20063,N_21883);
or UO_1905 (O_1905,N_21108,N_24857);
nand UO_1906 (O_1906,N_21141,N_20487);
nor UO_1907 (O_1907,N_20688,N_24895);
xor UO_1908 (O_1908,N_24303,N_23634);
nand UO_1909 (O_1909,N_20367,N_24367);
and UO_1910 (O_1910,N_20256,N_20087);
or UO_1911 (O_1911,N_21173,N_22141);
and UO_1912 (O_1912,N_21160,N_20359);
and UO_1913 (O_1913,N_22664,N_24904);
nand UO_1914 (O_1914,N_24167,N_23724);
or UO_1915 (O_1915,N_20402,N_20524);
and UO_1916 (O_1916,N_22490,N_21525);
xnor UO_1917 (O_1917,N_22140,N_22586);
nand UO_1918 (O_1918,N_20166,N_24495);
nand UO_1919 (O_1919,N_24938,N_23082);
nand UO_1920 (O_1920,N_24685,N_22614);
nand UO_1921 (O_1921,N_20714,N_20368);
nand UO_1922 (O_1922,N_24042,N_22432);
or UO_1923 (O_1923,N_24064,N_23121);
xor UO_1924 (O_1924,N_23943,N_21800);
nand UO_1925 (O_1925,N_20111,N_20734);
nand UO_1926 (O_1926,N_20764,N_21665);
xnor UO_1927 (O_1927,N_22784,N_22530);
and UO_1928 (O_1928,N_21322,N_23584);
and UO_1929 (O_1929,N_23524,N_21167);
nor UO_1930 (O_1930,N_24915,N_20802);
xnor UO_1931 (O_1931,N_21656,N_20318);
or UO_1932 (O_1932,N_23510,N_22858);
nand UO_1933 (O_1933,N_20181,N_24396);
nand UO_1934 (O_1934,N_21941,N_21679);
xnor UO_1935 (O_1935,N_24305,N_22137);
nand UO_1936 (O_1936,N_22224,N_22506);
nand UO_1937 (O_1937,N_22852,N_22395);
or UO_1938 (O_1938,N_24237,N_20457);
and UO_1939 (O_1939,N_24651,N_21105);
nor UO_1940 (O_1940,N_24070,N_20211);
nor UO_1941 (O_1941,N_24689,N_24478);
nor UO_1942 (O_1942,N_22551,N_20994);
or UO_1943 (O_1943,N_23325,N_22890);
nor UO_1944 (O_1944,N_24183,N_22905);
nand UO_1945 (O_1945,N_22927,N_20260);
xor UO_1946 (O_1946,N_20317,N_21125);
or UO_1947 (O_1947,N_22807,N_21977);
xor UO_1948 (O_1948,N_21786,N_23033);
xor UO_1949 (O_1949,N_21602,N_24397);
xor UO_1950 (O_1950,N_23769,N_21856);
nand UO_1951 (O_1951,N_22031,N_22666);
nand UO_1952 (O_1952,N_23666,N_22269);
nor UO_1953 (O_1953,N_20507,N_20574);
xor UO_1954 (O_1954,N_21671,N_22779);
nor UO_1955 (O_1955,N_21239,N_22992);
or UO_1956 (O_1956,N_23327,N_23113);
or UO_1957 (O_1957,N_22329,N_20254);
and UO_1958 (O_1958,N_24119,N_20916);
or UO_1959 (O_1959,N_23825,N_22120);
nor UO_1960 (O_1960,N_22228,N_23687);
nand UO_1961 (O_1961,N_23409,N_23411);
and UO_1962 (O_1962,N_24103,N_20493);
nor UO_1963 (O_1963,N_20777,N_21844);
and UO_1964 (O_1964,N_20370,N_24034);
or UO_1965 (O_1965,N_23850,N_22527);
xnor UO_1966 (O_1966,N_23536,N_23951);
or UO_1967 (O_1967,N_24328,N_20497);
and UO_1968 (O_1968,N_21633,N_23658);
nand UO_1969 (O_1969,N_23175,N_24977);
and UO_1970 (O_1970,N_23034,N_22471);
xor UO_1971 (O_1971,N_21204,N_20291);
nor UO_1972 (O_1972,N_22859,N_22918);
nand UO_1973 (O_1973,N_21682,N_20705);
xor UO_1974 (O_1974,N_21224,N_22741);
xnor UO_1975 (O_1975,N_22575,N_21117);
nand UO_1976 (O_1976,N_23902,N_20732);
and UO_1977 (O_1977,N_23167,N_23760);
or UO_1978 (O_1978,N_22363,N_23920);
nand UO_1979 (O_1979,N_20905,N_22326);
xnor UO_1980 (O_1980,N_22694,N_23288);
nor UO_1981 (O_1981,N_21659,N_22544);
or UO_1982 (O_1982,N_21654,N_20238);
or UO_1983 (O_1983,N_22841,N_24623);
nand UO_1984 (O_1984,N_23057,N_23765);
nand UO_1985 (O_1985,N_21028,N_24589);
and UO_1986 (O_1986,N_20881,N_21923);
or UO_1987 (O_1987,N_24299,N_21900);
and UO_1988 (O_1988,N_23801,N_22192);
nand UO_1989 (O_1989,N_22719,N_22932);
xnor UO_1990 (O_1990,N_21396,N_23995);
or UO_1991 (O_1991,N_24998,N_21984);
xor UO_1992 (O_1992,N_23376,N_24288);
nor UO_1993 (O_1993,N_23083,N_23931);
nor UO_1994 (O_1994,N_23197,N_22186);
or UO_1995 (O_1995,N_20825,N_24821);
nand UO_1996 (O_1996,N_22167,N_21884);
xor UO_1997 (O_1997,N_20586,N_22383);
nand UO_1998 (O_1998,N_21461,N_22392);
xor UO_1999 (O_1999,N_21657,N_21757);
nor UO_2000 (O_2000,N_23517,N_21632);
or UO_2001 (O_2001,N_23173,N_22906);
and UO_2002 (O_2002,N_22529,N_22844);
xnor UO_2003 (O_2003,N_21392,N_22683);
xor UO_2004 (O_2004,N_20275,N_20800);
nor UO_2005 (O_2005,N_22029,N_22017);
nor UO_2006 (O_2006,N_20353,N_21526);
nor UO_2007 (O_2007,N_22591,N_23863);
or UO_2008 (O_2008,N_21542,N_23293);
or UO_2009 (O_2009,N_23149,N_24038);
xor UO_2010 (O_2010,N_24592,N_24970);
xnor UO_2011 (O_2011,N_20727,N_20022);
nand UO_2012 (O_2012,N_24989,N_21347);
and UO_2013 (O_2013,N_22034,N_24078);
and UO_2014 (O_2014,N_20135,N_22040);
xnor UO_2015 (O_2015,N_24914,N_21030);
nor UO_2016 (O_2016,N_20573,N_21003);
nor UO_2017 (O_2017,N_21060,N_23467);
xnor UO_2018 (O_2018,N_24565,N_21087);
xnor UO_2019 (O_2019,N_21908,N_23186);
or UO_2020 (O_2020,N_23671,N_21344);
and UO_2021 (O_2021,N_23819,N_22928);
nand UO_2022 (O_2022,N_20776,N_23523);
nand UO_2023 (O_2023,N_24958,N_22219);
xor UO_2024 (O_2024,N_22580,N_21766);
nor UO_2025 (O_2025,N_24057,N_22917);
nor UO_2026 (O_2026,N_22832,N_22469);
or UO_2027 (O_2027,N_21823,N_22681);
xor UO_2028 (O_2028,N_20767,N_20049);
nand UO_2029 (O_2029,N_20590,N_20766);
nor UO_2030 (O_2030,N_21610,N_20074);
nor UO_2031 (O_2031,N_20428,N_22984);
nor UO_2032 (O_2032,N_22087,N_20578);
and UO_2033 (O_2033,N_21115,N_22870);
nand UO_2034 (O_2034,N_21491,N_22673);
nand UO_2035 (O_2035,N_24441,N_24492);
and UO_2036 (O_2036,N_24957,N_24020);
and UO_2037 (O_2037,N_20791,N_22996);
and UO_2038 (O_2038,N_21824,N_22686);
or UO_2039 (O_2039,N_21276,N_22537);
nor UO_2040 (O_2040,N_20615,N_23154);
nor UO_2041 (O_2041,N_22710,N_20807);
nor UO_2042 (O_2042,N_24981,N_24903);
and UO_2043 (O_2043,N_21096,N_20338);
or UO_2044 (O_2044,N_20719,N_22376);
nand UO_2045 (O_2045,N_23285,N_20816);
xor UO_2046 (O_2046,N_22324,N_21806);
or UO_2047 (O_2047,N_24745,N_24824);
xor UO_2048 (O_2048,N_24582,N_24466);
or UO_2049 (O_2049,N_22201,N_22067);
nor UO_2050 (O_2050,N_24089,N_20123);
and UO_2051 (O_2051,N_22748,N_23711);
or UO_2052 (O_2052,N_20456,N_21650);
or UO_2053 (O_2053,N_20170,N_21418);
or UO_2054 (O_2054,N_22306,N_24595);
nor UO_2055 (O_2055,N_23731,N_20975);
nand UO_2056 (O_2056,N_23515,N_23958);
or UO_2057 (O_2057,N_21902,N_22660);
and UO_2058 (O_2058,N_23143,N_22914);
and UO_2059 (O_2059,N_20213,N_20208);
xnor UO_2060 (O_2060,N_22340,N_24066);
nand UO_2061 (O_2061,N_20898,N_23384);
xnor UO_2062 (O_2062,N_20296,N_22788);
nor UO_2063 (O_2063,N_24204,N_23437);
nor UO_2064 (O_2064,N_22658,N_24956);
nor UO_2065 (O_2065,N_24546,N_24754);
xor UO_2066 (O_2066,N_23326,N_20871);
nor UO_2067 (O_2067,N_21399,N_23044);
xnor UO_2068 (O_2068,N_24973,N_24932);
and UO_2069 (O_2069,N_24625,N_23876);
nand UO_2070 (O_2070,N_23226,N_21051);
xor UO_2071 (O_2071,N_21057,N_24154);
nand UO_2072 (O_2072,N_20909,N_21797);
and UO_2073 (O_2073,N_24680,N_24647);
nand UO_2074 (O_2074,N_24952,N_22915);
xor UO_2075 (O_2075,N_23689,N_24665);
and UO_2076 (O_2076,N_20341,N_22499);
and UO_2077 (O_2077,N_22799,N_21285);
or UO_2078 (O_2078,N_24001,N_24075);
xnor UO_2079 (O_2079,N_21619,N_24276);
and UO_2080 (O_2080,N_23630,N_20165);
or UO_2081 (O_2081,N_23184,N_22670);
nand UO_2082 (O_2082,N_22736,N_23256);
xnor UO_2083 (O_2083,N_24405,N_24796);
or UO_2084 (O_2084,N_21848,N_23521);
xnor UO_2085 (O_2085,N_23320,N_23811);
and UO_2086 (O_2086,N_21181,N_20140);
nor UO_2087 (O_2087,N_20066,N_21449);
nand UO_2088 (O_2088,N_22330,N_24080);
or UO_2089 (O_2089,N_22153,N_21207);
and UO_2090 (O_2090,N_20454,N_21709);
nor UO_2091 (O_2091,N_23000,N_24165);
xnor UO_2092 (O_2092,N_21509,N_21514);
and UO_2093 (O_2093,N_24776,N_22292);
nand UO_2094 (O_2094,N_22175,N_23851);
nand UO_2095 (O_2095,N_20431,N_21987);
xnor UO_2096 (O_2096,N_22743,N_24268);
and UO_2097 (O_2097,N_21000,N_22423);
xnor UO_2098 (O_2098,N_23503,N_22682);
nand UO_2099 (O_2099,N_24831,N_24282);
nand UO_2100 (O_2100,N_23495,N_21886);
and UO_2101 (O_2101,N_21937,N_21221);
nor UO_2102 (O_2102,N_23845,N_24205);
and UO_2103 (O_2103,N_23993,N_22184);
and UO_2104 (O_2104,N_21649,N_21537);
nand UO_2105 (O_2105,N_21059,N_24523);
xor UO_2106 (O_2106,N_23405,N_21192);
xor UO_2107 (O_2107,N_21780,N_20201);
or UO_2108 (O_2108,N_22977,N_21021);
and UO_2109 (O_2109,N_21973,N_22631);
xor UO_2110 (O_2110,N_24509,N_23385);
or UO_2111 (O_2111,N_24010,N_24918);
and UO_2112 (O_2112,N_23305,N_20762);
xnor UO_2113 (O_2113,N_21244,N_21455);
xnor UO_2114 (O_2114,N_24208,N_23759);
nand UO_2115 (O_2115,N_20155,N_20445);
xor UO_2116 (O_2116,N_22181,N_22920);
nor UO_2117 (O_2117,N_22639,N_22221);
nand UO_2118 (O_2118,N_20215,N_21255);
and UO_2119 (O_2119,N_22532,N_22380);
nor UO_2120 (O_2120,N_24317,N_23162);
and UO_2121 (O_2121,N_20126,N_24607);
nor UO_2122 (O_2122,N_23303,N_23114);
nor UO_2123 (O_2123,N_21494,N_22838);
or UO_2124 (O_2124,N_23457,N_21327);
nor UO_2125 (O_2125,N_22690,N_24863);
xor UO_2126 (O_2126,N_24245,N_23386);
or UO_2127 (O_2127,N_23364,N_22105);
or UO_2128 (O_2128,N_21943,N_24415);
and UO_2129 (O_2129,N_20973,N_20511);
nor UO_2130 (O_2130,N_22885,N_24247);
nor UO_2131 (O_2131,N_22442,N_23712);
xnor UO_2132 (O_2132,N_22055,N_20604);
or UO_2133 (O_2133,N_23512,N_24050);
and UO_2134 (O_2134,N_21062,N_20489);
xor UO_2135 (O_2135,N_22038,N_21454);
or UO_2136 (O_2136,N_24178,N_23003);
nor UO_2137 (O_2137,N_24024,N_24873);
and UO_2138 (O_2138,N_24736,N_20625);
xor UO_2139 (O_2139,N_20947,N_21978);
nand UO_2140 (O_2140,N_24765,N_24273);
nand UO_2141 (O_2141,N_24322,N_22320);
or UO_2142 (O_2142,N_20012,N_21475);
nor UO_2143 (O_2143,N_20175,N_20530);
xnor UO_2144 (O_2144,N_24248,N_23938);
xnor UO_2145 (O_2145,N_22479,N_24350);
nand UO_2146 (O_2146,N_24329,N_20720);
and UO_2147 (O_2147,N_23311,N_21406);
and UO_2148 (O_2148,N_24637,N_23163);
nor UO_2149 (O_2149,N_23046,N_20080);
and UO_2150 (O_2150,N_22264,N_20710);
nor UO_2151 (O_2151,N_24556,N_21906);
xnor UO_2152 (O_2152,N_23458,N_20173);
xor UO_2153 (O_2153,N_24272,N_23700);
xor UO_2154 (O_2154,N_20894,N_22243);
and UO_2155 (O_2155,N_22912,N_22864);
and UO_2156 (O_2156,N_24624,N_24158);
or UO_2157 (O_2157,N_22173,N_20195);
nand UO_2158 (O_2158,N_23767,N_24975);
nor UO_2159 (O_2159,N_23810,N_23403);
nor UO_2160 (O_2160,N_20579,N_20017);
and UO_2161 (O_2161,N_22939,N_23764);
xor UO_2162 (O_2162,N_24708,N_24035);
nand UO_2163 (O_2163,N_22685,N_20193);
nor UO_2164 (O_2164,N_21077,N_24835);
nand UO_2165 (O_2165,N_23112,N_22245);
and UO_2166 (O_2166,N_23462,N_22513);
or UO_2167 (O_2167,N_21499,N_22652);
nor UO_2168 (O_2168,N_22738,N_24692);
nand UO_2169 (O_2169,N_21427,N_21297);
or UO_2170 (O_2170,N_24088,N_20284);
nor UO_2171 (O_2171,N_22750,N_20228);
nor UO_2172 (O_2172,N_21041,N_23009);
nand UO_2173 (O_2173,N_24480,N_22629);
nor UO_2174 (O_2174,N_20430,N_24908);
or UO_2175 (O_2175,N_23632,N_21642);
xor UO_2176 (O_2176,N_22158,N_23861);
or UO_2177 (O_2177,N_20078,N_21857);
and UO_2178 (O_2178,N_22542,N_23539);
or UO_2179 (O_2179,N_24160,N_21366);
or UO_2180 (O_2180,N_21124,N_21885);
or UO_2181 (O_2181,N_20651,N_21675);
nor UO_2182 (O_2182,N_24242,N_22866);
nand UO_2183 (O_2183,N_21247,N_21249);
xor UO_2184 (O_2184,N_21812,N_20669);
nor UO_2185 (O_2185,N_20427,N_21864);
nand UO_2186 (O_2186,N_20908,N_23001);
nor UO_2187 (O_2187,N_20189,N_23257);
and UO_2188 (O_2188,N_24614,N_22989);
nor UO_2189 (O_2189,N_21433,N_22332);
xor UO_2190 (O_2190,N_20488,N_20550);
or UO_2191 (O_2191,N_24439,N_21599);
nand UO_2192 (O_2192,N_24030,N_21953);
nor UO_2193 (O_2193,N_22481,N_20592);
nand UO_2194 (O_2194,N_24151,N_22887);
xnor UO_2195 (O_2195,N_24017,N_24356);
nand UO_2196 (O_2196,N_20419,N_24710);
nand UO_2197 (O_2197,N_22407,N_21252);
and UO_2198 (O_2198,N_21687,N_20141);
nand UO_2199 (O_2199,N_20706,N_21646);
or UO_2200 (O_2200,N_22805,N_20159);
nand UO_2201 (O_2201,N_21292,N_24300);
nand UO_2202 (O_2202,N_20537,N_20585);
xnor UO_2203 (O_2203,N_22012,N_21748);
nor UO_2204 (O_2204,N_23862,N_23417);
or UO_2205 (O_2205,N_23460,N_24068);
and UO_2206 (O_2206,N_23611,N_21855);
or UO_2207 (O_2207,N_21971,N_23773);
xnor UO_2208 (O_2208,N_24113,N_21972);
nor UO_2209 (O_2209,N_24095,N_20172);
and UO_2210 (O_2210,N_22746,N_20513);
nor UO_2211 (O_2211,N_20852,N_24476);
and UO_2212 (O_2212,N_24259,N_20399);
nor UO_2213 (O_2213,N_23022,N_24224);
nor UO_2214 (O_2214,N_20047,N_20931);
nor UO_2215 (O_2215,N_24675,N_21275);
xnor UO_2216 (O_2216,N_20668,N_24275);
nor UO_2217 (O_2217,N_24891,N_22817);
xnor UO_2218 (O_2218,N_23428,N_22378);
xor UO_2219 (O_2219,N_21861,N_21260);
and UO_2220 (O_2220,N_22951,N_20205);
nand UO_2221 (O_2221,N_21596,N_22894);
and UO_2222 (O_2222,N_20949,N_21217);
or UO_2223 (O_2223,N_23541,N_23722);
and UO_2224 (O_2224,N_22253,N_24354);
or UO_2225 (O_2225,N_24834,N_22956);
or UO_2226 (O_2226,N_22337,N_20413);
nor UO_2227 (O_2227,N_23021,N_23623);
and UO_2228 (O_2228,N_21046,N_23015);
or UO_2229 (O_2229,N_20944,N_24209);
nor UO_2230 (O_2230,N_21448,N_23172);
or UO_2231 (O_2231,N_22393,N_21145);
or UO_2232 (O_2232,N_24967,N_23620);
or UO_2233 (O_2233,N_24499,N_20890);
xor UO_2234 (O_2234,N_20874,N_24352);
or UO_2235 (O_2235,N_22521,N_24203);
nor UO_2236 (O_2236,N_22601,N_22628);
or UO_2237 (O_2237,N_22433,N_23537);
nand UO_2238 (O_2238,N_21541,N_22938);
xor UO_2239 (O_2239,N_20541,N_23490);
or UO_2240 (O_2240,N_20207,N_22006);
xnor UO_2241 (O_2241,N_24261,N_22848);
xnor UO_2242 (O_2242,N_20595,N_24836);
and UO_2243 (O_2243,N_23357,N_21483);
nand UO_2244 (O_2244,N_23625,N_20468);
or UO_2245 (O_2245,N_20678,N_22572);
and UO_2246 (O_2246,N_23838,N_22972);
and UO_2247 (O_2247,N_21422,N_21521);
nand UO_2248 (O_2248,N_23686,N_23968);
and UO_2249 (O_2249,N_22752,N_23854);
or UO_2250 (O_2250,N_23130,N_22934);
nor UO_2251 (O_2251,N_20831,N_21912);
nor UO_2252 (O_2252,N_24827,N_23146);
nand UO_2253 (O_2253,N_22833,N_20901);
or UO_2254 (O_2254,N_20304,N_21153);
or UO_2255 (O_2255,N_24574,N_21349);
nand UO_2256 (O_2256,N_24206,N_24983);
or UO_2257 (O_2257,N_24585,N_23637);
and UO_2258 (O_2258,N_24194,N_24712);
xor UO_2259 (O_2259,N_21996,N_21310);
nor UO_2260 (O_2260,N_22693,N_24522);
and UO_2261 (O_2261,N_23487,N_21866);
or UO_2262 (O_2262,N_21904,N_21256);
xnor UO_2263 (O_2263,N_20369,N_21601);
or UO_2264 (O_2264,N_23598,N_23269);
xor UO_2265 (O_2265,N_23766,N_21172);
nand UO_2266 (O_2266,N_20112,N_20935);
nand UO_2267 (O_2267,N_21997,N_23763);
nor UO_2268 (O_2268,N_23527,N_20648);
nor UO_2269 (O_2269,N_24528,N_24417);
and UO_2270 (O_2270,N_22418,N_22921);
nand UO_2271 (O_2271,N_20911,N_23006);
or UO_2272 (O_2272,N_23380,N_20665);
nor UO_2273 (O_2273,N_23672,N_20799);
nor UO_2274 (O_2274,N_24774,N_22554);
nor UO_2275 (O_2275,N_23281,N_24865);
and UO_2276 (O_2276,N_23776,N_20056);
nor UO_2277 (O_2277,N_20655,N_23651);
or UO_2278 (O_2278,N_23444,N_24598);
nor UO_2279 (O_2279,N_20357,N_21232);
nor UO_2280 (O_2280,N_23925,N_23497);
nand UO_2281 (O_2281,N_24741,N_23992);
nand UO_2282 (O_2282,N_20750,N_23050);
and UO_2283 (O_2283,N_21143,N_23084);
xnor UO_2284 (O_2284,N_21107,N_24302);
nand UO_2285 (O_2285,N_23250,N_24389);
nor UO_2286 (O_2286,N_22033,N_22346);
nand UO_2287 (O_2287,N_21880,N_20576);
or UO_2288 (O_2288,N_20040,N_23195);
xnor UO_2289 (O_2289,N_24539,N_21792);
and UO_2290 (O_2290,N_20783,N_20089);
xor UO_2291 (O_2291,N_23771,N_23841);
or UO_2292 (O_2292,N_22789,N_20637);
nor UO_2293 (O_2293,N_23761,N_24029);
or UO_2294 (O_2294,N_20638,N_21437);
xor UO_2295 (O_2295,N_21451,N_21928);
xor UO_2296 (O_2296,N_20561,N_22277);
and UO_2297 (O_2297,N_20255,N_20958);
xnor UO_2298 (O_2298,N_24635,N_24107);
or UO_2299 (O_2299,N_23805,N_21549);
nor UO_2300 (O_2300,N_21994,N_20996);
or UO_2301 (O_2301,N_23866,N_20034);
nand UO_2302 (O_2302,N_23744,N_21082);
xnor UO_2303 (O_2303,N_21872,N_21211);
or UO_2304 (O_2304,N_22108,N_23105);
and UO_2305 (O_2305,N_23734,N_20723);
nand UO_2306 (O_2306,N_22032,N_22134);
nor UO_2307 (O_2307,N_20865,N_24678);
xnor UO_2308 (O_2308,N_24169,N_21136);
and UO_2309 (O_2309,N_21151,N_22054);
nand UO_2310 (O_2310,N_20298,N_22343);
or UO_2311 (O_2311,N_23934,N_20408);
or UO_2312 (O_2312,N_21257,N_22000);
xor UO_2313 (O_2313,N_21611,N_20007);
xor UO_2314 (O_2314,N_20085,N_20115);
or UO_2315 (O_2315,N_23264,N_21609);
nor UO_2316 (O_2316,N_21644,N_23120);
xor UO_2317 (O_2317,N_21315,N_23905);
and UO_2318 (O_2318,N_20327,N_23058);
nand UO_2319 (O_2319,N_20998,N_23740);
xor UO_2320 (O_2320,N_23887,N_23572);
and UO_2321 (O_2321,N_24777,N_22611);
and UO_2322 (O_2322,N_21209,N_20779);
and UO_2323 (O_2323,N_20299,N_21429);
nor UO_2324 (O_2324,N_22007,N_20292);
nand UO_2325 (O_2325,N_24163,N_23471);
nor UO_2326 (O_2326,N_23282,N_24142);
nand UO_2327 (O_2327,N_22370,N_22025);
or UO_2328 (O_2328,N_22473,N_22699);
nand UO_2329 (O_2329,N_21843,N_23677);
and UO_2330 (O_2330,N_21808,N_22892);
and UO_2331 (O_2331,N_23451,N_24027);
xnor UO_2332 (O_2332,N_21111,N_21443);
xor UO_2333 (O_2333,N_23794,N_23133);
nor UO_2334 (O_2334,N_20840,N_21045);
xor UO_2335 (O_2335,N_21935,N_20449);
nor UO_2336 (O_2336,N_24366,N_20451);
and UO_2337 (O_2337,N_23504,N_23489);
nor UO_2338 (O_2338,N_21329,N_22643);
or UO_2339 (O_2339,N_20070,N_22118);
nand UO_2340 (O_2340,N_23170,N_24893);
xnor UO_2341 (O_2341,N_20384,N_21237);
xor UO_2342 (O_2342,N_24257,N_21554);
nand UO_2343 (O_2343,N_22516,N_22911);
xnor UO_2344 (O_2344,N_22641,N_20818);
or UO_2345 (O_2345,N_24347,N_23448);
nand UO_2346 (O_2346,N_22955,N_23589);
and UO_2347 (O_2347,N_21316,N_23638);
xor UO_2348 (O_2348,N_20051,N_23984);
and UO_2349 (O_2349,N_23063,N_23904);
xnor UO_2350 (O_2350,N_20914,N_24097);
nor UO_2351 (O_2351,N_22061,N_24788);
or UO_2352 (O_2352,N_22482,N_21495);
and UO_2353 (O_2353,N_20377,N_23660);
nor UO_2354 (O_2354,N_20919,N_21558);
xor UO_2355 (O_2355,N_24875,N_24783);
or UO_2356 (O_2356,N_22279,N_22913);
or UO_2357 (O_2357,N_20009,N_21270);
or UO_2358 (O_2358,N_20295,N_23928);
and UO_2359 (O_2359,N_23937,N_21034);
xnor UO_2360 (O_2360,N_24979,N_24723);
nand UO_2361 (O_2361,N_21183,N_20013);
and UO_2362 (O_2362,N_24368,N_23103);
nor UO_2363 (O_2363,N_20661,N_21934);
nor UO_2364 (O_2364,N_20042,N_21841);
xor UO_2365 (O_2365,N_20306,N_21006);
or UO_2366 (O_2366,N_20823,N_22589);
nand UO_2367 (O_2367,N_21647,N_20610);
nor UO_2368 (O_2368,N_22708,N_20851);
xor UO_2369 (O_2369,N_24153,N_21989);
and UO_2370 (O_2370,N_23259,N_22062);
nor UO_2371 (O_2371,N_23266,N_21768);
or UO_2372 (O_2372,N_20429,N_22868);
and UO_2373 (O_2373,N_24826,N_24934);
and UO_2374 (O_2374,N_22400,N_20226);
nand UO_2375 (O_2375,N_22287,N_23892);
xor UO_2376 (O_2376,N_24327,N_23148);
and UO_2377 (O_2377,N_22238,N_21661);
xor UO_2378 (O_2378,N_21109,N_23501);
or UO_2379 (O_2379,N_20930,N_21830);
and UO_2380 (O_2380,N_22797,N_22901);
nand UO_2381 (O_2381,N_20521,N_20539);
xor UO_2382 (O_2382,N_24111,N_24987);
nand UO_2383 (O_2383,N_24454,N_24563);
and UO_2384 (O_2384,N_20294,N_23528);
nor UO_2385 (O_2385,N_24428,N_23079);
and UO_2386 (O_2386,N_24239,N_22821);
and UO_2387 (O_2387,N_23783,N_23855);
nor UO_2388 (O_2388,N_23886,N_24586);
or UO_2389 (O_2389,N_20946,N_24198);
and UO_2390 (O_2390,N_24521,N_21913);
or UO_2391 (O_2391,N_21957,N_21720);
nor UO_2392 (O_2392,N_22950,N_21710);
and UO_2393 (O_2393,N_21803,N_21782);
and UO_2394 (O_2394,N_21393,N_24808);
and UO_2395 (O_2395,N_22028,N_20772);
nand UO_2396 (O_2396,N_23511,N_24552);
or UO_2397 (O_2397,N_21099,N_24561);
nand UO_2398 (O_2398,N_24087,N_22843);
nand UO_2399 (O_2399,N_22179,N_21336);
xor UO_2400 (O_2400,N_23675,N_23035);
nand UO_2401 (O_2401,N_21745,N_22248);
nor UO_2402 (O_2402,N_24148,N_23806);
and UO_2403 (O_2403,N_21026,N_21180);
or UO_2404 (O_2404,N_23865,N_22278);
or UO_2405 (O_2405,N_23155,N_22043);
and UO_2406 (O_2406,N_20789,N_21477);
or UO_2407 (O_2407,N_22701,N_23802);
nand UO_2408 (O_2408,N_24740,N_21504);
nor UO_2409 (O_2409,N_21732,N_23099);
nor UO_2410 (O_2410,N_22237,N_22526);
or UO_2411 (O_2411,N_24742,N_20664);
or UO_2412 (O_2412,N_23492,N_21189);
or UO_2413 (O_2413,N_23043,N_21191);
or UO_2414 (O_2414,N_22672,N_22360);
or UO_2415 (O_2415,N_21819,N_23418);
or UO_2416 (O_2416,N_22770,N_20697);
nand UO_2417 (O_2417,N_22494,N_21110);
and UO_2418 (O_2418,N_23260,N_23906);
and UO_2419 (O_2419,N_22903,N_23429);
or UO_2420 (O_2420,N_24429,N_21085);
nand UO_2421 (O_2421,N_22990,N_24128);
or UO_2422 (O_2422,N_21763,N_20412);
or UO_2423 (O_2423,N_22667,N_24800);
nand UO_2424 (O_2424,N_24296,N_23398);
nand UO_2425 (O_2425,N_23896,N_24946);
xor UO_2426 (O_2426,N_21185,N_21362);
nand UO_2427 (O_2427,N_22550,N_20752);
nor UO_2428 (O_2428,N_21802,N_21568);
xnor UO_2429 (O_2429,N_22372,N_24560);
nand UO_2430 (O_2430,N_21691,N_22813);
and UO_2431 (O_2431,N_23191,N_23977);
xor UO_2432 (O_2432,N_20522,N_22898);
nand UO_2433 (O_2433,N_24145,N_21039);
nor UO_2434 (O_2434,N_23337,N_21854);
nor UO_2435 (O_2435,N_22131,N_20945);
nand UO_2436 (O_2436,N_23071,N_24120);
nor UO_2437 (O_2437,N_21616,N_23869);
and UO_2438 (O_2438,N_21126,N_20325);
xnor UO_2439 (O_2439,N_24197,N_23323);
xor UO_2440 (O_2440,N_22114,N_21936);
and UO_2441 (O_2441,N_23908,N_23096);
and UO_2442 (O_2442,N_22534,N_21070);
xnor UO_2443 (O_2443,N_23339,N_23025);
or UO_2444 (O_2444,N_24059,N_24929);
nand UO_2445 (O_2445,N_20204,N_22319);
nand UO_2446 (O_2446,N_24847,N_20501);
or UO_2447 (O_2447,N_23434,N_20757);
nor UO_2448 (O_2448,N_22895,N_20966);
and UO_2449 (O_2449,N_21645,N_24880);
nand UO_2450 (O_2450,N_20139,N_24810);
nand UO_2451 (O_2451,N_24815,N_21795);
nand UO_2452 (O_2452,N_21438,N_21002);
xor UO_2453 (O_2453,N_22130,N_23073);
nand UO_2454 (O_2454,N_20176,N_22147);
nand UO_2455 (O_2455,N_23918,N_20127);
nor UO_2456 (O_2456,N_23959,N_24230);
nand UO_2457 (O_2457,N_21505,N_22185);
or UO_2458 (O_2458,N_22460,N_21919);
nor UO_2459 (O_2459,N_24411,N_20582);
or UO_2460 (O_2460,N_24668,N_22582);
nand UO_2461 (O_2461,N_20337,N_23081);
nor UO_2462 (O_2462,N_20855,N_20418);
nor UO_2463 (O_2463,N_21535,N_23754);
nand UO_2464 (O_2464,N_23561,N_20523);
and UO_2465 (O_2465,N_20955,N_20794);
or UO_2466 (O_2466,N_21212,N_24862);
nand UO_2467 (O_2467,N_20814,N_24830);
and UO_2468 (O_2468,N_22648,N_23750);
nand UO_2469 (O_2469,N_21326,N_21174);
nor UO_2470 (O_2470,N_22003,N_20689);
or UO_2471 (O_2471,N_23520,N_22583);
nor UO_2472 (O_2472,N_24813,N_21674);
nor UO_2473 (O_2473,N_24966,N_21995);
xor UO_2474 (O_2474,N_21580,N_20650);
or UO_2475 (O_2475,N_21202,N_23785);
or UO_2476 (O_2476,N_22974,N_23560);
nand UO_2477 (O_2477,N_24425,N_22644);
and UO_2478 (O_2478,N_22659,N_22080);
or UO_2479 (O_2479,N_22851,N_22632);
and UO_2480 (O_2480,N_23122,N_24964);
or UO_2481 (O_2481,N_22349,N_22993);
nand UO_2482 (O_2482,N_21985,N_22189);
nand UO_2483 (O_2483,N_22745,N_23247);
nand UO_2484 (O_2484,N_22492,N_24626);
nor UO_2485 (O_2485,N_22916,N_21652);
or UO_2486 (O_2486,N_23221,N_22758);
nand UO_2487 (O_2487,N_23587,N_22126);
nor UO_2488 (O_2488,N_21918,N_21029);
or UO_2489 (O_2489,N_24922,N_21825);
xor UO_2490 (O_2490,N_21954,N_20351);
nor UO_2491 (O_2491,N_22065,N_24342);
nand UO_2492 (O_2492,N_20694,N_20027);
nor UO_2493 (O_2493,N_21863,N_24076);
xor UO_2494 (O_2494,N_21607,N_22425);
xnor UO_2495 (O_2495,N_24040,N_24474);
and UO_2496 (O_2496,N_21955,N_20105);
nand UO_2497 (O_2497,N_22443,N_22435);
nand UO_2498 (O_2498,N_21828,N_23346);
nand UO_2499 (O_2499,N_22070,N_20364);
and UO_2500 (O_2500,N_23425,N_21543);
xor UO_2501 (O_2501,N_21548,N_21996);
nor UO_2502 (O_2502,N_20987,N_22219);
or UO_2503 (O_2503,N_20091,N_24120);
xor UO_2504 (O_2504,N_20401,N_24479);
nand UO_2505 (O_2505,N_20331,N_23551);
nor UO_2506 (O_2506,N_22672,N_24090);
nor UO_2507 (O_2507,N_21759,N_24544);
or UO_2508 (O_2508,N_20496,N_22520);
nor UO_2509 (O_2509,N_23116,N_24865);
and UO_2510 (O_2510,N_21214,N_24746);
or UO_2511 (O_2511,N_21645,N_23011);
or UO_2512 (O_2512,N_21197,N_24736);
nor UO_2513 (O_2513,N_23710,N_23881);
and UO_2514 (O_2514,N_22302,N_22776);
xnor UO_2515 (O_2515,N_23321,N_23679);
xnor UO_2516 (O_2516,N_24659,N_20323);
and UO_2517 (O_2517,N_20592,N_24677);
or UO_2518 (O_2518,N_22240,N_23479);
xor UO_2519 (O_2519,N_23755,N_24178);
nand UO_2520 (O_2520,N_22898,N_21378);
nand UO_2521 (O_2521,N_21660,N_21170);
xnor UO_2522 (O_2522,N_24525,N_21217);
nor UO_2523 (O_2523,N_22687,N_21685);
nand UO_2524 (O_2524,N_22258,N_21397);
xor UO_2525 (O_2525,N_24906,N_24400);
or UO_2526 (O_2526,N_23431,N_22297);
nor UO_2527 (O_2527,N_22751,N_20296);
xnor UO_2528 (O_2528,N_22551,N_23308);
nand UO_2529 (O_2529,N_21137,N_21415);
and UO_2530 (O_2530,N_24353,N_24659);
nand UO_2531 (O_2531,N_22856,N_23526);
or UO_2532 (O_2532,N_21657,N_23138);
xnor UO_2533 (O_2533,N_22911,N_21755);
or UO_2534 (O_2534,N_20583,N_23486);
nor UO_2535 (O_2535,N_20648,N_22058);
or UO_2536 (O_2536,N_20336,N_20086);
and UO_2537 (O_2537,N_20774,N_20535);
nand UO_2538 (O_2538,N_20979,N_22645);
or UO_2539 (O_2539,N_23442,N_23427);
nor UO_2540 (O_2540,N_23946,N_23231);
nand UO_2541 (O_2541,N_21141,N_20229);
xnor UO_2542 (O_2542,N_21681,N_24796);
and UO_2543 (O_2543,N_22059,N_20781);
nor UO_2544 (O_2544,N_22286,N_24718);
and UO_2545 (O_2545,N_21891,N_21185);
and UO_2546 (O_2546,N_24673,N_24604);
nor UO_2547 (O_2547,N_20834,N_24928);
or UO_2548 (O_2548,N_22869,N_23533);
nand UO_2549 (O_2549,N_24054,N_23629);
or UO_2550 (O_2550,N_21013,N_20277);
xor UO_2551 (O_2551,N_20938,N_24929);
nand UO_2552 (O_2552,N_23733,N_22895);
nor UO_2553 (O_2553,N_21285,N_24693);
nand UO_2554 (O_2554,N_22896,N_22781);
or UO_2555 (O_2555,N_23773,N_23736);
and UO_2556 (O_2556,N_23301,N_20935);
and UO_2557 (O_2557,N_24187,N_23678);
or UO_2558 (O_2558,N_24520,N_23890);
and UO_2559 (O_2559,N_23978,N_20827);
xnor UO_2560 (O_2560,N_23074,N_21088);
nor UO_2561 (O_2561,N_23798,N_22477);
nand UO_2562 (O_2562,N_23831,N_21072);
nor UO_2563 (O_2563,N_21655,N_20610);
and UO_2564 (O_2564,N_23561,N_20704);
and UO_2565 (O_2565,N_23025,N_24039);
nand UO_2566 (O_2566,N_23787,N_22472);
nand UO_2567 (O_2567,N_20480,N_20871);
nand UO_2568 (O_2568,N_20710,N_21618);
nor UO_2569 (O_2569,N_20230,N_24626);
nand UO_2570 (O_2570,N_21427,N_20189);
or UO_2571 (O_2571,N_23066,N_22925);
and UO_2572 (O_2572,N_23977,N_24726);
or UO_2573 (O_2573,N_23674,N_23213);
or UO_2574 (O_2574,N_23014,N_22356);
and UO_2575 (O_2575,N_22008,N_21618);
and UO_2576 (O_2576,N_24982,N_22299);
and UO_2577 (O_2577,N_23343,N_24886);
or UO_2578 (O_2578,N_24663,N_22535);
nor UO_2579 (O_2579,N_23084,N_23149);
or UO_2580 (O_2580,N_23943,N_23196);
xnor UO_2581 (O_2581,N_24875,N_20162);
xor UO_2582 (O_2582,N_20559,N_21957);
xor UO_2583 (O_2583,N_24540,N_21649);
nand UO_2584 (O_2584,N_21248,N_21028);
and UO_2585 (O_2585,N_21756,N_24925);
nand UO_2586 (O_2586,N_24326,N_20906);
nor UO_2587 (O_2587,N_22359,N_21378);
nor UO_2588 (O_2588,N_20758,N_22264);
xor UO_2589 (O_2589,N_23003,N_21348);
and UO_2590 (O_2590,N_22196,N_21927);
nor UO_2591 (O_2591,N_22342,N_24151);
nand UO_2592 (O_2592,N_24934,N_21879);
and UO_2593 (O_2593,N_23966,N_21042);
or UO_2594 (O_2594,N_24164,N_23770);
and UO_2595 (O_2595,N_20742,N_22807);
or UO_2596 (O_2596,N_22326,N_23029);
nand UO_2597 (O_2597,N_23783,N_23902);
nor UO_2598 (O_2598,N_24202,N_24569);
xnor UO_2599 (O_2599,N_24247,N_23086);
or UO_2600 (O_2600,N_24328,N_23019);
nand UO_2601 (O_2601,N_20535,N_20039);
or UO_2602 (O_2602,N_20564,N_21576);
and UO_2603 (O_2603,N_23582,N_23841);
xor UO_2604 (O_2604,N_20284,N_21890);
nand UO_2605 (O_2605,N_21388,N_24970);
or UO_2606 (O_2606,N_23314,N_20005);
xor UO_2607 (O_2607,N_20233,N_21177);
nand UO_2608 (O_2608,N_22725,N_20541);
and UO_2609 (O_2609,N_20147,N_23629);
and UO_2610 (O_2610,N_22680,N_24374);
and UO_2611 (O_2611,N_20831,N_23584);
xor UO_2612 (O_2612,N_24934,N_20026);
nor UO_2613 (O_2613,N_22202,N_24026);
nor UO_2614 (O_2614,N_24536,N_23287);
nor UO_2615 (O_2615,N_20064,N_21746);
nor UO_2616 (O_2616,N_24886,N_22408);
nor UO_2617 (O_2617,N_23151,N_23699);
nand UO_2618 (O_2618,N_20595,N_24059);
nand UO_2619 (O_2619,N_23590,N_24859);
or UO_2620 (O_2620,N_23251,N_21927);
or UO_2621 (O_2621,N_21682,N_23998);
and UO_2622 (O_2622,N_22160,N_24400);
and UO_2623 (O_2623,N_21525,N_23769);
xnor UO_2624 (O_2624,N_23157,N_20729);
nand UO_2625 (O_2625,N_23804,N_22611);
or UO_2626 (O_2626,N_24802,N_24124);
or UO_2627 (O_2627,N_24719,N_23585);
nand UO_2628 (O_2628,N_23073,N_21261);
or UO_2629 (O_2629,N_21384,N_20180);
nand UO_2630 (O_2630,N_23022,N_22504);
nand UO_2631 (O_2631,N_23337,N_24992);
or UO_2632 (O_2632,N_21672,N_23481);
nand UO_2633 (O_2633,N_22009,N_23480);
nor UO_2634 (O_2634,N_20365,N_20779);
or UO_2635 (O_2635,N_22497,N_22868);
xor UO_2636 (O_2636,N_20576,N_24033);
and UO_2637 (O_2637,N_20749,N_20775);
nand UO_2638 (O_2638,N_20920,N_23067);
xor UO_2639 (O_2639,N_20041,N_20817);
or UO_2640 (O_2640,N_23089,N_24762);
nand UO_2641 (O_2641,N_20644,N_23536);
nand UO_2642 (O_2642,N_23709,N_20930);
or UO_2643 (O_2643,N_22405,N_22693);
nor UO_2644 (O_2644,N_23616,N_21307);
and UO_2645 (O_2645,N_20638,N_20851);
xnor UO_2646 (O_2646,N_22077,N_22337);
xor UO_2647 (O_2647,N_23833,N_24070);
xor UO_2648 (O_2648,N_23006,N_22414);
nand UO_2649 (O_2649,N_21129,N_20085);
nor UO_2650 (O_2650,N_23258,N_20993);
nand UO_2651 (O_2651,N_24491,N_21499);
nor UO_2652 (O_2652,N_21500,N_22432);
xor UO_2653 (O_2653,N_20496,N_21298);
or UO_2654 (O_2654,N_20028,N_23881);
and UO_2655 (O_2655,N_23270,N_20155);
nand UO_2656 (O_2656,N_24955,N_21281);
nand UO_2657 (O_2657,N_23474,N_22521);
xnor UO_2658 (O_2658,N_21664,N_20202);
xor UO_2659 (O_2659,N_20303,N_21721);
xnor UO_2660 (O_2660,N_23886,N_20635);
and UO_2661 (O_2661,N_23776,N_20971);
xor UO_2662 (O_2662,N_23979,N_24682);
and UO_2663 (O_2663,N_24265,N_24558);
nand UO_2664 (O_2664,N_20519,N_22360);
or UO_2665 (O_2665,N_23124,N_23079);
xor UO_2666 (O_2666,N_22129,N_20823);
nand UO_2667 (O_2667,N_24866,N_20574);
and UO_2668 (O_2668,N_23667,N_23814);
xnor UO_2669 (O_2669,N_24476,N_22288);
xnor UO_2670 (O_2670,N_24868,N_20081);
nand UO_2671 (O_2671,N_21144,N_20549);
or UO_2672 (O_2672,N_24497,N_23944);
nand UO_2673 (O_2673,N_20804,N_24447);
nor UO_2674 (O_2674,N_21534,N_24026);
and UO_2675 (O_2675,N_21364,N_23961);
and UO_2676 (O_2676,N_20131,N_20339);
nor UO_2677 (O_2677,N_24559,N_21492);
or UO_2678 (O_2678,N_22587,N_24774);
or UO_2679 (O_2679,N_20697,N_22570);
nor UO_2680 (O_2680,N_22304,N_22051);
and UO_2681 (O_2681,N_24287,N_20760);
or UO_2682 (O_2682,N_23157,N_24976);
and UO_2683 (O_2683,N_24393,N_24478);
or UO_2684 (O_2684,N_20698,N_20846);
xor UO_2685 (O_2685,N_20400,N_21316);
nand UO_2686 (O_2686,N_20544,N_22714);
xnor UO_2687 (O_2687,N_22082,N_22627);
nor UO_2688 (O_2688,N_21302,N_21954);
xor UO_2689 (O_2689,N_21224,N_22824);
xnor UO_2690 (O_2690,N_20753,N_23492);
xor UO_2691 (O_2691,N_20810,N_24343);
or UO_2692 (O_2692,N_22318,N_23269);
xor UO_2693 (O_2693,N_22871,N_21413);
or UO_2694 (O_2694,N_21041,N_20945);
nand UO_2695 (O_2695,N_23449,N_24972);
nand UO_2696 (O_2696,N_21508,N_24951);
xor UO_2697 (O_2697,N_23182,N_21357);
and UO_2698 (O_2698,N_24662,N_21439);
and UO_2699 (O_2699,N_22410,N_24363);
nand UO_2700 (O_2700,N_24136,N_23601);
or UO_2701 (O_2701,N_20585,N_24512);
xnor UO_2702 (O_2702,N_22547,N_23827);
and UO_2703 (O_2703,N_23049,N_22715);
or UO_2704 (O_2704,N_24429,N_21845);
and UO_2705 (O_2705,N_20701,N_24600);
nor UO_2706 (O_2706,N_22654,N_20657);
xor UO_2707 (O_2707,N_24122,N_20565);
or UO_2708 (O_2708,N_23579,N_21918);
or UO_2709 (O_2709,N_20084,N_23448);
xor UO_2710 (O_2710,N_24335,N_22520);
nor UO_2711 (O_2711,N_21157,N_21021);
and UO_2712 (O_2712,N_22837,N_22450);
xor UO_2713 (O_2713,N_23335,N_24566);
and UO_2714 (O_2714,N_24427,N_23206);
xor UO_2715 (O_2715,N_21643,N_21123);
nor UO_2716 (O_2716,N_21973,N_23193);
nand UO_2717 (O_2717,N_21297,N_24935);
or UO_2718 (O_2718,N_22910,N_22943);
or UO_2719 (O_2719,N_24512,N_23832);
nand UO_2720 (O_2720,N_24193,N_20132);
and UO_2721 (O_2721,N_23254,N_22128);
and UO_2722 (O_2722,N_20656,N_22466);
xor UO_2723 (O_2723,N_24876,N_20852);
nand UO_2724 (O_2724,N_21246,N_23153);
nand UO_2725 (O_2725,N_20471,N_21621);
xnor UO_2726 (O_2726,N_20442,N_23748);
and UO_2727 (O_2727,N_21000,N_23128);
xor UO_2728 (O_2728,N_21147,N_20324);
nand UO_2729 (O_2729,N_23461,N_20936);
nand UO_2730 (O_2730,N_22386,N_20298);
xor UO_2731 (O_2731,N_21549,N_24039);
nand UO_2732 (O_2732,N_20065,N_22186);
xor UO_2733 (O_2733,N_23593,N_23938);
nor UO_2734 (O_2734,N_24341,N_22366);
nor UO_2735 (O_2735,N_21818,N_21084);
nand UO_2736 (O_2736,N_21497,N_20543);
nor UO_2737 (O_2737,N_20470,N_23264);
nor UO_2738 (O_2738,N_24007,N_24718);
nor UO_2739 (O_2739,N_21701,N_21956);
nor UO_2740 (O_2740,N_23140,N_21340);
nand UO_2741 (O_2741,N_22638,N_22326);
xor UO_2742 (O_2742,N_22007,N_22227);
nand UO_2743 (O_2743,N_22762,N_20514);
and UO_2744 (O_2744,N_20239,N_20942);
and UO_2745 (O_2745,N_22067,N_20770);
nand UO_2746 (O_2746,N_23737,N_22877);
nand UO_2747 (O_2747,N_23550,N_21471);
xor UO_2748 (O_2748,N_21884,N_21861);
nor UO_2749 (O_2749,N_24559,N_23682);
and UO_2750 (O_2750,N_20038,N_24639);
and UO_2751 (O_2751,N_24284,N_24412);
and UO_2752 (O_2752,N_24527,N_24054);
nand UO_2753 (O_2753,N_20624,N_23199);
and UO_2754 (O_2754,N_21106,N_21037);
and UO_2755 (O_2755,N_24498,N_24478);
and UO_2756 (O_2756,N_20572,N_23622);
and UO_2757 (O_2757,N_20145,N_20282);
or UO_2758 (O_2758,N_24054,N_22856);
xnor UO_2759 (O_2759,N_24603,N_21730);
nand UO_2760 (O_2760,N_20165,N_21092);
and UO_2761 (O_2761,N_21447,N_24227);
or UO_2762 (O_2762,N_20403,N_24130);
and UO_2763 (O_2763,N_22890,N_20437);
and UO_2764 (O_2764,N_21051,N_21587);
xor UO_2765 (O_2765,N_22205,N_23925);
nand UO_2766 (O_2766,N_23041,N_20044);
or UO_2767 (O_2767,N_21440,N_23807);
nor UO_2768 (O_2768,N_24084,N_21572);
nor UO_2769 (O_2769,N_21224,N_23803);
or UO_2770 (O_2770,N_21533,N_24282);
and UO_2771 (O_2771,N_23070,N_20542);
xor UO_2772 (O_2772,N_21762,N_24303);
and UO_2773 (O_2773,N_22176,N_22361);
nor UO_2774 (O_2774,N_22046,N_23350);
and UO_2775 (O_2775,N_20551,N_20713);
and UO_2776 (O_2776,N_24818,N_23732);
xor UO_2777 (O_2777,N_22348,N_24491);
nor UO_2778 (O_2778,N_23943,N_20491);
or UO_2779 (O_2779,N_20434,N_23457);
xor UO_2780 (O_2780,N_22336,N_23810);
xor UO_2781 (O_2781,N_22899,N_22308);
nor UO_2782 (O_2782,N_22737,N_21742);
nor UO_2783 (O_2783,N_21128,N_22167);
nor UO_2784 (O_2784,N_22693,N_21099);
or UO_2785 (O_2785,N_22717,N_23459);
xnor UO_2786 (O_2786,N_23083,N_24760);
or UO_2787 (O_2787,N_20524,N_20200);
or UO_2788 (O_2788,N_23878,N_24779);
or UO_2789 (O_2789,N_21242,N_20722);
and UO_2790 (O_2790,N_22571,N_24424);
nor UO_2791 (O_2791,N_22139,N_23468);
and UO_2792 (O_2792,N_22236,N_23233);
nor UO_2793 (O_2793,N_21417,N_23660);
xor UO_2794 (O_2794,N_22054,N_21729);
or UO_2795 (O_2795,N_24625,N_21283);
nor UO_2796 (O_2796,N_22887,N_21164);
nor UO_2797 (O_2797,N_22615,N_24476);
or UO_2798 (O_2798,N_20514,N_21506);
nor UO_2799 (O_2799,N_23063,N_23092);
xor UO_2800 (O_2800,N_22307,N_24856);
or UO_2801 (O_2801,N_20645,N_20342);
or UO_2802 (O_2802,N_23060,N_22579);
nor UO_2803 (O_2803,N_23007,N_22770);
and UO_2804 (O_2804,N_24356,N_23542);
nor UO_2805 (O_2805,N_24571,N_23923);
xor UO_2806 (O_2806,N_24452,N_23344);
nor UO_2807 (O_2807,N_21334,N_21603);
and UO_2808 (O_2808,N_20572,N_21486);
nor UO_2809 (O_2809,N_24131,N_20767);
and UO_2810 (O_2810,N_20555,N_21432);
or UO_2811 (O_2811,N_20033,N_24403);
and UO_2812 (O_2812,N_22934,N_24885);
nor UO_2813 (O_2813,N_24141,N_20517);
or UO_2814 (O_2814,N_22733,N_20354);
and UO_2815 (O_2815,N_20119,N_20011);
nand UO_2816 (O_2816,N_23622,N_21319);
xnor UO_2817 (O_2817,N_21943,N_23282);
nand UO_2818 (O_2818,N_24151,N_24876);
xnor UO_2819 (O_2819,N_21497,N_22551);
or UO_2820 (O_2820,N_22131,N_21969);
nor UO_2821 (O_2821,N_24192,N_22373);
or UO_2822 (O_2822,N_20939,N_23955);
nor UO_2823 (O_2823,N_24968,N_21049);
nor UO_2824 (O_2824,N_20255,N_22262);
and UO_2825 (O_2825,N_21222,N_23352);
nor UO_2826 (O_2826,N_22692,N_22217);
and UO_2827 (O_2827,N_21869,N_21940);
nand UO_2828 (O_2828,N_23038,N_22174);
and UO_2829 (O_2829,N_24567,N_23763);
nor UO_2830 (O_2830,N_21834,N_23035);
and UO_2831 (O_2831,N_23907,N_23486);
or UO_2832 (O_2832,N_23464,N_23637);
nor UO_2833 (O_2833,N_22440,N_20247);
nand UO_2834 (O_2834,N_24365,N_23094);
nor UO_2835 (O_2835,N_20289,N_24236);
xnor UO_2836 (O_2836,N_23994,N_24424);
nand UO_2837 (O_2837,N_24853,N_21184);
or UO_2838 (O_2838,N_23292,N_21742);
nand UO_2839 (O_2839,N_22996,N_21146);
nor UO_2840 (O_2840,N_23984,N_23567);
and UO_2841 (O_2841,N_24557,N_20856);
or UO_2842 (O_2842,N_21518,N_22163);
or UO_2843 (O_2843,N_20867,N_22885);
and UO_2844 (O_2844,N_24010,N_21838);
nand UO_2845 (O_2845,N_21948,N_20392);
xor UO_2846 (O_2846,N_20808,N_23907);
nand UO_2847 (O_2847,N_21667,N_21508);
and UO_2848 (O_2848,N_23296,N_23112);
nor UO_2849 (O_2849,N_20730,N_22399);
nor UO_2850 (O_2850,N_21985,N_20823);
and UO_2851 (O_2851,N_24339,N_21259);
nor UO_2852 (O_2852,N_20536,N_20631);
nor UO_2853 (O_2853,N_22633,N_22813);
or UO_2854 (O_2854,N_20181,N_24862);
and UO_2855 (O_2855,N_23798,N_20293);
nor UO_2856 (O_2856,N_21179,N_22113);
xnor UO_2857 (O_2857,N_24318,N_21353);
xnor UO_2858 (O_2858,N_23534,N_23483);
or UO_2859 (O_2859,N_23358,N_22043);
or UO_2860 (O_2860,N_24407,N_20120);
xor UO_2861 (O_2861,N_20161,N_21219);
nor UO_2862 (O_2862,N_20104,N_23362);
or UO_2863 (O_2863,N_23852,N_24737);
and UO_2864 (O_2864,N_24387,N_22785);
or UO_2865 (O_2865,N_20495,N_21761);
nand UO_2866 (O_2866,N_23312,N_23511);
nand UO_2867 (O_2867,N_24905,N_22501);
xnor UO_2868 (O_2868,N_23184,N_20760);
or UO_2869 (O_2869,N_24617,N_21011);
nand UO_2870 (O_2870,N_24252,N_22582);
and UO_2871 (O_2871,N_23463,N_24453);
nor UO_2872 (O_2872,N_21294,N_24776);
or UO_2873 (O_2873,N_24070,N_24804);
or UO_2874 (O_2874,N_22854,N_23988);
or UO_2875 (O_2875,N_21881,N_22376);
and UO_2876 (O_2876,N_21344,N_20822);
xnor UO_2877 (O_2877,N_23907,N_20584);
nand UO_2878 (O_2878,N_24331,N_24177);
or UO_2879 (O_2879,N_20682,N_24830);
xor UO_2880 (O_2880,N_21112,N_20172);
xnor UO_2881 (O_2881,N_22530,N_21998);
nand UO_2882 (O_2882,N_20623,N_23503);
nand UO_2883 (O_2883,N_24531,N_21610);
nand UO_2884 (O_2884,N_22179,N_23148);
nand UO_2885 (O_2885,N_22276,N_22484);
xnor UO_2886 (O_2886,N_24217,N_21578);
and UO_2887 (O_2887,N_23122,N_23622);
and UO_2888 (O_2888,N_24276,N_23778);
or UO_2889 (O_2889,N_24743,N_21944);
and UO_2890 (O_2890,N_22731,N_22244);
nand UO_2891 (O_2891,N_23644,N_22934);
nand UO_2892 (O_2892,N_21077,N_20326);
nand UO_2893 (O_2893,N_23368,N_23288);
or UO_2894 (O_2894,N_23653,N_23084);
nor UO_2895 (O_2895,N_22048,N_23112);
or UO_2896 (O_2896,N_20564,N_21788);
nand UO_2897 (O_2897,N_24874,N_22786);
nand UO_2898 (O_2898,N_23307,N_22649);
xor UO_2899 (O_2899,N_24300,N_20024);
and UO_2900 (O_2900,N_20484,N_21358);
nand UO_2901 (O_2901,N_23667,N_23373);
nor UO_2902 (O_2902,N_22692,N_21922);
nand UO_2903 (O_2903,N_21308,N_24113);
nor UO_2904 (O_2904,N_23657,N_20101);
xnor UO_2905 (O_2905,N_20132,N_20216);
and UO_2906 (O_2906,N_21749,N_20828);
nor UO_2907 (O_2907,N_20654,N_22682);
and UO_2908 (O_2908,N_24139,N_24519);
and UO_2909 (O_2909,N_22619,N_24910);
nor UO_2910 (O_2910,N_23421,N_23152);
or UO_2911 (O_2911,N_24059,N_23240);
or UO_2912 (O_2912,N_20769,N_20871);
nor UO_2913 (O_2913,N_20258,N_21922);
or UO_2914 (O_2914,N_21553,N_22643);
or UO_2915 (O_2915,N_23036,N_23113);
and UO_2916 (O_2916,N_24175,N_23282);
xnor UO_2917 (O_2917,N_24638,N_23021);
and UO_2918 (O_2918,N_22209,N_23579);
nand UO_2919 (O_2919,N_23627,N_24410);
nand UO_2920 (O_2920,N_23462,N_20877);
xnor UO_2921 (O_2921,N_24252,N_21779);
or UO_2922 (O_2922,N_20063,N_22577);
nand UO_2923 (O_2923,N_22461,N_22478);
or UO_2924 (O_2924,N_20010,N_21006);
nand UO_2925 (O_2925,N_24786,N_22863);
nor UO_2926 (O_2926,N_21967,N_24395);
or UO_2927 (O_2927,N_24311,N_21199);
xnor UO_2928 (O_2928,N_21930,N_24615);
and UO_2929 (O_2929,N_24111,N_23419);
and UO_2930 (O_2930,N_24451,N_23854);
nand UO_2931 (O_2931,N_20452,N_24656);
xnor UO_2932 (O_2932,N_24143,N_20236);
and UO_2933 (O_2933,N_22927,N_24186);
xnor UO_2934 (O_2934,N_23828,N_20960);
or UO_2935 (O_2935,N_22407,N_23691);
and UO_2936 (O_2936,N_24666,N_24729);
and UO_2937 (O_2937,N_20985,N_23371);
nand UO_2938 (O_2938,N_21093,N_22814);
nand UO_2939 (O_2939,N_24335,N_21929);
xor UO_2940 (O_2940,N_20361,N_20179);
nand UO_2941 (O_2941,N_22663,N_24521);
nand UO_2942 (O_2942,N_22116,N_21814);
nor UO_2943 (O_2943,N_20017,N_24426);
xor UO_2944 (O_2944,N_24762,N_22978);
nand UO_2945 (O_2945,N_21256,N_23498);
and UO_2946 (O_2946,N_21378,N_23443);
and UO_2947 (O_2947,N_23339,N_21073);
or UO_2948 (O_2948,N_24224,N_22188);
nor UO_2949 (O_2949,N_23063,N_23647);
or UO_2950 (O_2950,N_20430,N_24714);
nor UO_2951 (O_2951,N_20105,N_22680);
or UO_2952 (O_2952,N_22481,N_22286);
nor UO_2953 (O_2953,N_24900,N_24123);
xor UO_2954 (O_2954,N_20373,N_24157);
nand UO_2955 (O_2955,N_23417,N_23226);
nand UO_2956 (O_2956,N_20220,N_20811);
nor UO_2957 (O_2957,N_20897,N_22338);
and UO_2958 (O_2958,N_21155,N_22615);
and UO_2959 (O_2959,N_21698,N_20380);
xnor UO_2960 (O_2960,N_24045,N_21216);
nor UO_2961 (O_2961,N_21051,N_24991);
or UO_2962 (O_2962,N_23893,N_21337);
xor UO_2963 (O_2963,N_20797,N_23744);
or UO_2964 (O_2964,N_20684,N_21555);
nand UO_2965 (O_2965,N_20705,N_23840);
xor UO_2966 (O_2966,N_23534,N_20272);
nor UO_2967 (O_2967,N_22657,N_20902);
xnor UO_2968 (O_2968,N_23226,N_23080);
and UO_2969 (O_2969,N_22493,N_22216);
nand UO_2970 (O_2970,N_24029,N_22328);
and UO_2971 (O_2971,N_21672,N_20918);
xor UO_2972 (O_2972,N_20652,N_24101);
and UO_2973 (O_2973,N_23446,N_23806);
nand UO_2974 (O_2974,N_23781,N_20409);
and UO_2975 (O_2975,N_21126,N_23736);
or UO_2976 (O_2976,N_20388,N_20434);
nor UO_2977 (O_2977,N_23547,N_20798);
or UO_2978 (O_2978,N_21647,N_20482);
and UO_2979 (O_2979,N_24841,N_21891);
nor UO_2980 (O_2980,N_24975,N_24720);
nand UO_2981 (O_2981,N_23173,N_20923);
xor UO_2982 (O_2982,N_21623,N_22435);
nand UO_2983 (O_2983,N_21423,N_23916);
and UO_2984 (O_2984,N_22929,N_24819);
xnor UO_2985 (O_2985,N_21499,N_22125);
or UO_2986 (O_2986,N_23310,N_22895);
xor UO_2987 (O_2987,N_24313,N_22835);
and UO_2988 (O_2988,N_22675,N_20853);
xor UO_2989 (O_2989,N_20864,N_21093);
and UO_2990 (O_2990,N_24428,N_20121);
nand UO_2991 (O_2991,N_23849,N_21971);
and UO_2992 (O_2992,N_24288,N_20345);
and UO_2993 (O_2993,N_20964,N_21497);
nand UO_2994 (O_2994,N_20334,N_21723);
xnor UO_2995 (O_2995,N_20352,N_24338);
nand UO_2996 (O_2996,N_20210,N_24174);
or UO_2997 (O_2997,N_24053,N_23462);
nand UO_2998 (O_2998,N_23017,N_21315);
or UO_2999 (O_2999,N_24554,N_24399);
endmodule