module basic_500_3000_500_40_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_61,In_133);
nand U1 (N_1,In_150,In_41);
nor U2 (N_2,In_155,In_270);
or U3 (N_3,In_399,In_23);
nand U4 (N_4,In_295,In_205);
nor U5 (N_5,In_254,In_354);
nor U6 (N_6,In_117,In_186);
or U7 (N_7,In_65,In_175);
and U8 (N_8,In_457,In_43);
or U9 (N_9,In_404,In_160);
and U10 (N_10,In_57,In_176);
nand U11 (N_11,In_441,In_313);
and U12 (N_12,In_11,In_20);
nand U13 (N_13,In_344,In_263);
nor U14 (N_14,In_67,In_109);
nor U15 (N_15,In_421,In_467);
nand U16 (N_16,In_290,In_286);
nor U17 (N_17,In_233,In_50);
nand U18 (N_18,In_104,In_89);
and U19 (N_19,In_15,In_82);
nor U20 (N_20,In_314,In_164);
or U21 (N_21,In_243,In_495);
and U22 (N_22,In_278,In_27);
nor U23 (N_23,In_106,In_272);
nor U24 (N_24,In_18,In_14);
nand U25 (N_25,In_203,In_283);
or U26 (N_26,In_232,In_4);
nand U27 (N_27,In_269,In_139);
nor U28 (N_28,In_339,In_137);
or U29 (N_29,In_22,In_180);
nand U30 (N_30,In_84,In_474);
nor U31 (N_31,In_154,In_494);
and U32 (N_32,In_102,In_173);
nor U33 (N_33,In_51,In_294);
and U34 (N_34,In_93,In_382);
nand U35 (N_35,In_287,In_265);
nand U36 (N_36,In_210,In_490);
nand U37 (N_37,In_236,In_140);
nand U38 (N_38,In_324,In_416);
nor U39 (N_39,In_152,In_85);
or U40 (N_40,In_182,In_128);
nand U41 (N_41,In_56,In_429);
xor U42 (N_42,In_248,In_466);
and U43 (N_43,In_410,In_480);
nand U44 (N_44,In_240,In_482);
and U45 (N_45,In_40,In_190);
nor U46 (N_46,In_464,In_45);
nand U47 (N_47,In_326,In_499);
or U48 (N_48,In_259,In_379);
nor U49 (N_49,In_491,In_385);
nand U50 (N_50,In_52,In_262);
nand U51 (N_51,In_308,In_195);
nor U52 (N_52,In_252,In_397);
nor U53 (N_53,In_479,In_200);
nand U54 (N_54,In_275,In_260);
nor U55 (N_55,In_289,In_181);
or U56 (N_56,In_322,In_422);
nor U57 (N_57,In_111,In_73);
nand U58 (N_58,In_121,In_298);
and U59 (N_59,In_369,In_25);
and U60 (N_60,In_432,In_235);
and U61 (N_61,In_336,In_485);
or U62 (N_62,In_273,In_250);
or U63 (N_63,In_493,In_215);
nand U64 (N_64,In_189,In_148);
or U65 (N_65,In_388,In_446);
or U66 (N_66,In_194,In_115);
or U67 (N_67,In_403,In_55);
and U68 (N_68,In_129,In_319);
and U69 (N_69,In_35,In_311);
or U70 (N_70,In_202,In_86);
nor U71 (N_71,In_361,In_219);
nor U72 (N_72,In_1,In_374);
nor U73 (N_73,In_384,In_221);
nand U74 (N_74,In_212,In_271);
or U75 (N_75,In_280,In_33);
nand U76 (N_76,In_419,In_224);
or U77 (N_77,In_373,In_151);
nand U78 (N_78,In_257,In_381);
or U79 (N_79,In_284,In_193);
nand U80 (N_80,In_341,In_332);
and U81 (N_81,In_213,In_321);
or U82 (N_82,In_112,N_9);
or U83 (N_83,In_301,In_185);
nor U84 (N_84,In_476,In_188);
or U85 (N_85,In_62,N_55);
or U86 (N_86,In_279,In_108);
nand U87 (N_87,In_145,In_393);
nor U88 (N_88,N_34,In_497);
nor U89 (N_89,In_299,In_348);
nor U90 (N_90,In_216,In_444);
and U91 (N_91,In_101,In_435);
nand U92 (N_92,In_402,In_208);
nand U93 (N_93,In_12,N_45);
nor U94 (N_94,In_391,In_120);
nand U95 (N_95,N_56,In_66);
and U96 (N_96,In_103,N_11);
nor U97 (N_97,In_231,In_118);
or U98 (N_98,In_445,In_87);
nand U99 (N_99,In_414,In_304);
nand U100 (N_100,In_383,In_206);
nand U101 (N_101,In_47,In_242);
and U102 (N_102,In_296,In_302);
nor U103 (N_103,N_23,In_222);
or U104 (N_104,In_163,N_35);
nand U105 (N_105,In_199,In_471);
or U106 (N_106,N_1,N_33);
and U107 (N_107,In_187,In_458);
nor U108 (N_108,In_484,N_41);
nor U109 (N_109,N_29,In_83);
and U110 (N_110,In_114,In_98);
nor U111 (N_111,N_30,In_335);
and U112 (N_112,In_415,In_398);
or U113 (N_113,In_229,In_309);
nor U114 (N_114,In_498,In_94);
or U115 (N_115,In_358,In_307);
or U116 (N_116,N_64,In_126);
or U117 (N_117,In_405,In_7);
or U118 (N_118,N_18,In_331);
and U119 (N_119,In_238,In_179);
and U120 (N_120,N_25,In_423);
and U121 (N_121,In_5,In_401);
and U122 (N_122,In_478,N_40);
or U123 (N_123,N_50,In_472);
and U124 (N_124,In_327,N_47);
or U125 (N_125,N_12,In_24);
nand U126 (N_126,In_333,In_95);
or U127 (N_127,In_127,N_67);
nor U128 (N_128,In_487,In_178);
or U129 (N_129,N_74,In_303);
and U130 (N_130,N_51,In_357);
nand U131 (N_131,In_267,In_44);
and U132 (N_132,In_315,In_375);
nor U133 (N_133,In_424,In_355);
and U134 (N_134,In_395,In_153);
nand U135 (N_135,N_8,In_468);
or U136 (N_136,In_400,In_367);
nor U137 (N_137,N_0,In_264);
or U138 (N_138,N_69,In_300);
nor U139 (N_139,N_61,In_197);
nor U140 (N_140,In_149,In_184);
nor U141 (N_141,In_244,In_266);
nor U142 (N_142,In_97,N_71);
and U143 (N_143,In_125,In_253);
nor U144 (N_144,In_438,N_14);
nor U145 (N_145,In_165,In_430);
nor U146 (N_146,In_337,In_318);
or U147 (N_147,In_192,In_486);
nand U148 (N_148,In_207,In_345);
xor U149 (N_149,In_31,N_32);
nand U150 (N_150,In_274,N_143);
or U151 (N_151,In_0,N_94);
nor U152 (N_152,N_115,In_91);
and U153 (N_153,In_352,In_167);
nand U154 (N_154,In_48,In_225);
and U155 (N_155,In_483,In_159);
and U156 (N_156,In_447,In_157);
nand U157 (N_157,In_59,N_83);
and U158 (N_158,N_147,In_63);
nor U159 (N_159,N_38,In_46);
nand U160 (N_160,In_123,In_366);
and U161 (N_161,N_26,In_170);
nor U162 (N_162,N_106,In_53);
nor U163 (N_163,N_52,N_15);
nor U164 (N_164,In_370,N_77);
nor U165 (N_165,N_107,In_171);
or U166 (N_166,In_439,In_147);
nor U167 (N_167,In_451,N_43);
or U168 (N_168,In_144,In_426);
xnor U169 (N_169,In_17,In_470);
nor U170 (N_170,N_53,In_79);
nand U171 (N_171,In_122,In_38);
and U172 (N_172,In_378,N_135);
nor U173 (N_173,N_48,N_130);
or U174 (N_174,In_277,In_177);
and U175 (N_175,N_136,N_7);
nand U176 (N_176,In_360,In_29);
nand U177 (N_177,In_368,N_90);
and U178 (N_178,In_459,In_362);
nand U179 (N_179,N_134,In_390);
nand U180 (N_180,In_246,In_10);
nand U181 (N_181,In_42,N_20);
nor U182 (N_182,N_146,N_99);
nand U183 (N_183,N_111,In_347);
nand U184 (N_184,N_120,In_136);
and U185 (N_185,N_84,In_473);
nor U186 (N_186,In_396,In_436);
nor U187 (N_187,In_54,In_19);
nand U188 (N_188,In_131,In_481);
nand U189 (N_189,N_97,In_312);
and U190 (N_190,In_161,In_392);
nand U191 (N_191,In_36,N_2);
or U192 (N_192,In_317,N_78);
or U193 (N_193,In_58,N_140);
and U194 (N_194,N_58,N_109);
or U195 (N_195,In_305,N_42);
nand U196 (N_196,In_174,In_228);
nand U197 (N_197,N_98,In_28);
nand U198 (N_198,In_60,N_44);
and U199 (N_199,In_310,In_359);
and U200 (N_200,In_316,In_99);
nand U201 (N_201,N_60,N_121);
nand U202 (N_202,In_387,In_32);
xor U203 (N_203,In_211,In_88);
nand U204 (N_204,In_349,In_442);
nand U205 (N_205,N_31,In_492);
and U206 (N_206,In_110,N_149);
and U207 (N_207,In_76,In_288);
nor U208 (N_208,In_105,In_256);
and U209 (N_209,In_389,In_30);
or U210 (N_210,In_70,N_36);
and U211 (N_211,In_418,In_34);
and U212 (N_212,In_406,In_453);
nand U213 (N_213,N_104,N_49);
and U214 (N_214,N_46,In_230);
nor U215 (N_215,In_132,In_239);
nand U216 (N_216,In_477,In_223);
nand U217 (N_217,N_73,N_129);
nand U218 (N_218,In_9,N_75);
or U219 (N_219,In_320,In_141);
xor U220 (N_220,N_39,In_124);
or U221 (N_221,In_49,N_89);
or U222 (N_222,In_37,In_434);
nor U223 (N_223,In_469,In_386);
and U224 (N_224,In_168,In_363);
nand U225 (N_225,In_465,In_143);
or U226 (N_226,In_96,In_169);
nand U227 (N_227,N_22,N_194);
nor U228 (N_228,In_78,N_186);
and U229 (N_229,In_191,In_245);
nor U230 (N_230,N_166,In_2);
nor U231 (N_231,In_356,N_80);
and U232 (N_232,N_62,N_70);
or U233 (N_233,In_365,N_195);
or U234 (N_234,In_16,N_37);
or U235 (N_235,N_196,N_126);
nor U236 (N_236,In_100,N_210);
or U237 (N_237,N_66,In_72);
and U238 (N_238,In_346,In_292);
or U239 (N_239,In_276,N_217);
or U240 (N_240,N_3,N_204);
and U241 (N_241,In_196,N_137);
and U242 (N_242,In_217,In_407);
nor U243 (N_243,In_218,N_152);
or U244 (N_244,N_223,N_132);
or U245 (N_245,In_443,In_90);
nor U246 (N_246,N_221,N_224);
nor U247 (N_247,N_213,N_161);
and U248 (N_248,N_116,N_118);
nand U249 (N_249,N_119,In_255);
and U250 (N_250,In_460,N_160);
and U251 (N_251,N_165,N_114);
and U252 (N_252,In_394,In_251);
nor U253 (N_253,In_226,In_220);
nand U254 (N_254,In_351,In_413);
and U255 (N_255,In_249,In_297);
nor U256 (N_256,In_74,N_5);
nand U257 (N_257,In_68,In_433);
nor U258 (N_258,In_158,N_105);
or U259 (N_259,N_198,N_154);
or U260 (N_260,In_237,N_82);
nand U261 (N_261,In_156,N_189);
or U262 (N_262,N_185,N_215);
and U263 (N_263,N_79,In_488);
nor U264 (N_264,N_68,N_218);
and U265 (N_265,N_142,N_128);
or U266 (N_266,In_372,N_10);
nor U267 (N_267,N_102,In_291);
xor U268 (N_268,N_4,In_411);
and U269 (N_269,In_412,In_342);
or U270 (N_270,In_227,N_199);
nand U271 (N_271,In_440,In_285);
nand U272 (N_272,In_329,N_123);
nand U273 (N_273,In_6,In_247);
and U274 (N_274,In_282,N_214);
and U275 (N_275,In_462,In_475);
or U276 (N_276,N_108,In_380);
or U277 (N_277,N_212,N_208);
and U278 (N_278,N_180,N_145);
and U279 (N_279,In_119,N_169);
and U280 (N_280,In_69,N_24);
nand U281 (N_281,N_131,N_222);
or U282 (N_282,N_162,In_456);
nor U283 (N_283,N_113,In_71);
nor U284 (N_284,N_171,N_85);
and U285 (N_285,In_328,N_101);
nor U286 (N_286,In_496,N_88);
nor U287 (N_287,In_408,In_234);
and U288 (N_288,In_420,N_95);
nor U289 (N_289,N_197,N_155);
and U290 (N_290,In_452,In_142);
nor U291 (N_291,In_130,In_75);
nand U292 (N_292,In_13,N_167);
or U293 (N_293,N_156,N_164);
nor U294 (N_294,N_81,N_100);
nor U295 (N_295,In_198,N_124);
nor U296 (N_296,N_168,In_489);
and U297 (N_297,N_63,In_330);
and U298 (N_298,N_190,In_146);
and U299 (N_299,N_176,N_202);
nor U300 (N_300,N_54,N_264);
and U301 (N_301,In_323,N_209);
nor U302 (N_302,N_252,N_271);
or U303 (N_303,In_353,N_286);
nand U304 (N_304,N_19,N_281);
and U305 (N_305,N_283,N_297);
nor U306 (N_306,N_241,In_463);
or U307 (N_307,In_81,In_450);
nand U308 (N_308,N_294,N_253);
or U309 (N_309,N_211,N_59);
and U310 (N_310,In_162,N_182);
nand U311 (N_311,N_117,In_214);
and U312 (N_312,N_243,N_279);
and U313 (N_313,N_262,N_261);
and U314 (N_314,N_259,N_228);
nor U315 (N_315,N_87,N_284);
and U316 (N_316,N_287,N_141);
and U317 (N_317,In_268,N_103);
nand U318 (N_318,N_278,N_174);
nor U319 (N_319,N_163,N_257);
nor U320 (N_320,In_343,N_298);
and U321 (N_321,In_26,N_150);
or U322 (N_322,N_249,N_157);
nand U323 (N_323,N_175,N_268);
or U324 (N_324,N_92,N_285);
and U325 (N_325,In_376,N_288);
and U326 (N_326,N_28,N_230);
nor U327 (N_327,In_425,N_200);
nand U328 (N_328,N_207,N_240);
nor U329 (N_329,N_256,N_219);
nand U330 (N_330,N_151,N_292);
nand U331 (N_331,N_234,In_364);
nor U332 (N_332,N_289,N_269);
nand U333 (N_333,In_258,N_184);
or U334 (N_334,N_265,N_138);
nor U335 (N_335,N_290,In_135);
nand U336 (N_336,In_371,N_96);
or U337 (N_337,N_255,In_64);
nor U338 (N_338,In_427,In_334);
nor U339 (N_339,N_191,N_72);
nand U340 (N_340,N_170,N_277);
nor U341 (N_341,In_431,N_133);
nor U342 (N_342,N_244,In_261);
or U343 (N_343,N_173,In_338);
or U344 (N_344,In_3,N_267);
and U345 (N_345,N_177,In_92);
nand U346 (N_346,N_57,N_205);
and U347 (N_347,In_77,N_276);
nor U348 (N_348,N_188,N_158);
nor U349 (N_349,N_251,N_127);
and U350 (N_350,N_206,N_225);
nand U351 (N_351,In_201,In_39);
nor U352 (N_352,In_306,N_229);
nand U353 (N_353,In_448,N_144);
nand U354 (N_354,N_258,N_293);
and U355 (N_355,In_80,N_227);
or U356 (N_356,In_325,In_437);
nand U357 (N_357,N_27,N_291);
nand U358 (N_358,N_270,N_148);
nor U359 (N_359,N_216,N_295);
and U360 (N_360,N_266,N_275);
nor U361 (N_361,N_93,N_112);
or U362 (N_362,N_242,N_263);
and U363 (N_363,N_179,In_340);
nand U364 (N_364,N_181,N_250);
nand U365 (N_365,N_236,N_299);
nor U366 (N_366,N_226,N_16);
and U367 (N_367,N_220,In_209);
and U368 (N_368,In_293,In_172);
and U369 (N_369,In_454,N_172);
nand U370 (N_370,In_107,N_272);
and U371 (N_371,N_139,N_13);
nor U372 (N_372,N_125,N_187);
or U373 (N_373,In_377,In_417);
and U374 (N_374,N_248,N_231);
and U375 (N_375,N_364,N_363);
nor U376 (N_376,In_21,N_358);
or U377 (N_377,N_339,N_193);
nand U378 (N_378,N_233,N_246);
nand U379 (N_379,N_300,N_178);
nand U380 (N_380,N_322,N_235);
and U381 (N_381,N_260,N_332);
nor U382 (N_382,N_159,N_340);
nand U383 (N_383,N_374,N_341);
nand U384 (N_384,N_351,N_346);
and U385 (N_385,N_357,N_356);
nor U386 (N_386,N_347,In_166);
or U387 (N_387,N_371,N_305);
nor U388 (N_388,N_368,N_274);
nand U389 (N_389,In_241,N_320);
and U390 (N_390,N_6,N_317);
or U391 (N_391,N_336,N_370);
nor U392 (N_392,N_306,N_203);
and U393 (N_393,In_428,N_254);
nand U394 (N_394,N_321,N_307);
or U395 (N_395,N_330,In_449);
or U396 (N_396,N_309,N_192);
nand U397 (N_397,N_238,N_282);
nor U398 (N_398,N_318,N_327);
nor U399 (N_399,N_302,N_304);
nor U400 (N_400,N_153,N_373);
nand U401 (N_401,N_369,N_329);
or U402 (N_402,In_350,N_280);
or U403 (N_403,N_315,N_349);
and U404 (N_404,N_360,N_343);
nand U405 (N_405,N_367,N_323);
nor U406 (N_406,N_76,N_338);
and U407 (N_407,In_134,N_201);
or U408 (N_408,N_345,N_296);
nor U409 (N_409,N_355,N_350);
nor U410 (N_410,N_91,N_326);
and U411 (N_411,N_313,In_409);
and U412 (N_412,N_352,N_110);
nor U413 (N_413,N_314,N_324);
nand U414 (N_414,In_281,In_204);
and U415 (N_415,In_183,N_245);
and U416 (N_416,N_334,N_310);
or U417 (N_417,N_337,In_113);
nand U418 (N_418,In_455,N_372);
nor U419 (N_419,N_247,N_17);
or U420 (N_420,N_359,N_303);
nor U421 (N_421,In_138,N_344);
and U422 (N_422,N_86,N_21);
nor U423 (N_423,N_362,N_311);
or U424 (N_424,N_325,N_319);
or U425 (N_425,N_122,In_116);
and U426 (N_426,N_342,N_331);
and U427 (N_427,N_301,In_8);
nand U428 (N_428,N_328,N_273);
or U429 (N_429,N_333,N_354);
nand U430 (N_430,N_65,N_348);
nor U431 (N_431,N_239,N_308);
or U432 (N_432,N_335,N_365);
or U433 (N_433,N_232,N_316);
nor U434 (N_434,N_183,N_353);
nand U435 (N_435,In_461,N_237);
and U436 (N_436,N_312,N_361);
nand U437 (N_437,N_366,N_308);
or U438 (N_438,N_337,N_76);
or U439 (N_439,N_342,N_233);
nand U440 (N_440,N_273,N_280);
nor U441 (N_441,N_305,N_233);
and U442 (N_442,N_21,N_254);
nand U443 (N_443,N_203,N_337);
or U444 (N_444,N_345,N_330);
nor U445 (N_445,N_296,N_305);
nand U446 (N_446,N_353,N_338);
or U447 (N_447,N_303,In_21);
nor U448 (N_448,In_8,N_183);
and U449 (N_449,N_21,N_367);
nand U450 (N_450,N_427,N_435);
and U451 (N_451,N_401,N_447);
or U452 (N_452,N_416,N_404);
or U453 (N_453,N_395,N_449);
and U454 (N_454,N_380,N_379);
nor U455 (N_455,N_425,N_394);
nand U456 (N_456,N_405,N_437);
nor U457 (N_457,N_396,N_387);
nor U458 (N_458,N_412,N_444);
and U459 (N_459,N_389,N_418);
and U460 (N_460,N_411,N_388);
nor U461 (N_461,N_410,N_408);
and U462 (N_462,N_436,N_428);
or U463 (N_463,N_377,N_423);
or U464 (N_464,N_403,N_434);
nor U465 (N_465,N_413,N_448);
and U466 (N_466,N_392,N_430);
nor U467 (N_467,N_424,N_421);
nand U468 (N_468,N_400,N_406);
or U469 (N_469,N_390,N_375);
nor U470 (N_470,N_440,N_432);
nand U471 (N_471,N_381,N_420);
nor U472 (N_472,N_397,N_417);
nor U473 (N_473,N_426,N_398);
and U474 (N_474,N_415,N_378);
nor U475 (N_475,N_393,N_438);
nand U476 (N_476,N_382,N_399);
or U477 (N_477,N_409,N_433);
nand U478 (N_478,N_386,N_385);
and U479 (N_479,N_445,N_407);
and U480 (N_480,N_376,N_384);
or U481 (N_481,N_414,N_441);
or U482 (N_482,N_439,N_429);
nand U483 (N_483,N_422,N_431);
or U484 (N_484,N_442,N_391);
or U485 (N_485,N_419,N_446);
and U486 (N_486,N_383,N_443);
nand U487 (N_487,N_402,N_414);
nor U488 (N_488,N_396,N_410);
nor U489 (N_489,N_441,N_384);
nand U490 (N_490,N_431,N_394);
and U491 (N_491,N_385,N_394);
and U492 (N_492,N_387,N_418);
or U493 (N_493,N_393,N_405);
and U494 (N_494,N_382,N_400);
and U495 (N_495,N_415,N_410);
nor U496 (N_496,N_425,N_421);
nand U497 (N_497,N_436,N_390);
and U498 (N_498,N_382,N_430);
nand U499 (N_499,N_432,N_405);
nand U500 (N_500,N_407,N_396);
nor U501 (N_501,N_442,N_377);
nor U502 (N_502,N_415,N_421);
and U503 (N_503,N_449,N_403);
nor U504 (N_504,N_437,N_377);
nor U505 (N_505,N_406,N_429);
and U506 (N_506,N_402,N_445);
nand U507 (N_507,N_428,N_378);
or U508 (N_508,N_389,N_380);
and U509 (N_509,N_404,N_394);
or U510 (N_510,N_385,N_387);
or U511 (N_511,N_418,N_449);
nor U512 (N_512,N_419,N_425);
nand U513 (N_513,N_386,N_448);
or U514 (N_514,N_439,N_425);
and U515 (N_515,N_401,N_400);
nand U516 (N_516,N_422,N_399);
or U517 (N_517,N_407,N_420);
nor U518 (N_518,N_404,N_419);
nor U519 (N_519,N_397,N_381);
nand U520 (N_520,N_403,N_423);
nor U521 (N_521,N_377,N_400);
nand U522 (N_522,N_375,N_380);
and U523 (N_523,N_393,N_417);
nor U524 (N_524,N_425,N_443);
nand U525 (N_525,N_477,N_469);
nand U526 (N_526,N_523,N_478);
nand U527 (N_527,N_517,N_522);
or U528 (N_528,N_510,N_462);
nor U529 (N_529,N_464,N_475);
and U530 (N_530,N_461,N_482);
or U531 (N_531,N_458,N_452);
nand U532 (N_532,N_521,N_473);
nand U533 (N_533,N_455,N_519);
nand U534 (N_534,N_512,N_516);
or U535 (N_535,N_503,N_515);
nor U536 (N_536,N_485,N_508);
or U537 (N_537,N_501,N_460);
nand U538 (N_538,N_498,N_489);
nand U539 (N_539,N_456,N_465);
and U540 (N_540,N_454,N_506);
and U541 (N_541,N_513,N_453);
nand U542 (N_542,N_494,N_468);
nand U543 (N_543,N_467,N_520);
nand U544 (N_544,N_480,N_492);
nand U545 (N_545,N_511,N_466);
or U546 (N_546,N_472,N_504);
and U547 (N_547,N_496,N_463);
and U548 (N_548,N_499,N_484);
and U549 (N_549,N_488,N_495);
or U550 (N_550,N_490,N_451);
or U551 (N_551,N_471,N_476);
or U552 (N_552,N_509,N_486);
nand U553 (N_553,N_507,N_505);
nand U554 (N_554,N_524,N_470);
or U555 (N_555,N_500,N_497);
nor U556 (N_556,N_479,N_483);
nor U557 (N_557,N_491,N_474);
nor U558 (N_558,N_518,N_459);
nand U559 (N_559,N_481,N_457);
xor U560 (N_560,N_502,N_487);
or U561 (N_561,N_493,N_514);
nand U562 (N_562,N_450,N_461);
nand U563 (N_563,N_518,N_512);
and U564 (N_564,N_519,N_465);
and U565 (N_565,N_520,N_517);
nand U566 (N_566,N_487,N_524);
nand U567 (N_567,N_479,N_487);
and U568 (N_568,N_492,N_511);
or U569 (N_569,N_472,N_516);
nor U570 (N_570,N_517,N_501);
and U571 (N_571,N_503,N_466);
nand U572 (N_572,N_464,N_517);
or U573 (N_573,N_498,N_501);
or U574 (N_574,N_481,N_465);
and U575 (N_575,N_479,N_467);
nor U576 (N_576,N_500,N_462);
nand U577 (N_577,N_501,N_507);
and U578 (N_578,N_498,N_510);
nor U579 (N_579,N_516,N_494);
nand U580 (N_580,N_494,N_520);
nor U581 (N_581,N_470,N_483);
or U582 (N_582,N_516,N_463);
and U583 (N_583,N_520,N_465);
nor U584 (N_584,N_512,N_466);
or U585 (N_585,N_522,N_505);
and U586 (N_586,N_489,N_508);
nand U587 (N_587,N_454,N_485);
and U588 (N_588,N_461,N_478);
nor U589 (N_589,N_457,N_498);
and U590 (N_590,N_519,N_471);
nor U591 (N_591,N_488,N_481);
and U592 (N_592,N_499,N_497);
and U593 (N_593,N_517,N_474);
and U594 (N_594,N_462,N_497);
and U595 (N_595,N_491,N_494);
and U596 (N_596,N_471,N_486);
or U597 (N_597,N_518,N_451);
nor U598 (N_598,N_508,N_513);
nor U599 (N_599,N_456,N_460);
or U600 (N_600,N_560,N_575);
nand U601 (N_601,N_576,N_593);
nand U602 (N_602,N_550,N_577);
or U603 (N_603,N_527,N_540);
nand U604 (N_604,N_590,N_557);
nand U605 (N_605,N_525,N_594);
and U606 (N_606,N_538,N_587);
and U607 (N_607,N_555,N_569);
and U608 (N_608,N_559,N_533);
and U609 (N_609,N_561,N_545);
and U610 (N_610,N_537,N_536);
and U611 (N_611,N_556,N_553);
nor U612 (N_612,N_549,N_597);
or U613 (N_613,N_554,N_591);
nor U614 (N_614,N_578,N_547);
and U615 (N_615,N_546,N_589);
or U616 (N_616,N_571,N_563);
and U617 (N_617,N_579,N_535);
nor U618 (N_618,N_534,N_552);
and U619 (N_619,N_543,N_528);
nand U620 (N_620,N_592,N_548);
and U621 (N_621,N_566,N_567);
or U622 (N_622,N_531,N_599);
nand U623 (N_623,N_584,N_564);
nor U624 (N_624,N_595,N_532);
nand U625 (N_625,N_573,N_544);
and U626 (N_626,N_542,N_529);
nand U627 (N_627,N_586,N_551);
nor U628 (N_628,N_583,N_582);
or U629 (N_629,N_526,N_562);
or U630 (N_630,N_572,N_558);
and U631 (N_631,N_585,N_574);
or U632 (N_632,N_581,N_598);
nor U633 (N_633,N_568,N_596);
nor U634 (N_634,N_539,N_570);
and U635 (N_635,N_530,N_588);
or U636 (N_636,N_541,N_565);
nand U637 (N_637,N_580,N_540);
or U638 (N_638,N_595,N_544);
or U639 (N_639,N_533,N_596);
nand U640 (N_640,N_529,N_584);
nand U641 (N_641,N_573,N_562);
or U642 (N_642,N_553,N_573);
nand U643 (N_643,N_561,N_598);
nand U644 (N_644,N_562,N_546);
nand U645 (N_645,N_547,N_551);
nor U646 (N_646,N_531,N_570);
and U647 (N_647,N_573,N_583);
nor U648 (N_648,N_566,N_585);
nor U649 (N_649,N_539,N_568);
nand U650 (N_650,N_555,N_597);
or U651 (N_651,N_573,N_591);
nor U652 (N_652,N_577,N_556);
nor U653 (N_653,N_550,N_582);
or U654 (N_654,N_590,N_598);
nor U655 (N_655,N_556,N_579);
nand U656 (N_656,N_583,N_555);
or U657 (N_657,N_575,N_583);
nand U658 (N_658,N_581,N_560);
or U659 (N_659,N_525,N_574);
nand U660 (N_660,N_571,N_564);
or U661 (N_661,N_583,N_539);
nand U662 (N_662,N_595,N_570);
nand U663 (N_663,N_575,N_546);
nand U664 (N_664,N_558,N_528);
nand U665 (N_665,N_577,N_589);
nand U666 (N_666,N_589,N_561);
or U667 (N_667,N_541,N_574);
nor U668 (N_668,N_596,N_530);
and U669 (N_669,N_573,N_567);
and U670 (N_670,N_536,N_590);
nand U671 (N_671,N_571,N_538);
and U672 (N_672,N_598,N_557);
nand U673 (N_673,N_597,N_533);
or U674 (N_674,N_531,N_533);
nor U675 (N_675,N_653,N_604);
xnor U676 (N_676,N_660,N_610);
or U677 (N_677,N_616,N_608);
and U678 (N_678,N_669,N_673);
or U679 (N_679,N_623,N_664);
or U680 (N_680,N_636,N_649);
or U681 (N_681,N_658,N_638);
nand U682 (N_682,N_641,N_633);
or U683 (N_683,N_671,N_635);
nand U684 (N_684,N_628,N_615);
or U685 (N_685,N_609,N_631);
and U686 (N_686,N_662,N_611);
nand U687 (N_687,N_626,N_629);
nand U688 (N_688,N_674,N_652);
nand U689 (N_689,N_666,N_650);
nand U690 (N_690,N_601,N_670);
nand U691 (N_691,N_643,N_625);
nor U692 (N_692,N_613,N_654);
nor U693 (N_693,N_672,N_640);
and U694 (N_694,N_630,N_655);
nor U695 (N_695,N_634,N_620);
nor U696 (N_696,N_612,N_637);
or U697 (N_697,N_602,N_606);
nor U698 (N_698,N_665,N_644);
or U699 (N_699,N_651,N_645);
or U700 (N_700,N_624,N_607);
nor U701 (N_701,N_639,N_605);
nor U702 (N_702,N_614,N_663);
nand U703 (N_703,N_659,N_600);
and U704 (N_704,N_668,N_622);
nand U705 (N_705,N_656,N_617);
and U706 (N_706,N_603,N_642);
xnor U707 (N_707,N_619,N_648);
nand U708 (N_708,N_661,N_647);
nor U709 (N_709,N_632,N_646);
or U710 (N_710,N_657,N_618);
xnor U711 (N_711,N_621,N_627);
nor U712 (N_712,N_667,N_625);
and U713 (N_713,N_650,N_606);
nor U714 (N_714,N_627,N_618);
nor U715 (N_715,N_601,N_613);
nor U716 (N_716,N_620,N_618);
or U717 (N_717,N_654,N_658);
nand U718 (N_718,N_618,N_640);
or U719 (N_719,N_625,N_653);
and U720 (N_720,N_619,N_667);
nor U721 (N_721,N_643,N_644);
and U722 (N_722,N_650,N_643);
nand U723 (N_723,N_616,N_603);
nor U724 (N_724,N_610,N_638);
or U725 (N_725,N_635,N_663);
nand U726 (N_726,N_612,N_618);
or U727 (N_727,N_613,N_626);
and U728 (N_728,N_647,N_665);
and U729 (N_729,N_649,N_667);
or U730 (N_730,N_611,N_671);
nand U731 (N_731,N_644,N_604);
nor U732 (N_732,N_643,N_638);
nand U733 (N_733,N_657,N_615);
or U734 (N_734,N_600,N_646);
nor U735 (N_735,N_605,N_658);
nor U736 (N_736,N_612,N_638);
nand U737 (N_737,N_636,N_639);
and U738 (N_738,N_672,N_641);
nand U739 (N_739,N_674,N_646);
or U740 (N_740,N_600,N_603);
or U741 (N_741,N_669,N_674);
and U742 (N_742,N_619,N_614);
nand U743 (N_743,N_637,N_617);
nor U744 (N_744,N_634,N_614);
nand U745 (N_745,N_602,N_613);
or U746 (N_746,N_625,N_614);
or U747 (N_747,N_626,N_608);
and U748 (N_748,N_632,N_633);
nor U749 (N_749,N_649,N_617);
or U750 (N_750,N_685,N_729);
nor U751 (N_751,N_721,N_703);
nor U752 (N_752,N_708,N_707);
nor U753 (N_753,N_675,N_700);
xnor U754 (N_754,N_726,N_690);
and U755 (N_755,N_680,N_710);
nor U756 (N_756,N_738,N_722);
nor U757 (N_757,N_683,N_749);
nand U758 (N_758,N_720,N_747);
and U759 (N_759,N_678,N_702);
nor U760 (N_760,N_712,N_695);
nor U761 (N_761,N_734,N_711);
or U762 (N_762,N_744,N_716);
or U763 (N_763,N_731,N_706);
or U764 (N_764,N_684,N_713);
nand U765 (N_765,N_688,N_677);
and U766 (N_766,N_686,N_730);
nor U767 (N_767,N_692,N_705);
nor U768 (N_768,N_717,N_724);
or U769 (N_769,N_741,N_733);
nand U770 (N_770,N_736,N_740);
nand U771 (N_771,N_709,N_701);
or U772 (N_772,N_693,N_714);
nand U773 (N_773,N_746,N_748);
nand U774 (N_774,N_704,N_681);
xnor U775 (N_775,N_745,N_715);
and U776 (N_776,N_728,N_723);
or U777 (N_777,N_739,N_698);
and U778 (N_778,N_687,N_737);
or U779 (N_779,N_679,N_676);
and U780 (N_780,N_694,N_742);
and U781 (N_781,N_727,N_732);
or U782 (N_782,N_718,N_735);
nor U783 (N_783,N_699,N_696);
and U784 (N_784,N_743,N_689);
or U785 (N_785,N_725,N_682);
and U786 (N_786,N_691,N_697);
and U787 (N_787,N_719,N_740);
and U788 (N_788,N_749,N_735);
xnor U789 (N_789,N_717,N_695);
nand U790 (N_790,N_745,N_724);
or U791 (N_791,N_683,N_737);
nor U792 (N_792,N_735,N_682);
or U793 (N_793,N_694,N_738);
nand U794 (N_794,N_692,N_677);
or U795 (N_795,N_704,N_745);
nor U796 (N_796,N_681,N_700);
or U797 (N_797,N_680,N_746);
nor U798 (N_798,N_675,N_727);
nor U799 (N_799,N_727,N_733);
nand U800 (N_800,N_700,N_745);
and U801 (N_801,N_702,N_730);
nor U802 (N_802,N_699,N_728);
and U803 (N_803,N_702,N_679);
and U804 (N_804,N_704,N_723);
or U805 (N_805,N_713,N_689);
or U806 (N_806,N_744,N_713);
nor U807 (N_807,N_686,N_699);
and U808 (N_808,N_682,N_709);
and U809 (N_809,N_696,N_706);
or U810 (N_810,N_701,N_707);
nand U811 (N_811,N_693,N_745);
or U812 (N_812,N_695,N_699);
and U813 (N_813,N_724,N_740);
or U814 (N_814,N_720,N_704);
nor U815 (N_815,N_707,N_679);
nor U816 (N_816,N_738,N_748);
or U817 (N_817,N_732,N_723);
or U818 (N_818,N_727,N_739);
and U819 (N_819,N_710,N_686);
nand U820 (N_820,N_696,N_683);
nor U821 (N_821,N_698,N_722);
or U822 (N_822,N_717,N_746);
or U823 (N_823,N_731,N_694);
nor U824 (N_824,N_706,N_683);
or U825 (N_825,N_793,N_763);
or U826 (N_826,N_760,N_798);
nor U827 (N_827,N_768,N_816);
nand U828 (N_828,N_755,N_777);
or U829 (N_829,N_783,N_810);
or U830 (N_830,N_797,N_773);
and U831 (N_831,N_778,N_779);
nand U832 (N_832,N_750,N_786);
nor U833 (N_833,N_800,N_769);
nor U834 (N_834,N_788,N_789);
nor U835 (N_835,N_822,N_807);
nor U836 (N_836,N_784,N_776);
and U837 (N_837,N_795,N_753);
nor U838 (N_838,N_820,N_787);
nand U839 (N_839,N_764,N_811);
or U840 (N_840,N_767,N_815);
or U841 (N_841,N_794,N_821);
and U842 (N_842,N_808,N_809);
and U843 (N_843,N_824,N_802);
and U844 (N_844,N_772,N_806);
and U845 (N_845,N_792,N_790);
nand U846 (N_846,N_775,N_774);
and U847 (N_847,N_770,N_766);
nor U848 (N_848,N_781,N_817);
nor U849 (N_849,N_752,N_804);
nand U850 (N_850,N_812,N_805);
nor U851 (N_851,N_780,N_813);
or U852 (N_852,N_823,N_762);
nor U853 (N_853,N_771,N_782);
nand U854 (N_854,N_761,N_803);
nand U855 (N_855,N_759,N_796);
and U856 (N_856,N_799,N_785);
nor U857 (N_857,N_756,N_819);
nor U858 (N_858,N_814,N_801);
nand U859 (N_859,N_818,N_765);
or U860 (N_860,N_751,N_791);
nand U861 (N_861,N_757,N_758);
nor U862 (N_862,N_754,N_760);
nand U863 (N_863,N_809,N_759);
nor U864 (N_864,N_807,N_763);
nor U865 (N_865,N_787,N_809);
nor U866 (N_866,N_802,N_761);
nor U867 (N_867,N_751,N_808);
nor U868 (N_868,N_751,N_815);
and U869 (N_869,N_802,N_758);
nand U870 (N_870,N_776,N_754);
or U871 (N_871,N_771,N_784);
or U872 (N_872,N_820,N_796);
nand U873 (N_873,N_763,N_762);
nand U874 (N_874,N_772,N_800);
nor U875 (N_875,N_805,N_788);
and U876 (N_876,N_811,N_801);
or U877 (N_877,N_811,N_822);
and U878 (N_878,N_777,N_779);
nor U879 (N_879,N_780,N_799);
nor U880 (N_880,N_774,N_776);
or U881 (N_881,N_818,N_805);
nand U882 (N_882,N_816,N_774);
nand U883 (N_883,N_759,N_804);
nor U884 (N_884,N_768,N_786);
nand U885 (N_885,N_777,N_786);
or U886 (N_886,N_783,N_784);
and U887 (N_887,N_755,N_770);
or U888 (N_888,N_789,N_779);
nand U889 (N_889,N_771,N_823);
nor U890 (N_890,N_770,N_758);
nor U891 (N_891,N_792,N_753);
nand U892 (N_892,N_760,N_755);
or U893 (N_893,N_752,N_795);
or U894 (N_894,N_801,N_802);
or U895 (N_895,N_785,N_819);
and U896 (N_896,N_817,N_818);
and U897 (N_897,N_768,N_757);
and U898 (N_898,N_776,N_794);
nand U899 (N_899,N_760,N_751);
or U900 (N_900,N_828,N_854);
or U901 (N_901,N_827,N_869);
nand U902 (N_902,N_836,N_832);
nor U903 (N_903,N_833,N_899);
nor U904 (N_904,N_826,N_852);
nand U905 (N_905,N_835,N_850);
nand U906 (N_906,N_845,N_890);
nand U907 (N_907,N_840,N_881);
or U908 (N_908,N_863,N_837);
nor U909 (N_909,N_887,N_853);
and U910 (N_910,N_864,N_848);
nor U911 (N_911,N_862,N_865);
nor U912 (N_912,N_880,N_896);
or U913 (N_913,N_866,N_860);
or U914 (N_914,N_898,N_851);
or U915 (N_915,N_859,N_868);
and U916 (N_916,N_849,N_886);
or U917 (N_917,N_882,N_858);
and U918 (N_918,N_897,N_876);
or U919 (N_919,N_861,N_844);
nand U920 (N_920,N_834,N_885);
nand U921 (N_921,N_889,N_838);
nor U922 (N_922,N_847,N_894);
or U923 (N_923,N_884,N_857);
or U924 (N_924,N_893,N_839);
or U925 (N_925,N_878,N_856);
or U926 (N_926,N_830,N_855);
nor U927 (N_927,N_825,N_891);
nor U928 (N_928,N_874,N_883);
or U929 (N_929,N_892,N_841);
nand U930 (N_930,N_843,N_873);
or U931 (N_931,N_870,N_831);
nand U932 (N_932,N_829,N_875);
nand U933 (N_933,N_867,N_895);
and U934 (N_934,N_879,N_871);
and U935 (N_935,N_842,N_846);
nor U936 (N_936,N_888,N_872);
and U937 (N_937,N_877,N_896);
nor U938 (N_938,N_856,N_832);
nor U939 (N_939,N_891,N_887);
nand U940 (N_940,N_842,N_861);
and U941 (N_941,N_857,N_850);
or U942 (N_942,N_849,N_879);
and U943 (N_943,N_858,N_889);
and U944 (N_944,N_856,N_855);
nand U945 (N_945,N_852,N_833);
nand U946 (N_946,N_885,N_841);
and U947 (N_947,N_834,N_835);
and U948 (N_948,N_874,N_846);
nor U949 (N_949,N_880,N_868);
nand U950 (N_950,N_846,N_859);
nor U951 (N_951,N_899,N_830);
and U952 (N_952,N_830,N_865);
or U953 (N_953,N_839,N_845);
nand U954 (N_954,N_856,N_853);
nand U955 (N_955,N_835,N_891);
or U956 (N_956,N_872,N_882);
and U957 (N_957,N_871,N_840);
nor U958 (N_958,N_889,N_841);
nor U959 (N_959,N_861,N_849);
and U960 (N_960,N_897,N_884);
or U961 (N_961,N_851,N_877);
and U962 (N_962,N_829,N_885);
nand U963 (N_963,N_852,N_876);
nor U964 (N_964,N_858,N_877);
and U965 (N_965,N_887,N_845);
nor U966 (N_966,N_848,N_836);
or U967 (N_967,N_839,N_826);
nor U968 (N_968,N_899,N_856);
or U969 (N_969,N_856,N_854);
nand U970 (N_970,N_850,N_831);
nand U971 (N_971,N_860,N_862);
nor U972 (N_972,N_868,N_863);
or U973 (N_973,N_859,N_873);
and U974 (N_974,N_828,N_869);
nor U975 (N_975,N_934,N_938);
nor U976 (N_976,N_946,N_922);
or U977 (N_977,N_963,N_929);
nor U978 (N_978,N_957,N_917);
nor U979 (N_979,N_926,N_940);
nor U980 (N_980,N_918,N_936);
nor U981 (N_981,N_939,N_967);
or U982 (N_982,N_949,N_928);
xnor U983 (N_983,N_916,N_974);
nor U984 (N_984,N_943,N_962);
nor U985 (N_985,N_951,N_968);
nor U986 (N_986,N_956,N_921);
nand U987 (N_987,N_901,N_900);
nand U988 (N_988,N_955,N_958);
or U989 (N_989,N_903,N_902);
or U990 (N_990,N_920,N_945);
and U991 (N_991,N_964,N_947);
nor U992 (N_992,N_919,N_966);
nand U993 (N_993,N_930,N_971);
nor U994 (N_994,N_914,N_935);
nand U995 (N_995,N_909,N_954);
and U996 (N_996,N_944,N_904);
nand U997 (N_997,N_965,N_959);
nor U998 (N_998,N_931,N_913);
and U999 (N_999,N_960,N_911);
or U1000 (N_1000,N_933,N_953);
nor U1001 (N_1001,N_961,N_923);
nor U1002 (N_1002,N_969,N_941);
nand U1003 (N_1003,N_924,N_932);
nor U1004 (N_1004,N_937,N_912);
or U1005 (N_1005,N_910,N_973);
and U1006 (N_1006,N_952,N_942);
and U1007 (N_1007,N_906,N_950);
or U1008 (N_1008,N_925,N_948);
nand U1009 (N_1009,N_908,N_970);
nor U1010 (N_1010,N_907,N_927);
nor U1011 (N_1011,N_905,N_972);
nor U1012 (N_1012,N_915,N_920);
and U1013 (N_1013,N_942,N_967);
or U1014 (N_1014,N_911,N_944);
and U1015 (N_1015,N_967,N_917);
nor U1016 (N_1016,N_901,N_954);
or U1017 (N_1017,N_924,N_965);
and U1018 (N_1018,N_907,N_913);
nand U1019 (N_1019,N_921,N_938);
or U1020 (N_1020,N_953,N_949);
nor U1021 (N_1021,N_903,N_932);
and U1022 (N_1022,N_946,N_957);
nand U1023 (N_1023,N_963,N_956);
nand U1024 (N_1024,N_960,N_916);
nand U1025 (N_1025,N_918,N_970);
or U1026 (N_1026,N_937,N_953);
nand U1027 (N_1027,N_958,N_910);
nand U1028 (N_1028,N_903,N_951);
or U1029 (N_1029,N_906,N_939);
xnor U1030 (N_1030,N_911,N_916);
nor U1031 (N_1031,N_945,N_939);
nor U1032 (N_1032,N_908,N_959);
or U1033 (N_1033,N_967,N_956);
nand U1034 (N_1034,N_926,N_920);
nand U1035 (N_1035,N_921,N_957);
and U1036 (N_1036,N_966,N_905);
or U1037 (N_1037,N_939,N_942);
and U1038 (N_1038,N_954,N_939);
and U1039 (N_1039,N_970,N_906);
and U1040 (N_1040,N_954,N_968);
nor U1041 (N_1041,N_964,N_914);
nor U1042 (N_1042,N_909,N_972);
or U1043 (N_1043,N_966,N_915);
nand U1044 (N_1044,N_928,N_914);
nand U1045 (N_1045,N_932,N_906);
or U1046 (N_1046,N_944,N_946);
and U1047 (N_1047,N_907,N_955);
nor U1048 (N_1048,N_920,N_961);
or U1049 (N_1049,N_937,N_936);
or U1050 (N_1050,N_1029,N_999);
and U1051 (N_1051,N_1018,N_1033);
and U1052 (N_1052,N_1048,N_1049);
or U1053 (N_1053,N_1013,N_1035);
nor U1054 (N_1054,N_978,N_1043);
and U1055 (N_1055,N_998,N_985);
and U1056 (N_1056,N_1017,N_1000);
and U1057 (N_1057,N_981,N_980);
or U1058 (N_1058,N_1001,N_1028);
or U1059 (N_1059,N_982,N_984);
nor U1060 (N_1060,N_1002,N_1004);
nand U1061 (N_1061,N_992,N_989);
and U1062 (N_1062,N_1036,N_1006);
nand U1063 (N_1063,N_1020,N_1009);
nand U1064 (N_1064,N_1044,N_1015);
nand U1065 (N_1065,N_983,N_979);
or U1066 (N_1066,N_1024,N_1026);
and U1067 (N_1067,N_1007,N_977);
or U1068 (N_1068,N_976,N_1039);
nor U1069 (N_1069,N_993,N_1019);
nor U1070 (N_1070,N_991,N_1038);
nand U1071 (N_1071,N_1037,N_995);
nor U1072 (N_1072,N_990,N_1023);
or U1073 (N_1073,N_1008,N_1032);
and U1074 (N_1074,N_975,N_1010);
nor U1075 (N_1075,N_1041,N_1025);
xnor U1076 (N_1076,N_1045,N_994);
or U1077 (N_1077,N_1042,N_1027);
or U1078 (N_1078,N_1040,N_1034);
or U1079 (N_1079,N_1022,N_996);
or U1080 (N_1080,N_1014,N_1012);
nand U1081 (N_1081,N_1047,N_1031);
nor U1082 (N_1082,N_987,N_988);
nor U1083 (N_1083,N_986,N_997);
nand U1084 (N_1084,N_1005,N_1021);
nand U1085 (N_1085,N_1046,N_1030);
nor U1086 (N_1086,N_1003,N_1011);
and U1087 (N_1087,N_1016,N_997);
or U1088 (N_1088,N_982,N_990);
or U1089 (N_1089,N_990,N_975);
or U1090 (N_1090,N_1005,N_1030);
and U1091 (N_1091,N_1002,N_1035);
nor U1092 (N_1092,N_1033,N_1026);
and U1093 (N_1093,N_1021,N_998);
and U1094 (N_1094,N_995,N_1020);
and U1095 (N_1095,N_1024,N_1033);
nor U1096 (N_1096,N_1016,N_1011);
or U1097 (N_1097,N_979,N_991);
nor U1098 (N_1098,N_993,N_994);
or U1099 (N_1099,N_992,N_1007);
nor U1100 (N_1100,N_989,N_1013);
nor U1101 (N_1101,N_1011,N_978);
or U1102 (N_1102,N_991,N_1021);
and U1103 (N_1103,N_1022,N_1006);
nor U1104 (N_1104,N_1020,N_1033);
xnor U1105 (N_1105,N_1000,N_982);
nor U1106 (N_1106,N_1030,N_975);
or U1107 (N_1107,N_1030,N_1012);
nor U1108 (N_1108,N_990,N_1027);
or U1109 (N_1109,N_976,N_1010);
nor U1110 (N_1110,N_1042,N_989);
nor U1111 (N_1111,N_1019,N_978);
or U1112 (N_1112,N_995,N_1048);
nor U1113 (N_1113,N_995,N_987);
or U1114 (N_1114,N_1037,N_1031);
and U1115 (N_1115,N_1031,N_977);
nand U1116 (N_1116,N_1014,N_1022);
and U1117 (N_1117,N_1029,N_1049);
xor U1118 (N_1118,N_1032,N_986);
nor U1119 (N_1119,N_1039,N_1019);
or U1120 (N_1120,N_976,N_1042);
or U1121 (N_1121,N_1044,N_1013);
or U1122 (N_1122,N_1026,N_982);
nand U1123 (N_1123,N_1022,N_1042);
or U1124 (N_1124,N_1006,N_1021);
nand U1125 (N_1125,N_1074,N_1095);
nor U1126 (N_1126,N_1111,N_1070);
nand U1127 (N_1127,N_1098,N_1094);
or U1128 (N_1128,N_1101,N_1088);
and U1129 (N_1129,N_1081,N_1115);
or U1130 (N_1130,N_1113,N_1075);
nand U1131 (N_1131,N_1112,N_1064);
nor U1132 (N_1132,N_1053,N_1103);
or U1133 (N_1133,N_1071,N_1073);
and U1134 (N_1134,N_1124,N_1080);
nand U1135 (N_1135,N_1086,N_1120);
or U1136 (N_1136,N_1057,N_1051);
or U1137 (N_1137,N_1052,N_1059);
nor U1138 (N_1138,N_1092,N_1060);
nor U1139 (N_1139,N_1105,N_1078);
nand U1140 (N_1140,N_1106,N_1056);
nand U1141 (N_1141,N_1109,N_1087);
nor U1142 (N_1142,N_1099,N_1076);
or U1143 (N_1143,N_1114,N_1108);
nor U1144 (N_1144,N_1055,N_1072);
nand U1145 (N_1145,N_1079,N_1066);
nand U1146 (N_1146,N_1091,N_1118);
nand U1147 (N_1147,N_1062,N_1117);
or U1148 (N_1148,N_1083,N_1107);
or U1149 (N_1149,N_1082,N_1093);
nor U1150 (N_1150,N_1054,N_1084);
nand U1151 (N_1151,N_1069,N_1061);
nand U1152 (N_1152,N_1100,N_1085);
and U1153 (N_1153,N_1089,N_1116);
nor U1154 (N_1154,N_1077,N_1058);
nand U1155 (N_1155,N_1110,N_1123);
nand U1156 (N_1156,N_1104,N_1121);
nand U1157 (N_1157,N_1065,N_1063);
nand U1158 (N_1158,N_1096,N_1097);
nand U1159 (N_1159,N_1068,N_1050);
or U1160 (N_1160,N_1067,N_1122);
or U1161 (N_1161,N_1102,N_1119);
nand U1162 (N_1162,N_1090,N_1072);
and U1163 (N_1163,N_1071,N_1106);
and U1164 (N_1164,N_1078,N_1068);
nor U1165 (N_1165,N_1085,N_1054);
or U1166 (N_1166,N_1081,N_1052);
and U1167 (N_1167,N_1091,N_1102);
nor U1168 (N_1168,N_1075,N_1062);
and U1169 (N_1169,N_1096,N_1120);
or U1170 (N_1170,N_1053,N_1089);
nand U1171 (N_1171,N_1091,N_1076);
nand U1172 (N_1172,N_1088,N_1054);
nor U1173 (N_1173,N_1089,N_1119);
and U1174 (N_1174,N_1123,N_1096);
and U1175 (N_1175,N_1116,N_1062);
or U1176 (N_1176,N_1075,N_1076);
or U1177 (N_1177,N_1054,N_1097);
and U1178 (N_1178,N_1090,N_1076);
or U1179 (N_1179,N_1114,N_1062);
or U1180 (N_1180,N_1069,N_1055);
nand U1181 (N_1181,N_1105,N_1077);
nor U1182 (N_1182,N_1085,N_1050);
and U1183 (N_1183,N_1122,N_1066);
nor U1184 (N_1184,N_1085,N_1073);
or U1185 (N_1185,N_1059,N_1099);
or U1186 (N_1186,N_1072,N_1118);
xnor U1187 (N_1187,N_1061,N_1067);
or U1188 (N_1188,N_1104,N_1051);
nor U1189 (N_1189,N_1082,N_1109);
nand U1190 (N_1190,N_1065,N_1060);
nand U1191 (N_1191,N_1102,N_1120);
nand U1192 (N_1192,N_1084,N_1073);
nand U1193 (N_1193,N_1057,N_1114);
nor U1194 (N_1194,N_1080,N_1099);
and U1195 (N_1195,N_1109,N_1095);
nand U1196 (N_1196,N_1055,N_1105);
nand U1197 (N_1197,N_1098,N_1084);
nand U1198 (N_1198,N_1089,N_1050);
and U1199 (N_1199,N_1100,N_1078);
or U1200 (N_1200,N_1134,N_1171);
or U1201 (N_1201,N_1127,N_1177);
nor U1202 (N_1202,N_1142,N_1180);
and U1203 (N_1203,N_1149,N_1150);
nor U1204 (N_1204,N_1182,N_1199);
nor U1205 (N_1205,N_1170,N_1187);
or U1206 (N_1206,N_1144,N_1139);
nor U1207 (N_1207,N_1190,N_1135);
nor U1208 (N_1208,N_1140,N_1146);
or U1209 (N_1209,N_1175,N_1188);
or U1210 (N_1210,N_1183,N_1186);
nand U1211 (N_1211,N_1198,N_1130);
nand U1212 (N_1212,N_1158,N_1131);
or U1213 (N_1213,N_1189,N_1191);
nor U1214 (N_1214,N_1197,N_1185);
nor U1215 (N_1215,N_1152,N_1128);
nand U1216 (N_1216,N_1161,N_1181);
or U1217 (N_1217,N_1153,N_1166);
xnor U1218 (N_1218,N_1138,N_1163);
nand U1219 (N_1219,N_1143,N_1145);
and U1220 (N_1220,N_1169,N_1174);
or U1221 (N_1221,N_1164,N_1132);
and U1222 (N_1222,N_1172,N_1194);
nor U1223 (N_1223,N_1156,N_1184);
nand U1224 (N_1224,N_1195,N_1193);
nor U1225 (N_1225,N_1155,N_1179);
nor U1226 (N_1226,N_1129,N_1159);
and U1227 (N_1227,N_1157,N_1196);
or U1228 (N_1228,N_1192,N_1165);
nand U1229 (N_1229,N_1148,N_1133);
or U1230 (N_1230,N_1126,N_1136);
nand U1231 (N_1231,N_1154,N_1162);
or U1232 (N_1232,N_1173,N_1141);
nor U1233 (N_1233,N_1160,N_1176);
nor U1234 (N_1234,N_1151,N_1147);
nand U1235 (N_1235,N_1167,N_1178);
and U1236 (N_1236,N_1125,N_1168);
nand U1237 (N_1237,N_1137,N_1183);
nand U1238 (N_1238,N_1161,N_1178);
nor U1239 (N_1239,N_1140,N_1176);
and U1240 (N_1240,N_1171,N_1184);
nor U1241 (N_1241,N_1133,N_1168);
and U1242 (N_1242,N_1170,N_1131);
nand U1243 (N_1243,N_1160,N_1192);
xnor U1244 (N_1244,N_1161,N_1154);
and U1245 (N_1245,N_1125,N_1166);
or U1246 (N_1246,N_1173,N_1133);
and U1247 (N_1247,N_1166,N_1191);
and U1248 (N_1248,N_1141,N_1195);
and U1249 (N_1249,N_1170,N_1181);
nand U1250 (N_1250,N_1189,N_1183);
or U1251 (N_1251,N_1176,N_1188);
or U1252 (N_1252,N_1195,N_1159);
nand U1253 (N_1253,N_1140,N_1150);
nand U1254 (N_1254,N_1134,N_1183);
or U1255 (N_1255,N_1151,N_1186);
nor U1256 (N_1256,N_1136,N_1164);
nor U1257 (N_1257,N_1151,N_1175);
nand U1258 (N_1258,N_1147,N_1173);
or U1259 (N_1259,N_1132,N_1133);
or U1260 (N_1260,N_1172,N_1153);
or U1261 (N_1261,N_1175,N_1196);
and U1262 (N_1262,N_1157,N_1165);
or U1263 (N_1263,N_1173,N_1153);
nand U1264 (N_1264,N_1182,N_1180);
nor U1265 (N_1265,N_1184,N_1195);
or U1266 (N_1266,N_1190,N_1164);
and U1267 (N_1267,N_1136,N_1150);
nor U1268 (N_1268,N_1147,N_1172);
nand U1269 (N_1269,N_1143,N_1141);
xnor U1270 (N_1270,N_1152,N_1178);
or U1271 (N_1271,N_1139,N_1161);
nand U1272 (N_1272,N_1193,N_1125);
or U1273 (N_1273,N_1161,N_1136);
nand U1274 (N_1274,N_1156,N_1197);
or U1275 (N_1275,N_1273,N_1251);
or U1276 (N_1276,N_1258,N_1272);
nor U1277 (N_1277,N_1266,N_1222);
and U1278 (N_1278,N_1229,N_1243);
or U1279 (N_1279,N_1238,N_1225);
and U1280 (N_1280,N_1201,N_1226);
or U1281 (N_1281,N_1255,N_1202);
nor U1282 (N_1282,N_1260,N_1211);
nor U1283 (N_1283,N_1264,N_1268);
or U1284 (N_1284,N_1246,N_1271);
nor U1285 (N_1285,N_1207,N_1205);
or U1286 (N_1286,N_1249,N_1269);
or U1287 (N_1287,N_1237,N_1233);
xnor U1288 (N_1288,N_1239,N_1256);
nor U1289 (N_1289,N_1245,N_1247);
nor U1290 (N_1290,N_1230,N_1223);
and U1291 (N_1291,N_1244,N_1265);
nor U1292 (N_1292,N_1234,N_1210);
and U1293 (N_1293,N_1216,N_1212);
xnor U1294 (N_1294,N_1270,N_1267);
nor U1295 (N_1295,N_1263,N_1227);
nor U1296 (N_1296,N_1209,N_1203);
nand U1297 (N_1297,N_1218,N_1206);
or U1298 (N_1298,N_1231,N_1252);
nor U1299 (N_1299,N_1214,N_1242);
or U1300 (N_1300,N_1254,N_1228);
or U1301 (N_1301,N_1215,N_1217);
nand U1302 (N_1302,N_1208,N_1261);
nor U1303 (N_1303,N_1262,N_1224);
and U1304 (N_1304,N_1248,N_1241);
or U1305 (N_1305,N_1200,N_1219);
and U1306 (N_1306,N_1220,N_1259);
and U1307 (N_1307,N_1250,N_1213);
nand U1308 (N_1308,N_1204,N_1240);
nor U1309 (N_1309,N_1236,N_1221);
nor U1310 (N_1310,N_1235,N_1253);
nand U1311 (N_1311,N_1274,N_1232);
nand U1312 (N_1312,N_1257,N_1219);
nand U1313 (N_1313,N_1255,N_1201);
and U1314 (N_1314,N_1228,N_1223);
or U1315 (N_1315,N_1236,N_1271);
nor U1316 (N_1316,N_1250,N_1270);
nand U1317 (N_1317,N_1204,N_1272);
or U1318 (N_1318,N_1272,N_1212);
and U1319 (N_1319,N_1266,N_1215);
or U1320 (N_1320,N_1220,N_1200);
and U1321 (N_1321,N_1249,N_1204);
nand U1322 (N_1322,N_1202,N_1272);
nand U1323 (N_1323,N_1200,N_1208);
or U1324 (N_1324,N_1242,N_1205);
nor U1325 (N_1325,N_1237,N_1213);
nand U1326 (N_1326,N_1228,N_1214);
nor U1327 (N_1327,N_1212,N_1262);
and U1328 (N_1328,N_1273,N_1215);
nor U1329 (N_1329,N_1259,N_1252);
nor U1330 (N_1330,N_1220,N_1256);
or U1331 (N_1331,N_1260,N_1257);
nand U1332 (N_1332,N_1207,N_1235);
nor U1333 (N_1333,N_1237,N_1216);
nor U1334 (N_1334,N_1230,N_1201);
nand U1335 (N_1335,N_1250,N_1268);
or U1336 (N_1336,N_1263,N_1238);
and U1337 (N_1337,N_1211,N_1231);
or U1338 (N_1338,N_1210,N_1207);
or U1339 (N_1339,N_1259,N_1236);
nor U1340 (N_1340,N_1201,N_1222);
and U1341 (N_1341,N_1242,N_1266);
and U1342 (N_1342,N_1231,N_1219);
and U1343 (N_1343,N_1230,N_1202);
nor U1344 (N_1344,N_1239,N_1272);
and U1345 (N_1345,N_1203,N_1272);
or U1346 (N_1346,N_1207,N_1263);
or U1347 (N_1347,N_1272,N_1245);
nand U1348 (N_1348,N_1266,N_1214);
or U1349 (N_1349,N_1246,N_1201);
or U1350 (N_1350,N_1319,N_1326);
nor U1351 (N_1351,N_1317,N_1310);
and U1352 (N_1352,N_1345,N_1299);
nand U1353 (N_1353,N_1331,N_1278);
xor U1354 (N_1354,N_1304,N_1302);
or U1355 (N_1355,N_1292,N_1307);
nand U1356 (N_1356,N_1281,N_1330);
or U1357 (N_1357,N_1327,N_1286);
or U1358 (N_1358,N_1334,N_1347);
and U1359 (N_1359,N_1283,N_1335);
nand U1360 (N_1360,N_1322,N_1296);
or U1361 (N_1361,N_1341,N_1287);
nand U1362 (N_1362,N_1294,N_1324);
and U1363 (N_1363,N_1314,N_1289);
nand U1364 (N_1364,N_1343,N_1291);
and U1365 (N_1365,N_1320,N_1306);
nor U1366 (N_1366,N_1311,N_1333);
nor U1367 (N_1367,N_1346,N_1280);
nor U1368 (N_1368,N_1329,N_1305);
or U1369 (N_1369,N_1275,N_1279);
xor U1370 (N_1370,N_1316,N_1309);
and U1371 (N_1371,N_1321,N_1290);
nor U1372 (N_1372,N_1318,N_1312);
or U1373 (N_1373,N_1338,N_1323);
xor U1374 (N_1374,N_1297,N_1298);
nand U1375 (N_1375,N_1340,N_1313);
nor U1376 (N_1376,N_1293,N_1288);
and U1377 (N_1377,N_1277,N_1339);
nand U1378 (N_1378,N_1308,N_1349);
and U1379 (N_1379,N_1328,N_1337);
nand U1380 (N_1380,N_1301,N_1344);
and U1381 (N_1381,N_1284,N_1325);
nor U1382 (N_1382,N_1285,N_1315);
nand U1383 (N_1383,N_1276,N_1303);
and U1384 (N_1384,N_1336,N_1348);
or U1385 (N_1385,N_1300,N_1295);
or U1386 (N_1386,N_1332,N_1282);
nand U1387 (N_1387,N_1342,N_1312);
and U1388 (N_1388,N_1329,N_1324);
nand U1389 (N_1389,N_1338,N_1307);
nand U1390 (N_1390,N_1309,N_1349);
nand U1391 (N_1391,N_1316,N_1283);
nor U1392 (N_1392,N_1316,N_1339);
nand U1393 (N_1393,N_1328,N_1314);
nand U1394 (N_1394,N_1310,N_1299);
or U1395 (N_1395,N_1276,N_1345);
and U1396 (N_1396,N_1312,N_1336);
or U1397 (N_1397,N_1319,N_1308);
and U1398 (N_1398,N_1283,N_1293);
or U1399 (N_1399,N_1277,N_1343);
and U1400 (N_1400,N_1329,N_1340);
nor U1401 (N_1401,N_1329,N_1286);
and U1402 (N_1402,N_1299,N_1342);
nor U1403 (N_1403,N_1285,N_1342);
and U1404 (N_1404,N_1314,N_1339);
nand U1405 (N_1405,N_1349,N_1334);
nor U1406 (N_1406,N_1295,N_1297);
or U1407 (N_1407,N_1320,N_1338);
nor U1408 (N_1408,N_1328,N_1318);
or U1409 (N_1409,N_1296,N_1328);
and U1410 (N_1410,N_1284,N_1324);
nor U1411 (N_1411,N_1331,N_1321);
nand U1412 (N_1412,N_1278,N_1300);
nor U1413 (N_1413,N_1278,N_1316);
or U1414 (N_1414,N_1344,N_1318);
or U1415 (N_1415,N_1282,N_1306);
or U1416 (N_1416,N_1307,N_1329);
or U1417 (N_1417,N_1307,N_1275);
and U1418 (N_1418,N_1348,N_1292);
nor U1419 (N_1419,N_1299,N_1280);
and U1420 (N_1420,N_1283,N_1286);
and U1421 (N_1421,N_1325,N_1296);
or U1422 (N_1422,N_1337,N_1311);
nor U1423 (N_1423,N_1278,N_1297);
nand U1424 (N_1424,N_1317,N_1279);
or U1425 (N_1425,N_1369,N_1422);
or U1426 (N_1426,N_1378,N_1421);
nor U1427 (N_1427,N_1408,N_1368);
nand U1428 (N_1428,N_1400,N_1403);
and U1429 (N_1429,N_1398,N_1383);
nor U1430 (N_1430,N_1373,N_1379);
or U1431 (N_1431,N_1364,N_1393);
and U1432 (N_1432,N_1399,N_1370);
or U1433 (N_1433,N_1394,N_1380);
and U1434 (N_1434,N_1356,N_1375);
or U1435 (N_1435,N_1423,N_1365);
or U1436 (N_1436,N_1376,N_1396);
nand U1437 (N_1437,N_1377,N_1412);
nor U1438 (N_1438,N_1414,N_1417);
nand U1439 (N_1439,N_1374,N_1361);
nand U1440 (N_1440,N_1415,N_1387);
nor U1441 (N_1441,N_1418,N_1351);
and U1442 (N_1442,N_1366,N_1367);
nor U1443 (N_1443,N_1363,N_1388);
nand U1444 (N_1444,N_1359,N_1409);
nor U1445 (N_1445,N_1372,N_1362);
or U1446 (N_1446,N_1401,N_1410);
nor U1447 (N_1447,N_1371,N_1352);
and U1448 (N_1448,N_1402,N_1407);
and U1449 (N_1449,N_1353,N_1355);
nor U1450 (N_1450,N_1420,N_1360);
or U1451 (N_1451,N_1385,N_1358);
nand U1452 (N_1452,N_1397,N_1386);
nor U1453 (N_1453,N_1419,N_1390);
nor U1454 (N_1454,N_1389,N_1413);
nor U1455 (N_1455,N_1350,N_1406);
nor U1456 (N_1456,N_1354,N_1391);
nand U1457 (N_1457,N_1411,N_1404);
and U1458 (N_1458,N_1381,N_1382);
and U1459 (N_1459,N_1405,N_1416);
and U1460 (N_1460,N_1424,N_1357);
nor U1461 (N_1461,N_1395,N_1384);
and U1462 (N_1462,N_1392,N_1388);
nor U1463 (N_1463,N_1367,N_1419);
nor U1464 (N_1464,N_1362,N_1417);
and U1465 (N_1465,N_1389,N_1419);
nor U1466 (N_1466,N_1387,N_1382);
nor U1467 (N_1467,N_1381,N_1395);
nand U1468 (N_1468,N_1404,N_1367);
nand U1469 (N_1469,N_1356,N_1415);
xnor U1470 (N_1470,N_1376,N_1361);
or U1471 (N_1471,N_1404,N_1380);
and U1472 (N_1472,N_1379,N_1415);
nor U1473 (N_1473,N_1390,N_1382);
and U1474 (N_1474,N_1412,N_1352);
or U1475 (N_1475,N_1361,N_1397);
or U1476 (N_1476,N_1421,N_1389);
nor U1477 (N_1477,N_1421,N_1394);
nand U1478 (N_1478,N_1393,N_1361);
and U1479 (N_1479,N_1369,N_1377);
and U1480 (N_1480,N_1390,N_1408);
nor U1481 (N_1481,N_1364,N_1419);
nand U1482 (N_1482,N_1412,N_1395);
nor U1483 (N_1483,N_1357,N_1422);
nand U1484 (N_1484,N_1366,N_1382);
nor U1485 (N_1485,N_1368,N_1366);
nor U1486 (N_1486,N_1373,N_1354);
nand U1487 (N_1487,N_1381,N_1407);
nor U1488 (N_1488,N_1350,N_1391);
and U1489 (N_1489,N_1367,N_1394);
or U1490 (N_1490,N_1423,N_1363);
nand U1491 (N_1491,N_1366,N_1413);
nor U1492 (N_1492,N_1403,N_1399);
or U1493 (N_1493,N_1410,N_1376);
nor U1494 (N_1494,N_1400,N_1368);
nand U1495 (N_1495,N_1377,N_1374);
or U1496 (N_1496,N_1394,N_1388);
nand U1497 (N_1497,N_1360,N_1419);
or U1498 (N_1498,N_1401,N_1391);
and U1499 (N_1499,N_1398,N_1387);
or U1500 (N_1500,N_1434,N_1463);
or U1501 (N_1501,N_1447,N_1499);
or U1502 (N_1502,N_1481,N_1487);
and U1503 (N_1503,N_1427,N_1438);
nor U1504 (N_1504,N_1443,N_1457);
or U1505 (N_1505,N_1453,N_1454);
and U1506 (N_1506,N_1440,N_1477);
nor U1507 (N_1507,N_1426,N_1444);
nand U1508 (N_1508,N_1436,N_1435);
or U1509 (N_1509,N_1471,N_1425);
or U1510 (N_1510,N_1466,N_1489);
and U1511 (N_1511,N_1482,N_1461);
and U1512 (N_1512,N_1468,N_1429);
and U1513 (N_1513,N_1448,N_1492);
and U1514 (N_1514,N_1475,N_1498);
nor U1515 (N_1515,N_1451,N_1437);
or U1516 (N_1516,N_1449,N_1470);
and U1517 (N_1517,N_1464,N_1491);
or U1518 (N_1518,N_1497,N_1459);
nand U1519 (N_1519,N_1479,N_1467);
and U1520 (N_1520,N_1476,N_1432);
and U1521 (N_1521,N_1460,N_1495);
or U1522 (N_1522,N_1465,N_1452);
nor U1523 (N_1523,N_1490,N_1469);
nor U1524 (N_1524,N_1456,N_1493);
nor U1525 (N_1525,N_1484,N_1439);
or U1526 (N_1526,N_1446,N_1433);
nand U1527 (N_1527,N_1483,N_1472);
or U1528 (N_1528,N_1441,N_1428);
or U1529 (N_1529,N_1480,N_1473);
and U1530 (N_1530,N_1442,N_1450);
nor U1531 (N_1531,N_1474,N_1478);
or U1532 (N_1532,N_1486,N_1458);
xor U1533 (N_1533,N_1462,N_1445);
and U1534 (N_1534,N_1496,N_1430);
nand U1535 (N_1535,N_1494,N_1488);
nand U1536 (N_1536,N_1431,N_1455);
nand U1537 (N_1537,N_1485,N_1492);
nor U1538 (N_1538,N_1447,N_1426);
nand U1539 (N_1539,N_1481,N_1459);
nor U1540 (N_1540,N_1477,N_1456);
and U1541 (N_1541,N_1430,N_1482);
or U1542 (N_1542,N_1445,N_1430);
nor U1543 (N_1543,N_1498,N_1495);
and U1544 (N_1544,N_1464,N_1490);
nand U1545 (N_1545,N_1480,N_1434);
and U1546 (N_1546,N_1481,N_1478);
nand U1547 (N_1547,N_1444,N_1484);
nand U1548 (N_1548,N_1470,N_1474);
nand U1549 (N_1549,N_1499,N_1451);
and U1550 (N_1550,N_1487,N_1486);
and U1551 (N_1551,N_1427,N_1453);
or U1552 (N_1552,N_1457,N_1442);
nand U1553 (N_1553,N_1467,N_1440);
and U1554 (N_1554,N_1433,N_1436);
nor U1555 (N_1555,N_1490,N_1467);
and U1556 (N_1556,N_1446,N_1472);
or U1557 (N_1557,N_1470,N_1489);
nor U1558 (N_1558,N_1441,N_1438);
nor U1559 (N_1559,N_1490,N_1448);
nor U1560 (N_1560,N_1449,N_1451);
nor U1561 (N_1561,N_1445,N_1425);
or U1562 (N_1562,N_1454,N_1465);
nand U1563 (N_1563,N_1456,N_1484);
and U1564 (N_1564,N_1430,N_1441);
nand U1565 (N_1565,N_1497,N_1484);
and U1566 (N_1566,N_1443,N_1451);
and U1567 (N_1567,N_1475,N_1478);
nor U1568 (N_1568,N_1458,N_1482);
and U1569 (N_1569,N_1425,N_1489);
or U1570 (N_1570,N_1497,N_1429);
or U1571 (N_1571,N_1462,N_1449);
nor U1572 (N_1572,N_1498,N_1477);
and U1573 (N_1573,N_1471,N_1495);
and U1574 (N_1574,N_1440,N_1448);
nand U1575 (N_1575,N_1509,N_1503);
nor U1576 (N_1576,N_1513,N_1567);
nor U1577 (N_1577,N_1540,N_1520);
nor U1578 (N_1578,N_1544,N_1512);
nor U1579 (N_1579,N_1572,N_1510);
or U1580 (N_1580,N_1505,N_1531);
or U1581 (N_1581,N_1500,N_1501);
nand U1582 (N_1582,N_1553,N_1534);
nor U1583 (N_1583,N_1557,N_1573);
or U1584 (N_1584,N_1564,N_1537);
nor U1585 (N_1585,N_1522,N_1547);
nand U1586 (N_1586,N_1527,N_1511);
nand U1587 (N_1587,N_1515,N_1551);
nor U1588 (N_1588,N_1539,N_1568);
nand U1589 (N_1589,N_1570,N_1523);
or U1590 (N_1590,N_1514,N_1525);
or U1591 (N_1591,N_1552,N_1566);
or U1592 (N_1592,N_1518,N_1508);
or U1593 (N_1593,N_1550,N_1536);
nand U1594 (N_1594,N_1563,N_1526);
or U1595 (N_1595,N_1565,N_1530);
and U1596 (N_1596,N_1554,N_1504);
and U1597 (N_1597,N_1546,N_1524);
and U1598 (N_1598,N_1556,N_1533);
nand U1599 (N_1599,N_1528,N_1562);
nor U1600 (N_1600,N_1569,N_1506);
nor U1601 (N_1601,N_1574,N_1532);
and U1602 (N_1602,N_1502,N_1548);
nand U1603 (N_1603,N_1558,N_1561);
or U1604 (N_1604,N_1521,N_1545);
nor U1605 (N_1605,N_1555,N_1516);
or U1606 (N_1606,N_1541,N_1507);
and U1607 (N_1607,N_1519,N_1560);
and U1608 (N_1608,N_1535,N_1549);
nor U1609 (N_1609,N_1517,N_1529);
nand U1610 (N_1610,N_1542,N_1571);
or U1611 (N_1611,N_1559,N_1543);
nor U1612 (N_1612,N_1538,N_1551);
and U1613 (N_1613,N_1514,N_1521);
and U1614 (N_1614,N_1507,N_1571);
nor U1615 (N_1615,N_1568,N_1549);
nand U1616 (N_1616,N_1512,N_1540);
or U1617 (N_1617,N_1559,N_1520);
nand U1618 (N_1618,N_1515,N_1506);
or U1619 (N_1619,N_1574,N_1572);
and U1620 (N_1620,N_1532,N_1542);
and U1621 (N_1621,N_1538,N_1545);
nand U1622 (N_1622,N_1540,N_1522);
nor U1623 (N_1623,N_1505,N_1507);
xnor U1624 (N_1624,N_1537,N_1531);
nand U1625 (N_1625,N_1559,N_1566);
or U1626 (N_1626,N_1506,N_1517);
or U1627 (N_1627,N_1506,N_1563);
or U1628 (N_1628,N_1516,N_1528);
nor U1629 (N_1629,N_1544,N_1533);
or U1630 (N_1630,N_1544,N_1557);
nand U1631 (N_1631,N_1503,N_1534);
nor U1632 (N_1632,N_1519,N_1544);
and U1633 (N_1633,N_1514,N_1524);
nor U1634 (N_1634,N_1502,N_1517);
nand U1635 (N_1635,N_1509,N_1553);
and U1636 (N_1636,N_1566,N_1500);
nor U1637 (N_1637,N_1521,N_1502);
nor U1638 (N_1638,N_1517,N_1501);
or U1639 (N_1639,N_1507,N_1533);
and U1640 (N_1640,N_1542,N_1502);
nand U1641 (N_1641,N_1545,N_1564);
or U1642 (N_1642,N_1539,N_1551);
nor U1643 (N_1643,N_1568,N_1538);
nand U1644 (N_1644,N_1569,N_1566);
or U1645 (N_1645,N_1566,N_1506);
nand U1646 (N_1646,N_1542,N_1556);
or U1647 (N_1647,N_1509,N_1563);
nor U1648 (N_1648,N_1568,N_1574);
nor U1649 (N_1649,N_1545,N_1515);
nand U1650 (N_1650,N_1640,N_1586);
and U1651 (N_1651,N_1649,N_1577);
nor U1652 (N_1652,N_1608,N_1625);
nor U1653 (N_1653,N_1589,N_1618);
nand U1654 (N_1654,N_1639,N_1592);
nand U1655 (N_1655,N_1588,N_1576);
nand U1656 (N_1656,N_1609,N_1591);
nor U1657 (N_1657,N_1648,N_1634);
nand U1658 (N_1658,N_1602,N_1644);
or U1659 (N_1659,N_1616,N_1647);
and U1660 (N_1660,N_1624,N_1642);
nor U1661 (N_1661,N_1580,N_1581);
nand U1662 (N_1662,N_1621,N_1632);
nor U1663 (N_1663,N_1627,N_1575);
nand U1664 (N_1664,N_1617,N_1637);
xnor U1665 (N_1665,N_1645,N_1596);
or U1666 (N_1666,N_1643,N_1610);
nand U1667 (N_1667,N_1604,N_1638);
and U1668 (N_1668,N_1614,N_1623);
or U1669 (N_1669,N_1612,N_1629);
nor U1670 (N_1670,N_1628,N_1585);
nand U1671 (N_1671,N_1626,N_1594);
or U1672 (N_1672,N_1598,N_1606);
nor U1673 (N_1673,N_1600,N_1605);
nor U1674 (N_1674,N_1597,N_1619);
nand U1675 (N_1675,N_1584,N_1613);
nand U1676 (N_1676,N_1615,N_1646);
nand U1677 (N_1677,N_1590,N_1607);
and U1678 (N_1678,N_1603,N_1595);
nand U1679 (N_1679,N_1611,N_1635);
nand U1680 (N_1680,N_1641,N_1578);
and U1681 (N_1681,N_1579,N_1593);
nand U1682 (N_1682,N_1631,N_1620);
nand U1683 (N_1683,N_1582,N_1622);
or U1684 (N_1684,N_1633,N_1587);
and U1685 (N_1685,N_1583,N_1636);
and U1686 (N_1686,N_1630,N_1601);
and U1687 (N_1687,N_1599,N_1623);
nand U1688 (N_1688,N_1596,N_1578);
and U1689 (N_1689,N_1646,N_1600);
and U1690 (N_1690,N_1578,N_1592);
and U1691 (N_1691,N_1641,N_1598);
nand U1692 (N_1692,N_1633,N_1595);
nand U1693 (N_1693,N_1632,N_1588);
nor U1694 (N_1694,N_1610,N_1611);
nor U1695 (N_1695,N_1581,N_1588);
nor U1696 (N_1696,N_1627,N_1582);
or U1697 (N_1697,N_1618,N_1576);
or U1698 (N_1698,N_1631,N_1628);
and U1699 (N_1699,N_1634,N_1621);
nor U1700 (N_1700,N_1648,N_1633);
or U1701 (N_1701,N_1648,N_1646);
nor U1702 (N_1702,N_1646,N_1585);
nor U1703 (N_1703,N_1612,N_1584);
or U1704 (N_1704,N_1647,N_1598);
or U1705 (N_1705,N_1625,N_1648);
xnor U1706 (N_1706,N_1616,N_1587);
or U1707 (N_1707,N_1613,N_1643);
and U1708 (N_1708,N_1620,N_1640);
and U1709 (N_1709,N_1636,N_1595);
nor U1710 (N_1710,N_1637,N_1579);
or U1711 (N_1711,N_1603,N_1619);
or U1712 (N_1712,N_1605,N_1602);
and U1713 (N_1713,N_1593,N_1600);
nor U1714 (N_1714,N_1582,N_1617);
nor U1715 (N_1715,N_1635,N_1598);
or U1716 (N_1716,N_1649,N_1610);
nand U1717 (N_1717,N_1579,N_1610);
and U1718 (N_1718,N_1630,N_1643);
and U1719 (N_1719,N_1624,N_1583);
or U1720 (N_1720,N_1648,N_1631);
or U1721 (N_1721,N_1628,N_1643);
and U1722 (N_1722,N_1596,N_1589);
or U1723 (N_1723,N_1638,N_1587);
nor U1724 (N_1724,N_1606,N_1619);
nand U1725 (N_1725,N_1652,N_1708);
and U1726 (N_1726,N_1707,N_1724);
nor U1727 (N_1727,N_1692,N_1690);
and U1728 (N_1728,N_1660,N_1676);
nand U1729 (N_1729,N_1683,N_1681);
or U1730 (N_1730,N_1656,N_1658);
or U1731 (N_1731,N_1667,N_1661);
or U1732 (N_1732,N_1653,N_1675);
nor U1733 (N_1733,N_1696,N_1678);
nand U1734 (N_1734,N_1688,N_1682);
and U1735 (N_1735,N_1709,N_1717);
nand U1736 (N_1736,N_1670,N_1684);
or U1737 (N_1737,N_1662,N_1712);
nand U1738 (N_1738,N_1715,N_1685);
or U1739 (N_1739,N_1654,N_1666);
nand U1740 (N_1740,N_1689,N_1665);
nand U1741 (N_1741,N_1664,N_1713);
nor U1742 (N_1742,N_1651,N_1719);
or U1743 (N_1743,N_1716,N_1677);
nand U1744 (N_1744,N_1705,N_1702);
and U1745 (N_1745,N_1674,N_1691);
nand U1746 (N_1746,N_1704,N_1671);
nor U1747 (N_1747,N_1714,N_1698);
and U1748 (N_1748,N_1703,N_1720);
nand U1749 (N_1749,N_1655,N_1694);
nor U1750 (N_1750,N_1695,N_1659);
nand U1751 (N_1751,N_1650,N_1687);
nand U1752 (N_1752,N_1663,N_1706);
nor U1753 (N_1753,N_1679,N_1668);
nor U1754 (N_1754,N_1700,N_1697);
nor U1755 (N_1755,N_1657,N_1711);
or U1756 (N_1756,N_1672,N_1680);
nand U1757 (N_1757,N_1721,N_1710);
nand U1758 (N_1758,N_1718,N_1723);
nor U1759 (N_1759,N_1669,N_1686);
or U1760 (N_1760,N_1699,N_1693);
nand U1761 (N_1761,N_1673,N_1701);
nand U1762 (N_1762,N_1722,N_1694);
or U1763 (N_1763,N_1690,N_1664);
or U1764 (N_1764,N_1667,N_1665);
and U1765 (N_1765,N_1692,N_1695);
and U1766 (N_1766,N_1695,N_1690);
nand U1767 (N_1767,N_1660,N_1658);
or U1768 (N_1768,N_1722,N_1693);
or U1769 (N_1769,N_1684,N_1698);
nand U1770 (N_1770,N_1655,N_1687);
nand U1771 (N_1771,N_1654,N_1717);
nand U1772 (N_1772,N_1694,N_1673);
and U1773 (N_1773,N_1670,N_1722);
nand U1774 (N_1774,N_1702,N_1713);
or U1775 (N_1775,N_1678,N_1684);
and U1776 (N_1776,N_1654,N_1676);
nand U1777 (N_1777,N_1701,N_1699);
nand U1778 (N_1778,N_1682,N_1664);
nor U1779 (N_1779,N_1720,N_1681);
or U1780 (N_1780,N_1707,N_1678);
nor U1781 (N_1781,N_1675,N_1711);
and U1782 (N_1782,N_1724,N_1723);
and U1783 (N_1783,N_1672,N_1699);
or U1784 (N_1784,N_1709,N_1707);
nor U1785 (N_1785,N_1690,N_1659);
and U1786 (N_1786,N_1715,N_1714);
or U1787 (N_1787,N_1670,N_1702);
nor U1788 (N_1788,N_1660,N_1683);
nor U1789 (N_1789,N_1716,N_1724);
and U1790 (N_1790,N_1720,N_1650);
nand U1791 (N_1791,N_1694,N_1703);
nand U1792 (N_1792,N_1674,N_1710);
or U1793 (N_1793,N_1707,N_1697);
or U1794 (N_1794,N_1698,N_1656);
or U1795 (N_1795,N_1723,N_1694);
and U1796 (N_1796,N_1674,N_1706);
or U1797 (N_1797,N_1674,N_1715);
nor U1798 (N_1798,N_1657,N_1698);
nand U1799 (N_1799,N_1676,N_1715);
nand U1800 (N_1800,N_1746,N_1753);
or U1801 (N_1801,N_1738,N_1768);
and U1802 (N_1802,N_1789,N_1757);
and U1803 (N_1803,N_1796,N_1773);
nand U1804 (N_1804,N_1776,N_1747);
and U1805 (N_1805,N_1728,N_1760);
and U1806 (N_1806,N_1729,N_1793);
nor U1807 (N_1807,N_1756,N_1769);
or U1808 (N_1808,N_1727,N_1790);
or U1809 (N_1809,N_1788,N_1754);
or U1810 (N_1810,N_1791,N_1745);
nor U1811 (N_1811,N_1743,N_1742);
or U1812 (N_1812,N_1736,N_1731);
xor U1813 (N_1813,N_1784,N_1767);
nor U1814 (N_1814,N_1759,N_1752);
and U1815 (N_1815,N_1772,N_1787);
and U1816 (N_1816,N_1732,N_1779);
and U1817 (N_1817,N_1771,N_1778);
and U1818 (N_1818,N_1761,N_1799);
nor U1819 (N_1819,N_1763,N_1781);
or U1820 (N_1820,N_1726,N_1730);
or U1821 (N_1821,N_1764,N_1739);
and U1822 (N_1822,N_1785,N_1751);
nor U1823 (N_1823,N_1758,N_1786);
and U1824 (N_1824,N_1733,N_1794);
nand U1825 (N_1825,N_1735,N_1797);
nor U1826 (N_1826,N_1770,N_1782);
nand U1827 (N_1827,N_1795,N_1734);
and U1828 (N_1828,N_1777,N_1798);
or U1829 (N_1829,N_1741,N_1755);
or U1830 (N_1830,N_1780,N_1765);
or U1831 (N_1831,N_1774,N_1749);
and U1832 (N_1832,N_1792,N_1766);
nor U1833 (N_1833,N_1740,N_1762);
and U1834 (N_1834,N_1775,N_1748);
xnor U1835 (N_1835,N_1744,N_1737);
nand U1836 (N_1836,N_1725,N_1750);
nand U1837 (N_1837,N_1783,N_1735);
nor U1838 (N_1838,N_1788,N_1760);
nand U1839 (N_1839,N_1750,N_1742);
nor U1840 (N_1840,N_1777,N_1783);
nand U1841 (N_1841,N_1740,N_1757);
nand U1842 (N_1842,N_1750,N_1797);
or U1843 (N_1843,N_1729,N_1751);
nor U1844 (N_1844,N_1784,N_1725);
and U1845 (N_1845,N_1727,N_1757);
and U1846 (N_1846,N_1788,N_1732);
or U1847 (N_1847,N_1740,N_1734);
or U1848 (N_1848,N_1737,N_1768);
nand U1849 (N_1849,N_1762,N_1727);
nor U1850 (N_1850,N_1750,N_1741);
nand U1851 (N_1851,N_1741,N_1768);
or U1852 (N_1852,N_1767,N_1736);
or U1853 (N_1853,N_1748,N_1746);
and U1854 (N_1854,N_1757,N_1765);
nand U1855 (N_1855,N_1774,N_1726);
or U1856 (N_1856,N_1751,N_1788);
nand U1857 (N_1857,N_1762,N_1751);
nand U1858 (N_1858,N_1725,N_1738);
and U1859 (N_1859,N_1781,N_1754);
or U1860 (N_1860,N_1751,N_1770);
or U1861 (N_1861,N_1757,N_1728);
and U1862 (N_1862,N_1779,N_1770);
and U1863 (N_1863,N_1756,N_1736);
nor U1864 (N_1864,N_1789,N_1797);
nand U1865 (N_1865,N_1768,N_1788);
nand U1866 (N_1866,N_1792,N_1733);
nand U1867 (N_1867,N_1784,N_1774);
or U1868 (N_1868,N_1734,N_1743);
or U1869 (N_1869,N_1744,N_1770);
nor U1870 (N_1870,N_1790,N_1749);
nand U1871 (N_1871,N_1763,N_1786);
nand U1872 (N_1872,N_1755,N_1743);
and U1873 (N_1873,N_1765,N_1737);
or U1874 (N_1874,N_1773,N_1737);
nand U1875 (N_1875,N_1865,N_1802);
nand U1876 (N_1876,N_1821,N_1800);
nand U1877 (N_1877,N_1809,N_1843);
and U1878 (N_1878,N_1801,N_1845);
and U1879 (N_1879,N_1805,N_1833);
nand U1880 (N_1880,N_1839,N_1818);
and U1881 (N_1881,N_1873,N_1869);
nand U1882 (N_1882,N_1852,N_1834);
and U1883 (N_1883,N_1830,N_1861);
or U1884 (N_1884,N_1829,N_1838);
or U1885 (N_1885,N_1840,N_1870);
nor U1886 (N_1886,N_1806,N_1808);
or U1887 (N_1887,N_1846,N_1860);
or U1888 (N_1888,N_1841,N_1804);
nor U1889 (N_1889,N_1863,N_1813);
or U1890 (N_1890,N_1824,N_1814);
nand U1891 (N_1891,N_1850,N_1867);
and U1892 (N_1892,N_1857,N_1848);
and U1893 (N_1893,N_1816,N_1836);
or U1894 (N_1894,N_1864,N_1825);
or U1895 (N_1895,N_1822,N_1837);
nor U1896 (N_1896,N_1866,N_1859);
nor U1897 (N_1897,N_1820,N_1811);
nor U1898 (N_1898,N_1842,N_1844);
nor U1899 (N_1899,N_1819,N_1823);
or U1900 (N_1900,N_1817,N_1831);
nor U1901 (N_1901,N_1812,N_1815);
nor U1902 (N_1902,N_1855,N_1858);
and U1903 (N_1903,N_1856,N_1827);
nor U1904 (N_1904,N_1851,N_1872);
and U1905 (N_1905,N_1853,N_1835);
or U1906 (N_1906,N_1871,N_1826);
nor U1907 (N_1907,N_1807,N_1810);
and U1908 (N_1908,N_1862,N_1849);
nand U1909 (N_1909,N_1832,N_1847);
nand U1910 (N_1910,N_1874,N_1868);
or U1911 (N_1911,N_1803,N_1854);
and U1912 (N_1912,N_1828,N_1856);
nand U1913 (N_1913,N_1840,N_1864);
or U1914 (N_1914,N_1858,N_1829);
and U1915 (N_1915,N_1830,N_1810);
nand U1916 (N_1916,N_1852,N_1816);
and U1917 (N_1917,N_1873,N_1827);
and U1918 (N_1918,N_1839,N_1855);
or U1919 (N_1919,N_1856,N_1817);
and U1920 (N_1920,N_1838,N_1874);
and U1921 (N_1921,N_1826,N_1872);
nand U1922 (N_1922,N_1833,N_1844);
nand U1923 (N_1923,N_1832,N_1833);
nor U1924 (N_1924,N_1803,N_1860);
nand U1925 (N_1925,N_1822,N_1812);
and U1926 (N_1926,N_1800,N_1872);
nor U1927 (N_1927,N_1870,N_1830);
and U1928 (N_1928,N_1866,N_1844);
nor U1929 (N_1929,N_1849,N_1842);
or U1930 (N_1930,N_1817,N_1864);
and U1931 (N_1931,N_1831,N_1838);
or U1932 (N_1932,N_1848,N_1854);
nor U1933 (N_1933,N_1840,N_1828);
nand U1934 (N_1934,N_1858,N_1818);
and U1935 (N_1935,N_1805,N_1862);
nor U1936 (N_1936,N_1835,N_1822);
nor U1937 (N_1937,N_1846,N_1825);
or U1938 (N_1938,N_1866,N_1836);
or U1939 (N_1939,N_1811,N_1852);
or U1940 (N_1940,N_1840,N_1856);
or U1941 (N_1941,N_1849,N_1815);
or U1942 (N_1942,N_1805,N_1804);
and U1943 (N_1943,N_1857,N_1827);
nor U1944 (N_1944,N_1842,N_1835);
or U1945 (N_1945,N_1823,N_1809);
or U1946 (N_1946,N_1802,N_1800);
nor U1947 (N_1947,N_1816,N_1872);
and U1948 (N_1948,N_1805,N_1822);
and U1949 (N_1949,N_1852,N_1843);
and U1950 (N_1950,N_1880,N_1904);
nand U1951 (N_1951,N_1877,N_1941);
nor U1952 (N_1952,N_1912,N_1919);
or U1953 (N_1953,N_1922,N_1910);
and U1954 (N_1954,N_1920,N_1939);
or U1955 (N_1955,N_1949,N_1916);
or U1956 (N_1956,N_1909,N_1948);
nand U1957 (N_1957,N_1928,N_1944);
nor U1958 (N_1958,N_1908,N_1926);
or U1959 (N_1959,N_1892,N_1901);
nor U1960 (N_1960,N_1913,N_1878);
nor U1961 (N_1961,N_1917,N_1911);
and U1962 (N_1962,N_1890,N_1887);
nor U1963 (N_1963,N_1930,N_1879);
and U1964 (N_1964,N_1885,N_1947);
nand U1965 (N_1965,N_1905,N_1897);
nand U1966 (N_1966,N_1927,N_1935);
and U1967 (N_1967,N_1883,N_1891);
or U1968 (N_1968,N_1893,N_1924);
nor U1969 (N_1969,N_1921,N_1915);
nand U1970 (N_1970,N_1906,N_1931);
or U1971 (N_1971,N_1943,N_1918);
or U1972 (N_1972,N_1940,N_1923);
nor U1973 (N_1973,N_1900,N_1899);
nand U1974 (N_1974,N_1942,N_1936);
and U1975 (N_1975,N_1902,N_1882);
and U1976 (N_1976,N_1929,N_1895);
nand U1977 (N_1977,N_1938,N_1881);
nand U1978 (N_1978,N_1896,N_1933);
and U1979 (N_1979,N_1945,N_1914);
or U1980 (N_1980,N_1889,N_1898);
nand U1981 (N_1981,N_1925,N_1894);
and U1982 (N_1982,N_1937,N_1946);
and U1983 (N_1983,N_1886,N_1934);
or U1984 (N_1984,N_1903,N_1932);
nand U1985 (N_1985,N_1888,N_1884);
nor U1986 (N_1986,N_1907,N_1876);
and U1987 (N_1987,N_1875,N_1909);
or U1988 (N_1988,N_1913,N_1939);
nor U1989 (N_1989,N_1928,N_1918);
nor U1990 (N_1990,N_1891,N_1930);
and U1991 (N_1991,N_1947,N_1886);
nand U1992 (N_1992,N_1914,N_1947);
or U1993 (N_1993,N_1884,N_1876);
and U1994 (N_1994,N_1907,N_1879);
nor U1995 (N_1995,N_1928,N_1896);
or U1996 (N_1996,N_1929,N_1881);
nand U1997 (N_1997,N_1940,N_1922);
nor U1998 (N_1998,N_1946,N_1908);
and U1999 (N_1999,N_1920,N_1900);
or U2000 (N_2000,N_1889,N_1947);
nand U2001 (N_2001,N_1937,N_1942);
nor U2002 (N_2002,N_1889,N_1933);
nand U2003 (N_2003,N_1887,N_1914);
nor U2004 (N_2004,N_1877,N_1911);
or U2005 (N_2005,N_1906,N_1911);
or U2006 (N_2006,N_1875,N_1945);
and U2007 (N_2007,N_1880,N_1884);
nor U2008 (N_2008,N_1904,N_1926);
and U2009 (N_2009,N_1944,N_1926);
or U2010 (N_2010,N_1927,N_1928);
and U2011 (N_2011,N_1884,N_1914);
and U2012 (N_2012,N_1878,N_1904);
and U2013 (N_2013,N_1879,N_1914);
and U2014 (N_2014,N_1934,N_1949);
and U2015 (N_2015,N_1902,N_1913);
or U2016 (N_2016,N_1904,N_1930);
nand U2017 (N_2017,N_1876,N_1926);
and U2018 (N_2018,N_1938,N_1883);
and U2019 (N_2019,N_1911,N_1921);
nor U2020 (N_2020,N_1890,N_1945);
and U2021 (N_2021,N_1887,N_1942);
nor U2022 (N_2022,N_1909,N_1927);
or U2023 (N_2023,N_1884,N_1886);
or U2024 (N_2024,N_1903,N_1906);
nand U2025 (N_2025,N_1997,N_2007);
or U2026 (N_2026,N_1954,N_2019);
and U2027 (N_2027,N_1953,N_1989);
nand U2028 (N_2028,N_1985,N_2006);
or U2029 (N_2029,N_2002,N_1964);
or U2030 (N_2030,N_1990,N_1980);
or U2031 (N_2031,N_1984,N_1959);
or U2032 (N_2032,N_2005,N_1976);
nor U2033 (N_2033,N_2020,N_2004);
nand U2034 (N_2034,N_1966,N_1951);
or U2035 (N_2035,N_2014,N_1999);
nand U2036 (N_2036,N_1987,N_1958);
nand U2037 (N_2037,N_1983,N_1982);
nand U2038 (N_2038,N_1957,N_1992);
and U2039 (N_2039,N_1963,N_1991);
or U2040 (N_2040,N_1974,N_1988);
or U2041 (N_2041,N_1977,N_1955);
nand U2042 (N_2042,N_2008,N_2010);
and U2043 (N_2043,N_1996,N_1970);
and U2044 (N_2044,N_1978,N_2001);
or U2045 (N_2045,N_1993,N_2011);
nand U2046 (N_2046,N_2021,N_2024);
and U2047 (N_2047,N_2016,N_1994);
nor U2048 (N_2048,N_2022,N_1971);
or U2049 (N_2049,N_2018,N_1950);
xnor U2050 (N_2050,N_1961,N_1956);
nor U2051 (N_2051,N_1981,N_2000);
or U2052 (N_2052,N_2017,N_1995);
nor U2053 (N_2053,N_1979,N_1973);
or U2054 (N_2054,N_2012,N_1952);
nor U2055 (N_2055,N_1972,N_1968);
nand U2056 (N_2056,N_2013,N_1986);
nand U2057 (N_2057,N_1962,N_1998);
nor U2058 (N_2058,N_2015,N_1965);
nor U2059 (N_2059,N_1960,N_2023);
or U2060 (N_2060,N_1967,N_2009);
and U2061 (N_2061,N_1975,N_2003);
nor U2062 (N_2062,N_1969,N_1952);
nor U2063 (N_2063,N_1983,N_1968);
and U2064 (N_2064,N_1950,N_1961);
nor U2065 (N_2065,N_2001,N_1969);
nor U2066 (N_2066,N_1981,N_1983);
nand U2067 (N_2067,N_2008,N_2014);
nand U2068 (N_2068,N_2022,N_1986);
and U2069 (N_2069,N_1981,N_1952);
nand U2070 (N_2070,N_2018,N_1955);
and U2071 (N_2071,N_1979,N_1974);
nand U2072 (N_2072,N_2018,N_2023);
or U2073 (N_2073,N_2024,N_1989);
and U2074 (N_2074,N_1978,N_1951);
nand U2075 (N_2075,N_1970,N_1960);
nor U2076 (N_2076,N_1954,N_2022);
nor U2077 (N_2077,N_1965,N_2021);
or U2078 (N_2078,N_1958,N_2021);
nand U2079 (N_2079,N_1995,N_1987);
and U2080 (N_2080,N_2009,N_2002);
nand U2081 (N_2081,N_2015,N_1998);
or U2082 (N_2082,N_1962,N_1977);
or U2083 (N_2083,N_2009,N_1984);
and U2084 (N_2084,N_2010,N_1998);
and U2085 (N_2085,N_2003,N_2008);
or U2086 (N_2086,N_2004,N_1991);
nor U2087 (N_2087,N_1958,N_2008);
and U2088 (N_2088,N_2010,N_2002);
and U2089 (N_2089,N_2020,N_1958);
nand U2090 (N_2090,N_2014,N_1972);
and U2091 (N_2091,N_1956,N_2005);
nand U2092 (N_2092,N_1997,N_1963);
or U2093 (N_2093,N_1957,N_1971);
nand U2094 (N_2094,N_2015,N_1977);
nand U2095 (N_2095,N_1962,N_2002);
nor U2096 (N_2096,N_1995,N_1975);
or U2097 (N_2097,N_2019,N_1999);
and U2098 (N_2098,N_1964,N_1972);
or U2099 (N_2099,N_1996,N_1999);
and U2100 (N_2100,N_2037,N_2026);
or U2101 (N_2101,N_2062,N_2075);
or U2102 (N_2102,N_2059,N_2091);
nand U2103 (N_2103,N_2029,N_2088);
nor U2104 (N_2104,N_2045,N_2086);
nand U2105 (N_2105,N_2057,N_2041);
or U2106 (N_2106,N_2087,N_2089);
xor U2107 (N_2107,N_2027,N_2058);
nand U2108 (N_2108,N_2097,N_2094);
nand U2109 (N_2109,N_2090,N_2053);
nand U2110 (N_2110,N_2032,N_2072);
nor U2111 (N_2111,N_2028,N_2083);
or U2112 (N_2112,N_2073,N_2080);
or U2113 (N_2113,N_2048,N_2033);
and U2114 (N_2114,N_2076,N_2098);
or U2115 (N_2115,N_2055,N_2042);
nor U2116 (N_2116,N_2056,N_2060);
nor U2117 (N_2117,N_2025,N_2038);
nand U2118 (N_2118,N_2082,N_2085);
nor U2119 (N_2119,N_2051,N_2054);
and U2120 (N_2120,N_2031,N_2095);
nand U2121 (N_2121,N_2092,N_2069);
or U2122 (N_2122,N_2052,N_2081);
nand U2123 (N_2123,N_2039,N_2079);
nor U2124 (N_2124,N_2063,N_2096);
nor U2125 (N_2125,N_2049,N_2030);
nand U2126 (N_2126,N_2067,N_2077);
nand U2127 (N_2127,N_2064,N_2047);
nand U2128 (N_2128,N_2078,N_2034);
nor U2129 (N_2129,N_2071,N_2074);
and U2130 (N_2130,N_2068,N_2084);
and U2131 (N_2131,N_2043,N_2044);
or U2132 (N_2132,N_2061,N_2036);
nand U2133 (N_2133,N_2070,N_2065);
or U2134 (N_2134,N_2066,N_2093);
nand U2135 (N_2135,N_2050,N_2099);
nand U2136 (N_2136,N_2046,N_2035);
and U2137 (N_2137,N_2040,N_2047);
nand U2138 (N_2138,N_2063,N_2082);
or U2139 (N_2139,N_2052,N_2080);
nor U2140 (N_2140,N_2030,N_2091);
nor U2141 (N_2141,N_2043,N_2028);
nor U2142 (N_2142,N_2048,N_2070);
xnor U2143 (N_2143,N_2072,N_2084);
nand U2144 (N_2144,N_2067,N_2042);
or U2145 (N_2145,N_2055,N_2056);
nor U2146 (N_2146,N_2075,N_2079);
nor U2147 (N_2147,N_2073,N_2096);
nor U2148 (N_2148,N_2095,N_2037);
and U2149 (N_2149,N_2063,N_2066);
or U2150 (N_2150,N_2086,N_2064);
or U2151 (N_2151,N_2052,N_2067);
or U2152 (N_2152,N_2070,N_2039);
nor U2153 (N_2153,N_2095,N_2035);
or U2154 (N_2154,N_2052,N_2049);
and U2155 (N_2155,N_2027,N_2040);
nand U2156 (N_2156,N_2097,N_2027);
nor U2157 (N_2157,N_2085,N_2095);
nor U2158 (N_2158,N_2080,N_2043);
nor U2159 (N_2159,N_2096,N_2048);
or U2160 (N_2160,N_2071,N_2038);
or U2161 (N_2161,N_2041,N_2081);
or U2162 (N_2162,N_2081,N_2062);
nor U2163 (N_2163,N_2064,N_2091);
nand U2164 (N_2164,N_2079,N_2068);
and U2165 (N_2165,N_2041,N_2099);
nand U2166 (N_2166,N_2042,N_2091);
and U2167 (N_2167,N_2052,N_2084);
and U2168 (N_2168,N_2054,N_2041);
nand U2169 (N_2169,N_2056,N_2072);
or U2170 (N_2170,N_2075,N_2026);
nand U2171 (N_2171,N_2079,N_2086);
and U2172 (N_2172,N_2063,N_2043);
xor U2173 (N_2173,N_2056,N_2063);
or U2174 (N_2174,N_2035,N_2059);
or U2175 (N_2175,N_2104,N_2106);
nand U2176 (N_2176,N_2124,N_2159);
nand U2177 (N_2177,N_2135,N_2130);
and U2178 (N_2178,N_2162,N_2133);
nor U2179 (N_2179,N_2129,N_2119);
and U2180 (N_2180,N_2168,N_2157);
nand U2181 (N_2181,N_2116,N_2152);
nand U2182 (N_2182,N_2167,N_2102);
and U2183 (N_2183,N_2120,N_2156);
and U2184 (N_2184,N_2142,N_2145);
or U2185 (N_2185,N_2118,N_2143);
xnor U2186 (N_2186,N_2149,N_2160);
or U2187 (N_2187,N_2103,N_2163);
nand U2188 (N_2188,N_2153,N_2125);
nor U2189 (N_2189,N_2154,N_2140);
nand U2190 (N_2190,N_2141,N_2132);
nand U2191 (N_2191,N_2139,N_2161);
and U2192 (N_2192,N_2150,N_2128);
or U2193 (N_2193,N_2138,N_2115);
and U2194 (N_2194,N_2110,N_2137);
and U2195 (N_2195,N_2169,N_2174);
or U2196 (N_2196,N_2172,N_2123);
nor U2197 (N_2197,N_2136,N_2134);
or U2198 (N_2198,N_2148,N_2101);
or U2199 (N_2199,N_2131,N_2146);
nand U2200 (N_2200,N_2155,N_2121);
nor U2201 (N_2201,N_2111,N_2109);
and U2202 (N_2202,N_2112,N_2108);
nand U2203 (N_2203,N_2170,N_2151);
nor U2204 (N_2204,N_2107,N_2173);
or U2205 (N_2205,N_2100,N_2144);
nand U2206 (N_2206,N_2117,N_2171);
or U2207 (N_2207,N_2113,N_2166);
nor U2208 (N_2208,N_2164,N_2147);
or U2209 (N_2209,N_2105,N_2165);
and U2210 (N_2210,N_2158,N_2126);
or U2211 (N_2211,N_2127,N_2122);
and U2212 (N_2212,N_2114,N_2144);
nand U2213 (N_2213,N_2108,N_2149);
and U2214 (N_2214,N_2169,N_2116);
nor U2215 (N_2215,N_2131,N_2116);
and U2216 (N_2216,N_2156,N_2127);
nand U2217 (N_2217,N_2166,N_2145);
or U2218 (N_2218,N_2149,N_2147);
nand U2219 (N_2219,N_2132,N_2152);
nor U2220 (N_2220,N_2148,N_2127);
or U2221 (N_2221,N_2103,N_2116);
nand U2222 (N_2222,N_2142,N_2130);
nand U2223 (N_2223,N_2111,N_2122);
and U2224 (N_2224,N_2139,N_2142);
nand U2225 (N_2225,N_2107,N_2163);
and U2226 (N_2226,N_2147,N_2106);
nor U2227 (N_2227,N_2111,N_2145);
nor U2228 (N_2228,N_2133,N_2110);
and U2229 (N_2229,N_2132,N_2148);
nor U2230 (N_2230,N_2117,N_2133);
and U2231 (N_2231,N_2157,N_2121);
and U2232 (N_2232,N_2131,N_2115);
nand U2233 (N_2233,N_2129,N_2157);
nor U2234 (N_2234,N_2161,N_2106);
and U2235 (N_2235,N_2142,N_2123);
nor U2236 (N_2236,N_2113,N_2116);
and U2237 (N_2237,N_2172,N_2147);
and U2238 (N_2238,N_2141,N_2128);
and U2239 (N_2239,N_2160,N_2108);
or U2240 (N_2240,N_2105,N_2152);
nor U2241 (N_2241,N_2113,N_2174);
and U2242 (N_2242,N_2110,N_2124);
or U2243 (N_2243,N_2147,N_2168);
or U2244 (N_2244,N_2148,N_2161);
nor U2245 (N_2245,N_2111,N_2102);
and U2246 (N_2246,N_2171,N_2144);
nand U2247 (N_2247,N_2166,N_2144);
nor U2248 (N_2248,N_2125,N_2143);
or U2249 (N_2249,N_2131,N_2147);
nor U2250 (N_2250,N_2244,N_2178);
and U2251 (N_2251,N_2229,N_2193);
and U2252 (N_2252,N_2208,N_2216);
and U2253 (N_2253,N_2202,N_2191);
or U2254 (N_2254,N_2214,N_2239);
or U2255 (N_2255,N_2235,N_2213);
or U2256 (N_2256,N_2197,N_2240);
nand U2257 (N_2257,N_2184,N_2226);
nand U2258 (N_2258,N_2194,N_2225);
nor U2259 (N_2259,N_2176,N_2181);
and U2260 (N_2260,N_2245,N_2238);
and U2261 (N_2261,N_2177,N_2217);
nand U2262 (N_2262,N_2222,N_2249);
or U2263 (N_2263,N_2175,N_2203);
nor U2264 (N_2264,N_2221,N_2182);
nand U2265 (N_2265,N_2207,N_2185);
and U2266 (N_2266,N_2243,N_2209);
or U2267 (N_2267,N_2180,N_2198);
and U2268 (N_2268,N_2210,N_2241);
nor U2269 (N_2269,N_2228,N_2204);
or U2270 (N_2270,N_2246,N_2233);
nand U2271 (N_2271,N_2192,N_2218);
and U2272 (N_2272,N_2232,N_2236);
nand U2273 (N_2273,N_2179,N_2201);
nand U2274 (N_2274,N_2183,N_2200);
nand U2275 (N_2275,N_2190,N_2219);
and U2276 (N_2276,N_2220,N_2187);
nand U2277 (N_2277,N_2247,N_2231);
nand U2278 (N_2278,N_2248,N_2234);
or U2279 (N_2279,N_2206,N_2195);
or U2280 (N_2280,N_2227,N_2205);
or U2281 (N_2281,N_2199,N_2215);
and U2282 (N_2282,N_2188,N_2212);
nor U2283 (N_2283,N_2237,N_2230);
and U2284 (N_2284,N_2186,N_2189);
nor U2285 (N_2285,N_2196,N_2242);
nand U2286 (N_2286,N_2211,N_2223);
and U2287 (N_2287,N_2224,N_2229);
nand U2288 (N_2288,N_2229,N_2206);
nor U2289 (N_2289,N_2237,N_2227);
and U2290 (N_2290,N_2206,N_2245);
and U2291 (N_2291,N_2204,N_2209);
and U2292 (N_2292,N_2212,N_2225);
nand U2293 (N_2293,N_2240,N_2244);
or U2294 (N_2294,N_2204,N_2239);
and U2295 (N_2295,N_2208,N_2177);
nor U2296 (N_2296,N_2227,N_2200);
or U2297 (N_2297,N_2229,N_2191);
or U2298 (N_2298,N_2193,N_2231);
nand U2299 (N_2299,N_2211,N_2236);
nand U2300 (N_2300,N_2226,N_2221);
and U2301 (N_2301,N_2187,N_2239);
or U2302 (N_2302,N_2225,N_2247);
or U2303 (N_2303,N_2192,N_2205);
nand U2304 (N_2304,N_2208,N_2191);
and U2305 (N_2305,N_2207,N_2194);
nand U2306 (N_2306,N_2249,N_2184);
nand U2307 (N_2307,N_2188,N_2196);
nand U2308 (N_2308,N_2246,N_2248);
nand U2309 (N_2309,N_2198,N_2209);
and U2310 (N_2310,N_2179,N_2235);
nor U2311 (N_2311,N_2199,N_2238);
and U2312 (N_2312,N_2198,N_2181);
nand U2313 (N_2313,N_2178,N_2242);
nand U2314 (N_2314,N_2189,N_2242);
and U2315 (N_2315,N_2227,N_2234);
nand U2316 (N_2316,N_2191,N_2201);
or U2317 (N_2317,N_2191,N_2188);
or U2318 (N_2318,N_2186,N_2192);
and U2319 (N_2319,N_2209,N_2233);
and U2320 (N_2320,N_2248,N_2233);
or U2321 (N_2321,N_2218,N_2177);
nor U2322 (N_2322,N_2175,N_2191);
or U2323 (N_2323,N_2204,N_2221);
nor U2324 (N_2324,N_2224,N_2233);
or U2325 (N_2325,N_2310,N_2306);
and U2326 (N_2326,N_2318,N_2270);
and U2327 (N_2327,N_2273,N_2312);
nor U2328 (N_2328,N_2250,N_2311);
nand U2329 (N_2329,N_2259,N_2301);
and U2330 (N_2330,N_2295,N_2266);
nand U2331 (N_2331,N_2279,N_2265);
nor U2332 (N_2332,N_2252,N_2253);
and U2333 (N_2333,N_2257,N_2280);
nor U2334 (N_2334,N_2293,N_2272);
or U2335 (N_2335,N_2274,N_2267);
or U2336 (N_2336,N_2302,N_2286);
nand U2337 (N_2337,N_2261,N_2317);
and U2338 (N_2338,N_2316,N_2323);
nor U2339 (N_2339,N_2297,N_2320);
nand U2340 (N_2340,N_2289,N_2305);
and U2341 (N_2341,N_2308,N_2304);
and U2342 (N_2342,N_2258,N_2268);
or U2343 (N_2343,N_2291,N_2294);
or U2344 (N_2344,N_2255,N_2300);
and U2345 (N_2345,N_2275,N_2307);
nand U2346 (N_2346,N_2324,N_2263);
nand U2347 (N_2347,N_2276,N_2260);
and U2348 (N_2348,N_2292,N_2321);
and U2349 (N_2349,N_2251,N_2288);
nand U2350 (N_2350,N_2313,N_2283);
and U2351 (N_2351,N_2278,N_2277);
and U2352 (N_2352,N_2314,N_2299);
or U2353 (N_2353,N_2285,N_2269);
nor U2354 (N_2354,N_2264,N_2287);
or U2355 (N_2355,N_2254,N_2309);
nor U2356 (N_2356,N_2303,N_2290);
and U2357 (N_2357,N_2271,N_2319);
nor U2358 (N_2358,N_2284,N_2322);
nor U2359 (N_2359,N_2281,N_2315);
nand U2360 (N_2360,N_2296,N_2298);
nor U2361 (N_2361,N_2256,N_2262);
or U2362 (N_2362,N_2282,N_2306);
or U2363 (N_2363,N_2260,N_2265);
or U2364 (N_2364,N_2314,N_2277);
or U2365 (N_2365,N_2260,N_2309);
nand U2366 (N_2366,N_2251,N_2320);
and U2367 (N_2367,N_2276,N_2313);
nor U2368 (N_2368,N_2314,N_2267);
nor U2369 (N_2369,N_2274,N_2311);
nand U2370 (N_2370,N_2307,N_2285);
nand U2371 (N_2371,N_2323,N_2268);
and U2372 (N_2372,N_2306,N_2321);
nand U2373 (N_2373,N_2283,N_2264);
nor U2374 (N_2374,N_2309,N_2252);
and U2375 (N_2375,N_2301,N_2277);
nor U2376 (N_2376,N_2273,N_2290);
nor U2377 (N_2377,N_2265,N_2286);
nor U2378 (N_2378,N_2275,N_2290);
nor U2379 (N_2379,N_2277,N_2320);
nor U2380 (N_2380,N_2308,N_2292);
or U2381 (N_2381,N_2265,N_2323);
or U2382 (N_2382,N_2293,N_2303);
or U2383 (N_2383,N_2257,N_2289);
nor U2384 (N_2384,N_2309,N_2256);
nor U2385 (N_2385,N_2302,N_2304);
and U2386 (N_2386,N_2265,N_2278);
or U2387 (N_2387,N_2267,N_2306);
nor U2388 (N_2388,N_2297,N_2264);
and U2389 (N_2389,N_2265,N_2256);
nor U2390 (N_2390,N_2288,N_2312);
nor U2391 (N_2391,N_2281,N_2268);
and U2392 (N_2392,N_2322,N_2321);
nor U2393 (N_2393,N_2263,N_2270);
or U2394 (N_2394,N_2284,N_2307);
nor U2395 (N_2395,N_2289,N_2282);
and U2396 (N_2396,N_2317,N_2283);
and U2397 (N_2397,N_2318,N_2273);
or U2398 (N_2398,N_2308,N_2310);
nand U2399 (N_2399,N_2268,N_2285);
nor U2400 (N_2400,N_2352,N_2354);
nand U2401 (N_2401,N_2394,N_2380);
or U2402 (N_2402,N_2339,N_2355);
or U2403 (N_2403,N_2376,N_2345);
and U2404 (N_2404,N_2337,N_2382);
xor U2405 (N_2405,N_2386,N_2356);
nand U2406 (N_2406,N_2327,N_2353);
nor U2407 (N_2407,N_2363,N_2391);
and U2408 (N_2408,N_2332,N_2385);
and U2409 (N_2409,N_2390,N_2342);
or U2410 (N_2410,N_2370,N_2328);
nor U2411 (N_2411,N_2344,N_2350);
nor U2412 (N_2412,N_2366,N_2362);
nand U2413 (N_2413,N_2387,N_2351);
or U2414 (N_2414,N_2378,N_2333);
or U2415 (N_2415,N_2389,N_2349);
and U2416 (N_2416,N_2365,N_2381);
or U2417 (N_2417,N_2325,N_2375);
and U2418 (N_2418,N_2379,N_2334);
nand U2419 (N_2419,N_2346,N_2326);
and U2420 (N_2420,N_2360,N_2329);
or U2421 (N_2421,N_2373,N_2377);
nor U2422 (N_2422,N_2397,N_2384);
nand U2423 (N_2423,N_2398,N_2399);
nor U2424 (N_2424,N_2371,N_2372);
nand U2425 (N_2425,N_2383,N_2388);
nand U2426 (N_2426,N_2361,N_2343);
nor U2427 (N_2427,N_2368,N_2357);
or U2428 (N_2428,N_2340,N_2336);
or U2429 (N_2429,N_2330,N_2374);
or U2430 (N_2430,N_2331,N_2341);
nand U2431 (N_2431,N_2367,N_2358);
or U2432 (N_2432,N_2369,N_2395);
or U2433 (N_2433,N_2338,N_2335);
or U2434 (N_2434,N_2359,N_2392);
and U2435 (N_2435,N_2393,N_2364);
nand U2436 (N_2436,N_2347,N_2348);
or U2437 (N_2437,N_2396,N_2377);
nor U2438 (N_2438,N_2393,N_2395);
and U2439 (N_2439,N_2345,N_2327);
nor U2440 (N_2440,N_2354,N_2388);
or U2441 (N_2441,N_2361,N_2329);
and U2442 (N_2442,N_2349,N_2362);
nand U2443 (N_2443,N_2379,N_2351);
nor U2444 (N_2444,N_2398,N_2357);
nor U2445 (N_2445,N_2329,N_2398);
and U2446 (N_2446,N_2396,N_2340);
nand U2447 (N_2447,N_2325,N_2338);
nor U2448 (N_2448,N_2377,N_2370);
nand U2449 (N_2449,N_2335,N_2358);
nor U2450 (N_2450,N_2372,N_2327);
and U2451 (N_2451,N_2339,N_2356);
nand U2452 (N_2452,N_2398,N_2384);
nand U2453 (N_2453,N_2368,N_2327);
nor U2454 (N_2454,N_2342,N_2373);
nor U2455 (N_2455,N_2395,N_2348);
and U2456 (N_2456,N_2362,N_2345);
nor U2457 (N_2457,N_2343,N_2368);
and U2458 (N_2458,N_2363,N_2332);
nor U2459 (N_2459,N_2330,N_2353);
and U2460 (N_2460,N_2331,N_2375);
nor U2461 (N_2461,N_2387,N_2366);
or U2462 (N_2462,N_2332,N_2352);
xnor U2463 (N_2463,N_2337,N_2376);
or U2464 (N_2464,N_2366,N_2352);
and U2465 (N_2465,N_2328,N_2390);
nand U2466 (N_2466,N_2343,N_2385);
or U2467 (N_2467,N_2343,N_2333);
nand U2468 (N_2468,N_2365,N_2330);
nand U2469 (N_2469,N_2397,N_2345);
nor U2470 (N_2470,N_2327,N_2357);
nand U2471 (N_2471,N_2356,N_2388);
nor U2472 (N_2472,N_2382,N_2397);
nor U2473 (N_2473,N_2352,N_2389);
and U2474 (N_2474,N_2339,N_2396);
and U2475 (N_2475,N_2405,N_2425);
and U2476 (N_2476,N_2471,N_2455);
and U2477 (N_2477,N_2402,N_2418);
and U2478 (N_2478,N_2434,N_2459);
and U2479 (N_2479,N_2457,N_2442);
and U2480 (N_2480,N_2414,N_2468);
and U2481 (N_2481,N_2444,N_2421);
nand U2482 (N_2482,N_2469,N_2420);
and U2483 (N_2483,N_2473,N_2464);
or U2484 (N_2484,N_2431,N_2461);
or U2485 (N_2485,N_2441,N_2423);
and U2486 (N_2486,N_2426,N_2403);
or U2487 (N_2487,N_2447,N_2417);
nor U2488 (N_2488,N_2429,N_2410);
and U2489 (N_2489,N_2424,N_2430);
nor U2490 (N_2490,N_2443,N_2406);
and U2491 (N_2491,N_2466,N_2416);
and U2492 (N_2492,N_2458,N_2438);
nor U2493 (N_2493,N_2448,N_2415);
nor U2494 (N_2494,N_2440,N_2454);
or U2495 (N_2495,N_2428,N_2407);
and U2496 (N_2496,N_2470,N_2449);
nand U2497 (N_2497,N_2456,N_2419);
or U2498 (N_2498,N_2401,N_2422);
or U2499 (N_2499,N_2453,N_2404);
or U2500 (N_2500,N_2463,N_2433);
nand U2501 (N_2501,N_2451,N_2432);
nand U2502 (N_2502,N_2439,N_2474);
nand U2503 (N_2503,N_2408,N_2427);
and U2504 (N_2504,N_2465,N_2446);
and U2505 (N_2505,N_2450,N_2462);
or U2506 (N_2506,N_2460,N_2435);
or U2507 (N_2507,N_2452,N_2412);
nand U2508 (N_2508,N_2436,N_2400);
nor U2509 (N_2509,N_2467,N_2411);
nand U2510 (N_2510,N_2409,N_2472);
nor U2511 (N_2511,N_2445,N_2437);
nand U2512 (N_2512,N_2413,N_2412);
or U2513 (N_2513,N_2435,N_2457);
and U2514 (N_2514,N_2434,N_2433);
and U2515 (N_2515,N_2409,N_2412);
nor U2516 (N_2516,N_2413,N_2428);
or U2517 (N_2517,N_2461,N_2416);
and U2518 (N_2518,N_2469,N_2467);
nand U2519 (N_2519,N_2420,N_2452);
and U2520 (N_2520,N_2454,N_2418);
and U2521 (N_2521,N_2451,N_2457);
and U2522 (N_2522,N_2459,N_2420);
and U2523 (N_2523,N_2429,N_2427);
or U2524 (N_2524,N_2426,N_2441);
nand U2525 (N_2525,N_2409,N_2425);
and U2526 (N_2526,N_2464,N_2462);
nand U2527 (N_2527,N_2422,N_2468);
nor U2528 (N_2528,N_2433,N_2461);
or U2529 (N_2529,N_2416,N_2448);
and U2530 (N_2530,N_2453,N_2444);
nand U2531 (N_2531,N_2465,N_2400);
or U2532 (N_2532,N_2462,N_2427);
nand U2533 (N_2533,N_2415,N_2437);
nand U2534 (N_2534,N_2428,N_2442);
and U2535 (N_2535,N_2409,N_2438);
nor U2536 (N_2536,N_2402,N_2410);
nand U2537 (N_2537,N_2456,N_2404);
nand U2538 (N_2538,N_2446,N_2400);
nand U2539 (N_2539,N_2431,N_2457);
nand U2540 (N_2540,N_2420,N_2424);
or U2541 (N_2541,N_2429,N_2433);
nor U2542 (N_2542,N_2425,N_2419);
or U2543 (N_2543,N_2418,N_2421);
nand U2544 (N_2544,N_2473,N_2425);
nand U2545 (N_2545,N_2423,N_2474);
nand U2546 (N_2546,N_2429,N_2452);
or U2547 (N_2547,N_2403,N_2431);
and U2548 (N_2548,N_2407,N_2433);
and U2549 (N_2549,N_2443,N_2439);
or U2550 (N_2550,N_2517,N_2513);
nor U2551 (N_2551,N_2509,N_2533);
and U2552 (N_2552,N_2477,N_2529);
nand U2553 (N_2553,N_2495,N_2482);
nand U2554 (N_2554,N_2489,N_2480);
nand U2555 (N_2555,N_2491,N_2481);
and U2556 (N_2556,N_2531,N_2542);
nand U2557 (N_2557,N_2537,N_2492);
or U2558 (N_2558,N_2514,N_2544);
and U2559 (N_2559,N_2538,N_2527);
nand U2560 (N_2560,N_2530,N_2545);
or U2561 (N_2561,N_2476,N_2512);
and U2562 (N_2562,N_2534,N_2522);
nor U2563 (N_2563,N_2496,N_2502);
or U2564 (N_2564,N_2540,N_2547);
nor U2565 (N_2565,N_2515,N_2494);
and U2566 (N_2566,N_2528,N_2526);
nor U2567 (N_2567,N_2520,N_2504);
and U2568 (N_2568,N_2493,N_2498);
or U2569 (N_2569,N_2536,N_2523);
nand U2570 (N_2570,N_2524,N_2506);
or U2571 (N_2571,N_2484,N_2511);
and U2572 (N_2572,N_2521,N_2549);
nor U2573 (N_2573,N_2532,N_2510);
nor U2574 (N_2574,N_2485,N_2501);
nor U2575 (N_2575,N_2518,N_2535);
or U2576 (N_2576,N_2486,N_2519);
or U2577 (N_2577,N_2539,N_2546);
nor U2578 (N_2578,N_2503,N_2483);
and U2579 (N_2579,N_2499,N_2543);
and U2580 (N_2580,N_2497,N_2487);
nand U2581 (N_2581,N_2548,N_2541);
nand U2582 (N_2582,N_2525,N_2505);
and U2583 (N_2583,N_2488,N_2475);
nor U2584 (N_2584,N_2479,N_2490);
nor U2585 (N_2585,N_2508,N_2507);
nor U2586 (N_2586,N_2478,N_2500);
nor U2587 (N_2587,N_2516,N_2508);
and U2588 (N_2588,N_2479,N_2501);
or U2589 (N_2589,N_2535,N_2538);
nand U2590 (N_2590,N_2526,N_2503);
or U2591 (N_2591,N_2504,N_2526);
nor U2592 (N_2592,N_2532,N_2503);
nor U2593 (N_2593,N_2536,N_2529);
or U2594 (N_2594,N_2536,N_2501);
nor U2595 (N_2595,N_2540,N_2520);
nand U2596 (N_2596,N_2479,N_2487);
xor U2597 (N_2597,N_2500,N_2526);
nand U2598 (N_2598,N_2534,N_2492);
and U2599 (N_2599,N_2533,N_2482);
nor U2600 (N_2600,N_2475,N_2546);
nand U2601 (N_2601,N_2487,N_2517);
and U2602 (N_2602,N_2526,N_2538);
and U2603 (N_2603,N_2527,N_2513);
and U2604 (N_2604,N_2516,N_2504);
or U2605 (N_2605,N_2498,N_2522);
and U2606 (N_2606,N_2546,N_2516);
nand U2607 (N_2607,N_2489,N_2525);
and U2608 (N_2608,N_2547,N_2507);
and U2609 (N_2609,N_2508,N_2522);
nand U2610 (N_2610,N_2536,N_2482);
or U2611 (N_2611,N_2541,N_2516);
nand U2612 (N_2612,N_2491,N_2546);
nor U2613 (N_2613,N_2490,N_2544);
nor U2614 (N_2614,N_2534,N_2507);
nor U2615 (N_2615,N_2504,N_2536);
and U2616 (N_2616,N_2526,N_2546);
or U2617 (N_2617,N_2524,N_2500);
and U2618 (N_2618,N_2548,N_2524);
and U2619 (N_2619,N_2549,N_2520);
nand U2620 (N_2620,N_2512,N_2546);
nand U2621 (N_2621,N_2520,N_2525);
nand U2622 (N_2622,N_2477,N_2487);
or U2623 (N_2623,N_2503,N_2523);
and U2624 (N_2624,N_2487,N_2534);
and U2625 (N_2625,N_2553,N_2584);
or U2626 (N_2626,N_2572,N_2573);
nor U2627 (N_2627,N_2558,N_2599);
or U2628 (N_2628,N_2586,N_2600);
and U2629 (N_2629,N_2554,N_2582);
xor U2630 (N_2630,N_2555,N_2618);
nor U2631 (N_2631,N_2561,N_2552);
nand U2632 (N_2632,N_2617,N_2611);
nor U2633 (N_2633,N_2585,N_2612);
nand U2634 (N_2634,N_2551,N_2566);
and U2635 (N_2635,N_2622,N_2620);
or U2636 (N_2636,N_2563,N_2594);
and U2637 (N_2637,N_2619,N_2579);
and U2638 (N_2638,N_2574,N_2568);
nor U2639 (N_2639,N_2597,N_2575);
nor U2640 (N_2640,N_2570,N_2608);
nand U2641 (N_2641,N_2610,N_2605);
and U2642 (N_2642,N_2609,N_2577);
or U2643 (N_2643,N_2621,N_2567);
and U2644 (N_2644,N_2588,N_2593);
or U2645 (N_2645,N_2606,N_2557);
nor U2646 (N_2646,N_2595,N_2613);
nand U2647 (N_2647,N_2564,N_2560);
nor U2648 (N_2648,N_2576,N_2614);
or U2649 (N_2649,N_2590,N_2592);
and U2650 (N_2650,N_2602,N_2624);
xor U2651 (N_2651,N_2556,N_2607);
or U2652 (N_2652,N_2616,N_2565);
nand U2653 (N_2653,N_2583,N_2559);
and U2654 (N_2654,N_2604,N_2589);
and U2655 (N_2655,N_2580,N_2601);
nand U2656 (N_2656,N_2550,N_2571);
nand U2657 (N_2657,N_2569,N_2581);
or U2658 (N_2658,N_2562,N_2578);
or U2659 (N_2659,N_2587,N_2596);
and U2660 (N_2660,N_2591,N_2615);
nand U2661 (N_2661,N_2623,N_2598);
and U2662 (N_2662,N_2603,N_2619);
and U2663 (N_2663,N_2559,N_2558);
and U2664 (N_2664,N_2612,N_2572);
and U2665 (N_2665,N_2595,N_2569);
nand U2666 (N_2666,N_2601,N_2619);
or U2667 (N_2667,N_2619,N_2611);
nor U2668 (N_2668,N_2603,N_2611);
or U2669 (N_2669,N_2564,N_2611);
nor U2670 (N_2670,N_2605,N_2556);
xor U2671 (N_2671,N_2600,N_2580);
nand U2672 (N_2672,N_2593,N_2579);
nand U2673 (N_2673,N_2617,N_2574);
and U2674 (N_2674,N_2616,N_2570);
nand U2675 (N_2675,N_2579,N_2617);
or U2676 (N_2676,N_2611,N_2581);
or U2677 (N_2677,N_2573,N_2604);
nand U2678 (N_2678,N_2594,N_2611);
nor U2679 (N_2679,N_2593,N_2560);
or U2680 (N_2680,N_2559,N_2553);
or U2681 (N_2681,N_2569,N_2566);
and U2682 (N_2682,N_2567,N_2565);
nor U2683 (N_2683,N_2587,N_2609);
or U2684 (N_2684,N_2550,N_2599);
or U2685 (N_2685,N_2577,N_2553);
nand U2686 (N_2686,N_2571,N_2619);
or U2687 (N_2687,N_2609,N_2608);
or U2688 (N_2688,N_2624,N_2596);
nor U2689 (N_2689,N_2551,N_2559);
nand U2690 (N_2690,N_2597,N_2603);
and U2691 (N_2691,N_2594,N_2550);
nor U2692 (N_2692,N_2601,N_2550);
or U2693 (N_2693,N_2616,N_2600);
or U2694 (N_2694,N_2615,N_2568);
and U2695 (N_2695,N_2585,N_2582);
xor U2696 (N_2696,N_2604,N_2555);
nand U2697 (N_2697,N_2607,N_2564);
or U2698 (N_2698,N_2617,N_2577);
nand U2699 (N_2699,N_2605,N_2555);
nor U2700 (N_2700,N_2651,N_2682);
nor U2701 (N_2701,N_2653,N_2692);
nor U2702 (N_2702,N_2659,N_2673);
and U2703 (N_2703,N_2697,N_2683);
nand U2704 (N_2704,N_2665,N_2685);
nor U2705 (N_2705,N_2628,N_2663);
nor U2706 (N_2706,N_2649,N_2639);
nor U2707 (N_2707,N_2662,N_2677);
and U2708 (N_2708,N_2696,N_2629);
and U2709 (N_2709,N_2654,N_2636);
or U2710 (N_2710,N_2640,N_2657);
nand U2711 (N_2711,N_2660,N_2686);
and U2712 (N_2712,N_2668,N_2658);
and U2713 (N_2713,N_2694,N_2647);
and U2714 (N_2714,N_2635,N_2644);
or U2715 (N_2715,N_2632,N_2643);
nor U2716 (N_2716,N_2650,N_2691);
nor U2717 (N_2717,N_2638,N_2648);
and U2718 (N_2718,N_2689,N_2678);
and U2719 (N_2719,N_2627,N_2633);
and U2720 (N_2720,N_2675,N_2652);
and U2721 (N_2721,N_2642,N_2674);
or U2722 (N_2722,N_2661,N_2680);
and U2723 (N_2723,N_2679,N_2630);
and U2724 (N_2724,N_2669,N_2634);
nor U2725 (N_2725,N_2664,N_2688);
nand U2726 (N_2726,N_2666,N_2681);
and U2727 (N_2727,N_2699,N_2670);
or U2728 (N_2728,N_2626,N_2631);
nand U2729 (N_2729,N_2646,N_2693);
nand U2730 (N_2730,N_2687,N_2645);
nand U2731 (N_2731,N_2695,N_2667);
and U2732 (N_2732,N_2698,N_2672);
nand U2733 (N_2733,N_2690,N_2656);
nor U2734 (N_2734,N_2641,N_2676);
nor U2735 (N_2735,N_2655,N_2684);
nand U2736 (N_2736,N_2625,N_2671);
nand U2737 (N_2737,N_2637,N_2699);
nand U2738 (N_2738,N_2641,N_2669);
and U2739 (N_2739,N_2648,N_2641);
or U2740 (N_2740,N_2675,N_2647);
and U2741 (N_2741,N_2666,N_2659);
nor U2742 (N_2742,N_2690,N_2645);
nor U2743 (N_2743,N_2666,N_2658);
and U2744 (N_2744,N_2661,N_2650);
nor U2745 (N_2745,N_2648,N_2649);
nand U2746 (N_2746,N_2647,N_2670);
xnor U2747 (N_2747,N_2661,N_2676);
and U2748 (N_2748,N_2674,N_2640);
and U2749 (N_2749,N_2659,N_2688);
and U2750 (N_2750,N_2686,N_2682);
nand U2751 (N_2751,N_2670,N_2691);
xor U2752 (N_2752,N_2686,N_2633);
nor U2753 (N_2753,N_2688,N_2666);
nor U2754 (N_2754,N_2671,N_2668);
and U2755 (N_2755,N_2676,N_2651);
nand U2756 (N_2756,N_2661,N_2665);
or U2757 (N_2757,N_2658,N_2655);
nand U2758 (N_2758,N_2681,N_2657);
and U2759 (N_2759,N_2658,N_2663);
or U2760 (N_2760,N_2682,N_2634);
and U2761 (N_2761,N_2672,N_2696);
or U2762 (N_2762,N_2670,N_2644);
nor U2763 (N_2763,N_2643,N_2634);
nand U2764 (N_2764,N_2661,N_2664);
or U2765 (N_2765,N_2648,N_2693);
nor U2766 (N_2766,N_2666,N_2649);
or U2767 (N_2767,N_2686,N_2638);
or U2768 (N_2768,N_2672,N_2665);
nor U2769 (N_2769,N_2663,N_2685);
or U2770 (N_2770,N_2675,N_2664);
nor U2771 (N_2771,N_2678,N_2662);
or U2772 (N_2772,N_2691,N_2644);
and U2773 (N_2773,N_2646,N_2690);
nand U2774 (N_2774,N_2663,N_2642);
nor U2775 (N_2775,N_2713,N_2735);
or U2776 (N_2776,N_2736,N_2704);
or U2777 (N_2777,N_2742,N_2769);
and U2778 (N_2778,N_2745,N_2755);
nand U2779 (N_2779,N_2748,N_2743);
xnor U2780 (N_2780,N_2707,N_2711);
or U2781 (N_2781,N_2740,N_2701);
or U2782 (N_2782,N_2708,N_2723);
nor U2783 (N_2783,N_2709,N_2761);
nor U2784 (N_2784,N_2726,N_2724);
and U2785 (N_2785,N_2729,N_2758);
or U2786 (N_2786,N_2749,N_2751);
or U2787 (N_2787,N_2753,N_2770);
or U2788 (N_2788,N_2714,N_2722);
nor U2789 (N_2789,N_2765,N_2746);
nand U2790 (N_2790,N_2717,N_2763);
and U2791 (N_2791,N_2773,N_2762);
nor U2792 (N_2792,N_2731,N_2771);
nand U2793 (N_2793,N_2710,N_2721);
nor U2794 (N_2794,N_2718,N_2767);
or U2795 (N_2795,N_2702,N_2741);
nand U2796 (N_2796,N_2720,N_2730);
nand U2797 (N_2797,N_2757,N_2738);
nand U2798 (N_2798,N_2715,N_2732);
nor U2799 (N_2799,N_2706,N_2760);
and U2800 (N_2800,N_2739,N_2737);
nor U2801 (N_2801,N_2766,N_2768);
nand U2802 (N_2802,N_2764,N_2744);
nor U2803 (N_2803,N_2703,N_2754);
or U2804 (N_2804,N_2725,N_2734);
or U2805 (N_2805,N_2719,N_2759);
nand U2806 (N_2806,N_2747,N_2756);
or U2807 (N_2807,N_2716,N_2774);
and U2808 (N_2808,N_2728,N_2772);
nor U2809 (N_2809,N_2727,N_2705);
and U2810 (N_2810,N_2700,N_2750);
or U2811 (N_2811,N_2712,N_2752);
or U2812 (N_2812,N_2733,N_2719);
or U2813 (N_2813,N_2713,N_2736);
nand U2814 (N_2814,N_2723,N_2718);
or U2815 (N_2815,N_2758,N_2726);
nand U2816 (N_2816,N_2704,N_2767);
and U2817 (N_2817,N_2756,N_2750);
and U2818 (N_2818,N_2764,N_2747);
and U2819 (N_2819,N_2744,N_2763);
and U2820 (N_2820,N_2736,N_2742);
and U2821 (N_2821,N_2723,N_2722);
nor U2822 (N_2822,N_2763,N_2748);
nor U2823 (N_2823,N_2759,N_2734);
or U2824 (N_2824,N_2730,N_2731);
nor U2825 (N_2825,N_2723,N_2750);
xor U2826 (N_2826,N_2731,N_2700);
and U2827 (N_2827,N_2723,N_2761);
and U2828 (N_2828,N_2756,N_2759);
and U2829 (N_2829,N_2706,N_2719);
nor U2830 (N_2830,N_2727,N_2702);
and U2831 (N_2831,N_2727,N_2746);
nand U2832 (N_2832,N_2764,N_2720);
nand U2833 (N_2833,N_2712,N_2762);
nand U2834 (N_2834,N_2722,N_2730);
nand U2835 (N_2835,N_2726,N_2774);
and U2836 (N_2836,N_2701,N_2774);
or U2837 (N_2837,N_2703,N_2751);
nand U2838 (N_2838,N_2701,N_2773);
nor U2839 (N_2839,N_2706,N_2764);
nor U2840 (N_2840,N_2716,N_2746);
nand U2841 (N_2841,N_2764,N_2773);
or U2842 (N_2842,N_2719,N_2707);
nand U2843 (N_2843,N_2739,N_2709);
and U2844 (N_2844,N_2713,N_2747);
or U2845 (N_2845,N_2759,N_2739);
nand U2846 (N_2846,N_2706,N_2772);
and U2847 (N_2847,N_2719,N_2746);
and U2848 (N_2848,N_2753,N_2762);
nor U2849 (N_2849,N_2757,N_2726);
and U2850 (N_2850,N_2844,N_2793);
nand U2851 (N_2851,N_2847,N_2837);
nor U2852 (N_2852,N_2807,N_2829);
nand U2853 (N_2853,N_2806,N_2832);
and U2854 (N_2854,N_2800,N_2827);
or U2855 (N_2855,N_2839,N_2787);
and U2856 (N_2856,N_2836,N_2782);
and U2857 (N_2857,N_2786,N_2828);
nor U2858 (N_2858,N_2838,N_2830);
and U2859 (N_2859,N_2815,N_2789);
nand U2860 (N_2860,N_2824,N_2825);
and U2861 (N_2861,N_2791,N_2808);
nor U2862 (N_2862,N_2783,N_2831);
and U2863 (N_2863,N_2814,N_2790);
or U2864 (N_2864,N_2809,N_2820);
nand U2865 (N_2865,N_2792,N_2810);
or U2866 (N_2866,N_2797,N_2817);
nand U2867 (N_2867,N_2802,N_2812);
nor U2868 (N_2868,N_2846,N_2799);
or U2869 (N_2869,N_2780,N_2834);
nor U2870 (N_2870,N_2796,N_2778);
and U2871 (N_2871,N_2826,N_2805);
and U2872 (N_2872,N_2801,N_2798);
nor U2873 (N_2873,N_2803,N_2819);
nand U2874 (N_2874,N_2848,N_2804);
or U2875 (N_2875,N_2822,N_2795);
and U2876 (N_2876,N_2788,N_2794);
or U2877 (N_2877,N_2775,N_2823);
nand U2878 (N_2878,N_2785,N_2842);
nor U2879 (N_2879,N_2818,N_2777);
or U2880 (N_2880,N_2821,N_2833);
and U2881 (N_2881,N_2845,N_2784);
and U2882 (N_2882,N_2840,N_2813);
or U2883 (N_2883,N_2816,N_2843);
and U2884 (N_2884,N_2835,N_2811);
or U2885 (N_2885,N_2841,N_2849);
nand U2886 (N_2886,N_2776,N_2781);
xor U2887 (N_2887,N_2779,N_2837);
and U2888 (N_2888,N_2821,N_2785);
and U2889 (N_2889,N_2823,N_2815);
or U2890 (N_2890,N_2800,N_2810);
nor U2891 (N_2891,N_2836,N_2822);
nor U2892 (N_2892,N_2837,N_2841);
and U2893 (N_2893,N_2812,N_2822);
and U2894 (N_2894,N_2832,N_2784);
nand U2895 (N_2895,N_2807,N_2801);
nor U2896 (N_2896,N_2794,N_2790);
and U2897 (N_2897,N_2807,N_2816);
and U2898 (N_2898,N_2832,N_2844);
or U2899 (N_2899,N_2843,N_2836);
nor U2900 (N_2900,N_2834,N_2802);
nand U2901 (N_2901,N_2808,N_2832);
or U2902 (N_2902,N_2821,N_2777);
and U2903 (N_2903,N_2785,N_2780);
nand U2904 (N_2904,N_2826,N_2819);
and U2905 (N_2905,N_2825,N_2841);
nor U2906 (N_2906,N_2837,N_2776);
nor U2907 (N_2907,N_2825,N_2842);
or U2908 (N_2908,N_2784,N_2781);
xor U2909 (N_2909,N_2775,N_2837);
and U2910 (N_2910,N_2843,N_2801);
nor U2911 (N_2911,N_2843,N_2830);
nand U2912 (N_2912,N_2846,N_2779);
nand U2913 (N_2913,N_2784,N_2791);
and U2914 (N_2914,N_2818,N_2847);
or U2915 (N_2915,N_2836,N_2807);
or U2916 (N_2916,N_2823,N_2832);
or U2917 (N_2917,N_2791,N_2829);
or U2918 (N_2918,N_2840,N_2848);
nand U2919 (N_2919,N_2785,N_2822);
or U2920 (N_2920,N_2789,N_2781);
nand U2921 (N_2921,N_2835,N_2819);
nand U2922 (N_2922,N_2788,N_2829);
or U2923 (N_2923,N_2822,N_2828);
or U2924 (N_2924,N_2834,N_2821);
nand U2925 (N_2925,N_2892,N_2851);
or U2926 (N_2926,N_2923,N_2867);
nor U2927 (N_2927,N_2913,N_2854);
and U2928 (N_2928,N_2895,N_2871);
nand U2929 (N_2929,N_2893,N_2904);
nand U2930 (N_2930,N_2869,N_2908);
nor U2931 (N_2931,N_2890,N_2879);
and U2932 (N_2932,N_2922,N_2857);
nor U2933 (N_2933,N_2919,N_2873);
nand U2934 (N_2934,N_2898,N_2917);
nand U2935 (N_2935,N_2911,N_2905);
nand U2936 (N_2936,N_2915,N_2852);
nor U2937 (N_2937,N_2921,N_2862);
and U2938 (N_2938,N_2860,N_2878);
nor U2939 (N_2939,N_2868,N_2876);
nor U2940 (N_2940,N_2907,N_2906);
nor U2941 (N_2941,N_2853,N_2896);
and U2942 (N_2942,N_2875,N_2891);
or U2943 (N_2943,N_2889,N_2912);
and U2944 (N_2944,N_2859,N_2901);
and U2945 (N_2945,N_2864,N_2863);
or U2946 (N_2946,N_2888,N_2902);
nand U2947 (N_2947,N_2856,N_2866);
nor U2948 (N_2948,N_2918,N_2855);
nand U2949 (N_2949,N_2870,N_2924);
nand U2950 (N_2950,N_2850,N_2897);
nand U2951 (N_2951,N_2880,N_2920);
nor U2952 (N_2952,N_2887,N_2872);
nand U2953 (N_2953,N_2883,N_2909);
or U2954 (N_2954,N_2858,N_2916);
or U2955 (N_2955,N_2861,N_2882);
or U2956 (N_2956,N_2885,N_2900);
or U2957 (N_2957,N_2877,N_2884);
nor U2958 (N_2958,N_2886,N_2894);
and U2959 (N_2959,N_2914,N_2865);
nand U2960 (N_2960,N_2899,N_2874);
and U2961 (N_2961,N_2903,N_2910);
or U2962 (N_2962,N_2881,N_2895);
nor U2963 (N_2963,N_2869,N_2872);
nand U2964 (N_2964,N_2874,N_2914);
and U2965 (N_2965,N_2919,N_2851);
or U2966 (N_2966,N_2906,N_2901);
nand U2967 (N_2967,N_2861,N_2893);
or U2968 (N_2968,N_2924,N_2916);
nand U2969 (N_2969,N_2913,N_2857);
and U2970 (N_2970,N_2896,N_2903);
or U2971 (N_2971,N_2897,N_2906);
nand U2972 (N_2972,N_2887,N_2877);
or U2973 (N_2973,N_2900,N_2890);
or U2974 (N_2974,N_2867,N_2896);
nand U2975 (N_2975,N_2904,N_2854);
and U2976 (N_2976,N_2918,N_2864);
or U2977 (N_2977,N_2911,N_2921);
and U2978 (N_2978,N_2914,N_2901);
nor U2979 (N_2979,N_2884,N_2924);
nand U2980 (N_2980,N_2871,N_2859);
or U2981 (N_2981,N_2898,N_2915);
nor U2982 (N_2982,N_2919,N_2857);
and U2983 (N_2983,N_2887,N_2899);
and U2984 (N_2984,N_2924,N_2868);
and U2985 (N_2985,N_2905,N_2879);
or U2986 (N_2986,N_2904,N_2899);
nor U2987 (N_2987,N_2909,N_2850);
nand U2988 (N_2988,N_2921,N_2859);
and U2989 (N_2989,N_2903,N_2905);
nor U2990 (N_2990,N_2893,N_2903);
nor U2991 (N_2991,N_2900,N_2908);
or U2992 (N_2992,N_2888,N_2894);
or U2993 (N_2993,N_2875,N_2884);
or U2994 (N_2994,N_2921,N_2902);
nor U2995 (N_2995,N_2891,N_2905);
nand U2996 (N_2996,N_2850,N_2871);
and U2997 (N_2997,N_2889,N_2915);
or U2998 (N_2998,N_2903,N_2873);
nand U2999 (N_2999,N_2860,N_2868);
nand UO_0 (O_0,N_2967,N_2927);
and UO_1 (O_1,N_2943,N_2962);
xor UO_2 (O_2,N_2998,N_2931);
nor UO_3 (O_3,N_2982,N_2949);
and UO_4 (O_4,N_2957,N_2939);
and UO_5 (O_5,N_2950,N_2969);
nor UO_6 (O_6,N_2988,N_2926);
or UO_7 (O_7,N_2940,N_2958);
and UO_8 (O_8,N_2997,N_2933);
nor UO_9 (O_9,N_2947,N_2941);
and UO_10 (O_10,N_2964,N_2970);
nand UO_11 (O_11,N_2928,N_2990);
nor UO_12 (O_12,N_2960,N_2983);
and UO_13 (O_13,N_2942,N_2948);
nand UO_14 (O_14,N_2959,N_2961);
nor UO_15 (O_15,N_2991,N_2979);
or UO_16 (O_16,N_2966,N_2937);
or UO_17 (O_17,N_2992,N_2994);
nand UO_18 (O_18,N_2934,N_2978);
nand UO_19 (O_19,N_2945,N_2930);
nand UO_20 (O_20,N_2996,N_2985);
or UO_21 (O_21,N_2956,N_2980);
and UO_22 (O_22,N_2993,N_2981);
and UO_23 (O_23,N_2999,N_2936);
nor UO_24 (O_24,N_2955,N_2986);
nor UO_25 (O_25,N_2965,N_2932);
xor UO_26 (O_26,N_2954,N_2976);
nor UO_27 (O_27,N_2952,N_2971);
or UO_28 (O_28,N_2984,N_2935);
and UO_29 (O_29,N_2972,N_2995);
nor UO_30 (O_30,N_2963,N_2944);
or UO_31 (O_31,N_2929,N_2951);
nor UO_32 (O_32,N_2974,N_2968);
nand UO_33 (O_33,N_2977,N_2946);
and UO_34 (O_34,N_2987,N_2989);
xnor UO_35 (O_35,N_2938,N_2953);
or UO_36 (O_36,N_2975,N_2925);
nor UO_37 (O_37,N_2973,N_2974);
nand UO_38 (O_38,N_2992,N_2974);
and UO_39 (O_39,N_2977,N_2972);
and UO_40 (O_40,N_2932,N_2947);
or UO_41 (O_41,N_2962,N_2985);
and UO_42 (O_42,N_2983,N_2925);
or UO_43 (O_43,N_2953,N_2950);
or UO_44 (O_44,N_2964,N_2980);
nand UO_45 (O_45,N_2960,N_2927);
nor UO_46 (O_46,N_2936,N_2940);
nand UO_47 (O_47,N_2931,N_2989);
nand UO_48 (O_48,N_2983,N_2964);
nand UO_49 (O_49,N_2930,N_2980);
or UO_50 (O_50,N_2990,N_2930);
nor UO_51 (O_51,N_2955,N_2961);
nor UO_52 (O_52,N_2978,N_2932);
and UO_53 (O_53,N_2999,N_2985);
nor UO_54 (O_54,N_2977,N_2969);
and UO_55 (O_55,N_2934,N_2935);
nand UO_56 (O_56,N_2987,N_2954);
nand UO_57 (O_57,N_2962,N_2998);
or UO_58 (O_58,N_2981,N_2942);
and UO_59 (O_59,N_2993,N_2957);
or UO_60 (O_60,N_2963,N_2925);
and UO_61 (O_61,N_2979,N_2965);
nand UO_62 (O_62,N_2986,N_2985);
and UO_63 (O_63,N_2929,N_2933);
and UO_64 (O_64,N_2960,N_2952);
xnor UO_65 (O_65,N_2927,N_2928);
nor UO_66 (O_66,N_2967,N_2995);
nor UO_67 (O_67,N_2978,N_2928);
or UO_68 (O_68,N_2952,N_2951);
nand UO_69 (O_69,N_2968,N_2984);
nand UO_70 (O_70,N_2930,N_2972);
nor UO_71 (O_71,N_2954,N_2969);
nand UO_72 (O_72,N_2962,N_2987);
or UO_73 (O_73,N_2934,N_2928);
and UO_74 (O_74,N_2954,N_2982);
nand UO_75 (O_75,N_2974,N_2964);
or UO_76 (O_76,N_2980,N_2948);
nand UO_77 (O_77,N_2992,N_2948);
or UO_78 (O_78,N_2983,N_2980);
nor UO_79 (O_79,N_2929,N_2961);
and UO_80 (O_80,N_2950,N_2957);
or UO_81 (O_81,N_2953,N_2933);
nand UO_82 (O_82,N_2963,N_2989);
nand UO_83 (O_83,N_2997,N_2927);
and UO_84 (O_84,N_2947,N_2959);
nand UO_85 (O_85,N_2983,N_2992);
and UO_86 (O_86,N_2925,N_2950);
and UO_87 (O_87,N_2954,N_2936);
nand UO_88 (O_88,N_2929,N_2943);
nor UO_89 (O_89,N_2972,N_2955);
nand UO_90 (O_90,N_2947,N_2962);
nor UO_91 (O_91,N_2989,N_2998);
nor UO_92 (O_92,N_2952,N_2942);
and UO_93 (O_93,N_2952,N_2987);
and UO_94 (O_94,N_2942,N_2990);
xor UO_95 (O_95,N_2998,N_2978);
or UO_96 (O_96,N_2972,N_2987);
or UO_97 (O_97,N_2938,N_2957);
nor UO_98 (O_98,N_2958,N_2962);
nor UO_99 (O_99,N_2935,N_2926);
or UO_100 (O_100,N_2996,N_2945);
nor UO_101 (O_101,N_2958,N_2981);
or UO_102 (O_102,N_2979,N_2970);
nor UO_103 (O_103,N_2940,N_2989);
and UO_104 (O_104,N_2958,N_2948);
or UO_105 (O_105,N_2999,N_2966);
nand UO_106 (O_106,N_2994,N_2981);
and UO_107 (O_107,N_2989,N_2969);
and UO_108 (O_108,N_2951,N_2982);
nor UO_109 (O_109,N_2936,N_2987);
nor UO_110 (O_110,N_2986,N_2954);
or UO_111 (O_111,N_2956,N_2997);
and UO_112 (O_112,N_2928,N_2998);
nand UO_113 (O_113,N_2972,N_2969);
and UO_114 (O_114,N_2939,N_2963);
nor UO_115 (O_115,N_2949,N_2955);
or UO_116 (O_116,N_2936,N_2968);
and UO_117 (O_117,N_2946,N_2951);
nor UO_118 (O_118,N_2961,N_2944);
and UO_119 (O_119,N_2986,N_2999);
nor UO_120 (O_120,N_2956,N_2983);
or UO_121 (O_121,N_2984,N_2957);
nor UO_122 (O_122,N_2973,N_2927);
and UO_123 (O_123,N_2993,N_2984);
and UO_124 (O_124,N_2979,N_2937);
and UO_125 (O_125,N_2999,N_2983);
nand UO_126 (O_126,N_2975,N_2938);
nand UO_127 (O_127,N_2981,N_2949);
nand UO_128 (O_128,N_2976,N_2993);
nor UO_129 (O_129,N_2941,N_2974);
nor UO_130 (O_130,N_2992,N_2950);
nand UO_131 (O_131,N_2965,N_2972);
or UO_132 (O_132,N_2972,N_2979);
nand UO_133 (O_133,N_2986,N_2971);
nor UO_134 (O_134,N_2939,N_2990);
nor UO_135 (O_135,N_2991,N_2967);
nand UO_136 (O_136,N_2982,N_2945);
nor UO_137 (O_137,N_2941,N_2946);
nor UO_138 (O_138,N_2983,N_2974);
or UO_139 (O_139,N_2939,N_2950);
or UO_140 (O_140,N_2995,N_2938);
nand UO_141 (O_141,N_2937,N_2995);
or UO_142 (O_142,N_2942,N_2966);
nand UO_143 (O_143,N_2986,N_2952);
nor UO_144 (O_144,N_2999,N_2928);
or UO_145 (O_145,N_2926,N_2978);
or UO_146 (O_146,N_2988,N_2983);
and UO_147 (O_147,N_2927,N_2950);
and UO_148 (O_148,N_2944,N_2972);
nor UO_149 (O_149,N_2968,N_2950);
and UO_150 (O_150,N_2945,N_2983);
nand UO_151 (O_151,N_2931,N_2994);
and UO_152 (O_152,N_2954,N_2997);
and UO_153 (O_153,N_2934,N_2964);
nand UO_154 (O_154,N_2949,N_2975);
or UO_155 (O_155,N_2975,N_2929);
or UO_156 (O_156,N_2975,N_2998);
or UO_157 (O_157,N_2925,N_2936);
nand UO_158 (O_158,N_2960,N_2982);
and UO_159 (O_159,N_2948,N_2972);
nor UO_160 (O_160,N_2939,N_2974);
nor UO_161 (O_161,N_2940,N_2955);
nand UO_162 (O_162,N_2938,N_2973);
nand UO_163 (O_163,N_2960,N_2997);
or UO_164 (O_164,N_2931,N_2978);
or UO_165 (O_165,N_2937,N_2956);
or UO_166 (O_166,N_2990,N_2967);
nor UO_167 (O_167,N_2980,N_2943);
and UO_168 (O_168,N_2932,N_2940);
nor UO_169 (O_169,N_2947,N_2980);
nor UO_170 (O_170,N_2938,N_2960);
and UO_171 (O_171,N_2934,N_2931);
nor UO_172 (O_172,N_2964,N_2989);
and UO_173 (O_173,N_2971,N_2966);
nand UO_174 (O_174,N_2940,N_2978);
nand UO_175 (O_175,N_2981,N_2953);
nand UO_176 (O_176,N_2970,N_2995);
and UO_177 (O_177,N_2929,N_2972);
nor UO_178 (O_178,N_2957,N_2986);
nand UO_179 (O_179,N_2935,N_2945);
nor UO_180 (O_180,N_2969,N_2955);
nor UO_181 (O_181,N_2925,N_2980);
or UO_182 (O_182,N_2997,N_2929);
nand UO_183 (O_183,N_2994,N_2939);
and UO_184 (O_184,N_2925,N_2984);
or UO_185 (O_185,N_2940,N_2928);
and UO_186 (O_186,N_2953,N_2985);
nand UO_187 (O_187,N_2995,N_2971);
and UO_188 (O_188,N_2983,N_2944);
nand UO_189 (O_189,N_2968,N_2942);
and UO_190 (O_190,N_2947,N_2998);
nor UO_191 (O_191,N_2992,N_2975);
nand UO_192 (O_192,N_2928,N_2933);
nor UO_193 (O_193,N_2942,N_2949);
or UO_194 (O_194,N_2988,N_2963);
and UO_195 (O_195,N_2983,N_2971);
nor UO_196 (O_196,N_2925,N_2927);
or UO_197 (O_197,N_2945,N_2940);
nand UO_198 (O_198,N_2978,N_2966);
nor UO_199 (O_199,N_2933,N_2999);
nand UO_200 (O_200,N_2967,N_2940);
and UO_201 (O_201,N_2963,N_2994);
and UO_202 (O_202,N_2929,N_2947);
or UO_203 (O_203,N_2939,N_2985);
nor UO_204 (O_204,N_2972,N_2953);
or UO_205 (O_205,N_2951,N_2940);
and UO_206 (O_206,N_2987,N_2943);
or UO_207 (O_207,N_2960,N_2934);
or UO_208 (O_208,N_2998,N_2996);
nor UO_209 (O_209,N_2956,N_2970);
nand UO_210 (O_210,N_2938,N_2985);
nor UO_211 (O_211,N_2939,N_2949);
or UO_212 (O_212,N_2992,N_2969);
or UO_213 (O_213,N_2991,N_2962);
and UO_214 (O_214,N_2954,N_2983);
and UO_215 (O_215,N_2995,N_2930);
and UO_216 (O_216,N_2938,N_2933);
xnor UO_217 (O_217,N_2942,N_2955);
nor UO_218 (O_218,N_2928,N_2944);
or UO_219 (O_219,N_2967,N_2956);
or UO_220 (O_220,N_2953,N_2957);
nor UO_221 (O_221,N_2951,N_2956);
nor UO_222 (O_222,N_2997,N_2998);
nand UO_223 (O_223,N_2959,N_2967);
or UO_224 (O_224,N_2958,N_2969);
xnor UO_225 (O_225,N_2965,N_2968);
and UO_226 (O_226,N_2965,N_2984);
and UO_227 (O_227,N_2965,N_2962);
or UO_228 (O_228,N_2975,N_2970);
or UO_229 (O_229,N_2943,N_2968);
or UO_230 (O_230,N_2970,N_2941);
nand UO_231 (O_231,N_2974,N_2950);
or UO_232 (O_232,N_2991,N_2959);
or UO_233 (O_233,N_2954,N_2966);
or UO_234 (O_234,N_2929,N_2970);
or UO_235 (O_235,N_2937,N_2991);
nor UO_236 (O_236,N_2957,N_2971);
or UO_237 (O_237,N_2958,N_2939);
or UO_238 (O_238,N_2996,N_2980);
or UO_239 (O_239,N_2934,N_2991);
nor UO_240 (O_240,N_2958,N_2997);
nand UO_241 (O_241,N_2941,N_2936);
or UO_242 (O_242,N_2976,N_2995);
or UO_243 (O_243,N_2951,N_2997);
nor UO_244 (O_244,N_2957,N_2977);
or UO_245 (O_245,N_2979,N_2964);
and UO_246 (O_246,N_2995,N_2975);
nand UO_247 (O_247,N_2935,N_2997);
nand UO_248 (O_248,N_2969,N_2979);
and UO_249 (O_249,N_2991,N_2963);
nand UO_250 (O_250,N_2972,N_2980);
nor UO_251 (O_251,N_2990,N_2991);
or UO_252 (O_252,N_2995,N_2962);
or UO_253 (O_253,N_2994,N_2986);
and UO_254 (O_254,N_2983,N_2989);
or UO_255 (O_255,N_2975,N_2982);
and UO_256 (O_256,N_2953,N_2937);
and UO_257 (O_257,N_2996,N_2942);
or UO_258 (O_258,N_2990,N_2946);
nor UO_259 (O_259,N_2928,N_2966);
nor UO_260 (O_260,N_2988,N_2962);
nor UO_261 (O_261,N_2939,N_2973);
xnor UO_262 (O_262,N_2970,N_2973);
or UO_263 (O_263,N_2992,N_2970);
nor UO_264 (O_264,N_2957,N_2970);
nor UO_265 (O_265,N_2990,N_2972);
nor UO_266 (O_266,N_2968,N_2946);
and UO_267 (O_267,N_2955,N_2957);
and UO_268 (O_268,N_2938,N_2948);
nor UO_269 (O_269,N_2957,N_2966);
nor UO_270 (O_270,N_2963,N_2964);
and UO_271 (O_271,N_2938,N_2929);
nor UO_272 (O_272,N_2972,N_2968);
nor UO_273 (O_273,N_2940,N_2966);
and UO_274 (O_274,N_2935,N_2942);
or UO_275 (O_275,N_2963,N_2984);
and UO_276 (O_276,N_2980,N_2979);
nor UO_277 (O_277,N_2944,N_2990);
and UO_278 (O_278,N_2942,N_2985);
nor UO_279 (O_279,N_2973,N_2956);
nand UO_280 (O_280,N_2998,N_2958);
and UO_281 (O_281,N_2998,N_2988);
or UO_282 (O_282,N_2937,N_2981);
nor UO_283 (O_283,N_2974,N_2991);
nand UO_284 (O_284,N_2967,N_2943);
nor UO_285 (O_285,N_2925,N_2992);
and UO_286 (O_286,N_2935,N_2978);
xnor UO_287 (O_287,N_2996,N_2973);
or UO_288 (O_288,N_2949,N_2974);
nor UO_289 (O_289,N_2968,N_2955);
nand UO_290 (O_290,N_2944,N_2959);
and UO_291 (O_291,N_2962,N_2997);
and UO_292 (O_292,N_2994,N_2996);
and UO_293 (O_293,N_2932,N_2966);
or UO_294 (O_294,N_2946,N_2943);
or UO_295 (O_295,N_2925,N_2952);
nor UO_296 (O_296,N_2960,N_2929);
or UO_297 (O_297,N_2946,N_2983);
and UO_298 (O_298,N_2942,N_2995);
xnor UO_299 (O_299,N_2935,N_2933);
or UO_300 (O_300,N_2988,N_2980);
nand UO_301 (O_301,N_2988,N_2937);
or UO_302 (O_302,N_2938,N_2972);
and UO_303 (O_303,N_2987,N_2942);
nand UO_304 (O_304,N_2933,N_2985);
nor UO_305 (O_305,N_2959,N_2977);
and UO_306 (O_306,N_2927,N_2972);
or UO_307 (O_307,N_2974,N_2932);
and UO_308 (O_308,N_2955,N_2933);
and UO_309 (O_309,N_2961,N_2986);
nor UO_310 (O_310,N_2980,N_2997);
and UO_311 (O_311,N_2947,N_2978);
nand UO_312 (O_312,N_2983,N_2993);
and UO_313 (O_313,N_2992,N_2929);
and UO_314 (O_314,N_2995,N_2961);
nand UO_315 (O_315,N_2973,N_2925);
and UO_316 (O_316,N_2978,N_2955);
nand UO_317 (O_317,N_2956,N_2996);
nand UO_318 (O_318,N_2934,N_2992);
nand UO_319 (O_319,N_2942,N_2977);
nor UO_320 (O_320,N_2963,N_2973);
or UO_321 (O_321,N_2989,N_2978);
xnor UO_322 (O_322,N_2965,N_2973);
and UO_323 (O_323,N_2946,N_2944);
nand UO_324 (O_324,N_2985,N_2993);
or UO_325 (O_325,N_2947,N_2997);
or UO_326 (O_326,N_2939,N_2984);
nand UO_327 (O_327,N_2952,N_2955);
or UO_328 (O_328,N_2982,N_2950);
nor UO_329 (O_329,N_2954,N_2933);
nor UO_330 (O_330,N_2993,N_2928);
or UO_331 (O_331,N_2956,N_2989);
and UO_332 (O_332,N_2928,N_2969);
nand UO_333 (O_333,N_2989,N_2959);
and UO_334 (O_334,N_2926,N_2957);
or UO_335 (O_335,N_2928,N_2963);
nand UO_336 (O_336,N_2949,N_2961);
nand UO_337 (O_337,N_2966,N_2953);
xor UO_338 (O_338,N_2929,N_2935);
nand UO_339 (O_339,N_2950,N_2946);
and UO_340 (O_340,N_2955,N_2965);
nand UO_341 (O_341,N_2949,N_2945);
and UO_342 (O_342,N_2935,N_2991);
or UO_343 (O_343,N_2938,N_2932);
and UO_344 (O_344,N_2979,N_2944);
nor UO_345 (O_345,N_2937,N_2942);
nand UO_346 (O_346,N_2985,N_2977);
nor UO_347 (O_347,N_2989,N_2966);
or UO_348 (O_348,N_2958,N_2952);
nand UO_349 (O_349,N_2945,N_2941);
nand UO_350 (O_350,N_2934,N_2997);
and UO_351 (O_351,N_2961,N_2940);
or UO_352 (O_352,N_2992,N_2952);
or UO_353 (O_353,N_2950,N_2931);
nor UO_354 (O_354,N_2932,N_2963);
nor UO_355 (O_355,N_2985,N_2925);
and UO_356 (O_356,N_2946,N_2959);
or UO_357 (O_357,N_2943,N_2960);
nor UO_358 (O_358,N_2970,N_2960);
nand UO_359 (O_359,N_2959,N_2994);
nor UO_360 (O_360,N_2990,N_2971);
and UO_361 (O_361,N_2950,N_2964);
nor UO_362 (O_362,N_2986,N_2926);
or UO_363 (O_363,N_2968,N_2932);
and UO_364 (O_364,N_2993,N_2975);
nor UO_365 (O_365,N_2989,N_2932);
and UO_366 (O_366,N_2975,N_2940);
and UO_367 (O_367,N_2926,N_2943);
nor UO_368 (O_368,N_2966,N_2979);
nor UO_369 (O_369,N_2973,N_2955);
or UO_370 (O_370,N_2956,N_2950);
and UO_371 (O_371,N_2976,N_2994);
nor UO_372 (O_372,N_2986,N_2938);
nand UO_373 (O_373,N_2971,N_2955);
or UO_374 (O_374,N_2944,N_2994);
nor UO_375 (O_375,N_2956,N_2976);
or UO_376 (O_376,N_2952,N_2949);
nand UO_377 (O_377,N_2928,N_2995);
and UO_378 (O_378,N_2943,N_2961);
or UO_379 (O_379,N_2984,N_2930);
or UO_380 (O_380,N_2959,N_2999);
nor UO_381 (O_381,N_2971,N_2982);
and UO_382 (O_382,N_2945,N_2984);
and UO_383 (O_383,N_2988,N_2930);
nor UO_384 (O_384,N_2989,N_2977);
nor UO_385 (O_385,N_2996,N_2931);
or UO_386 (O_386,N_2929,N_2949);
or UO_387 (O_387,N_2997,N_2932);
or UO_388 (O_388,N_2937,N_2987);
and UO_389 (O_389,N_2934,N_2958);
nand UO_390 (O_390,N_2968,N_2953);
or UO_391 (O_391,N_2994,N_2954);
and UO_392 (O_392,N_2975,N_2948);
nor UO_393 (O_393,N_2928,N_2945);
or UO_394 (O_394,N_2954,N_2967);
xnor UO_395 (O_395,N_2975,N_2991);
nand UO_396 (O_396,N_2969,N_2975);
xnor UO_397 (O_397,N_2944,N_2968);
or UO_398 (O_398,N_2948,N_2936);
nand UO_399 (O_399,N_2942,N_2941);
nor UO_400 (O_400,N_2925,N_2953);
or UO_401 (O_401,N_2986,N_2965);
or UO_402 (O_402,N_2975,N_2983);
and UO_403 (O_403,N_2925,N_2962);
and UO_404 (O_404,N_2966,N_2982);
nor UO_405 (O_405,N_2950,N_2985);
and UO_406 (O_406,N_2977,N_2961);
and UO_407 (O_407,N_2975,N_2954);
and UO_408 (O_408,N_2993,N_2986);
nand UO_409 (O_409,N_2961,N_2925);
and UO_410 (O_410,N_2951,N_2985);
nor UO_411 (O_411,N_2977,N_2932);
and UO_412 (O_412,N_2951,N_2960);
nor UO_413 (O_413,N_2982,N_2937);
or UO_414 (O_414,N_2936,N_2957);
and UO_415 (O_415,N_2928,N_2976);
nor UO_416 (O_416,N_2997,N_2989);
nand UO_417 (O_417,N_2935,N_2963);
or UO_418 (O_418,N_2941,N_2971);
nor UO_419 (O_419,N_2928,N_2991);
nor UO_420 (O_420,N_2990,N_2951);
nand UO_421 (O_421,N_2978,N_2927);
nand UO_422 (O_422,N_2965,N_2935);
nor UO_423 (O_423,N_2954,N_2927);
or UO_424 (O_424,N_2971,N_2968);
or UO_425 (O_425,N_2937,N_2957);
xnor UO_426 (O_426,N_2972,N_2981);
or UO_427 (O_427,N_2983,N_2949);
nor UO_428 (O_428,N_2983,N_2936);
nand UO_429 (O_429,N_2962,N_2946);
nand UO_430 (O_430,N_2951,N_2961);
nor UO_431 (O_431,N_2977,N_2971);
or UO_432 (O_432,N_2977,N_2966);
or UO_433 (O_433,N_2957,N_2974);
nand UO_434 (O_434,N_2943,N_2932);
nor UO_435 (O_435,N_2943,N_2963);
nor UO_436 (O_436,N_2945,N_2978);
or UO_437 (O_437,N_2984,N_2971);
and UO_438 (O_438,N_2925,N_2974);
nand UO_439 (O_439,N_2940,N_2985);
and UO_440 (O_440,N_2970,N_2959);
nand UO_441 (O_441,N_2959,N_2936);
nor UO_442 (O_442,N_2962,N_2975);
and UO_443 (O_443,N_2926,N_2925);
nor UO_444 (O_444,N_2945,N_2997);
nand UO_445 (O_445,N_2981,N_2948);
and UO_446 (O_446,N_2965,N_2976);
nand UO_447 (O_447,N_2941,N_2926);
nor UO_448 (O_448,N_2964,N_2975);
or UO_449 (O_449,N_2964,N_2967);
nand UO_450 (O_450,N_2976,N_2975);
or UO_451 (O_451,N_2960,N_2966);
and UO_452 (O_452,N_2944,N_2982);
or UO_453 (O_453,N_2992,N_2960);
or UO_454 (O_454,N_2933,N_2947);
or UO_455 (O_455,N_2967,N_2951);
nand UO_456 (O_456,N_2979,N_2929);
nand UO_457 (O_457,N_2956,N_2933);
and UO_458 (O_458,N_2938,N_2959);
nor UO_459 (O_459,N_2931,N_2937);
and UO_460 (O_460,N_2966,N_2985);
and UO_461 (O_461,N_2991,N_2996);
and UO_462 (O_462,N_2937,N_2986);
nor UO_463 (O_463,N_2935,N_2998);
nor UO_464 (O_464,N_2992,N_2926);
or UO_465 (O_465,N_2983,N_2985);
nor UO_466 (O_466,N_2984,N_2934);
and UO_467 (O_467,N_2988,N_2973);
and UO_468 (O_468,N_2950,N_2952);
and UO_469 (O_469,N_2945,N_2985);
and UO_470 (O_470,N_2932,N_2995);
and UO_471 (O_471,N_2988,N_2941);
and UO_472 (O_472,N_2980,N_2991);
and UO_473 (O_473,N_2952,N_2979);
nand UO_474 (O_474,N_2938,N_2946);
or UO_475 (O_475,N_2986,N_2953);
nor UO_476 (O_476,N_2962,N_2937);
and UO_477 (O_477,N_2936,N_2964);
nand UO_478 (O_478,N_2935,N_2938);
nand UO_479 (O_479,N_2930,N_2985);
or UO_480 (O_480,N_2939,N_2938);
and UO_481 (O_481,N_2964,N_2971);
nor UO_482 (O_482,N_2970,N_2947);
nor UO_483 (O_483,N_2971,N_2958);
nor UO_484 (O_484,N_2980,N_2927);
nand UO_485 (O_485,N_2965,N_2958);
and UO_486 (O_486,N_2929,N_2941);
nor UO_487 (O_487,N_2978,N_2951);
or UO_488 (O_488,N_2928,N_2984);
and UO_489 (O_489,N_2982,N_2936);
or UO_490 (O_490,N_2978,N_2982);
and UO_491 (O_491,N_2993,N_2974);
and UO_492 (O_492,N_2937,N_2955);
nor UO_493 (O_493,N_2979,N_2940);
or UO_494 (O_494,N_2959,N_2962);
or UO_495 (O_495,N_2947,N_2938);
nand UO_496 (O_496,N_2933,N_2931);
and UO_497 (O_497,N_2948,N_2932);
or UO_498 (O_498,N_2964,N_2982);
or UO_499 (O_499,N_2925,N_2965);
endmodule