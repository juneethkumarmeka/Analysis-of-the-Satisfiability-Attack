module basic_500_3000_500_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_37,In_107);
xor U1 (N_1,In_66,In_257);
nor U2 (N_2,In_485,In_175);
nand U3 (N_3,In_378,In_111);
nor U4 (N_4,In_92,In_80);
and U5 (N_5,In_360,In_142);
nor U6 (N_6,In_299,In_252);
and U7 (N_7,In_91,In_179);
nand U8 (N_8,In_258,In_14);
and U9 (N_9,In_165,In_251);
and U10 (N_10,In_269,In_127);
nand U11 (N_11,In_375,In_152);
nor U12 (N_12,In_6,In_319);
and U13 (N_13,In_355,In_496);
nand U14 (N_14,In_470,In_163);
and U15 (N_15,In_157,In_172);
and U16 (N_16,In_329,In_481);
xnor U17 (N_17,In_291,In_51);
nand U18 (N_18,In_483,In_106);
or U19 (N_19,In_90,In_144);
or U20 (N_20,In_387,In_495);
nand U21 (N_21,In_168,In_399);
nand U22 (N_22,In_373,In_323);
nor U23 (N_23,In_44,In_223);
nand U24 (N_24,In_148,In_290);
nand U25 (N_25,In_285,In_454);
and U26 (N_26,In_377,In_166);
nand U27 (N_27,In_292,In_449);
or U28 (N_28,In_262,In_53);
and U29 (N_29,In_42,In_105);
nand U30 (N_30,In_3,In_13);
nand U31 (N_31,In_126,In_88);
nand U32 (N_32,In_52,In_209);
or U33 (N_33,In_345,In_203);
and U34 (N_34,In_115,In_18);
nor U35 (N_35,In_185,In_327);
nor U36 (N_36,In_2,In_190);
or U37 (N_37,In_410,In_86);
nand U38 (N_38,In_308,In_491);
and U39 (N_39,In_171,In_353);
nand U40 (N_40,In_429,In_322);
nor U41 (N_41,In_247,In_189);
and U42 (N_42,In_181,In_186);
and U43 (N_43,In_73,In_121);
xor U44 (N_44,In_57,In_309);
nor U45 (N_45,In_374,In_476);
nand U46 (N_46,In_216,In_89);
or U47 (N_47,In_248,In_242);
and U48 (N_48,In_154,In_241);
xnor U49 (N_49,In_452,In_182);
or U50 (N_50,In_219,In_297);
or U51 (N_51,In_320,In_259);
or U52 (N_52,In_253,In_184);
and U53 (N_53,In_16,In_418);
and U54 (N_54,In_32,In_364);
and U55 (N_55,In_250,In_498);
nor U56 (N_56,In_408,In_124);
and U57 (N_57,In_25,In_348);
nand U58 (N_58,In_255,In_56);
or U59 (N_59,In_420,In_103);
xnor U60 (N_60,In_49,In_101);
or U61 (N_61,In_426,In_240);
and U62 (N_62,In_391,In_439);
nand U63 (N_63,In_451,In_150);
or U64 (N_64,In_278,In_445);
nand U65 (N_65,In_45,In_78);
nand U66 (N_66,In_300,In_233);
or U67 (N_67,In_74,In_493);
or U68 (N_68,In_95,In_135);
nor U69 (N_69,In_433,In_371);
and U70 (N_70,In_112,In_158);
and U71 (N_71,In_415,In_8);
xnor U72 (N_72,In_0,In_275);
nand U73 (N_73,In_384,In_314);
nor U74 (N_74,In_204,In_38);
or U75 (N_75,In_318,In_405);
nand U76 (N_76,In_134,In_153);
nor U77 (N_77,In_447,In_287);
and U78 (N_78,In_283,In_390);
nand U79 (N_79,In_43,In_335);
or U80 (N_80,In_354,In_392);
and U81 (N_81,In_407,In_465);
nor U82 (N_82,In_412,In_60);
xnor U83 (N_83,In_497,In_346);
nor U84 (N_84,In_211,In_347);
and U85 (N_85,In_351,In_382);
nor U86 (N_86,In_272,In_224);
nor U87 (N_87,In_487,In_201);
nor U88 (N_88,In_340,In_471);
or U89 (N_89,In_475,In_331);
nor U90 (N_90,In_232,In_243);
nor U91 (N_91,In_396,In_9);
nor U92 (N_92,In_381,In_443);
or U93 (N_93,In_468,In_486);
and U94 (N_94,In_302,In_450);
or U95 (N_95,In_194,In_427);
nand U96 (N_96,In_467,In_361);
nor U97 (N_97,In_169,In_424);
nand U98 (N_98,In_96,In_17);
and U99 (N_99,In_67,In_30);
or U100 (N_100,In_288,In_23);
or U101 (N_101,In_270,In_62);
nand U102 (N_102,In_342,In_197);
nand U103 (N_103,In_76,In_245);
nor U104 (N_104,In_440,In_130);
nand U105 (N_105,In_432,In_296);
and U106 (N_106,In_212,In_70);
nand U107 (N_107,In_389,In_28);
and U108 (N_108,In_466,In_341);
and U109 (N_109,In_231,In_114);
and U110 (N_110,In_33,In_457);
and U111 (N_111,In_456,In_100);
and U112 (N_112,In_178,In_227);
or U113 (N_113,In_305,In_406);
xor U114 (N_114,In_65,In_138);
nor U115 (N_115,In_210,In_455);
and U116 (N_116,In_409,In_221);
nor U117 (N_117,In_20,In_132);
nand U118 (N_118,In_237,In_330);
xor U119 (N_119,In_268,In_68);
xor U120 (N_120,In_98,In_417);
nand U121 (N_121,In_131,In_116);
or U122 (N_122,In_82,In_239);
or U123 (N_123,In_469,In_123);
and U124 (N_124,In_238,In_265);
xnor U125 (N_125,In_385,In_306);
and U126 (N_126,In_122,In_79);
nand U127 (N_127,In_128,In_192);
xor U128 (N_128,In_274,In_289);
and U129 (N_129,In_277,In_164);
or U130 (N_130,In_48,In_31);
or U131 (N_131,In_349,In_294);
xnor U132 (N_132,In_254,In_328);
and U133 (N_133,In_226,In_304);
and U134 (N_134,In_369,In_41);
and U135 (N_135,In_458,In_21);
nor U136 (N_136,In_206,In_11);
xor U137 (N_137,In_271,In_448);
or U138 (N_138,In_15,In_282);
and U139 (N_139,In_404,In_85);
or U140 (N_140,In_444,In_372);
and U141 (N_141,In_393,In_370);
nand U142 (N_142,In_359,In_50);
or U143 (N_143,In_125,In_273);
nand U144 (N_144,In_482,In_388);
xnor U145 (N_145,In_357,In_207);
nand U146 (N_146,In_477,In_149);
or U147 (N_147,In_325,In_441);
and U148 (N_148,In_380,In_379);
nor U149 (N_149,In_160,In_438);
xor U150 (N_150,In_386,In_198);
nand U151 (N_151,In_71,In_460);
nand U152 (N_152,In_94,In_326);
xor U153 (N_153,In_199,In_474);
nand U154 (N_154,In_208,In_337);
nand U155 (N_155,In_365,In_397);
nor U156 (N_156,In_4,In_222);
nand U157 (N_157,In_453,In_145);
nand U158 (N_158,In_193,In_110);
or U159 (N_159,In_244,In_431);
xor U160 (N_160,In_118,In_75);
nand U161 (N_161,In_58,In_298);
nand U162 (N_162,In_229,In_293);
and U163 (N_163,In_155,In_368);
or U164 (N_164,In_202,In_140);
xnor U165 (N_165,In_358,In_264);
or U166 (N_166,In_220,In_363);
and U167 (N_167,In_109,In_461);
nand U168 (N_168,In_214,In_217);
nand U169 (N_169,In_435,In_414);
nand U170 (N_170,In_27,In_416);
and U171 (N_171,In_108,In_77);
or U172 (N_172,In_421,In_307);
and U173 (N_173,In_187,In_81);
and U174 (N_174,In_36,In_263);
nor U175 (N_175,In_484,In_437);
nor U176 (N_176,In_200,In_464);
nor U177 (N_177,In_170,In_176);
nand U178 (N_178,In_225,In_183);
or U179 (N_179,In_488,In_246);
and U180 (N_180,In_195,In_10);
nand U181 (N_181,In_472,In_34);
and U182 (N_182,In_425,In_419);
and U183 (N_183,In_402,In_338);
nor U184 (N_184,In_312,In_156);
or U185 (N_185,In_230,In_494);
xnor U186 (N_186,In_411,In_301);
and U187 (N_187,In_234,In_343);
and U188 (N_188,In_54,In_40);
nand U189 (N_189,In_139,In_280);
or U190 (N_190,In_1,In_395);
nand U191 (N_191,In_12,In_260);
and U192 (N_192,In_339,In_310);
nand U193 (N_193,In_46,In_490);
nor U194 (N_194,In_26,In_167);
or U195 (N_195,In_434,In_22);
nand U196 (N_196,In_336,In_430);
or U197 (N_197,In_69,In_117);
nor U198 (N_198,In_311,In_266);
nand U199 (N_199,In_235,In_261);
nand U200 (N_200,In_303,In_356);
and U201 (N_201,In_147,In_84);
and U202 (N_202,In_236,In_191);
or U203 (N_203,In_281,In_442);
or U204 (N_204,In_120,In_492);
xnor U205 (N_205,In_141,In_332);
nand U206 (N_206,In_174,In_119);
or U207 (N_207,In_321,In_334);
or U208 (N_208,In_35,In_267);
xor U209 (N_209,In_83,In_480);
nor U210 (N_210,In_188,In_72);
and U211 (N_211,In_59,In_422);
and U212 (N_212,In_376,In_64);
and U213 (N_213,In_63,In_93);
nand U214 (N_214,In_459,In_398);
and U215 (N_215,In_413,In_143);
or U216 (N_216,In_104,In_344);
or U217 (N_217,In_394,In_102);
xnor U218 (N_218,In_436,In_446);
nand U219 (N_219,In_161,In_366);
xnor U220 (N_220,In_362,In_213);
nor U221 (N_221,In_249,In_177);
xor U222 (N_222,In_129,In_403);
nand U223 (N_223,In_173,In_317);
nand U224 (N_224,In_55,In_99);
and U225 (N_225,In_7,In_29);
and U226 (N_226,In_39,In_428);
and U227 (N_227,In_462,In_463);
and U228 (N_228,In_136,In_19);
nor U229 (N_229,In_499,In_61);
nand U230 (N_230,In_162,In_286);
or U231 (N_231,In_367,In_316);
nand U232 (N_232,In_313,In_324);
nor U233 (N_233,In_218,In_151);
nor U234 (N_234,In_205,In_489);
nand U235 (N_235,In_228,In_383);
nor U236 (N_236,In_113,In_276);
and U237 (N_237,In_479,In_47);
nand U238 (N_238,In_473,In_180);
and U239 (N_239,In_5,In_400);
nor U240 (N_240,In_401,In_196);
nand U241 (N_241,In_97,In_159);
and U242 (N_242,In_295,In_215);
xor U243 (N_243,In_87,In_315);
and U244 (N_244,In_423,In_146);
or U245 (N_245,In_284,In_279);
or U246 (N_246,In_133,In_478);
and U247 (N_247,In_24,In_137);
and U248 (N_248,In_256,In_350);
nor U249 (N_249,In_352,In_333);
or U250 (N_250,In_211,In_58);
or U251 (N_251,In_275,In_49);
and U252 (N_252,In_98,In_173);
or U253 (N_253,In_116,In_382);
nor U254 (N_254,In_122,In_260);
or U255 (N_255,In_169,In_324);
or U256 (N_256,In_169,In_189);
or U257 (N_257,In_162,In_220);
nand U258 (N_258,In_145,In_75);
and U259 (N_259,In_385,In_256);
or U260 (N_260,In_342,In_242);
nor U261 (N_261,In_43,In_413);
and U262 (N_262,In_142,In_334);
or U263 (N_263,In_253,In_32);
nor U264 (N_264,In_84,In_359);
and U265 (N_265,In_140,In_375);
nand U266 (N_266,In_192,In_313);
and U267 (N_267,In_490,In_259);
nand U268 (N_268,In_34,In_122);
or U269 (N_269,In_296,In_153);
nand U270 (N_270,In_430,In_363);
nor U271 (N_271,In_448,In_31);
nor U272 (N_272,In_421,In_423);
nor U273 (N_273,In_438,In_334);
and U274 (N_274,In_136,In_196);
nand U275 (N_275,In_337,In_273);
or U276 (N_276,In_261,In_6);
or U277 (N_277,In_69,In_374);
nand U278 (N_278,In_64,In_410);
or U279 (N_279,In_435,In_404);
xnor U280 (N_280,In_224,In_106);
nor U281 (N_281,In_183,In_281);
xor U282 (N_282,In_164,In_104);
and U283 (N_283,In_245,In_493);
or U284 (N_284,In_123,In_326);
or U285 (N_285,In_188,In_141);
and U286 (N_286,In_411,In_73);
nor U287 (N_287,In_16,In_13);
nand U288 (N_288,In_381,In_286);
and U289 (N_289,In_406,In_140);
nor U290 (N_290,In_371,In_427);
nand U291 (N_291,In_6,In_177);
and U292 (N_292,In_343,In_81);
and U293 (N_293,In_479,In_443);
nand U294 (N_294,In_4,In_336);
or U295 (N_295,In_145,In_203);
nand U296 (N_296,In_362,In_291);
and U297 (N_297,In_233,In_10);
nand U298 (N_298,In_228,In_46);
and U299 (N_299,In_367,In_177);
and U300 (N_300,In_82,In_480);
or U301 (N_301,In_49,In_245);
xnor U302 (N_302,In_476,In_58);
nand U303 (N_303,In_443,In_374);
and U304 (N_304,In_465,In_267);
nand U305 (N_305,In_241,In_447);
or U306 (N_306,In_344,In_117);
nand U307 (N_307,In_491,In_427);
nand U308 (N_308,In_37,In_462);
nand U309 (N_309,In_436,In_327);
nor U310 (N_310,In_90,In_29);
or U311 (N_311,In_258,In_295);
and U312 (N_312,In_402,In_237);
nor U313 (N_313,In_254,In_55);
and U314 (N_314,In_483,In_332);
and U315 (N_315,In_383,In_33);
nor U316 (N_316,In_95,In_216);
xnor U317 (N_317,In_297,In_364);
xor U318 (N_318,In_252,In_157);
and U319 (N_319,In_165,In_436);
nand U320 (N_320,In_241,In_301);
or U321 (N_321,In_255,In_429);
nand U322 (N_322,In_291,In_207);
nor U323 (N_323,In_57,In_126);
or U324 (N_324,In_97,In_61);
nor U325 (N_325,In_173,In_455);
nand U326 (N_326,In_431,In_418);
or U327 (N_327,In_194,In_310);
and U328 (N_328,In_477,In_252);
nor U329 (N_329,In_196,In_391);
nor U330 (N_330,In_492,In_401);
or U331 (N_331,In_175,In_136);
or U332 (N_332,In_325,In_339);
nor U333 (N_333,In_40,In_300);
and U334 (N_334,In_80,In_113);
xor U335 (N_335,In_253,In_78);
xor U336 (N_336,In_431,In_465);
xnor U337 (N_337,In_457,In_241);
and U338 (N_338,In_94,In_220);
and U339 (N_339,In_417,In_4);
nor U340 (N_340,In_70,In_259);
nand U341 (N_341,In_108,In_387);
nor U342 (N_342,In_185,In_451);
or U343 (N_343,In_304,In_67);
and U344 (N_344,In_157,In_122);
nor U345 (N_345,In_281,In_146);
xnor U346 (N_346,In_83,In_134);
nor U347 (N_347,In_189,In_473);
nand U348 (N_348,In_457,In_287);
and U349 (N_349,In_240,In_141);
nand U350 (N_350,In_302,In_462);
xor U351 (N_351,In_110,In_190);
nor U352 (N_352,In_346,In_357);
or U353 (N_353,In_78,In_377);
or U354 (N_354,In_79,In_110);
xnor U355 (N_355,In_115,In_263);
nand U356 (N_356,In_157,In_300);
nand U357 (N_357,In_325,In_288);
or U358 (N_358,In_122,In_117);
nand U359 (N_359,In_61,In_38);
or U360 (N_360,In_213,In_267);
or U361 (N_361,In_375,In_172);
nor U362 (N_362,In_72,In_288);
nor U363 (N_363,In_462,In_342);
and U364 (N_364,In_251,In_105);
nor U365 (N_365,In_328,In_373);
nand U366 (N_366,In_143,In_146);
xnor U367 (N_367,In_213,In_388);
nor U368 (N_368,In_284,In_442);
nand U369 (N_369,In_318,In_290);
nor U370 (N_370,In_232,In_484);
or U371 (N_371,In_164,In_143);
and U372 (N_372,In_446,In_234);
nor U373 (N_373,In_493,In_469);
nor U374 (N_374,In_76,In_113);
and U375 (N_375,In_359,In_323);
nand U376 (N_376,In_383,In_415);
and U377 (N_377,In_336,In_382);
xnor U378 (N_378,In_8,In_141);
or U379 (N_379,In_150,In_395);
or U380 (N_380,In_138,In_231);
nor U381 (N_381,In_379,In_58);
or U382 (N_382,In_473,In_293);
nand U383 (N_383,In_24,In_268);
nor U384 (N_384,In_59,In_72);
or U385 (N_385,In_237,In_340);
or U386 (N_386,In_322,In_399);
nor U387 (N_387,In_471,In_238);
or U388 (N_388,In_358,In_383);
nor U389 (N_389,In_349,In_57);
or U390 (N_390,In_169,In_367);
and U391 (N_391,In_250,In_457);
and U392 (N_392,In_164,In_28);
nand U393 (N_393,In_156,In_386);
nand U394 (N_394,In_125,In_281);
xnor U395 (N_395,In_299,In_376);
and U396 (N_396,In_208,In_240);
or U397 (N_397,In_301,In_473);
xnor U398 (N_398,In_449,In_263);
or U399 (N_399,In_252,In_165);
nand U400 (N_400,In_194,In_375);
nor U401 (N_401,In_405,In_11);
xnor U402 (N_402,In_86,In_263);
and U403 (N_403,In_458,In_199);
and U404 (N_404,In_381,In_55);
and U405 (N_405,In_11,In_133);
nand U406 (N_406,In_67,In_76);
nor U407 (N_407,In_400,In_25);
xor U408 (N_408,In_69,In_7);
nor U409 (N_409,In_1,In_398);
xnor U410 (N_410,In_389,In_1);
nor U411 (N_411,In_214,In_179);
or U412 (N_412,In_171,In_156);
nand U413 (N_413,In_469,In_384);
nand U414 (N_414,In_467,In_427);
and U415 (N_415,In_346,In_462);
nor U416 (N_416,In_44,In_414);
nor U417 (N_417,In_216,In_209);
xor U418 (N_418,In_422,In_420);
or U419 (N_419,In_401,In_279);
nand U420 (N_420,In_48,In_173);
nand U421 (N_421,In_245,In_463);
or U422 (N_422,In_27,In_330);
or U423 (N_423,In_349,In_84);
or U424 (N_424,In_254,In_130);
nor U425 (N_425,In_454,In_479);
xnor U426 (N_426,In_119,In_281);
xor U427 (N_427,In_207,In_432);
xnor U428 (N_428,In_173,In_74);
or U429 (N_429,In_462,In_152);
nor U430 (N_430,In_106,In_345);
nor U431 (N_431,In_56,In_479);
xnor U432 (N_432,In_82,In_323);
xnor U433 (N_433,In_46,In_76);
or U434 (N_434,In_496,In_194);
nor U435 (N_435,In_496,In_31);
xnor U436 (N_436,In_17,In_58);
or U437 (N_437,In_173,In_482);
xnor U438 (N_438,In_30,In_145);
and U439 (N_439,In_338,In_225);
and U440 (N_440,In_49,In_331);
xnor U441 (N_441,In_183,In_292);
nand U442 (N_442,In_441,In_292);
or U443 (N_443,In_193,In_173);
nand U444 (N_444,In_153,In_492);
and U445 (N_445,In_129,In_317);
nor U446 (N_446,In_8,In_226);
nor U447 (N_447,In_391,In_338);
xor U448 (N_448,In_311,In_264);
and U449 (N_449,In_206,In_443);
and U450 (N_450,In_41,In_8);
xnor U451 (N_451,In_100,In_444);
xor U452 (N_452,In_150,In_53);
and U453 (N_453,In_462,In_348);
and U454 (N_454,In_457,In_140);
and U455 (N_455,In_28,In_470);
and U456 (N_456,In_321,In_317);
nor U457 (N_457,In_154,In_136);
or U458 (N_458,In_441,In_188);
and U459 (N_459,In_228,In_201);
nand U460 (N_460,In_52,In_242);
nor U461 (N_461,In_412,In_93);
nor U462 (N_462,In_70,In_181);
nand U463 (N_463,In_443,In_110);
nand U464 (N_464,In_153,In_54);
and U465 (N_465,In_234,In_422);
or U466 (N_466,In_271,In_4);
nand U467 (N_467,In_363,In_420);
nand U468 (N_468,In_337,In_123);
nand U469 (N_469,In_43,In_129);
nand U470 (N_470,In_162,In_456);
and U471 (N_471,In_112,In_278);
or U472 (N_472,In_350,In_481);
xor U473 (N_473,In_272,In_107);
nor U474 (N_474,In_352,In_200);
xor U475 (N_475,In_488,In_438);
nor U476 (N_476,In_346,In_240);
or U477 (N_477,In_39,In_234);
xnor U478 (N_478,In_276,In_29);
xor U479 (N_479,In_371,In_413);
or U480 (N_480,In_77,In_468);
and U481 (N_481,In_254,In_494);
nand U482 (N_482,In_446,In_382);
nand U483 (N_483,In_159,In_487);
nand U484 (N_484,In_166,In_423);
xor U485 (N_485,In_470,In_475);
or U486 (N_486,In_394,In_480);
and U487 (N_487,In_409,In_488);
xor U488 (N_488,In_12,In_462);
nor U489 (N_489,In_245,In_369);
nor U490 (N_490,In_259,In_215);
nor U491 (N_491,In_236,In_144);
and U492 (N_492,In_406,In_301);
nor U493 (N_493,In_442,In_98);
nand U494 (N_494,In_272,In_140);
xor U495 (N_495,In_139,In_474);
nor U496 (N_496,In_79,In_344);
and U497 (N_497,In_84,In_49);
and U498 (N_498,In_11,In_395);
nor U499 (N_499,In_339,In_108);
nand U500 (N_500,In_355,In_33);
nand U501 (N_501,In_37,In_33);
xnor U502 (N_502,In_456,In_175);
nand U503 (N_503,In_277,In_247);
or U504 (N_504,In_234,In_493);
nand U505 (N_505,In_394,In_31);
or U506 (N_506,In_286,In_435);
nor U507 (N_507,In_364,In_29);
xnor U508 (N_508,In_428,In_255);
and U509 (N_509,In_293,In_445);
nor U510 (N_510,In_35,In_444);
and U511 (N_511,In_52,In_447);
and U512 (N_512,In_278,In_486);
or U513 (N_513,In_349,In_342);
or U514 (N_514,In_357,In_156);
and U515 (N_515,In_13,In_268);
nand U516 (N_516,In_491,In_189);
and U517 (N_517,In_416,In_471);
or U518 (N_518,In_52,In_117);
nor U519 (N_519,In_312,In_447);
nor U520 (N_520,In_118,In_112);
or U521 (N_521,In_452,In_348);
and U522 (N_522,In_481,In_229);
xor U523 (N_523,In_74,In_411);
xnor U524 (N_524,In_186,In_486);
nand U525 (N_525,In_103,In_129);
or U526 (N_526,In_235,In_306);
nand U527 (N_527,In_315,In_166);
nand U528 (N_528,In_197,In_164);
or U529 (N_529,In_310,In_372);
nand U530 (N_530,In_206,In_427);
nor U531 (N_531,In_188,In_318);
and U532 (N_532,In_439,In_237);
xor U533 (N_533,In_274,In_66);
nor U534 (N_534,In_385,In_421);
or U535 (N_535,In_364,In_220);
nor U536 (N_536,In_100,In_25);
nand U537 (N_537,In_285,In_334);
nor U538 (N_538,In_337,In_253);
nand U539 (N_539,In_455,In_413);
or U540 (N_540,In_414,In_71);
xor U541 (N_541,In_385,In_240);
nand U542 (N_542,In_164,In_456);
nand U543 (N_543,In_242,In_193);
and U544 (N_544,In_358,In_36);
nand U545 (N_545,In_384,In_375);
nand U546 (N_546,In_394,In_296);
or U547 (N_547,In_367,In_497);
xnor U548 (N_548,In_494,In_264);
nor U549 (N_549,In_122,In_255);
or U550 (N_550,In_232,In_26);
and U551 (N_551,In_80,In_319);
or U552 (N_552,In_22,In_260);
nor U553 (N_553,In_328,In_111);
and U554 (N_554,In_460,In_349);
nor U555 (N_555,In_69,In_17);
nor U556 (N_556,In_359,In_203);
and U557 (N_557,In_250,In_473);
xnor U558 (N_558,In_227,In_96);
nand U559 (N_559,In_28,In_486);
nand U560 (N_560,In_288,In_271);
nor U561 (N_561,In_200,In_433);
nor U562 (N_562,In_148,In_398);
and U563 (N_563,In_82,In_354);
nand U564 (N_564,In_452,In_449);
nand U565 (N_565,In_47,In_182);
nor U566 (N_566,In_69,In_491);
nand U567 (N_567,In_300,In_304);
xor U568 (N_568,In_483,In_343);
and U569 (N_569,In_19,In_206);
or U570 (N_570,In_426,In_100);
nand U571 (N_571,In_301,In_7);
nand U572 (N_572,In_156,In_84);
nor U573 (N_573,In_191,In_168);
and U574 (N_574,In_259,In_179);
and U575 (N_575,In_216,In_227);
and U576 (N_576,In_358,In_435);
nor U577 (N_577,In_296,In_186);
nand U578 (N_578,In_244,In_234);
or U579 (N_579,In_270,In_223);
nor U580 (N_580,In_265,In_131);
nor U581 (N_581,In_211,In_263);
and U582 (N_582,In_195,In_271);
nor U583 (N_583,In_19,In_70);
and U584 (N_584,In_400,In_79);
nand U585 (N_585,In_362,In_417);
or U586 (N_586,In_181,In_252);
or U587 (N_587,In_47,In_222);
nor U588 (N_588,In_364,In_287);
nor U589 (N_589,In_182,In_125);
and U590 (N_590,In_421,In_160);
and U591 (N_591,In_387,In_259);
nor U592 (N_592,In_143,In_67);
nor U593 (N_593,In_323,In_286);
nand U594 (N_594,In_199,In_163);
nand U595 (N_595,In_341,In_209);
nor U596 (N_596,In_306,In_301);
or U597 (N_597,In_318,In_87);
or U598 (N_598,In_33,In_400);
and U599 (N_599,In_165,In_82);
or U600 (N_600,N_559,N_539);
nor U601 (N_601,N_458,N_431);
nor U602 (N_602,N_482,N_134);
and U603 (N_603,N_288,N_466);
nor U604 (N_604,N_346,N_127);
or U605 (N_605,N_520,N_521);
xor U606 (N_606,N_102,N_473);
and U607 (N_607,N_506,N_548);
nand U608 (N_608,N_138,N_477);
or U609 (N_609,N_555,N_585);
nor U610 (N_610,N_315,N_461);
nor U611 (N_611,N_282,N_329);
nand U612 (N_612,N_440,N_434);
or U613 (N_613,N_25,N_170);
or U614 (N_614,N_422,N_536);
nor U615 (N_615,N_121,N_178);
and U616 (N_616,N_527,N_14);
xnor U617 (N_617,N_228,N_179);
xor U618 (N_618,N_216,N_165);
and U619 (N_619,N_50,N_151);
nor U620 (N_620,N_436,N_570);
nor U621 (N_621,N_441,N_38);
xnor U622 (N_622,N_572,N_129);
and U623 (N_623,N_556,N_567);
nor U624 (N_624,N_496,N_145);
nand U625 (N_625,N_10,N_388);
xor U626 (N_626,N_502,N_26);
nand U627 (N_627,N_116,N_15);
and U628 (N_628,N_231,N_428);
or U629 (N_629,N_375,N_300);
and U630 (N_630,N_190,N_4);
or U631 (N_631,N_381,N_128);
nand U632 (N_632,N_226,N_564);
or U633 (N_633,N_185,N_28);
nor U634 (N_634,N_443,N_135);
and U635 (N_635,N_132,N_297);
nor U636 (N_636,N_239,N_341);
nor U637 (N_637,N_211,N_480);
or U638 (N_638,N_513,N_435);
and U639 (N_639,N_212,N_317);
xor U640 (N_640,N_407,N_373);
nand U641 (N_641,N_318,N_319);
nor U642 (N_642,N_11,N_281);
and U643 (N_643,N_505,N_351);
nor U644 (N_644,N_68,N_543);
and U645 (N_645,N_425,N_159);
nor U646 (N_646,N_463,N_259);
and U647 (N_647,N_5,N_111);
nand U648 (N_648,N_308,N_143);
nor U649 (N_649,N_286,N_156);
nand U650 (N_650,N_194,N_336);
and U651 (N_651,N_123,N_574);
nand U652 (N_652,N_309,N_54);
nand U653 (N_653,N_568,N_538);
nor U654 (N_654,N_552,N_408);
nor U655 (N_655,N_331,N_219);
or U656 (N_656,N_485,N_540);
and U657 (N_657,N_354,N_587);
and U658 (N_658,N_217,N_209);
or U659 (N_659,N_291,N_472);
and U660 (N_660,N_376,N_1);
or U661 (N_661,N_389,N_563);
and U662 (N_662,N_426,N_530);
or U663 (N_663,N_130,N_36);
xor U664 (N_664,N_31,N_78);
nand U665 (N_665,N_84,N_204);
nor U666 (N_666,N_325,N_491);
xnor U667 (N_667,N_202,N_100);
nand U668 (N_668,N_122,N_504);
xor U669 (N_669,N_29,N_12);
nand U670 (N_670,N_531,N_87);
and U671 (N_671,N_0,N_30);
and U672 (N_672,N_103,N_582);
nor U673 (N_673,N_581,N_386);
nor U674 (N_674,N_283,N_23);
and U675 (N_675,N_478,N_141);
nor U676 (N_676,N_312,N_285);
xnor U677 (N_677,N_402,N_83);
or U678 (N_678,N_263,N_270);
or U679 (N_679,N_448,N_232);
or U680 (N_680,N_49,N_575);
or U681 (N_681,N_43,N_438);
and U682 (N_682,N_497,N_137);
nor U683 (N_683,N_119,N_313);
or U684 (N_684,N_230,N_61);
or U685 (N_685,N_526,N_363);
and U686 (N_686,N_278,N_79);
or U687 (N_687,N_105,N_411);
and U688 (N_688,N_593,N_366);
nor U689 (N_689,N_40,N_171);
nand U690 (N_690,N_13,N_189);
or U691 (N_691,N_72,N_580);
and U692 (N_692,N_592,N_522);
nand U693 (N_693,N_453,N_294);
or U694 (N_694,N_238,N_220);
and U695 (N_695,N_588,N_45);
nand U696 (N_696,N_335,N_508);
or U697 (N_697,N_409,N_410);
or U698 (N_698,N_140,N_390);
nor U699 (N_699,N_146,N_136);
and U700 (N_700,N_546,N_362);
or U701 (N_701,N_280,N_338);
and U702 (N_702,N_32,N_63);
nand U703 (N_703,N_21,N_17);
and U704 (N_704,N_305,N_579);
and U705 (N_705,N_244,N_553);
nand U706 (N_706,N_352,N_596);
and U707 (N_707,N_340,N_115);
nand U708 (N_708,N_598,N_88);
nor U709 (N_709,N_558,N_92);
nand U710 (N_710,N_457,N_406);
nand U711 (N_711,N_347,N_562);
or U712 (N_712,N_94,N_152);
nand U713 (N_713,N_258,N_494);
or U714 (N_714,N_333,N_166);
and U715 (N_715,N_423,N_169);
or U716 (N_716,N_233,N_549);
and U717 (N_717,N_70,N_157);
and U718 (N_718,N_235,N_284);
and U719 (N_719,N_243,N_515);
nor U720 (N_720,N_371,N_56);
nand U721 (N_721,N_184,N_274);
nand U722 (N_722,N_266,N_468);
nand U723 (N_723,N_516,N_39);
nor U724 (N_724,N_77,N_131);
nor U725 (N_725,N_348,N_501);
nand U726 (N_726,N_399,N_277);
nor U727 (N_727,N_566,N_193);
and U728 (N_728,N_203,N_481);
nor U729 (N_729,N_160,N_383);
nand U730 (N_730,N_427,N_551);
nand U731 (N_731,N_339,N_471);
and U732 (N_732,N_295,N_484);
nand U733 (N_733,N_330,N_58);
or U734 (N_734,N_20,N_89);
nor U735 (N_735,N_413,N_391);
and U736 (N_736,N_86,N_155);
nor U737 (N_737,N_392,N_377);
nor U738 (N_738,N_418,N_361);
and U739 (N_739,N_71,N_27);
and U740 (N_740,N_99,N_430);
or U741 (N_741,N_421,N_256);
or U742 (N_742,N_149,N_173);
and U743 (N_743,N_595,N_241);
nor U744 (N_744,N_469,N_349);
and U745 (N_745,N_55,N_483);
xor U746 (N_746,N_161,N_174);
nand U747 (N_747,N_343,N_344);
nor U748 (N_748,N_419,N_367);
xor U749 (N_749,N_52,N_442);
and U750 (N_750,N_37,N_359);
and U751 (N_751,N_60,N_205);
and U752 (N_752,N_109,N_208);
or U753 (N_753,N_251,N_187);
or U754 (N_754,N_275,N_69);
and U755 (N_755,N_192,N_240);
xnor U756 (N_756,N_493,N_433);
xor U757 (N_757,N_577,N_65);
or U758 (N_758,N_75,N_301);
nand U759 (N_759,N_142,N_401);
and U760 (N_760,N_7,N_268);
or U761 (N_761,N_269,N_215);
xnor U762 (N_762,N_287,N_307);
and U763 (N_763,N_133,N_565);
nor U764 (N_764,N_467,N_304);
nand U765 (N_765,N_112,N_255);
or U766 (N_766,N_517,N_227);
or U767 (N_767,N_372,N_544);
nor U768 (N_768,N_465,N_554);
or U769 (N_769,N_261,N_120);
nor U770 (N_770,N_221,N_511);
nor U771 (N_771,N_380,N_108);
and U772 (N_772,N_200,N_8);
and U773 (N_773,N_403,N_498);
nand U774 (N_774,N_198,N_486);
or U775 (N_775,N_162,N_42);
nor U776 (N_776,N_529,N_196);
nor U777 (N_777,N_455,N_487);
and U778 (N_778,N_85,N_124);
nor U779 (N_779,N_97,N_514);
xnor U780 (N_780,N_207,N_365);
nand U781 (N_781,N_289,N_404);
nor U782 (N_782,N_424,N_327);
nor U783 (N_783,N_569,N_345);
or U784 (N_784,N_46,N_334);
xor U785 (N_785,N_573,N_597);
or U786 (N_786,N_186,N_67);
nand U787 (N_787,N_394,N_57);
nand U788 (N_788,N_479,N_321);
nand U789 (N_789,N_512,N_523);
and U790 (N_790,N_534,N_48);
or U791 (N_791,N_254,N_107);
and U792 (N_792,N_492,N_265);
nor U793 (N_793,N_16,N_364);
and U794 (N_794,N_393,N_303);
nor U795 (N_795,N_62,N_414);
nand U796 (N_796,N_510,N_296);
nor U797 (N_797,N_550,N_326);
nor U798 (N_798,N_535,N_519);
nor U799 (N_799,N_81,N_398);
xnor U800 (N_800,N_495,N_248);
nand U801 (N_801,N_368,N_182);
and U802 (N_802,N_397,N_314);
nor U803 (N_803,N_576,N_450);
and U804 (N_804,N_74,N_118);
nor U805 (N_805,N_73,N_34);
nand U806 (N_806,N_452,N_3);
nand U807 (N_807,N_499,N_594);
nor U808 (N_808,N_279,N_311);
nor U809 (N_809,N_528,N_324);
nand U810 (N_810,N_474,N_415);
nand U811 (N_811,N_144,N_350);
xor U812 (N_812,N_267,N_489);
or U813 (N_813,N_545,N_584);
nand U814 (N_814,N_225,N_53);
nand U815 (N_815,N_395,N_176);
nor U816 (N_816,N_420,N_378);
and U817 (N_817,N_396,N_260);
nor U818 (N_818,N_306,N_101);
or U819 (N_819,N_412,N_249);
nand U820 (N_820,N_250,N_292);
or U821 (N_821,N_405,N_44);
nor U822 (N_822,N_560,N_387);
nor U823 (N_823,N_446,N_591);
xnor U824 (N_824,N_183,N_416);
nand U825 (N_825,N_51,N_172);
nor U826 (N_826,N_201,N_356);
nor U827 (N_827,N_518,N_195);
nand U828 (N_828,N_117,N_459);
or U829 (N_829,N_533,N_599);
and U830 (N_830,N_561,N_475);
or U831 (N_831,N_320,N_547);
and U832 (N_832,N_271,N_180);
nor U833 (N_833,N_328,N_525);
and U834 (N_834,N_299,N_444);
nor U835 (N_835,N_488,N_578);
nor U836 (N_836,N_242,N_106);
nor U837 (N_837,N_264,N_247);
xnor U838 (N_838,N_33,N_357);
nand U839 (N_839,N_589,N_91);
and U840 (N_840,N_384,N_47);
nor U841 (N_841,N_164,N_293);
and U842 (N_842,N_150,N_110);
or U843 (N_843,N_272,N_125);
nand U844 (N_844,N_24,N_358);
or U845 (N_845,N_234,N_210);
xor U846 (N_846,N_22,N_456);
or U847 (N_847,N_503,N_188);
or U848 (N_848,N_126,N_276);
nor U849 (N_849,N_9,N_18);
and U850 (N_850,N_175,N_590);
nand U851 (N_851,N_177,N_273);
and U852 (N_852,N_59,N_6);
and U853 (N_853,N_41,N_76);
nor U854 (N_854,N_237,N_332);
or U855 (N_855,N_439,N_337);
nand U856 (N_856,N_583,N_449);
nand U857 (N_857,N_429,N_500);
nor U858 (N_858,N_537,N_353);
or U859 (N_859,N_197,N_90);
or U860 (N_860,N_451,N_66);
and U861 (N_861,N_379,N_213);
or U862 (N_862,N_153,N_206);
and U863 (N_863,N_298,N_360);
nor U864 (N_864,N_342,N_586);
and U865 (N_865,N_432,N_222);
nor U866 (N_866,N_96,N_223);
nor U867 (N_867,N_382,N_95);
nor U868 (N_868,N_93,N_370);
nor U869 (N_869,N_437,N_236);
and U870 (N_870,N_104,N_400);
and U871 (N_871,N_158,N_218);
and U872 (N_872,N_252,N_509);
or U873 (N_873,N_417,N_524);
nor U874 (N_874,N_470,N_290);
xor U875 (N_875,N_245,N_355);
nor U876 (N_876,N_323,N_385);
nand U877 (N_877,N_229,N_82);
nor U878 (N_878,N_262,N_257);
nor U879 (N_879,N_181,N_316);
nand U880 (N_880,N_191,N_302);
nand U881 (N_881,N_445,N_310);
xor U882 (N_882,N_542,N_163);
or U883 (N_883,N_19,N_2);
xor U884 (N_884,N_447,N_168);
and U885 (N_885,N_64,N_253);
and U886 (N_886,N_139,N_148);
and U887 (N_887,N_454,N_541);
and U888 (N_888,N_113,N_246);
nor U889 (N_889,N_507,N_322);
nand U890 (N_890,N_224,N_464);
or U891 (N_891,N_476,N_490);
or U892 (N_892,N_460,N_80);
xnor U893 (N_893,N_114,N_167);
nand U894 (N_894,N_154,N_98);
nor U895 (N_895,N_199,N_369);
or U896 (N_896,N_147,N_214);
xnor U897 (N_897,N_571,N_532);
and U898 (N_898,N_557,N_35);
nor U899 (N_899,N_374,N_462);
or U900 (N_900,N_119,N_299);
nor U901 (N_901,N_406,N_99);
nand U902 (N_902,N_566,N_39);
and U903 (N_903,N_564,N_155);
nand U904 (N_904,N_203,N_83);
xor U905 (N_905,N_506,N_362);
and U906 (N_906,N_500,N_390);
nand U907 (N_907,N_137,N_255);
nor U908 (N_908,N_129,N_113);
or U909 (N_909,N_139,N_258);
xor U910 (N_910,N_53,N_253);
nand U911 (N_911,N_12,N_62);
nand U912 (N_912,N_314,N_421);
or U913 (N_913,N_64,N_390);
nor U914 (N_914,N_234,N_570);
and U915 (N_915,N_83,N_122);
or U916 (N_916,N_277,N_556);
nor U917 (N_917,N_261,N_11);
nor U918 (N_918,N_302,N_401);
xor U919 (N_919,N_0,N_329);
or U920 (N_920,N_417,N_74);
and U921 (N_921,N_19,N_453);
nand U922 (N_922,N_20,N_284);
or U923 (N_923,N_455,N_326);
and U924 (N_924,N_351,N_300);
or U925 (N_925,N_31,N_80);
and U926 (N_926,N_383,N_407);
or U927 (N_927,N_13,N_497);
nor U928 (N_928,N_462,N_335);
or U929 (N_929,N_532,N_462);
or U930 (N_930,N_523,N_210);
xnor U931 (N_931,N_530,N_498);
or U932 (N_932,N_11,N_274);
nor U933 (N_933,N_321,N_314);
and U934 (N_934,N_340,N_190);
and U935 (N_935,N_365,N_448);
or U936 (N_936,N_99,N_43);
xor U937 (N_937,N_260,N_287);
nor U938 (N_938,N_309,N_215);
nand U939 (N_939,N_413,N_466);
nand U940 (N_940,N_104,N_23);
nor U941 (N_941,N_469,N_450);
nor U942 (N_942,N_76,N_142);
nand U943 (N_943,N_12,N_572);
nand U944 (N_944,N_259,N_558);
or U945 (N_945,N_158,N_466);
and U946 (N_946,N_334,N_404);
and U947 (N_947,N_520,N_127);
nand U948 (N_948,N_487,N_231);
nor U949 (N_949,N_463,N_448);
xor U950 (N_950,N_441,N_175);
xnor U951 (N_951,N_73,N_590);
or U952 (N_952,N_574,N_24);
nor U953 (N_953,N_535,N_261);
or U954 (N_954,N_227,N_462);
and U955 (N_955,N_109,N_173);
or U956 (N_956,N_545,N_67);
or U957 (N_957,N_188,N_131);
nor U958 (N_958,N_76,N_177);
or U959 (N_959,N_132,N_358);
nand U960 (N_960,N_111,N_83);
or U961 (N_961,N_241,N_312);
or U962 (N_962,N_467,N_446);
and U963 (N_963,N_404,N_305);
nand U964 (N_964,N_160,N_173);
or U965 (N_965,N_358,N_444);
nor U966 (N_966,N_59,N_56);
and U967 (N_967,N_178,N_80);
nand U968 (N_968,N_206,N_340);
or U969 (N_969,N_395,N_82);
nor U970 (N_970,N_550,N_585);
nor U971 (N_971,N_568,N_172);
and U972 (N_972,N_128,N_524);
or U973 (N_973,N_305,N_385);
or U974 (N_974,N_199,N_570);
or U975 (N_975,N_584,N_212);
or U976 (N_976,N_257,N_432);
xor U977 (N_977,N_174,N_215);
nand U978 (N_978,N_592,N_263);
and U979 (N_979,N_568,N_169);
or U980 (N_980,N_281,N_556);
or U981 (N_981,N_264,N_495);
and U982 (N_982,N_533,N_156);
or U983 (N_983,N_305,N_148);
xor U984 (N_984,N_352,N_485);
nand U985 (N_985,N_576,N_282);
and U986 (N_986,N_427,N_199);
or U987 (N_987,N_254,N_546);
or U988 (N_988,N_3,N_94);
and U989 (N_989,N_6,N_252);
nand U990 (N_990,N_372,N_501);
and U991 (N_991,N_64,N_69);
nor U992 (N_992,N_244,N_520);
nand U993 (N_993,N_60,N_218);
and U994 (N_994,N_300,N_80);
nor U995 (N_995,N_252,N_177);
nand U996 (N_996,N_578,N_141);
nor U997 (N_997,N_127,N_195);
or U998 (N_998,N_522,N_231);
xnor U999 (N_999,N_389,N_451);
nor U1000 (N_1000,N_462,N_149);
xnor U1001 (N_1001,N_48,N_47);
nor U1002 (N_1002,N_79,N_582);
nor U1003 (N_1003,N_514,N_556);
and U1004 (N_1004,N_212,N_250);
and U1005 (N_1005,N_161,N_464);
or U1006 (N_1006,N_437,N_102);
xnor U1007 (N_1007,N_261,N_587);
or U1008 (N_1008,N_337,N_29);
nand U1009 (N_1009,N_235,N_84);
and U1010 (N_1010,N_276,N_291);
nor U1011 (N_1011,N_14,N_267);
or U1012 (N_1012,N_263,N_261);
nand U1013 (N_1013,N_218,N_554);
and U1014 (N_1014,N_475,N_130);
or U1015 (N_1015,N_355,N_140);
and U1016 (N_1016,N_414,N_387);
nor U1017 (N_1017,N_270,N_147);
and U1018 (N_1018,N_497,N_238);
xor U1019 (N_1019,N_183,N_18);
or U1020 (N_1020,N_543,N_26);
or U1021 (N_1021,N_369,N_249);
or U1022 (N_1022,N_99,N_354);
nor U1023 (N_1023,N_103,N_406);
and U1024 (N_1024,N_201,N_80);
or U1025 (N_1025,N_159,N_445);
nor U1026 (N_1026,N_118,N_571);
nand U1027 (N_1027,N_486,N_72);
nor U1028 (N_1028,N_161,N_572);
and U1029 (N_1029,N_56,N_475);
nand U1030 (N_1030,N_302,N_222);
nor U1031 (N_1031,N_100,N_159);
and U1032 (N_1032,N_298,N_436);
nand U1033 (N_1033,N_176,N_153);
or U1034 (N_1034,N_144,N_164);
nor U1035 (N_1035,N_575,N_172);
xor U1036 (N_1036,N_486,N_244);
xor U1037 (N_1037,N_242,N_457);
or U1038 (N_1038,N_410,N_224);
nor U1039 (N_1039,N_30,N_421);
xnor U1040 (N_1040,N_455,N_290);
nand U1041 (N_1041,N_238,N_477);
nand U1042 (N_1042,N_201,N_549);
nand U1043 (N_1043,N_305,N_493);
nand U1044 (N_1044,N_489,N_193);
or U1045 (N_1045,N_579,N_1);
nor U1046 (N_1046,N_202,N_336);
and U1047 (N_1047,N_9,N_436);
nand U1048 (N_1048,N_416,N_265);
nor U1049 (N_1049,N_560,N_124);
or U1050 (N_1050,N_353,N_146);
and U1051 (N_1051,N_393,N_147);
and U1052 (N_1052,N_585,N_27);
and U1053 (N_1053,N_364,N_383);
nor U1054 (N_1054,N_446,N_513);
nand U1055 (N_1055,N_153,N_256);
xor U1056 (N_1056,N_79,N_315);
and U1057 (N_1057,N_247,N_296);
nand U1058 (N_1058,N_380,N_220);
nand U1059 (N_1059,N_599,N_399);
nand U1060 (N_1060,N_168,N_246);
nor U1061 (N_1061,N_557,N_222);
or U1062 (N_1062,N_350,N_256);
nand U1063 (N_1063,N_481,N_116);
or U1064 (N_1064,N_461,N_434);
nand U1065 (N_1065,N_162,N_524);
nand U1066 (N_1066,N_512,N_425);
nor U1067 (N_1067,N_422,N_340);
nor U1068 (N_1068,N_204,N_210);
xnor U1069 (N_1069,N_238,N_479);
nand U1070 (N_1070,N_288,N_347);
nand U1071 (N_1071,N_583,N_520);
nand U1072 (N_1072,N_78,N_390);
or U1073 (N_1073,N_411,N_491);
and U1074 (N_1074,N_22,N_428);
or U1075 (N_1075,N_211,N_241);
and U1076 (N_1076,N_340,N_355);
nand U1077 (N_1077,N_23,N_551);
or U1078 (N_1078,N_152,N_248);
and U1079 (N_1079,N_464,N_440);
nor U1080 (N_1080,N_208,N_328);
nor U1081 (N_1081,N_409,N_170);
nor U1082 (N_1082,N_349,N_104);
nor U1083 (N_1083,N_244,N_576);
xor U1084 (N_1084,N_68,N_472);
nor U1085 (N_1085,N_456,N_282);
and U1086 (N_1086,N_271,N_307);
or U1087 (N_1087,N_234,N_22);
xnor U1088 (N_1088,N_492,N_546);
nand U1089 (N_1089,N_379,N_197);
nand U1090 (N_1090,N_335,N_502);
nand U1091 (N_1091,N_160,N_288);
xnor U1092 (N_1092,N_401,N_591);
nand U1093 (N_1093,N_370,N_55);
and U1094 (N_1094,N_286,N_323);
nor U1095 (N_1095,N_137,N_569);
and U1096 (N_1096,N_42,N_545);
nor U1097 (N_1097,N_511,N_525);
or U1098 (N_1098,N_547,N_46);
and U1099 (N_1099,N_473,N_323);
nor U1100 (N_1100,N_296,N_181);
nand U1101 (N_1101,N_469,N_333);
nor U1102 (N_1102,N_225,N_156);
and U1103 (N_1103,N_251,N_246);
nand U1104 (N_1104,N_17,N_27);
nand U1105 (N_1105,N_154,N_449);
or U1106 (N_1106,N_564,N_380);
and U1107 (N_1107,N_373,N_352);
nor U1108 (N_1108,N_36,N_351);
nor U1109 (N_1109,N_593,N_370);
or U1110 (N_1110,N_6,N_321);
nor U1111 (N_1111,N_240,N_440);
nand U1112 (N_1112,N_280,N_370);
nor U1113 (N_1113,N_377,N_320);
nand U1114 (N_1114,N_11,N_562);
xnor U1115 (N_1115,N_335,N_596);
and U1116 (N_1116,N_83,N_216);
nand U1117 (N_1117,N_164,N_591);
nor U1118 (N_1118,N_97,N_58);
or U1119 (N_1119,N_453,N_160);
nor U1120 (N_1120,N_56,N_132);
or U1121 (N_1121,N_572,N_241);
or U1122 (N_1122,N_409,N_43);
nand U1123 (N_1123,N_407,N_435);
or U1124 (N_1124,N_387,N_358);
nor U1125 (N_1125,N_243,N_575);
nand U1126 (N_1126,N_219,N_96);
nand U1127 (N_1127,N_296,N_538);
or U1128 (N_1128,N_442,N_46);
nand U1129 (N_1129,N_333,N_557);
nand U1130 (N_1130,N_413,N_147);
nor U1131 (N_1131,N_27,N_339);
and U1132 (N_1132,N_225,N_320);
nand U1133 (N_1133,N_336,N_190);
nand U1134 (N_1134,N_138,N_385);
nor U1135 (N_1135,N_584,N_216);
nand U1136 (N_1136,N_264,N_221);
and U1137 (N_1137,N_328,N_266);
or U1138 (N_1138,N_243,N_213);
or U1139 (N_1139,N_132,N_0);
or U1140 (N_1140,N_538,N_507);
nor U1141 (N_1141,N_409,N_535);
xnor U1142 (N_1142,N_149,N_160);
nand U1143 (N_1143,N_369,N_593);
nand U1144 (N_1144,N_8,N_591);
nor U1145 (N_1145,N_90,N_292);
nand U1146 (N_1146,N_588,N_593);
and U1147 (N_1147,N_245,N_289);
or U1148 (N_1148,N_378,N_259);
nor U1149 (N_1149,N_559,N_175);
and U1150 (N_1150,N_549,N_35);
nor U1151 (N_1151,N_383,N_453);
nand U1152 (N_1152,N_401,N_293);
or U1153 (N_1153,N_395,N_51);
or U1154 (N_1154,N_79,N_363);
nor U1155 (N_1155,N_185,N_457);
nor U1156 (N_1156,N_434,N_156);
and U1157 (N_1157,N_211,N_125);
and U1158 (N_1158,N_373,N_28);
nor U1159 (N_1159,N_81,N_355);
nand U1160 (N_1160,N_581,N_240);
nor U1161 (N_1161,N_11,N_417);
nand U1162 (N_1162,N_0,N_378);
nor U1163 (N_1163,N_305,N_228);
nor U1164 (N_1164,N_442,N_526);
or U1165 (N_1165,N_520,N_328);
nor U1166 (N_1166,N_110,N_302);
nor U1167 (N_1167,N_336,N_4);
or U1168 (N_1168,N_566,N_305);
xnor U1169 (N_1169,N_3,N_176);
or U1170 (N_1170,N_71,N_208);
nor U1171 (N_1171,N_521,N_108);
or U1172 (N_1172,N_463,N_450);
nand U1173 (N_1173,N_135,N_103);
xor U1174 (N_1174,N_143,N_586);
nand U1175 (N_1175,N_595,N_314);
xor U1176 (N_1176,N_102,N_52);
and U1177 (N_1177,N_344,N_445);
nand U1178 (N_1178,N_448,N_352);
and U1179 (N_1179,N_89,N_138);
nor U1180 (N_1180,N_351,N_192);
and U1181 (N_1181,N_487,N_187);
and U1182 (N_1182,N_29,N_398);
or U1183 (N_1183,N_439,N_186);
nor U1184 (N_1184,N_476,N_355);
or U1185 (N_1185,N_287,N_107);
and U1186 (N_1186,N_534,N_347);
xor U1187 (N_1187,N_547,N_408);
xor U1188 (N_1188,N_153,N_117);
nand U1189 (N_1189,N_388,N_159);
nand U1190 (N_1190,N_71,N_496);
or U1191 (N_1191,N_480,N_315);
nand U1192 (N_1192,N_505,N_166);
nor U1193 (N_1193,N_154,N_336);
and U1194 (N_1194,N_554,N_464);
or U1195 (N_1195,N_82,N_420);
and U1196 (N_1196,N_197,N_148);
nand U1197 (N_1197,N_539,N_28);
or U1198 (N_1198,N_238,N_119);
xor U1199 (N_1199,N_51,N_164);
nor U1200 (N_1200,N_686,N_659);
nand U1201 (N_1201,N_868,N_732);
xor U1202 (N_1202,N_694,N_925);
nand U1203 (N_1203,N_802,N_909);
or U1204 (N_1204,N_819,N_828);
nand U1205 (N_1205,N_1169,N_1117);
nor U1206 (N_1206,N_863,N_839);
and U1207 (N_1207,N_973,N_701);
nor U1208 (N_1208,N_1156,N_649);
nor U1209 (N_1209,N_616,N_1153);
nand U1210 (N_1210,N_789,N_1036);
and U1211 (N_1211,N_662,N_641);
and U1212 (N_1212,N_642,N_637);
xor U1213 (N_1213,N_1050,N_699);
or U1214 (N_1214,N_1178,N_869);
nand U1215 (N_1215,N_1171,N_1148);
nor U1216 (N_1216,N_1077,N_1186);
and U1217 (N_1217,N_823,N_874);
xnor U1218 (N_1218,N_1127,N_799);
or U1219 (N_1219,N_1170,N_896);
or U1220 (N_1220,N_1062,N_794);
nand U1221 (N_1221,N_1071,N_887);
or U1222 (N_1222,N_850,N_962);
nor U1223 (N_1223,N_1031,N_872);
and U1224 (N_1224,N_693,N_1033);
nand U1225 (N_1225,N_1003,N_740);
nand U1226 (N_1226,N_1124,N_1012);
nor U1227 (N_1227,N_646,N_861);
and U1228 (N_1228,N_716,N_947);
or U1229 (N_1229,N_747,N_1181);
and U1230 (N_1230,N_767,N_835);
or U1231 (N_1231,N_758,N_1191);
nor U1232 (N_1232,N_1000,N_972);
and U1233 (N_1233,N_1058,N_1111);
nand U1234 (N_1234,N_908,N_954);
xor U1235 (N_1235,N_1122,N_812);
nand U1236 (N_1236,N_911,N_1073);
or U1237 (N_1237,N_682,N_731);
nand U1238 (N_1238,N_772,N_854);
xor U1239 (N_1239,N_940,N_820);
and U1240 (N_1240,N_784,N_1080);
nor U1241 (N_1241,N_620,N_1149);
or U1242 (N_1242,N_933,N_907);
or U1243 (N_1243,N_991,N_1070);
nor U1244 (N_1244,N_1116,N_974);
nand U1245 (N_1245,N_1199,N_1079);
xnor U1246 (N_1246,N_1142,N_1189);
or U1247 (N_1247,N_664,N_999);
nand U1248 (N_1248,N_1106,N_929);
xnor U1249 (N_1249,N_916,N_622);
xnor U1250 (N_1250,N_844,N_808);
nor U1251 (N_1251,N_1087,N_845);
nand U1252 (N_1252,N_1167,N_1025);
nor U1253 (N_1253,N_827,N_853);
or U1254 (N_1254,N_702,N_866);
and U1255 (N_1255,N_1018,N_724);
nand U1256 (N_1256,N_1016,N_886);
nor U1257 (N_1257,N_696,N_1134);
or U1258 (N_1258,N_743,N_661);
and U1259 (N_1259,N_1023,N_735);
and U1260 (N_1260,N_993,N_1039);
nor U1261 (N_1261,N_1188,N_807);
nand U1262 (N_1262,N_782,N_1060);
nor U1263 (N_1263,N_1034,N_1193);
xnor U1264 (N_1264,N_793,N_1183);
and U1265 (N_1265,N_1173,N_1053);
nor U1266 (N_1266,N_904,N_1040);
nand U1267 (N_1267,N_1175,N_977);
or U1268 (N_1268,N_1104,N_707);
or U1269 (N_1269,N_848,N_779);
nand U1270 (N_1270,N_665,N_1126);
nand U1271 (N_1271,N_990,N_805);
nor U1272 (N_1272,N_912,N_1184);
nand U1273 (N_1273,N_858,N_697);
or U1274 (N_1274,N_674,N_618);
nand U1275 (N_1275,N_768,N_945);
and U1276 (N_1276,N_1054,N_870);
and U1277 (N_1277,N_1119,N_1030);
nor U1278 (N_1278,N_1125,N_836);
and U1279 (N_1279,N_915,N_856);
or U1280 (N_1280,N_1084,N_1051);
and U1281 (N_1281,N_1007,N_989);
nor U1282 (N_1282,N_725,N_1118);
nand U1283 (N_1283,N_1044,N_903);
nand U1284 (N_1284,N_838,N_1152);
or U1285 (N_1285,N_619,N_1158);
and U1286 (N_1286,N_1064,N_803);
nor U1287 (N_1287,N_1086,N_759);
nand U1288 (N_1288,N_749,N_917);
nand U1289 (N_1289,N_842,N_834);
and U1290 (N_1290,N_1081,N_656);
or U1291 (N_1291,N_624,N_713);
or U1292 (N_1292,N_780,N_944);
nor U1293 (N_1293,N_1174,N_1163);
nand U1294 (N_1294,N_1042,N_1093);
or U1295 (N_1295,N_613,N_718);
or U1296 (N_1296,N_652,N_660);
nor U1297 (N_1297,N_756,N_901);
or U1298 (N_1298,N_968,N_1105);
nand U1299 (N_1299,N_1066,N_636);
nand U1300 (N_1300,N_638,N_764);
nor U1301 (N_1301,N_643,N_817);
or U1302 (N_1302,N_971,N_942);
nor U1303 (N_1303,N_1147,N_683);
and U1304 (N_1304,N_985,N_918);
or U1305 (N_1305,N_1078,N_737);
or U1306 (N_1306,N_1197,N_634);
nand U1307 (N_1307,N_1021,N_1056);
nor U1308 (N_1308,N_964,N_1138);
nand U1309 (N_1309,N_607,N_988);
and U1310 (N_1310,N_1090,N_709);
or U1311 (N_1311,N_738,N_730);
or U1312 (N_1312,N_824,N_753);
or U1313 (N_1313,N_645,N_992);
nand U1314 (N_1314,N_966,N_891);
nand U1315 (N_1315,N_995,N_1097);
nand U1316 (N_1316,N_611,N_809);
nand U1317 (N_1317,N_935,N_1095);
xnor U1318 (N_1318,N_884,N_1008);
nor U1319 (N_1319,N_797,N_957);
or U1320 (N_1320,N_609,N_1146);
nor U1321 (N_1321,N_792,N_936);
nor U1322 (N_1322,N_913,N_1195);
or U1323 (N_1323,N_679,N_692);
and U1324 (N_1324,N_1168,N_1182);
and U1325 (N_1325,N_1075,N_1004);
or U1326 (N_1326,N_1143,N_1094);
and U1327 (N_1327,N_855,N_644);
nor U1328 (N_1328,N_762,N_804);
xor U1329 (N_1329,N_695,N_728);
nor U1330 (N_1330,N_841,N_606);
or U1331 (N_1331,N_996,N_905);
and U1332 (N_1332,N_705,N_932);
or U1333 (N_1333,N_1194,N_965);
nand U1334 (N_1334,N_734,N_859);
nand U1335 (N_1335,N_960,N_1096);
nor U1336 (N_1336,N_1068,N_847);
or U1337 (N_1337,N_1179,N_830);
nand U1338 (N_1338,N_640,N_885);
and U1339 (N_1339,N_748,N_1082);
or U1340 (N_1340,N_635,N_983);
xnor U1341 (N_1341,N_750,N_773);
nor U1342 (N_1342,N_1133,N_818);
nor U1343 (N_1343,N_938,N_941);
or U1344 (N_1344,N_744,N_951);
nand U1345 (N_1345,N_687,N_1061);
and U1346 (N_1346,N_895,N_790);
xnor U1347 (N_1347,N_976,N_733);
nor U1348 (N_1348,N_1135,N_787);
and U1349 (N_1349,N_608,N_1114);
or U1350 (N_1350,N_663,N_715);
nor U1351 (N_1351,N_684,N_952);
and U1352 (N_1352,N_603,N_1164);
nand U1353 (N_1353,N_771,N_956);
nor U1354 (N_1354,N_1043,N_722);
nand U1355 (N_1355,N_927,N_939);
nor U1356 (N_1356,N_751,N_979);
nor U1357 (N_1357,N_655,N_1067);
and U1358 (N_1358,N_876,N_1131);
and U1359 (N_1359,N_1045,N_857);
xor U1360 (N_1360,N_1128,N_1115);
and U1361 (N_1361,N_978,N_986);
nor U1362 (N_1362,N_1121,N_778);
nor U1363 (N_1363,N_760,N_926);
nand U1364 (N_1364,N_1102,N_680);
nor U1365 (N_1365,N_681,N_1047);
or U1366 (N_1366,N_1002,N_897);
and U1367 (N_1367,N_1177,N_628);
or U1368 (N_1368,N_610,N_651);
and U1369 (N_1369,N_1052,N_706);
nand U1370 (N_1370,N_967,N_955);
nand U1371 (N_1371,N_821,N_1013);
nor U1372 (N_1372,N_1091,N_1123);
and U1373 (N_1373,N_814,N_623);
and U1374 (N_1374,N_1072,N_658);
or U1375 (N_1375,N_1019,N_906);
and U1376 (N_1376,N_648,N_1162);
nor U1377 (N_1377,N_711,N_982);
or U1378 (N_1378,N_1176,N_948);
nand U1379 (N_1379,N_969,N_710);
or U1380 (N_1380,N_627,N_741);
or U1381 (N_1381,N_1166,N_1150);
or U1382 (N_1382,N_1109,N_1088);
nor U1383 (N_1383,N_796,N_1196);
or U1384 (N_1384,N_1057,N_1083);
and U1385 (N_1385,N_700,N_1159);
nand U1386 (N_1386,N_775,N_1038);
and U1387 (N_1387,N_677,N_883);
nand U1388 (N_1388,N_688,N_795);
or U1389 (N_1389,N_1139,N_825);
or U1390 (N_1390,N_840,N_879);
nor U1391 (N_1391,N_602,N_934);
nor U1392 (N_1392,N_647,N_852);
and U1393 (N_1393,N_1136,N_1157);
and U1394 (N_1394,N_1028,N_763);
xor U1395 (N_1395,N_1006,N_961);
and U1396 (N_1396,N_1035,N_777);
or U1397 (N_1397,N_984,N_980);
nand U1398 (N_1398,N_893,N_843);
xor U1399 (N_1399,N_987,N_630);
or U1400 (N_1400,N_1165,N_667);
and U1401 (N_1401,N_943,N_1132);
or U1402 (N_1402,N_832,N_846);
nand U1403 (N_1403,N_1112,N_1137);
or U1404 (N_1404,N_902,N_867);
and U1405 (N_1405,N_629,N_1048);
or U1406 (N_1406,N_785,N_921);
nand U1407 (N_1407,N_822,N_770);
nor U1408 (N_1408,N_754,N_1140);
and U1409 (N_1409,N_774,N_837);
nor U1410 (N_1410,N_1024,N_704);
and U1411 (N_1411,N_875,N_708);
xnor U1412 (N_1412,N_676,N_1198);
or U1413 (N_1413,N_1161,N_878);
xor U1414 (N_1414,N_626,N_765);
and U1415 (N_1415,N_949,N_1107);
nor U1416 (N_1416,N_877,N_1037);
nand U1417 (N_1417,N_650,N_757);
nand U1418 (N_1418,N_1049,N_761);
and U1419 (N_1419,N_1144,N_1145);
or U1420 (N_1420,N_1010,N_1085);
or U1421 (N_1421,N_1110,N_666);
or U1422 (N_1422,N_1022,N_1113);
nand U1423 (N_1423,N_1185,N_953);
nand U1424 (N_1424,N_1092,N_669);
nor U1425 (N_1425,N_865,N_691);
nand U1426 (N_1426,N_975,N_1026);
and U1427 (N_1427,N_899,N_752);
xnor U1428 (N_1428,N_849,N_690);
and U1429 (N_1429,N_717,N_970);
or U1430 (N_1430,N_633,N_673);
nand U1431 (N_1431,N_1020,N_798);
nor U1432 (N_1432,N_851,N_880);
nand U1433 (N_1433,N_721,N_654);
nand U1434 (N_1434,N_703,N_829);
and U1435 (N_1435,N_810,N_1059);
nor U1436 (N_1436,N_723,N_745);
and U1437 (N_1437,N_800,N_806);
xnor U1438 (N_1438,N_746,N_1017);
xnor U1439 (N_1439,N_727,N_922);
or U1440 (N_1440,N_1160,N_813);
nor U1441 (N_1441,N_924,N_882);
or U1442 (N_1442,N_1011,N_698);
xor U1443 (N_1443,N_788,N_889);
and U1444 (N_1444,N_689,N_1100);
or U1445 (N_1445,N_1190,N_1001);
and U1446 (N_1446,N_959,N_1055);
or U1447 (N_1447,N_950,N_1099);
nor U1448 (N_1448,N_958,N_726);
nand U1449 (N_1449,N_1172,N_675);
and U1450 (N_1450,N_930,N_900);
and U1451 (N_1451,N_712,N_781);
nor U1452 (N_1452,N_672,N_791);
and U1453 (N_1453,N_1154,N_631);
nor U1454 (N_1454,N_668,N_981);
xor U1455 (N_1455,N_1151,N_1108);
or U1456 (N_1456,N_1014,N_1141);
nor U1457 (N_1457,N_1129,N_1041);
and U1458 (N_1458,N_1032,N_671);
nand U1459 (N_1459,N_815,N_920);
xor U1460 (N_1460,N_625,N_621);
or U1461 (N_1461,N_605,N_720);
or U1462 (N_1462,N_1005,N_1009);
and U1463 (N_1463,N_614,N_657);
or U1464 (N_1464,N_1101,N_888);
nand U1465 (N_1465,N_881,N_776);
nand U1466 (N_1466,N_615,N_860);
nor U1467 (N_1467,N_601,N_862);
and U1468 (N_1468,N_714,N_739);
and U1469 (N_1469,N_1069,N_833);
nand U1470 (N_1470,N_914,N_1065);
and U1471 (N_1471,N_755,N_1155);
and U1472 (N_1472,N_1089,N_653);
nand U1473 (N_1473,N_963,N_617);
or U1474 (N_1474,N_811,N_719);
and U1475 (N_1475,N_890,N_604);
nor U1476 (N_1476,N_998,N_1074);
nand U1477 (N_1477,N_997,N_873);
nor U1478 (N_1478,N_1120,N_931);
and U1479 (N_1479,N_816,N_1103);
nor U1480 (N_1480,N_946,N_612);
nor U1481 (N_1481,N_678,N_729);
or U1482 (N_1482,N_1076,N_801);
and U1483 (N_1483,N_1015,N_632);
nor U1484 (N_1484,N_1192,N_831);
and U1485 (N_1485,N_766,N_1027);
nor U1486 (N_1486,N_994,N_1187);
and U1487 (N_1487,N_742,N_892);
xnor U1488 (N_1488,N_871,N_826);
or U1489 (N_1489,N_786,N_919);
and U1490 (N_1490,N_1029,N_670);
xnor U1491 (N_1491,N_769,N_783);
nand U1492 (N_1492,N_894,N_937);
xor U1493 (N_1493,N_1046,N_1098);
nor U1494 (N_1494,N_736,N_910);
or U1495 (N_1495,N_1180,N_864);
nor U1496 (N_1496,N_898,N_928);
xor U1497 (N_1497,N_923,N_639);
or U1498 (N_1498,N_1063,N_1130);
or U1499 (N_1499,N_685,N_600);
and U1500 (N_1500,N_738,N_854);
and U1501 (N_1501,N_877,N_827);
and U1502 (N_1502,N_999,N_876);
xnor U1503 (N_1503,N_612,N_1148);
or U1504 (N_1504,N_1170,N_658);
or U1505 (N_1505,N_962,N_986);
xor U1506 (N_1506,N_608,N_691);
and U1507 (N_1507,N_922,N_802);
or U1508 (N_1508,N_803,N_1021);
or U1509 (N_1509,N_1039,N_977);
nor U1510 (N_1510,N_905,N_838);
xor U1511 (N_1511,N_626,N_907);
and U1512 (N_1512,N_709,N_734);
or U1513 (N_1513,N_854,N_1048);
nor U1514 (N_1514,N_883,N_898);
and U1515 (N_1515,N_653,N_879);
or U1516 (N_1516,N_684,N_686);
nor U1517 (N_1517,N_845,N_776);
nor U1518 (N_1518,N_1018,N_765);
nand U1519 (N_1519,N_679,N_906);
and U1520 (N_1520,N_941,N_783);
or U1521 (N_1521,N_775,N_857);
and U1522 (N_1522,N_667,N_796);
nor U1523 (N_1523,N_1096,N_1107);
or U1524 (N_1524,N_640,N_755);
xor U1525 (N_1525,N_1037,N_1034);
and U1526 (N_1526,N_668,N_1050);
or U1527 (N_1527,N_1000,N_1128);
or U1528 (N_1528,N_1005,N_972);
nor U1529 (N_1529,N_897,N_764);
nand U1530 (N_1530,N_1103,N_821);
nor U1531 (N_1531,N_893,N_784);
and U1532 (N_1532,N_1130,N_1191);
and U1533 (N_1533,N_1103,N_854);
nand U1534 (N_1534,N_779,N_790);
or U1535 (N_1535,N_687,N_874);
or U1536 (N_1536,N_695,N_965);
xnor U1537 (N_1537,N_731,N_875);
nand U1538 (N_1538,N_913,N_834);
nor U1539 (N_1539,N_1095,N_798);
xnor U1540 (N_1540,N_706,N_1100);
nand U1541 (N_1541,N_713,N_1029);
and U1542 (N_1542,N_694,N_913);
nor U1543 (N_1543,N_906,N_794);
and U1544 (N_1544,N_1074,N_993);
nand U1545 (N_1545,N_1130,N_1068);
xor U1546 (N_1546,N_714,N_933);
or U1547 (N_1547,N_1134,N_753);
xnor U1548 (N_1548,N_1113,N_673);
and U1549 (N_1549,N_687,N_780);
nand U1550 (N_1550,N_1150,N_1035);
or U1551 (N_1551,N_1016,N_743);
nor U1552 (N_1552,N_1130,N_787);
nand U1553 (N_1553,N_1085,N_635);
or U1554 (N_1554,N_715,N_665);
nand U1555 (N_1555,N_702,N_779);
or U1556 (N_1556,N_670,N_854);
and U1557 (N_1557,N_1103,N_1147);
nand U1558 (N_1558,N_939,N_863);
and U1559 (N_1559,N_649,N_933);
nor U1560 (N_1560,N_923,N_637);
and U1561 (N_1561,N_709,N_1034);
nor U1562 (N_1562,N_1114,N_1069);
or U1563 (N_1563,N_798,N_990);
xnor U1564 (N_1564,N_907,N_937);
nand U1565 (N_1565,N_1114,N_1195);
and U1566 (N_1566,N_822,N_681);
or U1567 (N_1567,N_981,N_1054);
or U1568 (N_1568,N_696,N_1099);
nor U1569 (N_1569,N_1002,N_952);
nor U1570 (N_1570,N_1033,N_1029);
xor U1571 (N_1571,N_1144,N_1023);
or U1572 (N_1572,N_621,N_1192);
and U1573 (N_1573,N_633,N_606);
and U1574 (N_1574,N_1084,N_682);
xnor U1575 (N_1575,N_998,N_705);
or U1576 (N_1576,N_1137,N_1065);
nand U1577 (N_1577,N_1038,N_769);
xor U1578 (N_1578,N_1105,N_836);
nand U1579 (N_1579,N_741,N_873);
and U1580 (N_1580,N_977,N_1149);
xnor U1581 (N_1581,N_977,N_1005);
xnor U1582 (N_1582,N_1099,N_858);
nand U1583 (N_1583,N_859,N_1038);
and U1584 (N_1584,N_1139,N_774);
xnor U1585 (N_1585,N_854,N_1082);
and U1586 (N_1586,N_897,N_656);
nor U1587 (N_1587,N_844,N_675);
or U1588 (N_1588,N_975,N_1058);
or U1589 (N_1589,N_1021,N_827);
nor U1590 (N_1590,N_649,N_1000);
nand U1591 (N_1591,N_944,N_648);
and U1592 (N_1592,N_676,N_1121);
or U1593 (N_1593,N_842,N_884);
or U1594 (N_1594,N_628,N_1133);
xnor U1595 (N_1595,N_635,N_651);
nor U1596 (N_1596,N_872,N_1038);
and U1597 (N_1597,N_1051,N_979);
and U1598 (N_1598,N_782,N_708);
and U1599 (N_1599,N_950,N_683);
nand U1600 (N_1600,N_1004,N_1184);
and U1601 (N_1601,N_1193,N_1083);
nand U1602 (N_1602,N_757,N_791);
nor U1603 (N_1603,N_1139,N_917);
nor U1604 (N_1604,N_638,N_1056);
or U1605 (N_1605,N_1111,N_619);
xnor U1606 (N_1606,N_967,N_1177);
and U1607 (N_1607,N_968,N_681);
xnor U1608 (N_1608,N_955,N_768);
and U1609 (N_1609,N_644,N_678);
or U1610 (N_1610,N_704,N_1064);
or U1611 (N_1611,N_668,N_714);
and U1612 (N_1612,N_883,N_969);
or U1613 (N_1613,N_886,N_1185);
nor U1614 (N_1614,N_1040,N_1119);
nand U1615 (N_1615,N_663,N_728);
or U1616 (N_1616,N_707,N_1123);
or U1617 (N_1617,N_952,N_1062);
or U1618 (N_1618,N_825,N_927);
nor U1619 (N_1619,N_1078,N_664);
nand U1620 (N_1620,N_1141,N_1136);
nor U1621 (N_1621,N_787,N_988);
xnor U1622 (N_1622,N_974,N_889);
nor U1623 (N_1623,N_953,N_851);
nor U1624 (N_1624,N_1147,N_813);
nand U1625 (N_1625,N_670,N_709);
nor U1626 (N_1626,N_1193,N_724);
or U1627 (N_1627,N_1113,N_1068);
nand U1628 (N_1628,N_1152,N_1129);
or U1629 (N_1629,N_1086,N_617);
nand U1630 (N_1630,N_855,N_1188);
and U1631 (N_1631,N_882,N_863);
or U1632 (N_1632,N_812,N_1131);
nand U1633 (N_1633,N_1015,N_656);
and U1634 (N_1634,N_1198,N_852);
nor U1635 (N_1635,N_894,N_1198);
or U1636 (N_1636,N_1182,N_922);
or U1637 (N_1637,N_808,N_896);
nor U1638 (N_1638,N_1113,N_1069);
and U1639 (N_1639,N_1116,N_682);
nand U1640 (N_1640,N_670,N_693);
nor U1641 (N_1641,N_756,N_1106);
or U1642 (N_1642,N_935,N_1075);
or U1643 (N_1643,N_651,N_906);
or U1644 (N_1644,N_870,N_1109);
xnor U1645 (N_1645,N_805,N_979);
nor U1646 (N_1646,N_930,N_1168);
and U1647 (N_1647,N_984,N_798);
and U1648 (N_1648,N_1199,N_1034);
and U1649 (N_1649,N_696,N_1089);
nand U1650 (N_1650,N_950,N_1107);
and U1651 (N_1651,N_935,N_604);
nor U1652 (N_1652,N_1195,N_1160);
nor U1653 (N_1653,N_936,N_1078);
nor U1654 (N_1654,N_897,N_600);
nand U1655 (N_1655,N_789,N_1026);
and U1656 (N_1656,N_652,N_888);
or U1657 (N_1657,N_1168,N_977);
or U1658 (N_1658,N_1150,N_852);
nor U1659 (N_1659,N_1061,N_674);
or U1660 (N_1660,N_983,N_1085);
nand U1661 (N_1661,N_793,N_752);
nand U1662 (N_1662,N_722,N_1049);
or U1663 (N_1663,N_762,N_604);
and U1664 (N_1664,N_1137,N_769);
and U1665 (N_1665,N_625,N_1191);
and U1666 (N_1666,N_636,N_781);
or U1667 (N_1667,N_915,N_622);
or U1668 (N_1668,N_864,N_749);
and U1669 (N_1669,N_971,N_959);
nand U1670 (N_1670,N_994,N_1183);
nor U1671 (N_1671,N_773,N_623);
and U1672 (N_1672,N_604,N_994);
nor U1673 (N_1673,N_1131,N_783);
nand U1674 (N_1674,N_964,N_623);
nor U1675 (N_1675,N_729,N_638);
and U1676 (N_1676,N_610,N_1031);
nand U1677 (N_1677,N_761,N_1173);
xor U1678 (N_1678,N_633,N_950);
nor U1679 (N_1679,N_673,N_676);
nor U1680 (N_1680,N_1120,N_1103);
and U1681 (N_1681,N_1189,N_1136);
or U1682 (N_1682,N_819,N_1156);
xnor U1683 (N_1683,N_866,N_669);
or U1684 (N_1684,N_729,N_921);
or U1685 (N_1685,N_685,N_962);
nor U1686 (N_1686,N_1001,N_852);
nand U1687 (N_1687,N_670,N_781);
and U1688 (N_1688,N_914,N_847);
xor U1689 (N_1689,N_941,N_754);
or U1690 (N_1690,N_656,N_1041);
xor U1691 (N_1691,N_1118,N_894);
nor U1692 (N_1692,N_670,N_807);
or U1693 (N_1693,N_1166,N_753);
nor U1694 (N_1694,N_1132,N_970);
nand U1695 (N_1695,N_1075,N_722);
or U1696 (N_1696,N_964,N_970);
nand U1697 (N_1697,N_1136,N_1047);
or U1698 (N_1698,N_620,N_785);
and U1699 (N_1699,N_880,N_606);
and U1700 (N_1700,N_806,N_802);
nor U1701 (N_1701,N_858,N_834);
nand U1702 (N_1702,N_673,N_1087);
nand U1703 (N_1703,N_1019,N_850);
and U1704 (N_1704,N_863,N_1011);
and U1705 (N_1705,N_1077,N_676);
or U1706 (N_1706,N_604,N_833);
nor U1707 (N_1707,N_1190,N_928);
nor U1708 (N_1708,N_839,N_718);
and U1709 (N_1709,N_854,N_1145);
nand U1710 (N_1710,N_796,N_1159);
nor U1711 (N_1711,N_1170,N_1068);
or U1712 (N_1712,N_859,N_1190);
xor U1713 (N_1713,N_625,N_605);
and U1714 (N_1714,N_819,N_620);
or U1715 (N_1715,N_1118,N_682);
xnor U1716 (N_1716,N_740,N_1017);
nor U1717 (N_1717,N_1103,N_811);
and U1718 (N_1718,N_1154,N_647);
nor U1719 (N_1719,N_755,N_720);
or U1720 (N_1720,N_638,N_679);
nor U1721 (N_1721,N_654,N_836);
and U1722 (N_1722,N_1186,N_920);
nand U1723 (N_1723,N_1086,N_638);
nand U1724 (N_1724,N_812,N_975);
nor U1725 (N_1725,N_1042,N_913);
nand U1726 (N_1726,N_972,N_1178);
or U1727 (N_1727,N_1021,N_897);
and U1728 (N_1728,N_861,N_1042);
and U1729 (N_1729,N_990,N_977);
and U1730 (N_1730,N_775,N_911);
and U1731 (N_1731,N_1043,N_1106);
xor U1732 (N_1732,N_1199,N_1107);
or U1733 (N_1733,N_714,N_1094);
nor U1734 (N_1734,N_757,N_1183);
or U1735 (N_1735,N_1143,N_805);
and U1736 (N_1736,N_631,N_1106);
nor U1737 (N_1737,N_769,N_1168);
nor U1738 (N_1738,N_976,N_675);
or U1739 (N_1739,N_1009,N_1130);
nor U1740 (N_1740,N_614,N_775);
or U1741 (N_1741,N_1115,N_953);
or U1742 (N_1742,N_670,N_846);
nor U1743 (N_1743,N_841,N_1168);
xnor U1744 (N_1744,N_915,N_843);
nor U1745 (N_1745,N_922,N_878);
xnor U1746 (N_1746,N_1124,N_1006);
nor U1747 (N_1747,N_750,N_935);
nor U1748 (N_1748,N_749,N_942);
and U1749 (N_1749,N_1070,N_720);
and U1750 (N_1750,N_1154,N_868);
or U1751 (N_1751,N_909,N_924);
and U1752 (N_1752,N_888,N_717);
and U1753 (N_1753,N_1162,N_604);
and U1754 (N_1754,N_782,N_1015);
nor U1755 (N_1755,N_916,N_1053);
nand U1756 (N_1756,N_812,N_1018);
xor U1757 (N_1757,N_974,N_952);
nand U1758 (N_1758,N_730,N_1056);
nand U1759 (N_1759,N_604,N_693);
nand U1760 (N_1760,N_680,N_1104);
xor U1761 (N_1761,N_895,N_682);
and U1762 (N_1762,N_1087,N_1113);
or U1763 (N_1763,N_759,N_1103);
nor U1764 (N_1764,N_730,N_948);
nor U1765 (N_1765,N_876,N_671);
nor U1766 (N_1766,N_1009,N_742);
or U1767 (N_1767,N_673,N_900);
and U1768 (N_1768,N_670,N_999);
or U1769 (N_1769,N_1087,N_915);
and U1770 (N_1770,N_847,N_680);
nand U1771 (N_1771,N_1079,N_1156);
or U1772 (N_1772,N_974,N_885);
nor U1773 (N_1773,N_685,N_1022);
nor U1774 (N_1774,N_1033,N_852);
nor U1775 (N_1775,N_1078,N_646);
nor U1776 (N_1776,N_752,N_971);
and U1777 (N_1777,N_624,N_993);
or U1778 (N_1778,N_744,N_1032);
nor U1779 (N_1779,N_774,N_677);
and U1780 (N_1780,N_773,N_749);
or U1781 (N_1781,N_875,N_910);
nor U1782 (N_1782,N_1082,N_841);
nor U1783 (N_1783,N_735,N_1128);
and U1784 (N_1784,N_757,N_896);
nor U1785 (N_1785,N_1021,N_845);
nand U1786 (N_1786,N_936,N_933);
xor U1787 (N_1787,N_1163,N_1080);
xor U1788 (N_1788,N_1009,N_809);
nor U1789 (N_1789,N_752,N_1023);
and U1790 (N_1790,N_751,N_619);
xnor U1791 (N_1791,N_1080,N_958);
xnor U1792 (N_1792,N_962,N_738);
nand U1793 (N_1793,N_873,N_952);
and U1794 (N_1794,N_796,N_676);
xor U1795 (N_1795,N_955,N_1165);
or U1796 (N_1796,N_1182,N_982);
or U1797 (N_1797,N_877,N_809);
or U1798 (N_1798,N_633,N_1108);
or U1799 (N_1799,N_912,N_822);
and U1800 (N_1800,N_1641,N_1734);
and U1801 (N_1801,N_1787,N_1224);
nand U1802 (N_1802,N_1435,N_1769);
nor U1803 (N_1803,N_1572,N_1253);
xnor U1804 (N_1804,N_1430,N_1603);
nand U1805 (N_1805,N_1609,N_1447);
nand U1806 (N_1806,N_1379,N_1343);
nand U1807 (N_1807,N_1710,N_1776);
or U1808 (N_1808,N_1254,N_1522);
or U1809 (N_1809,N_1216,N_1271);
and U1810 (N_1810,N_1296,N_1506);
and U1811 (N_1811,N_1477,N_1546);
or U1812 (N_1812,N_1453,N_1606);
or U1813 (N_1813,N_1576,N_1735);
nand U1814 (N_1814,N_1708,N_1358);
and U1815 (N_1815,N_1528,N_1535);
xor U1816 (N_1816,N_1442,N_1539);
or U1817 (N_1817,N_1421,N_1246);
or U1818 (N_1818,N_1268,N_1459);
and U1819 (N_1819,N_1423,N_1542);
xnor U1820 (N_1820,N_1631,N_1645);
xor U1821 (N_1821,N_1479,N_1628);
and U1822 (N_1822,N_1327,N_1329);
nor U1823 (N_1823,N_1222,N_1277);
nor U1824 (N_1824,N_1719,N_1554);
xor U1825 (N_1825,N_1368,N_1771);
and U1826 (N_1826,N_1693,N_1515);
and U1827 (N_1827,N_1386,N_1387);
nand U1828 (N_1828,N_1591,N_1404);
nand U1829 (N_1829,N_1574,N_1629);
and U1830 (N_1830,N_1360,N_1309);
nand U1831 (N_1831,N_1491,N_1418);
xor U1832 (N_1832,N_1626,N_1793);
or U1833 (N_1833,N_1429,N_1310);
nor U1834 (N_1834,N_1208,N_1434);
xor U1835 (N_1835,N_1750,N_1560);
or U1836 (N_1836,N_1243,N_1478);
nand U1837 (N_1837,N_1403,N_1786);
and U1838 (N_1838,N_1215,N_1538);
nor U1839 (N_1839,N_1303,N_1685);
nor U1840 (N_1840,N_1739,N_1596);
or U1841 (N_1841,N_1751,N_1695);
xnor U1842 (N_1842,N_1394,N_1696);
nor U1843 (N_1843,N_1728,N_1266);
xor U1844 (N_1844,N_1627,N_1647);
and U1845 (N_1845,N_1231,N_1294);
nor U1846 (N_1846,N_1411,N_1683);
nor U1847 (N_1847,N_1748,N_1533);
xor U1848 (N_1848,N_1670,N_1264);
or U1849 (N_1849,N_1571,N_1514);
nor U1850 (N_1850,N_1233,N_1474);
nand U1851 (N_1851,N_1770,N_1798);
nor U1852 (N_1852,N_1331,N_1509);
or U1853 (N_1853,N_1284,N_1472);
nand U1854 (N_1854,N_1402,N_1413);
xnor U1855 (N_1855,N_1414,N_1427);
and U1856 (N_1856,N_1220,N_1649);
nand U1857 (N_1857,N_1541,N_1682);
nor U1858 (N_1858,N_1616,N_1729);
or U1859 (N_1859,N_1451,N_1741);
nor U1860 (N_1860,N_1717,N_1704);
and U1861 (N_1861,N_1740,N_1633);
nor U1862 (N_1862,N_1496,N_1230);
nand U1863 (N_1863,N_1356,N_1274);
xnor U1864 (N_1864,N_1625,N_1256);
and U1865 (N_1865,N_1621,N_1499);
nor U1866 (N_1866,N_1595,N_1565);
and U1867 (N_1867,N_1369,N_1476);
nand U1868 (N_1868,N_1531,N_1635);
nor U1869 (N_1869,N_1460,N_1723);
and U1870 (N_1870,N_1799,N_1619);
or U1871 (N_1871,N_1357,N_1273);
nor U1872 (N_1872,N_1382,N_1761);
nand U1873 (N_1873,N_1438,N_1305);
nand U1874 (N_1874,N_1431,N_1397);
and U1875 (N_1875,N_1237,N_1597);
nand U1876 (N_1876,N_1458,N_1601);
nor U1877 (N_1877,N_1433,N_1325);
or U1878 (N_1878,N_1784,N_1569);
nand U1879 (N_1879,N_1668,N_1275);
or U1880 (N_1880,N_1393,N_1241);
xor U1881 (N_1881,N_1406,N_1385);
nand U1882 (N_1882,N_1405,N_1390);
or U1883 (N_1883,N_1228,N_1760);
nor U1884 (N_1884,N_1753,N_1785);
or U1885 (N_1885,N_1267,N_1321);
nand U1886 (N_1886,N_1234,N_1529);
nand U1887 (N_1887,N_1745,N_1319);
and U1888 (N_1888,N_1507,N_1240);
or U1889 (N_1889,N_1440,N_1342);
nor U1890 (N_1890,N_1672,N_1518);
or U1891 (N_1891,N_1372,N_1444);
nor U1892 (N_1892,N_1422,N_1468);
nand U1893 (N_1893,N_1441,N_1485);
nor U1894 (N_1894,N_1756,N_1324);
nor U1895 (N_1895,N_1643,N_1494);
nor U1896 (N_1896,N_1791,N_1558);
and U1897 (N_1897,N_1346,N_1795);
xnor U1898 (N_1898,N_1295,N_1681);
nor U1899 (N_1899,N_1653,N_1260);
and U1900 (N_1900,N_1502,N_1248);
xnor U1901 (N_1901,N_1466,N_1646);
xor U1902 (N_1902,N_1450,N_1725);
nand U1903 (N_1903,N_1680,N_1280);
or U1904 (N_1904,N_1510,N_1252);
or U1905 (N_1905,N_1424,N_1408);
nor U1906 (N_1906,N_1209,N_1768);
and U1907 (N_1907,N_1512,N_1772);
nand U1908 (N_1908,N_1287,N_1634);
and U1909 (N_1909,N_1655,N_1376);
or U1910 (N_1910,N_1794,N_1561);
and U1911 (N_1911,N_1666,N_1698);
or U1912 (N_1912,N_1722,N_1437);
nand U1913 (N_1913,N_1604,N_1373);
nor U1914 (N_1914,N_1201,N_1553);
and U1915 (N_1915,N_1777,N_1480);
nor U1916 (N_1916,N_1232,N_1624);
or U1917 (N_1917,N_1694,N_1497);
or U1918 (N_1918,N_1333,N_1521);
nand U1919 (N_1919,N_1416,N_1299);
and U1920 (N_1920,N_1605,N_1773);
or U1921 (N_1921,N_1487,N_1742);
nor U1922 (N_1922,N_1720,N_1223);
nand U1923 (N_1923,N_1678,N_1545);
or U1924 (N_1924,N_1314,N_1524);
nor U1925 (N_1925,N_1270,N_1302);
nor U1926 (N_1926,N_1501,N_1613);
or U1927 (N_1927,N_1259,N_1242);
nor U1928 (N_1928,N_1712,N_1349);
or U1929 (N_1929,N_1570,N_1283);
or U1930 (N_1930,N_1548,N_1623);
nor U1931 (N_1931,N_1348,N_1426);
nor U1932 (N_1932,N_1486,N_1790);
nand U1933 (N_1933,N_1315,N_1263);
nor U1934 (N_1934,N_1508,N_1203);
and U1935 (N_1935,N_1205,N_1383);
or U1936 (N_1936,N_1513,N_1493);
nand U1937 (N_1937,N_1732,N_1339);
nor U1938 (N_1938,N_1419,N_1610);
or U1939 (N_1939,N_1550,N_1395);
or U1940 (N_1940,N_1318,N_1622);
nand U1941 (N_1941,N_1225,N_1367);
nand U1942 (N_1942,N_1279,N_1792);
or U1943 (N_1943,N_1443,N_1257);
nand U1944 (N_1944,N_1519,N_1779);
nand U1945 (N_1945,N_1557,N_1781);
and U1946 (N_1946,N_1488,N_1323);
or U1947 (N_1947,N_1640,N_1705);
nand U1948 (N_1948,N_1639,N_1612);
and U1949 (N_1949,N_1312,N_1286);
and U1950 (N_1950,N_1738,N_1330);
or U1951 (N_1951,N_1755,N_1638);
or U1952 (N_1952,N_1465,N_1620);
nand U1953 (N_1953,N_1552,N_1326);
and U1954 (N_1954,N_1446,N_1361);
nor U1955 (N_1955,N_1204,N_1445);
and U1956 (N_1956,N_1592,N_1229);
nand U1957 (N_1957,N_1463,N_1677);
xor U1958 (N_1958,N_1401,N_1316);
nand U1959 (N_1959,N_1285,N_1660);
nand U1960 (N_1960,N_1359,N_1389);
and U1961 (N_1961,N_1363,N_1354);
nand U1962 (N_1962,N_1311,N_1674);
or U1963 (N_1963,N_1365,N_1328);
or U1964 (N_1964,N_1600,N_1733);
and U1965 (N_1965,N_1731,N_1200);
nand U1966 (N_1966,N_1654,N_1530);
and U1967 (N_1967,N_1617,N_1543);
nor U1968 (N_1968,N_1308,N_1355);
or U1969 (N_1969,N_1532,N_1300);
or U1970 (N_1970,N_1523,N_1650);
nor U1971 (N_1971,N_1338,N_1218);
xnor U1972 (N_1972,N_1667,N_1227);
or U1973 (N_1973,N_1448,N_1239);
or U1974 (N_1974,N_1375,N_1526);
xor U1975 (N_1975,N_1797,N_1580);
xnor U1976 (N_1976,N_1614,N_1262);
nand U1977 (N_1977,N_1214,N_1636);
or U1978 (N_1978,N_1691,N_1258);
nor U1979 (N_1979,N_1737,N_1492);
or U1980 (N_1980,N_1454,N_1762);
nand U1981 (N_1981,N_1575,N_1747);
or U1982 (N_1982,N_1251,N_1377);
nor U1983 (N_1983,N_1727,N_1384);
nand U1984 (N_1984,N_1202,N_1744);
and U1985 (N_1985,N_1527,N_1743);
nand U1986 (N_1986,N_1707,N_1703);
nand U1987 (N_1987,N_1307,N_1481);
or U1988 (N_1988,N_1566,N_1313);
and U1989 (N_1989,N_1400,N_1767);
nor U1990 (N_1990,N_1412,N_1544);
or U1991 (N_1991,N_1334,N_1556);
xnor U1992 (N_1992,N_1632,N_1716);
xnor U1993 (N_1993,N_1503,N_1516);
nor U1994 (N_1994,N_1436,N_1581);
or U1995 (N_1995,N_1495,N_1352);
or U1996 (N_1996,N_1206,N_1505);
xor U1997 (N_1997,N_1297,N_1700);
and U1998 (N_1998,N_1415,N_1517);
xnor U1999 (N_1999,N_1238,N_1549);
nor U2000 (N_2000,N_1235,N_1362);
or U2001 (N_2001,N_1469,N_1679);
nor U2002 (N_2002,N_1726,N_1588);
and U2003 (N_2003,N_1461,N_1317);
nor U2004 (N_2004,N_1563,N_1226);
or U2005 (N_2005,N_1537,N_1462);
nor U2006 (N_2006,N_1714,N_1337);
or U2007 (N_2007,N_1380,N_1425);
nor U2008 (N_2008,N_1608,N_1378);
and U2009 (N_2009,N_1410,N_1336);
or U2010 (N_2010,N_1540,N_1483);
or U2011 (N_2011,N_1715,N_1599);
nor U2012 (N_2012,N_1269,N_1706);
or U2013 (N_2013,N_1536,N_1351);
nor U2014 (N_2014,N_1661,N_1290);
nor U2015 (N_2015,N_1702,N_1618);
or U2016 (N_2016,N_1675,N_1688);
nand U2017 (N_2017,N_1371,N_1511);
and U2018 (N_2018,N_1344,N_1607);
or U2019 (N_2019,N_1210,N_1250);
xor U2020 (N_2020,N_1292,N_1207);
nor U2021 (N_2021,N_1370,N_1345);
nor U2022 (N_2022,N_1759,N_1669);
nor U2023 (N_2023,N_1663,N_1432);
or U2024 (N_2024,N_1789,N_1244);
nand U2025 (N_2025,N_1775,N_1573);
xor U2026 (N_2026,N_1340,N_1579);
or U2027 (N_2027,N_1615,N_1288);
and U2028 (N_2028,N_1304,N_1651);
or U2029 (N_2029,N_1417,N_1648);
xor U2030 (N_2030,N_1664,N_1261);
or U2031 (N_2031,N_1709,N_1428);
nor U2032 (N_2032,N_1464,N_1322);
nand U2033 (N_2033,N_1455,N_1611);
nor U2034 (N_2034,N_1652,N_1746);
nor U2035 (N_2035,N_1347,N_1673);
nor U2036 (N_2036,N_1590,N_1467);
or U2037 (N_2037,N_1656,N_1765);
or U2038 (N_2038,N_1484,N_1594);
xnor U2039 (N_2039,N_1697,N_1212);
nand U2040 (N_2040,N_1783,N_1249);
xor U2041 (N_2041,N_1276,N_1724);
and U2042 (N_2042,N_1291,N_1452);
or U2043 (N_2043,N_1602,N_1713);
nor U2044 (N_2044,N_1551,N_1374);
nand U2045 (N_2045,N_1457,N_1490);
nand U2046 (N_2046,N_1657,N_1420);
nor U2047 (N_2047,N_1396,N_1350);
xor U2048 (N_2048,N_1564,N_1562);
or U2049 (N_2049,N_1236,N_1388);
or U2050 (N_2050,N_1585,N_1662);
nor U2051 (N_2051,N_1782,N_1578);
nand U2052 (N_2052,N_1439,N_1341);
or U2053 (N_2053,N_1278,N_1780);
nand U2054 (N_2054,N_1353,N_1763);
and U2055 (N_2055,N_1247,N_1301);
or U2056 (N_2056,N_1730,N_1520);
xor U2057 (N_2057,N_1534,N_1399);
nor U2058 (N_2058,N_1589,N_1407);
nor U2059 (N_2059,N_1475,N_1749);
nand U2060 (N_2060,N_1449,N_1699);
nor U2061 (N_2061,N_1686,N_1689);
nand U2062 (N_2062,N_1582,N_1593);
and U2063 (N_2063,N_1217,N_1473);
nand U2064 (N_2064,N_1676,N_1788);
or U2065 (N_2065,N_1255,N_1381);
or U2066 (N_2066,N_1711,N_1555);
and U2067 (N_2067,N_1721,N_1687);
and U2068 (N_2068,N_1754,N_1736);
nand U2069 (N_2069,N_1644,N_1659);
and U2070 (N_2070,N_1547,N_1690);
and U2071 (N_2071,N_1306,N_1364);
xor U2072 (N_2072,N_1586,N_1482);
nor U2073 (N_2073,N_1752,N_1692);
nand U2074 (N_2074,N_1525,N_1598);
nor U2075 (N_2075,N_1671,N_1587);
or U2076 (N_2076,N_1796,N_1245);
or U2077 (N_2077,N_1630,N_1366);
nand U2078 (N_2078,N_1642,N_1559);
nand U2079 (N_2079,N_1219,N_1658);
and U2080 (N_2080,N_1289,N_1398);
and U2081 (N_2081,N_1335,N_1211);
nor U2082 (N_2082,N_1213,N_1221);
xor U2083 (N_2083,N_1470,N_1504);
and U2084 (N_2084,N_1584,N_1684);
or U2085 (N_2085,N_1766,N_1332);
nor U2086 (N_2086,N_1583,N_1409);
nand U2087 (N_2087,N_1272,N_1778);
nor U2088 (N_2088,N_1282,N_1471);
xnor U2089 (N_2089,N_1701,N_1764);
or U2090 (N_2090,N_1718,N_1757);
nor U2091 (N_2091,N_1489,N_1391);
nor U2092 (N_2092,N_1298,N_1577);
nand U2093 (N_2093,N_1758,N_1392);
and U2094 (N_2094,N_1774,N_1281);
and U2095 (N_2095,N_1568,N_1293);
and U2096 (N_2096,N_1320,N_1567);
or U2097 (N_2097,N_1265,N_1498);
or U2098 (N_2098,N_1637,N_1456);
xor U2099 (N_2099,N_1665,N_1500);
nand U2100 (N_2100,N_1304,N_1604);
nand U2101 (N_2101,N_1670,N_1777);
or U2102 (N_2102,N_1596,N_1560);
or U2103 (N_2103,N_1687,N_1605);
xnor U2104 (N_2104,N_1254,N_1616);
and U2105 (N_2105,N_1795,N_1406);
nand U2106 (N_2106,N_1336,N_1279);
or U2107 (N_2107,N_1464,N_1503);
and U2108 (N_2108,N_1202,N_1221);
nor U2109 (N_2109,N_1250,N_1490);
nor U2110 (N_2110,N_1480,N_1608);
nor U2111 (N_2111,N_1785,N_1580);
xnor U2112 (N_2112,N_1390,N_1525);
nor U2113 (N_2113,N_1247,N_1296);
nor U2114 (N_2114,N_1214,N_1209);
xnor U2115 (N_2115,N_1296,N_1710);
and U2116 (N_2116,N_1727,N_1450);
nand U2117 (N_2117,N_1578,N_1419);
nand U2118 (N_2118,N_1222,N_1566);
and U2119 (N_2119,N_1343,N_1324);
and U2120 (N_2120,N_1712,N_1538);
or U2121 (N_2121,N_1702,N_1466);
nor U2122 (N_2122,N_1431,N_1511);
or U2123 (N_2123,N_1484,N_1637);
or U2124 (N_2124,N_1448,N_1451);
nor U2125 (N_2125,N_1364,N_1460);
and U2126 (N_2126,N_1502,N_1742);
nand U2127 (N_2127,N_1435,N_1207);
or U2128 (N_2128,N_1567,N_1325);
or U2129 (N_2129,N_1427,N_1685);
nand U2130 (N_2130,N_1221,N_1542);
nor U2131 (N_2131,N_1435,N_1487);
nor U2132 (N_2132,N_1248,N_1561);
and U2133 (N_2133,N_1449,N_1498);
or U2134 (N_2134,N_1772,N_1316);
or U2135 (N_2135,N_1361,N_1553);
or U2136 (N_2136,N_1380,N_1517);
nand U2137 (N_2137,N_1790,N_1379);
or U2138 (N_2138,N_1210,N_1430);
nand U2139 (N_2139,N_1340,N_1575);
nand U2140 (N_2140,N_1498,N_1595);
nor U2141 (N_2141,N_1549,N_1416);
nand U2142 (N_2142,N_1596,N_1480);
nand U2143 (N_2143,N_1228,N_1363);
nand U2144 (N_2144,N_1542,N_1734);
and U2145 (N_2145,N_1339,N_1207);
and U2146 (N_2146,N_1735,N_1554);
or U2147 (N_2147,N_1466,N_1242);
nor U2148 (N_2148,N_1633,N_1373);
nor U2149 (N_2149,N_1444,N_1433);
xor U2150 (N_2150,N_1240,N_1530);
nor U2151 (N_2151,N_1366,N_1783);
and U2152 (N_2152,N_1552,N_1507);
nand U2153 (N_2153,N_1799,N_1585);
nand U2154 (N_2154,N_1490,N_1508);
or U2155 (N_2155,N_1603,N_1512);
or U2156 (N_2156,N_1441,N_1685);
or U2157 (N_2157,N_1776,N_1638);
nor U2158 (N_2158,N_1724,N_1208);
xnor U2159 (N_2159,N_1513,N_1659);
xnor U2160 (N_2160,N_1593,N_1705);
xnor U2161 (N_2161,N_1645,N_1219);
or U2162 (N_2162,N_1413,N_1489);
xnor U2163 (N_2163,N_1346,N_1623);
nor U2164 (N_2164,N_1732,N_1420);
or U2165 (N_2165,N_1384,N_1226);
or U2166 (N_2166,N_1521,N_1447);
or U2167 (N_2167,N_1238,N_1594);
nor U2168 (N_2168,N_1338,N_1629);
and U2169 (N_2169,N_1736,N_1205);
or U2170 (N_2170,N_1503,N_1637);
nand U2171 (N_2171,N_1437,N_1625);
or U2172 (N_2172,N_1268,N_1688);
nor U2173 (N_2173,N_1445,N_1523);
or U2174 (N_2174,N_1603,N_1631);
or U2175 (N_2175,N_1288,N_1382);
and U2176 (N_2176,N_1282,N_1372);
and U2177 (N_2177,N_1789,N_1406);
or U2178 (N_2178,N_1422,N_1660);
nor U2179 (N_2179,N_1356,N_1487);
or U2180 (N_2180,N_1341,N_1289);
nand U2181 (N_2181,N_1733,N_1414);
and U2182 (N_2182,N_1769,N_1294);
and U2183 (N_2183,N_1626,N_1302);
and U2184 (N_2184,N_1237,N_1223);
nand U2185 (N_2185,N_1238,N_1525);
xnor U2186 (N_2186,N_1303,N_1427);
xnor U2187 (N_2187,N_1706,N_1227);
or U2188 (N_2188,N_1666,N_1251);
and U2189 (N_2189,N_1497,N_1376);
and U2190 (N_2190,N_1597,N_1484);
and U2191 (N_2191,N_1424,N_1248);
or U2192 (N_2192,N_1624,N_1616);
nand U2193 (N_2193,N_1608,N_1536);
nand U2194 (N_2194,N_1350,N_1225);
and U2195 (N_2195,N_1283,N_1453);
and U2196 (N_2196,N_1751,N_1682);
or U2197 (N_2197,N_1791,N_1636);
nor U2198 (N_2198,N_1798,N_1341);
nand U2199 (N_2199,N_1494,N_1653);
nand U2200 (N_2200,N_1602,N_1643);
or U2201 (N_2201,N_1263,N_1526);
nand U2202 (N_2202,N_1287,N_1260);
and U2203 (N_2203,N_1737,N_1418);
or U2204 (N_2204,N_1611,N_1433);
or U2205 (N_2205,N_1402,N_1569);
nand U2206 (N_2206,N_1349,N_1646);
nand U2207 (N_2207,N_1577,N_1456);
nand U2208 (N_2208,N_1393,N_1684);
or U2209 (N_2209,N_1433,N_1457);
or U2210 (N_2210,N_1429,N_1784);
or U2211 (N_2211,N_1572,N_1384);
xnor U2212 (N_2212,N_1691,N_1291);
or U2213 (N_2213,N_1561,N_1210);
nor U2214 (N_2214,N_1629,N_1217);
xor U2215 (N_2215,N_1555,N_1725);
nand U2216 (N_2216,N_1220,N_1522);
and U2217 (N_2217,N_1785,N_1730);
nand U2218 (N_2218,N_1446,N_1337);
nor U2219 (N_2219,N_1761,N_1646);
nand U2220 (N_2220,N_1759,N_1543);
xor U2221 (N_2221,N_1726,N_1350);
or U2222 (N_2222,N_1295,N_1793);
and U2223 (N_2223,N_1449,N_1331);
nand U2224 (N_2224,N_1422,N_1626);
or U2225 (N_2225,N_1272,N_1519);
and U2226 (N_2226,N_1281,N_1650);
nor U2227 (N_2227,N_1592,N_1679);
and U2228 (N_2228,N_1276,N_1342);
nor U2229 (N_2229,N_1395,N_1202);
and U2230 (N_2230,N_1502,N_1721);
nand U2231 (N_2231,N_1466,N_1344);
and U2232 (N_2232,N_1341,N_1469);
nand U2233 (N_2233,N_1207,N_1790);
or U2234 (N_2234,N_1641,N_1617);
xor U2235 (N_2235,N_1732,N_1440);
and U2236 (N_2236,N_1247,N_1311);
nor U2237 (N_2237,N_1350,N_1596);
and U2238 (N_2238,N_1655,N_1789);
nand U2239 (N_2239,N_1456,N_1563);
nand U2240 (N_2240,N_1657,N_1697);
or U2241 (N_2241,N_1701,N_1585);
nor U2242 (N_2242,N_1409,N_1627);
or U2243 (N_2243,N_1766,N_1389);
nand U2244 (N_2244,N_1240,N_1581);
and U2245 (N_2245,N_1627,N_1614);
xnor U2246 (N_2246,N_1646,N_1492);
or U2247 (N_2247,N_1727,N_1222);
nand U2248 (N_2248,N_1295,N_1527);
nand U2249 (N_2249,N_1736,N_1320);
nor U2250 (N_2250,N_1660,N_1333);
or U2251 (N_2251,N_1786,N_1730);
and U2252 (N_2252,N_1782,N_1743);
nor U2253 (N_2253,N_1494,N_1489);
or U2254 (N_2254,N_1297,N_1631);
nand U2255 (N_2255,N_1651,N_1760);
nand U2256 (N_2256,N_1403,N_1488);
or U2257 (N_2257,N_1234,N_1346);
and U2258 (N_2258,N_1693,N_1323);
or U2259 (N_2259,N_1435,N_1530);
and U2260 (N_2260,N_1273,N_1227);
or U2261 (N_2261,N_1338,N_1609);
nand U2262 (N_2262,N_1427,N_1366);
xor U2263 (N_2263,N_1585,N_1690);
or U2264 (N_2264,N_1201,N_1491);
nor U2265 (N_2265,N_1463,N_1316);
or U2266 (N_2266,N_1391,N_1333);
nand U2267 (N_2267,N_1613,N_1399);
or U2268 (N_2268,N_1789,N_1200);
and U2269 (N_2269,N_1669,N_1722);
nand U2270 (N_2270,N_1680,N_1759);
nand U2271 (N_2271,N_1555,N_1674);
nand U2272 (N_2272,N_1216,N_1642);
and U2273 (N_2273,N_1424,N_1745);
and U2274 (N_2274,N_1349,N_1565);
nor U2275 (N_2275,N_1500,N_1428);
nand U2276 (N_2276,N_1681,N_1298);
nand U2277 (N_2277,N_1368,N_1779);
or U2278 (N_2278,N_1346,N_1611);
and U2279 (N_2279,N_1682,N_1518);
and U2280 (N_2280,N_1782,N_1359);
or U2281 (N_2281,N_1567,N_1357);
and U2282 (N_2282,N_1346,N_1730);
nor U2283 (N_2283,N_1203,N_1376);
nand U2284 (N_2284,N_1498,N_1270);
xnor U2285 (N_2285,N_1760,N_1347);
xnor U2286 (N_2286,N_1471,N_1435);
and U2287 (N_2287,N_1312,N_1275);
nand U2288 (N_2288,N_1751,N_1309);
xor U2289 (N_2289,N_1776,N_1262);
nor U2290 (N_2290,N_1608,N_1760);
nand U2291 (N_2291,N_1658,N_1700);
and U2292 (N_2292,N_1287,N_1584);
xnor U2293 (N_2293,N_1242,N_1430);
and U2294 (N_2294,N_1722,N_1354);
xor U2295 (N_2295,N_1266,N_1462);
or U2296 (N_2296,N_1340,N_1516);
nand U2297 (N_2297,N_1742,N_1414);
nand U2298 (N_2298,N_1274,N_1642);
or U2299 (N_2299,N_1324,N_1617);
and U2300 (N_2300,N_1637,N_1698);
and U2301 (N_2301,N_1436,N_1768);
nand U2302 (N_2302,N_1764,N_1327);
nand U2303 (N_2303,N_1643,N_1736);
and U2304 (N_2304,N_1475,N_1557);
and U2305 (N_2305,N_1459,N_1700);
and U2306 (N_2306,N_1470,N_1503);
and U2307 (N_2307,N_1593,N_1432);
or U2308 (N_2308,N_1243,N_1618);
nor U2309 (N_2309,N_1368,N_1294);
nor U2310 (N_2310,N_1640,N_1716);
nor U2311 (N_2311,N_1385,N_1377);
or U2312 (N_2312,N_1362,N_1434);
nand U2313 (N_2313,N_1525,N_1728);
and U2314 (N_2314,N_1734,N_1599);
nor U2315 (N_2315,N_1418,N_1547);
xnor U2316 (N_2316,N_1278,N_1302);
and U2317 (N_2317,N_1565,N_1304);
nand U2318 (N_2318,N_1680,N_1219);
and U2319 (N_2319,N_1493,N_1520);
nor U2320 (N_2320,N_1614,N_1733);
and U2321 (N_2321,N_1284,N_1497);
nand U2322 (N_2322,N_1310,N_1296);
nor U2323 (N_2323,N_1354,N_1353);
nand U2324 (N_2324,N_1346,N_1443);
and U2325 (N_2325,N_1298,N_1307);
nor U2326 (N_2326,N_1555,N_1475);
nor U2327 (N_2327,N_1492,N_1756);
nand U2328 (N_2328,N_1637,N_1278);
nor U2329 (N_2329,N_1349,N_1428);
and U2330 (N_2330,N_1357,N_1506);
and U2331 (N_2331,N_1406,N_1386);
nand U2332 (N_2332,N_1237,N_1468);
or U2333 (N_2333,N_1524,N_1757);
or U2334 (N_2334,N_1590,N_1440);
nor U2335 (N_2335,N_1432,N_1761);
or U2336 (N_2336,N_1204,N_1705);
or U2337 (N_2337,N_1506,N_1424);
nor U2338 (N_2338,N_1467,N_1365);
xor U2339 (N_2339,N_1691,N_1536);
or U2340 (N_2340,N_1446,N_1758);
and U2341 (N_2341,N_1752,N_1368);
nand U2342 (N_2342,N_1592,N_1307);
and U2343 (N_2343,N_1241,N_1293);
xnor U2344 (N_2344,N_1277,N_1771);
nand U2345 (N_2345,N_1263,N_1376);
nand U2346 (N_2346,N_1256,N_1426);
and U2347 (N_2347,N_1490,N_1383);
nand U2348 (N_2348,N_1669,N_1791);
or U2349 (N_2349,N_1698,N_1216);
nand U2350 (N_2350,N_1470,N_1350);
and U2351 (N_2351,N_1732,N_1613);
or U2352 (N_2352,N_1482,N_1704);
xor U2353 (N_2353,N_1686,N_1350);
nand U2354 (N_2354,N_1448,N_1701);
or U2355 (N_2355,N_1353,N_1466);
or U2356 (N_2356,N_1782,N_1209);
nor U2357 (N_2357,N_1577,N_1278);
nor U2358 (N_2358,N_1422,N_1719);
nand U2359 (N_2359,N_1552,N_1600);
and U2360 (N_2360,N_1490,N_1225);
nor U2361 (N_2361,N_1370,N_1279);
nand U2362 (N_2362,N_1526,N_1460);
or U2363 (N_2363,N_1783,N_1724);
and U2364 (N_2364,N_1703,N_1255);
nand U2365 (N_2365,N_1753,N_1244);
nor U2366 (N_2366,N_1552,N_1484);
and U2367 (N_2367,N_1677,N_1548);
and U2368 (N_2368,N_1418,N_1666);
nor U2369 (N_2369,N_1499,N_1377);
or U2370 (N_2370,N_1722,N_1283);
or U2371 (N_2371,N_1316,N_1599);
nor U2372 (N_2372,N_1668,N_1749);
nand U2373 (N_2373,N_1646,N_1760);
nand U2374 (N_2374,N_1287,N_1606);
nor U2375 (N_2375,N_1265,N_1611);
or U2376 (N_2376,N_1786,N_1397);
and U2377 (N_2377,N_1628,N_1570);
and U2378 (N_2378,N_1692,N_1760);
nand U2379 (N_2379,N_1279,N_1377);
nor U2380 (N_2380,N_1537,N_1612);
xnor U2381 (N_2381,N_1404,N_1455);
nor U2382 (N_2382,N_1435,N_1359);
or U2383 (N_2383,N_1231,N_1296);
nor U2384 (N_2384,N_1361,N_1694);
nand U2385 (N_2385,N_1420,N_1210);
and U2386 (N_2386,N_1602,N_1775);
and U2387 (N_2387,N_1206,N_1327);
and U2388 (N_2388,N_1685,N_1265);
and U2389 (N_2389,N_1544,N_1268);
nand U2390 (N_2390,N_1476,N_1520);
nor U2391 (N_2391,N_1515,N_1499);
nand U2392 (N_2392,N_1302,N_1730);
or U2393 (N_2393,N_1236,N_1246);
nand U2394 (N_2394,N_1587,N_1685);
or U2395 (N_2395,N_1360,N_1741);
nor U2396 (N_2396,N_1790,N_1430);
and U2397 (N_2397,N_1379,N_1301);
nor U2398 (N_2398,N_1410,N_1433);
nand U2399 (N_2399,N_1660,N_1744);
and U2400 (N_2400,N_2331,N_2086);
xnor U2401 (N_2401,N_1808,N_2182);
nand U2402 (N_2402,N_1861,N_1908);
or U2403 (N_2403,N_2342,N_2002);
and U2404 (N_2404,N_1859,N_2313);
or U2405 (N_2405,N_2205,N_2030);
nor U2406 (N_2406,N_1932,N_2322);
nand U2407 (N_2407,N_1970,N_2260);
or U2408 (N_2408,N_2284,N_2223);
or U2409 (N_2409,N_2257,N_2363);
nand U2410 (N_2410,N_2184,N_2158);
nand U2411 (N_2411,N_2384,N_1941);
and U2412 (N_2412,N_1813,N_2147);
nand U2413 (N_2413,N_2349,N_2041);
or U2414 (N_2414,N_2169,N_2089);
or U2415 (N_2415,N_1802,N_2385);
or U2416 (N_2416,N_2154,N_2202);
nor U2417 (N_2417,N_1816,N_2161);
nand U2418 (N_2418,N_2321,N_1979);
nand U2419 (N_2419,N_2148,N_2338);
or U2420 (N_2420,N_1824,N_2017);
xnor U2421 (N_2421,N_1819,N_2370);
and U2422 (N_2422,N_2368,N_2299);
xnor U2423 (N_2423,N_1820,N_1878);
nand U2424 (N_2424,N_2249,N_2059);
nor U2425 (N_2425,N_2198,N_2176);
or U2426 (N_2426,N_2143,N_1942);
nor U2427 (N_2427,N_1851,N_2054);
nor U2428 (N_2428,N_1991,N_2354);
or U2429 (N_2429,N_1966,N_2206);
nand U2430 (N_2430,N_2092,N_1906);
or U2431 (N_2431,N_2314,N_2194);
nand U2432 (N_2432,N_1886,N_2173);
xor U2433 (N_2433,N_2282,N_2027);
xor U2434 (N_2434,N_1863,N_2247);
nand U2435 (N_2435,N_2311,N_2172);
nand U2436 (N_2436,N_2138,N_2300);
or U2437 (N_2437,N_1955,N_2372);
and U2438 (N_2438,N_2040,N_2269);
and U2439 (N_2439,N_2333,N_2026);
nand U2440 (N_2440,N_2188,N_2357);
nand U2441 (N_2441,N_1968,N_2035);
nor U2442 (N_2442,N_2341,N_2273);
nand U2443 (N_2443,N_2375,N_1917);
xor U2444 (N_2444,N_2265,N_2034);
and U2445 (N_2445,N_1843,N_2048);
nand U2446 (N_2446,N_2076,N_2068);
xor U2447 (N_2447,N_2009,N_1946);
nand U2448 (N_2448,N_2344,N_2125);
nor U2449 (N_2449,N_2355,N_2168);
or U2450 (N_2450,N_1922,N_2061);
and U2451 (N_2451,N_2398,N_1831);
nor U2452 (N_2452,N_2371,N_1903);
nor U2453 (N_2453,N_2107,N_1912);
or U2454 (N_2454,N_2013,N_1953);
and U2455 (N_2455,N_1977,N_1956);
or U2456 (N_2456,N_2327,N_1855);
nor U2457 (N_2457,N_1948,N_2139);
nor U2458 (N_2458,N_2256,N_1943);
nor U2459 (N_2459,N_2129,N_1891);
or U2460 (N_2460,N_2049,N_2011);
nor U2461 (N_2461,N_2018,N_2022);
nand U2462 (N_2462,N_1918,N_1865);
nand U2463 (N_2463,N_1880,N_2216);
nor U2464 (N_2464,N_2160,N_1974);
nand U2465 (N_2465,N_2175,N_2364);
nand U2466 (N_2466,N_2329,N_1998);
or U2467 (N_2467,N_2144,N_2225);
nor U2468 (N_2468,N_2283,N_2328);
and U2469 (N_2469,N_2276,N_2133);
and U2470 (N_2470,N_2196,N_2171);
xnor U2471 (N_2471,N_2153,N_1875);
nand U2472 (N_2472,N_2047,N_1829);
and U2473 (N_2473,N_1987,N_2072);
nand U2474 (N_2474,N_2248,N_2134);
and U2475 (N_2475,N_2152,N_2023);
or U2476 (N_2476,N_2395,N_1884);
and U2477 (N_2477,N_2108,N_2219);
or U2478 (N_2478,N_1925,N_1952);
and U2479 (N_2479,N_1934,N_1930);
nor U2480 (N_2480,N_2399,N_2008);
nor U2481 (N_2481,N_1904,N_1945);
and U2482 (N_2482,N_2119,N_2050);
nor U2483 (N_2483,N_1872,N_1835);
nor U2484 (N_2484,N_1993,N_2156);
xnor U2485 (N_2485,N_1984,N_1821);
nand U2486 (N_2486,N_1972,N_1990);
nand U2487 (N_2487,N_1992,N_2251);
and U2488 (N_2488,N_1848,N_2287);
and U2489 (N_2489,N_2288,N_2252);
nand U2490 (N_2490,N_2010,N_1804);
nand U2491 (N_2491,N_2359,N_2127);
nor U2492 (N_2492,N_2187,N_2128);
nand U2493 (N_2493,N_1857,N_2246);
xnor U2494 (N_2494,N_1837,N_1926);
and U2495 (N_2495,N_2084,N_2155);
nor U2496 (N_2496,N_1827,N_2056);
nor U2497 (N_2497,N_1988,N_2376);
nor U2498 (N_2498,N_2209,N_1995);
nor U2499 (N_2499,N_1898,N_2224);
xnor U2500 (N_2500,N_1889,N_2241);
or U2501 (N_2501,N_1919,N_2039);
xnor U2502 (N_2502,N_2220,N_2306);
nand U2503 (N_2503,N_2304,N_2240);
or U2504 (N_2504,N_2296,N_2393);
nor U2505 (N_2505,N_2270,N_2191);
xor U2506 (N_2506,N_1931,N_2290);
and U2507 (N_2507,N_1860,N_2316);
nor U2508 (N_2508,N_2294,N_2177);
or U2509 (N_2509,N_1928,N_2394);
nor U2510 (N_2510,N_2100,N_2070);
nor U2511 (N_2511,N_2345,N_2146);
xnor U2512 (N_2512,N_2232,N_1879);
nand U2513 (N_2513,N_2318,N_1964);
or U2514 (N_2514,N_2007,N_2149);
and U2515 (N_2515,N_1856,N_2014);
nor U2516 (N_2516,N_2136,N_2083);
and U2517 (N_2517,N_2235,N_2045);
nor U2518 (N_2518,N_2163,N_1805);
nand U2519 (N_2519,N_2062,N_1978);
and U2520 (N_2520,N_2382,N_1899);
and U2521 (N_2521,N_2190,N_1940);
or U2522 (N_2522,N_2337,N_2087);
nand U2523 (N_2523,N_2279,N_2101);
or U2524 (N_2524,N_2043,N_1938);
nand U2525 (N_2525,N_2356,N_2378);
nor U2526 (N_2526,N_1849,N_2347);
xnor U2527 (N_2527,N_1997,N_2025);
nor U2528 (N_2528,N_1927,N_1885);
xor U2529 (N_2529,N_2332,N_2093);
and U2530 (N_2530,N_2082,N_1989);
xnor U2531 (N_2531,N_1803,N_2080);
nand U2532 (N_2532,N_2366,N_2051);
nor U2533 (N_2533,N_2267,N_2373);
nand U2534 (N_2534,N_2113,N_1913);
nand U2535 (N_2535,N_2317,N_2073);
and U2536 (N_2536,N_2174,N_2181);
nor U2537 (N_2537,N_2186,N_2286);
nand U2538 (N_2538,N_2250,N_2320);
and U2539 (N_2539,N_2280,N_1905);
nand U2540 (N_2540,N_1870,N_2262);
or U2541 (N_2541,N_2033,N_1887);
xor U2542 (N_2542,N_1957,N_2388);
nand U2543 (N_2543,N_2391,N_1890);
nor U2544 (N_2544,N_1921,N_1876);
or U2545 (N_2545,N_2052,N_1975);
nor U2546 (N_2546,N_2104,N_1915);
nor U2547 (N_2547,N_2380,N_1840);
nand U2548 (N_2548,N_1902,N_2389);
nor U2549 (N_2549,N_2165,N_1935);
nor U2550 (N_2550,N_2397,N_1959);
xor U2551 (N_2551,N_1949,N_2263);
nor U2552 (N_2552,N_2227,N_2211);
nor U2553 (N_2553,N_2324,N_2374);
and U2554 (N_2554,N_1900,N_2095);
nand U2555 (N_2555,N_2193,N_2301);
nor U2556 (N_2556,N_2367,N_2180);
nand U2557 (N_2557,N_2110,N_2244);
and U2558 (N_2558,N_2131,N_1853);
nand U2559 (N_2559,N_2264,N_2336);
nand U2560 (N_2560,N_1967,N_2325);
nor U2561 (N_2561,N_2308,N_2207);
nand U2562 (N_2562,N_2255,N_2360);
and U2563 (N_2563,N_2330,N_1960);
or U2564 (N_2564,N_2189,N_2123);
or U2565 (N_2565,N_2310,N_2124);
nand U2566 (N_2566,N_2001,N_2326);
nor U2567 (N_2567,N_1866,N_2126);
xor U2568 (N_2568,N_2044,N_2141);
and U2569 (N_2569,N_1888,N_1814);
nand U2570 (N_2570,N_1937,N_2114);
nor U2571 (N_2571,N_2038,N_2130);
nor U2572 (N_2572,N_1973,N_2243);
and U2573 (N_2573,N_2096,N_2005);
xnor U2574 (N_2574,N_2230,N_1982);
nor U2575 (N_2575,N_1976,N_1910);
or U2576 (N_2576,N_2396,N_2069);
and U2577 (N_2577,N_2334,N_2120);
nand U2578 (N_2578,N_1999,N_2361);
and U2579 (N_2579,N_1936,N_2315);
and U2580 (N_2580,N_2004,N_2066);
nand U2581 (N_2581,N_2166,N_2271);
xor U2582 (N_2582,N_2132,N_2097);
nand U2583 (N_2583,N_1929,N_1845);
and U2584 (N_2584,N_2067,N_2032);
nor U2585 (N_2585,N_2098,N_2075);
xnor U2586 (N_2586,N_2064,N_1841);
or U2587 (N_2587,N_1939,N_1996);
nor U2588 (N_2588,N_2297,N_1817);
nor U2589 (N_2589,N_1895,N_1969);
nor U2590 (N_2590,N_2215,N_1911);
or U2591 (N_2591,N_2142,N_2293);
nand U2592 (N_2592,N_2029,N_2183);
nand U2593 (N_2593,N_2305,N_1844);
nand U2594 (N_2594,N_2003,N_1815);
nor U2595 (N_2595,N_1826,N_2091);
and U2596 (N_2596,N_2353,N_1862);
or U2597 (N_2597,N_2278,N_2150);
and U2598 (N_2598,N_1812,N_2238);
and U2599 (N_2599,N_2145,N_1801);
nand U2600 (N_2600,N_2259,N_1954);
nand U2601 (N_2601,N_2383,N_1830);
nor U2602 (N_2602,N_2339,N_2377);
nor U2603 (N_2603,N_2140,N_1950);
nand U2604 (N_2604,N_1892,N_2058);
and U2605 (N_2605,N_2028,N_1947);
nand U2606 (N_2606,N_2115,N_2019);
or U2607 (N_2607,N_1981,N_2106);
nor U2608 (N_2608,N_1916,N_2277);
and U2609 (N_2609,N_2178,N_2006);
nand U2610 (N_2610,N_1962,N_1896);
nor U2611 (N_2611,N_2112,N_2036);
nand U2612 (N_2612,N_2077,N_1807);
and U2613 (N_2613,N_2214,N_2135);
or U2614 (N_2614,N_1924,N_1822);
nor U2615 (N_2615,N_1832,N_2222);
or U2616 (N_2616,N_2351,N_2392);
or U2617 (N_2617,N_2057,N_2102);
nand U2618 (N_2618,N_2151,N_1834);
nand U2619 (N_2619,N_2268,N_1825);
nor U2620 (N_2620,N_2016,N_2309);
or U2621 (N_2621,N_1828,N_2281);
and U2622 (N_2622,N_1958,N_2063);
nor U2623 (N_2623,N_1980,N_2233);
nor U2624 (N_2624,N_1985,N_1839);
nor U2625 (N_2625,N_2218,N_2167);
or U2626 (N_2626,N_2362,N_2352);
nor U2627 (N_2627,N_2234,N_1811);
nand U2628 (N_2628,N_2099,N_1933);
nand U2629 (N_2629,N_2292,N_2346);
and U2630 (N_2630,N_1800,N_1854);
and U2631 (N_2631,N_2226,N_2229);
and U2632 (N_2632,N_2319,N_2195);
nor U2633 (N_2633,N_2302,N_1914);
nor U2634 (N_2634,N_2253,N_2053);
and U2635 (N_2635,N_1838,N_1818);
nand U2636 (N_2636,N_1850,N_1858);
and U2637 (N_2637,N_2021,N_1971);
or U2638 (N_2638,N_1809,N_1868);
nor U2639 (N_2639,N_1994,N_2254);
nand U2640 (N_2640,N_1907,N_2024);
or U2641 (N_2641,N_2242,N_1944);
nand U2642 (N_2642,N_2046,N_2261);
nand U2643 (N_2643,N_2210,N_2291);
or U2644 (N_2644,N_2071,N_2387);
nand U2645 (N_2645,N_2236,N_2031);
or U2646 (N_2646,N_2085,N_2090);
or U2647 (N_2647,N_2111,N_1836);
nor U2648 (N_2648,N_2258,N_2343);
or U2649 (N_2649,N_2078,N_2312);
or U2650 (N_2650,N_2159,N_2212);
nor U2651 (N_2651,N_1986,N_1810);
nor U2652 (N_2652,N_2358,N_1873);
and U2653 (N_2653,N_1961,N_2221);
nor U2654 (N_2654,N_2170,N_2369);
and U2655 (N_2655,N_2162,N_2199);
or U2656 (N_2656,N_2272,N_1901);
or U2657 (N_2657,N_2065,N_1923);
nand U2658 (N_2658,N_1909,N_1833);
and U2659 (N_2659,N_2094,N_1823);
nand U2660 (N_2660,N_2074,N_2060);
or U2661 (N_2661,N_2266,N_1893);
or U2662 (N_2662,N_2335,N_2379);
and U2663 (N_2663,N_2118,N_2012);
xnor U2664 (N_2664,N_2323,N_1864);
nor U2665 (N_2665,N_2348,N_1874);
and U2666 (N_2666,N_2185,N_2307);
or U2667 (N_2667,N_2037,N_2122);
and U2668 (N_2668,N_2350,N_2340);
or U2669 (N_2669,N_2245,N_2192);
or U2670 (N_2670,N_2117,N_2295);
and U2671 (N_2671,N_2116,N_2105);
and U2672 (N_2672,N_1882,N_2081);
nor U2673 (N_2673,N_2239,N_1894);
and U2674 (N_2674,N_2217,N_1869);
or U2675 (N_2675,N_1951,N_2103);
and U2676 (N_2676,N_2088,N_1867);
nand U2677 (N_2677,N_2390,N_1883);
nor U2678 (N_2678,N_2231,N_2386);
xnor U2679 (N_2679,N_2079,N_2179);
and U2680 (N_2680,N_2137,N_1920);
xnor U2681 (N_2681,N_2200,N_1877);
and U2682 (N_2682,N_2365,N_2197);
xnor U2683 (N_2683,N_2208,N_1847);
nand U2684 (N_2684,N_2015,N_2289);
or U2685 (N_2685,N_1897,N_1983);
nor U2686 (N_2686,N_1963,N_2164);
nor U2687 (N_2687,N_2228,N_1842);
and U2688 (N_2688,N_1965,N_2109);
nand U2689 (N_2689,N_2275,N_2020);
or U2690 (N_2690,N_1846,N_2237);
nor U2691 (N_2691,N_2055,N_2381);
and U2692 (N_2692,N_2121,N_2203);
nor U2693 (N_2693,N_2204,N_2285);
and U2694 (N_2694,N_1871,N_2303);
or U2695 (N_2695,N_2201,N_1852);
and U2696 (N_2696,N_2042,N_2298);
nand U2697 (N_2697,N_1881,N_1806);
xor U2698 (N_2698,N_2157,N_2274);
or U2699 (N_2699,N_2213,N_2000);
xnor U2700 (N_2700,N_2289,N_2293);
and U2701 (N_2701,N_2304,N_1968);
nor U2702 (N_2702,N_2179,N_1962);
or U2703 (N_2703,N_1845,N_1921);
nand U2704 (N_2704,N_2148,N_2069);
nor U2705 (N_2705,N_2268,N_2020);
nand U2706 (N_2706,N_2368,N_1810);
and U2707 (N_2707,N_1972,N_2341);
nor U2708 (N_2708,N_2095,N_1932);
or U2709 (N_2709,N_2293,N_1873);
and U2710 (N_2710,N_2367,N_2281);
or U2711 (N_2711,N_2093,N_2035);
or U2712 (N_2712,N_1911,N_2288);
and U2713 (N_2713,N_2086,N_2151);
nand U2714 (N_2714,N_2226,N_1971);
or U2715 (N_2715,N_2004,N_2171);
or U2716 (N_2716,N_2309,N_2377);
or U2717 (N_2717,N_2341,N_1811);
and U2718 (N_2718,N_2256,N_1883);
nand U2719 (N_2719,N_1861,N_2023);
and U2720 (N_2720,N_2125,N_2023);
and U2721 (N_2721,N_2393,N_2225);
or U2722 (N_2722,N_1827,N_2397);
xnor U2723 (N_2723,N_2224,N_2296);
nand U2724 (N_2724,N_2209,N_1992);
nor U2725 (N_2725,N_2113,N_1829);
and U2726 (N_2726,N_1936,N_2318);
and U2727 (N_2727,N_2033,N_2041);
or U2728 (N_2728,N_2130,N_1914);
nand U2729 (N_2729,N_2170,N_2143);
nand U2730 (N_2730,N_2119,N_2279);
and U2731 (N_2731,N_1965,N_2296);
nand U2732 (N_2732,N_2338,N_1919);
or U2733 (N_2733,N_1906,N_2201);
nor U2734 (N_2734,N_1850,N_2065);
nor U2735 (N_2735,N_1840,N_2304);
and U2736 (N_2736,N_1939,N_2093);
xnor U2737 (N_2737,N_1997,N_2218);
or U2738 (N_2738,N_1866,N_2286);
nand U2739 (N_2739,N_1966,N_2260);
nand U2740 (N_2740,N_2034,N_1970);
nand U2741 (N_2741,N_1823,N_1936);
xnor U2742 (N_2742,N_2086,N_1915);
and U2743 (N_2743,N_2250,N_2032);
nor U2744 (N_2744,N_1973,N_1823);
nor U2745 (N_2745,N_2102,N_1827);
nand U2746 (N_2746,N_2067,N_2106);
nand U2747 (N_2747,N_2005,N_2215);
xor U2748 (N_2748,N_2128,N_2367);
nor U2749 (N_2749,N_1972,N_2316);
nand U2750 (N_2750,N_2179,N_2310);
xnor U2751 (N_2751,N_2377,N_2316);
nor U2752 (N_2752,N_2198,N_2394);
or U2753 (N_2753,N_2136,N_1907);
or U2754 (N_2754,N_1936,N_2035);
or U2755 (N_2755,N_2084,N_2123);
or U2756 (N_2756,N_1995,N_1844);
xnor U2757 (N_2757,N_1959,N_2209);
xnor U2758 (N_2758,N_2168,N_2315);
and U2759 (N_2759,N_2374,N_2098);
or U2760 (N_2760,N_2247,N_2004);
and U2761 (N_2761,N_2020,N_1961);
or U2762 (N_2762,N_1846,N_2014);
or U2763 (N_2763,N_2163,N_2066);
nor U2764 (N_2764,N_1984,N_1805);
nand U2765 (N_2765,N_2227,N_1949);
nand U2766 (N_2766,N_1838,N_2210);
or U2767 (N_2767,N_2105,N_2084);
nand U2768 (N_2768,N_1829,N_1962);
or U2769 (N_2769,N_2222,N_1900);
nand U2770 (N_2770,N_2213,N_1951);
nand U2771 (N_2771,N_2373,N_2244);
and U2772 (N_2772,N_2217,N_1848);
xnor U2773 (N_2773,N_2288,N_1830);
and U2774 (N_2774,N_2231,N_2168);
nor U2775 (N_2775,N_2272,N_1812);
and U2776 (N_2776,N_2297,N_1957);
and U2777 (N_2777,N_2115,N_1876);
and U2778 (N_2778,N_2153,N_1994);
nand U2779 (N_2779,N_2078,N_2153);
or U2780 (N_2780,N_1940,N_1982);
and U2781 (N_2781,N_2296,N_2109);
and U2782 (N_2782,N_1851,N_1811);
xnor U2783 (N_2783,N_2389,N_2008);
or U2784 (N_2784,N_1981,N_2380);
and U2785 (N_2785,N_1810,N_1895);
nand U2786 (N_2786,N_1816,N_2212);
or U2787 (N_2787,N_1871,N_2023);
nand U2788 (N_2788,N_2036,N_2028);
xor U2789 (N_2789,N_1812,N_2046);
nand U2790 (N_2790,N_2006,N_2287);
nor U2791 (N_2791,N_2352,N_1955);
nand U2792 (N_2792,N_2005,N_2253);
nor U2793 (N_2793,N_2156,N_2187);
and U2794 (N_2794,N_1863,N_1983);
nand U2795 (N_2795,N_1976,N_2277);
and U2796 (N_2796,N_2288,N_2381);
xor U2797 (N_2797,N_2057,N_1999);
or U2798 (N_2798,N_2006,N_1864);
or U2799 (N_2799,N_2103,N_2169);
nor U2800 (N_2800,N_2124,N_2009);
and U2801 (N_2801,N_1929,N_2277);
nor U2802 (N_2802,N_1844,N_2112);
nor U2803 (N_2803,N_2108,N_2012);
or U2804 (N_2804,N_1843,N_2319);
and U2805 (N_2805,N_1895,N_1828);
or U2806 (N_2806,N_1940,N_1952);
nand U2807 (N_2807,N_1812,N_1811);
nand U2808 (N_2808,N_2191,N_1941);
and U2809 (N_2809,N_2064,N_2140);
and U2810 (N_2810,N_1938,N_1954);
or U2811 (N_2811,N_2068,N_2242);
or U2812 (N_2812,N_2269,N_2166);
and U2813 (N_2813,N_2326,N_2382);
xnor U2814 (N_2814,N_2227,N_1825);
nor U2815 (N_2815,N_2291,N_2072);
nor U2816 (N_2816,N_2175,N_2207);
or U2817 (N_2817,N_2130,N_2092);
xor U2818 (N_2818,N_2233,N_2136);
nor U2819 (N_2819,N_2238,N_1975);
nand U2820 (N_2820,N_2366,N_2329);
or U2821 (N_2821,N_1914,N_2152);
nor U2822 (N_2822,N_1940,N_1802);
and U2823 (N_2823,N_2214,N_1940);
nand U2824 (N_2824,N_1989,N_1914);
xnor U2825 (N_2825,N_2133,N_1905);
nand U2826 (N_2826,N_2251,N_2183);
nand U2827 (N_2827,N_2068,N_1921);
nor U2828 (N_2828,N_2383,N_2276);
and U2829 (N_2829,N_2240,N_2032);
or U2830 (N_2830,N_2204,N_2329);
nand U2831 (N_2831,N_2179,N_1854);
nor U2832 (N_2832,N_2251,N_1844);
or U2833 (N_2833,N_1833,N_1970);
nor U2834 (N_2834,N_2127,N_2352);
nor U2835 (N_2835,N_1987,N_2368);
nor U2836 (N_2836,N_1848,N_2254);
and U2837 (N_2837,N_1856,N_2210);
and U2838 (N_2838,N_2328,N_1804);
and U2839 (N_2839,N_2390,N_2084);
nand U2840 (N_2840,N_1893,N_1894);
nor U2841 (N_2841,N_2033,N_2038);
and U2842 (N_2842,N_2303,N_1816);
xor U2843 (N_2843,N_2171,N_2024);
nand U2844 (N_2844,N_2021,N_2084);
nand U2845 (N_2845,N_1844,N_2154);
nand U2846 (N_2846,N_2362,N_2148);
nand U2847 (N_2847,N_2387,N_2159);
and U2848 (N_2848,N_1881,N_1939);
nand U2849 (N_2849,N_2349,N_2392);
nand U2850 (N_2850,N_2045,N_2343);
nand U2851 (N_2851,N_1969,N_2066);
xor U2852 (N_2852,N_2371,N_2053);
or U2853 (N_2853,N_1832,N_1934);
and U2854 (N_2854,N_1988,N_1985);
and U2855 (N_2855,N_2054,N_2267);
nand U2856 (N_2856,N_2215,N_1904);
nor U2857 (N_2857,N_2157,N_2287);
or U2858 (N_2858,N_2038,N_2195);
nand U2859 (N_2859,N_2248,N_2269);
nand U2860 (N_2860,N_1991,N_2048);
nand U2861 (N_2861,N_1925,N_2048);
nand U2862 (N_2862,N_2155,N_1889);
or U2863 (N_2863,N_2334,N_2186);
or U2864 (N_2864,N_1871,N_1977);
or U2865 (N_2865,N_2190,N_2320);
and U2866 (N_2866,N_2246,N_1957);
nor U2867 (N_2867,N_2054,N_1889);
nand U2868 (N_2868,N_2164,N_2123);
nor U2869 (N_2869,N_1863,N_1982);
or U2870 (N_2870,N_2360,N_1881);
nand U2871 (N_2871,N_2184,N_2380);
or U2872 (N_2872,N_2126,N_2064);
nor U2873 (N_2873,N_1837,N_2019);
xnor U2874 (N_2874,N_1958,N_2015);
and U2875 (N_2875,N_2349,N_2300);
xnor U2876 (N_2876,N_2095,N_2291);
nand U2877 (N_2877,N_2392,N_1839);
or U2878 (N_2878,N_1936,N_2332);
nor U2879 (N_2879,N_2228,N_2236);
nand U2880 (N_2880,N_2209,N_1899);
and U2881 (N_2881,N_1855,N_1872);
nand U2882 (N_2882,N_2140,N_2366);
and U2883 (N_2883,N_2004,N_1870);
or U2884 (N_2884,N_2215,N_2374);
xor U2885 (N_2885,N_2186,N_2392);
and U2886 (N_2886,N_2376,N_2169);
nor U2887 (N_2887,N_1940,N_2083);
and U2888 (N_2888,N_2078,N_2173);
nor U2889 (N_2889,N_1855,N_1925);
nor U2890 (N_2890,N_2188,N_1889);
nand U2891 (N_2891,N_2327,N_2331);
nor U2892 (N_2892,N_2046,N_1999);
and U2893 (N_2893,N_1812,N_2137);
and U2894 (N_2894,N_2259,N_1810);
and U2895 (N_2895,N_2040,N_2115);
nand U2896 (N_2896,N_1869,N_2131);
and U2897 (N_2897,N_2190,N_2095);
xnor U2898 (N_2898,N_2340,N_2069);
or U2899 (N_2899,N_2351,N_2147);
and U2900 (N_2900,N_2084,N_2167);
nor U2901 (N_2901,N_2353,N_2272);
xor U2902 (N_2902,N_1965,N_2279);
nand U2903 (N_2903,N_2314,N_2255);
xor U2904 (N_2904,N_2380,N_2378);
or U2905 (N_2905,N_1874,N_2105);
or U2906 (N_2906,N_1894,N_2200);
or U2907 (N_2907,N_1925,N_2137);
or U2908 (N_2908,N_2391,N_2314);
nand U2909 (N_2909,N_2385,N_2257);
nand U2910 (N_2910,N_2368,N_2182);
and U2911 (N_2911,N_1943,N_2228);
and U2912 (N_2912,N_2096,N_1927);
or U2913 (N_2913,N_2354,N_2116);
nor U2914 (N_2914,N_2390,N_2232);
nand U2915 (N_2915,N_2046,N_2342);
nor U2916 (N_2916,N_2303,N_2348);
or U2917 (N_2917,N_2240,N_1895);
or U2918 (N_2918,N_2104,N_1811);
or U2919 (N_2919,N_2169,N_2036);
nor U2920 (N_2920,N_1959,N_1867);
nor U2921 (N_2921,N_1947,N_2102);
or U2922 (N_2922,N_2064,N_2322);
nand U2923 (N_2923,N_1845,N_2050);
and U2924 (N_2924,N_2067,N_1952);
nor U2925 (N_2925,N_2062,N_1841);
or U2926 (N_2926,N_2114,N_1928);
xor U2927 (N_2927,N_2236,N_2056);
nand U2928 (N_2928,N_2265,N_1922);
xor U2929 (N_2929,N_2073,N_2057);
or U2930 (N_2930,N_2221,N_2254);
nand U2931 (N_2931,N_1962,N_2284);
nand U2932 (N_2932,N_2375,N_2374);
xnor U2933 (N_2933,N_2215,N_2203);
nor U2934 (N_2934,N_2318,N_2199);
xor U2935 (N_2935,N_2270,N_2398);
nor U2936 (N_2936,N_2225,N_2058);
nor U2937 (N_2937,N_1869,N_2101);
nand U2938 (N_2938,N_1810,N_2107);
or U2939 (N_2939,N_2039,N_2235);
or U2940 (N_2940,N_1804,N_1819);
nand U2941 (N_2941,N_2138,N_1984);
nand U2942 (N_2942,N_2133,N_2216);
nand U2943 (N_2943,N_2027,N_2360);
or U2944 (N_2944,N_2322,N_1944);
or U2945 (N_2945,N_2017,N_2349);
nor U2946 (N_2946,N_2240,N_2390);
or U2947 (N_2947,N_1858,N_1847);
nor U2948 (N_2948,N_1985,N_2149);
or U2949 (N_2949,N_1909,N_2148);
nand U2950 (N_2950,N_2386,N_2353);
nand U2951 (N_2951,N_2125,N_2306);
and U2952 (N_2952,N_1883,N_2007);
xnor U2953 (N_2953,N_1836,N_1871);
nor U2954 (N_2954,N_2225,N_1928);
xnor U2955 (N_2955,N_2164,N_2024);
nor U2956 (N_2956,N_1974,N_2056);
nor U2957 (N_2957,N_1911,N_2228);
xor U2958 (N_2958,N_2056,N_1802);
and U2959 (N_2959,N_1829,N_1948);
or U2960 (N_2960,N_1940,N_1814);
nor U2961 (N_2961,N_2058,N_1860);
xor U2962 (N_2962,N_2232,N_1895);
xnor U2963 (N_2963,N_2272,N_2382);
or U2964 (N_2964,N_1955,N_1973);
xor U2965 (N_2965,N_2343,N_2156);
or U2966 (N_2966,N_1973,N_2327);
and U2967 (N_2967,N_1866,N_1969);
nor U2968 (N_2968,N_2134,N_1926);
xnor U2969 (N_2969,N_2242,N_2395);
and U2970 (N_2970,N_1899,N_1978);
and U2971 (N_2971,N_2220,N_2350);
or U2972 (N_2972,N_2323,N_2266);
or U2973 (N_2973,N_1856,N_2389);
nor U2974 (N_2974,N_1824,N_1921);
xor U2975 (N_2975,N_1861,N_1867);
and U2976 (N_2976,N_2354,N_2388);
xnor U2977 (N_2977,N_2160,N_2056);
nand U2978 (N_2978,N_1853,N_2336);
nand U2979 (N_2979,N_2072,N_1939);
nor U2980 (N_2980,N_1999,N_2259);
nor U2981 (N_2981,N_2036,N_1849);
nand U2982 (N_2982,N_1953,N_2369);
or U2983 (N_2983,N_1965,N_1839);
or U2984 (N_2984,N_2099,N_1878);
nor U2985 (N_2985,N_2039,N_2398);
and U2986 (N_2986,N_2127,N_2390);
nor U2987 (N_2987,N_2312,N_2372);
and U2988 (N_2988,N_2342,N_1815);
nand U2989 (N_2989,N_2014,N_1802);
or U2990 (N_2990,N_2208,N_2399);
or U2991 (N_2991,N_2371,N_2149);
and U2992 (N_2992,N_2206,N_2186);
and U2993 (N_2993,N_2113,N_2004);
nor U2994 (N_2994,N_2045,N_2283);
or U2995 (N_2995,N_2119,N_2331);
nand U2996 (N_2996,N_2223,N_1922);
nand U2997 (N_2997,N_2262,N_1838);
nand U2998 (N_2998,N_1808,N_1815);
or U2999 (N_2999,N_2087,N_2153);
or UO_0 (O_0,N_2703,N_2950);
or UO_1 (O_1,N_2575,N_2569);
nand UO_2 (O_2,N_2800,N_2947);
nand UO_3 (O_3,N_2746,N_2829);
nor UO_4 (O_4,N_2492,N_2914);
and UO_5 (O_5,N_2793,N_2493);
and UO_6 (O_6,N_2514,N_2517);
and UO_7 (O_7,N_2483,N_2423);
or UO_8 (O_8,N_2750,N_2741);
or UO_9 (O_9,N_2721,N_2874);
xor UO_10 (O_10,N_2515,N_2431);
nor UO_11 (O_11,N_2455,N_2811);
nor UO_12 (O_12,N_2581,N_2589);
nor UO_13 (O_13,N_2424,N_2406);
nor UO_14 (O_14,N_2419,N_2474);
nand UO_15 (O_15,N_2597,N_2679);
or UO_16 (O_16,N_2444,N_2845);
or UO_17 (O_17,N_2516,N_2662);
nor UO_18 (O_18,N_2963,N_2499);
and UO_19 (O_19,N_2883,N_2607);
xnor UO_20 (O_20,N_2526,N_2923);
and UO_21 (O_21,N_2549,N_2691);
and UO_22 (O_22,N_2990,N_2673);
or UO_23 (O_23,N_2951,N_2977);
nand UO_24 (O_24,N_2919,N_2877);
nand UO_25 (O_25,N_2468,N_2933);
and UO_26 (O_26,N_2988,N_2508);
or UO_27 (O_27,N_2825,N_2651);
and UO_28 (O_28,N_2677,N_2782);
nand UO_29 (O_29,N_2674,N_2412);
nor UO_30 (O_30,N_2924,N_2435);
or UO_31 (O_31,N_2828,N_2619);
nor UO_32 (O_32,N_2420,N_2823);
or UO_33 (O_33,N_2695,N_2718);
nand UO_34 (O_34,N_2660,N_2880);
or UO_35 (O_35,N_2475,N_2725);
nor UO_36 (O_36,N_2408,N_2458);
nand UO_37 (O_37,N_2798,N_2596);
and UO_38 (O_38,N_2533,N_2872);
or UO_39 (O_39,N_2489,N_2834);
nor UO_40 (O_40,N_2504,N_2649);
or UO_41 (O_41,N_2773,N_2661);
and UO_42 (O_42,N_2758,N_2779);
or UO_43 (O_43,N_2832,N_2745);
or UO_44 (O_44,N_2775,N_2970);
or UO_45 (O_45,N_2989,N_2663);
nor UO_46 (O_46,N_2638,N_2840);
nand UO_47 (O_47,N_2654,N_2585);
xor UO_48 (O_48,N_2764,N_2471);
or UO_49 (O_49,N_2598,N_2818);
xnor UO_50 (O_50,N_2503,N_2609);
nor UO_51 (O_51,N_2460,N_2694);
nand UO_52 (O_52,N_2814,N_2882);
xnor UO_53 (O_53,N_2652,N_2644);
nand UO_54 (O_54,N_2608,N_2860);
nor UO_55 (O_55,N_2894,N_2414);
and UO_56 (O_56,N_2647,N_2626);
nor UO_57 (O_57,N_2627,N_2720);
nor UO_58 (O_58,N_2805,N_2850);
nand UO_59 (O_59,N_2864,N_2437);
or UO_60 (O_60,N_2777,N_2646);
nand UO_61 (O_61,N_2731,N_2539);
xor UO_62 (O_62,N_2767,N_2891);
nand UO_63 (O_63,N_2885,N_2500);
or UO_64 (O_64,N_2965,N_2490);
nand UO_65 (O_65,N_2742,N_2620);
nor UO_66 (O_66,N_2804,N_2856);
nand UO_67 (O_67,N_2418,N_2407);
or UO_68 (O_68,N_2917,N_2579);
xnor UO_69 (O_69,N_2985,N_2612);
or UO_70 (O_70,N_2820,N_2562);
or UO_71 (O_71,N_2997,N_2634);
nor UO_72 (O_72,N_2712,N_2683);
xnor UO_73 (O_73,N_2540,N_2401);
nor UO_74 (O_74,N_2450,N_2920);
and UO_75 (O_75,N_2461,N_2484);
xor UO_76 (O_76,N_2429,N_2922);
and UO_77 (O_77,N_2893,N_2485);
and UO_78 (O_78,N_2439,N_2617);
xor UO_79 (O_79,N_2632,N_2687);
nand UO_80 (O_80,N_2568,N_2774);
and UO_81 (O_81,N_2888,N_2710);
nor UO_82 (O_82,N_2862,N_2563);
and UO_83 (O_83,N_2754,N_2521);
nand UO_84 (O_84,N_2719,N_2624);
nand UO_85 (O_85,N_2910,N_2852);
nor UO_86 (O_86,N_2451,N_2587);
or UO_87 (O_87,N_2837,N_2939);
nor UO_88 (O_88,N_2974,N_2570);
nor UO_89 (O_89,N_2670,N_2413);
or UO_90 (O_90,N_2921,N_2676);
and UO_91 (O_91,N_2494,N_2690);
or UO_92 (O_92,N_2941,N_2902);
nor UO_93 (O_93,N_2904,N_2509);
and UO_94 (O_94,N_2462,N_2978);
nand UO_95 (O_95,N_2622,N_2945);
and UO_96 (O_96,N_2467,N_2863);
or UO_97 (O_97,N_2696,N_2903);
nor UO_98 (O_98,N_2416,N_2841);
and UO_99 (O_99,N_2830,N_2421);
nand UO_100 (O_100,N_2497,N_2422);
or UO_101 (O_101,N_2479,N_2614);
nor UO_102 (O_102,N_2669,N_2826);
nor UO_103 (O_103,N_2964,N_2469);
nand UO_104 (O_104,N_2600,N_2572);
or UO_105 (O_105,N_2817,N_2992);
nor UO_106 (O_106,N_2534,N_2802);
nor UO_107 (O_107,N_2772,N_2459);
nor UO_108 (O_108,N_2524,N_2980);
and UO_109 (O_109,N_2987,N_2405);
xor UO_110 (O_110,N_2932,N_2452);
nand UO_111 (O_111,N_2957,N_2535);
or UO_112 (O_112,N_2955,N_2799);
nor UO_113 (O_113,N_2463,N_2803);
xor UO_114 (O_114,N_2928,N_2736);
or UO_115 (O_115,N_2954,N_2574);
or UO_116 (O_116,N_2833,N_2537);
and UO_117 (O_117,N_2870,N_2975);
nand UO_118 (O_118,N_2618,N_2749);
or UO_119 (O_119,N_2615,N_2576);
and UO_120 (O_120,N_2512,N_2771);
or UO_121 (O_121,N_2633,N_2428);
nand UO_122 (O_122,N_2756,N_2505);
nand UO_123 (O_123,N_2456,N_2876);
or UO_124 (O_124,N_2610,N_2507);
and UO_125 (O_125,N_2402,N_2605);
nor UO_126 (O_126,N_2763,N_2545);
nor UO_127 (O_127,N_2502,N_2556);
nand UO_128 (O_128,N_2664,N_2776);
nand UO_129 (O_129,N_2946,N_2592);
nor UO_130 (O_130,N_2487,N_2601);
nor UO_131 (O_131,N_2851,N_2409);
nand UO_132 (O_132,N_2853,N_2547);
and UO_133 (O_133,N_2795,N_2686);
nand UO_134 (O_134,N_2698,N_2470);
nand UO_135 (O_135,N_2527,N_2590);
nand UO_136 (O_136,N_2628,N_2982);
nand UO_137 (O_137,N_2541,N_2445);
and UO_138 (O_138,N_2960,N_2715);
or UO_139 (O_139,N_2453,N_2616);
nor UO_140 (O_140,N_2757,N_2723);
and UO_141 (O_141,N_2998,N_2659);
and UO_142 (O_142,N_2898,N_2865);
nand UO_143 (O_143,N_2498,N_2417);
and UO_144 (O_144,N_2641,N_2816);
or UO_145 (O_145,N_2681,N_2635);
or UO_146 (O_146,N_2753,N_2449);
nand UO_147 (O_147,N_2873,N_2430);
xor UO_148 (O_148,N_2740,N_2625);
xnor UO_149 (O_149,N_2476,N_2536);
nor UO_150 (O_150,N_2433,N_2979);
nor UO_151 (O_151,N_2699,N_2602);
nor UO_152 (O_152,N_2859,N_2636);
nand UO_153 (O_153,N_2656,N_2411);
and UO_154 (O_154,N_2611,N_2582);
or UO_155 (O_155,N_2953,N_2561);
xnor UO_156 (O_156,N_2734,N_2948);
nand UO_157 (O_157,N_2702,N_2836);
xor UO_158 (O_158,N_2890,N_2730);
nor UO_159 (O_159,N_2403,N_2613);
nand UO_160 (O_160,N_2966,N_2648);
xor UO_161 (O_161,N_2929,N_2680);
or UO_162 (O_162,N_2905,N_2808);
or UO_163 (O_163,N_2510,N_2743);
and UO_164 (O_164,N_2868,N_2558);
nand UO_165 (O_165,N_2454,N_2768);
and UO_166 (O_166,N_2520,N_2899);
nand UO_167 (O_167,N_2727,N_2496);
nand UO_168 (O_168,N_2684,N_2675);
and UO_169 (O_169,N_2724,N_2936);
nand UO_170 (O_170,N_2789,N_2956);
or UO_171 (O_171,N_2657,N_2784);
nand UO_172 (O_172,N_2495,N_2542);
nand UO_173 (O_173,N_2854,N_2847);
xnor UO_174 (O_174,N_2739,N_2713);
nand UO_175 (O_175,N_2786,N_2986);
nand UO_176 (O_176,N_2642,N_2551);
nor UO_177 (O_177,N_2869,N_2744);
or UO_178 (O_178,N_2543,N_2762);
or UO_179 (O_179,N_2571,N_2637);
nand UO_180 (O_180,N_2538,N_2708);
xor UO_181 (O_181,N_2518,N_2448);
nand UO_182 (O_182,N_2918,N_2806);
xnor UO_183 (O_183,N_2650,N_2916);
and UO_184 (O_184,N_2544,N_2706);
or UO_185 (O_185,N_2728,N_2546);
and UO_186 (O_186,N_2831,N_2961);
and UO_187 (O_187,N_2927,N_2791);
nor UO_188 (O_188,N_2915,N_2770);
and UO_189 (O_189,N_2577,N_2925);
or UO_190 (O_190,N_2682,N_2844);
xor UO_191 (O_191,N_2911,N_2566);
or UO_192 (O_192,N_2580,N_2665);
nand UO_193 (O_193,N_2881,N_2879);
or UO_194 (O_194,N_2511,N_2410);
and UO_195 (O_195,N_2578,N_2591);
and UO_196 (O_196,N_2550,N_2588);
nor UO_197 (O_197,N_2942,N_2857);
or UO_198 (O_198,N_2848,N_2810);
nand UO_199 (O_199,N_2678,N_2866);
nand UO_200 (O_200,N_2871,N_2972);
nand UO_201 (O_201,N_2486,N_2630);
nor UO_202 (O_202,N_2959,N_2564);
and UO_203 (O_203,N_2735,N_2701);
nor UO_204 (O_204,N_2884,N_2688);
nor UO_205 (O_205,N_2465,N_2755);
nand UO_206 (O_206,N_2595,N_2747);
or UO_207 (O_207,N_2969,N_2722);
nor UO_208 (O_208,N_2714,N_2631);
nand UO_209 (O_209,N_2685,N_2567);
nand UO_210 (O_210,N_2968,N_2704);
and UO_211 (O_211,N_2937,N_2967);
or UO_212 (O_212,N_2573,N_2586);
and UO_213 (O_213,N_2931,N_2886);
and UO_214 (O_214,N_2892,N_2643);
or UO_215 (O_215,N_2944,N_2559);
or UO_216 (O_216,N_2478,N_2788);
xnor UO_217 (O_217,N_2838,N_2809);
and UO_218 (O_218,N_2751,N_2934);
nand UO_219 (O_219,N_2813,N_2792);
or UO_220 (O_220,N_2790,N_2621);
and UO_221 (O_221,N_2781,N_2787);
and UO_222 (O_222,N_2835,N_2812);
or UO_223 (O_223,N_2738,N_2482);
and UO_224 (O_224,N_2949,N_2693);
or UO_225 (O_225,N_2464,N_2935);
or UO_226 (O_226,N_2709,N_2716);
nor UO_227 (O_227,N_2639,N_2442);
nor UO_228 (O_228,N_2842,N_2522);
and UO_229 (O_229,N_2603,N_2432);
nor UO_230 (O_230,N_2801,N_2958);
or UO_231 (O_231,N_2640,N_2553);
and UO_232 (O_232,N_2446,N_2440);
nor UO_233 (O_233,N_2671,N_2697);
or UO_234 (O_234,N_2952,N_2584);
or UO_235 (O_235,N_2425,N_2488);
or UO_236 (O_236,N_2473,N_2729);
nand UO_237 (O_237,N_2689,N_2973);
nor UO_238 (O_238,N_2783,N_2769);
nor UO_239 (O_239,N_2895,N_2976);
xor UO_240 (O_240,N_2707,N_2532);
or UO_241 (O_241,N_2778,N_2447);
or UO_242 (O_242,N_2438,N_2824);
or UO_243 (O_243,N_2480,N_2995);
and UO_244 (O_244,N_2996,N_2560);
xnor UO_245 (O_245,N_2906,N_2692);
nand UO_246 (O_246,N_2993,N_2896);
and UO_247 (O_247,N_2761,N_2552);
xor UO_248 (O_248,N_2875,N_2858);
or UO_249 (O_249,N_2759,N_2913);
and UO_250 (O_250,N_2481,N_2593);
nand UO_251 (O_251,N_2984,N_2519);
or UO_252 (O_252,N_2983,N_2604);
nor UO_253 (O_253,N_2994,N_2821);
nor UO_254 (O_254,N_2807,N_2666);
nand UO_255 (O_255,N_2780,N_2427);
or UO_256 (O_256,N_2765,N_2907);
or UO_257 (O_257,N_2441,N_2849);
nand UO_258 (O_258,N_2827,N_2938);
xnor UO_259 (O_259,N_2599,N_2565);
nand UO_260 (O_260,N_2717,N_2861);
nor UO_261 (O_261,N_2846,N_2843);
nand UO_262 (O_262,N_2940,N_2733);
nand UO_263 (O_263,N_2796,N_2606);
and UO_264 (O_264,N_2436,N_2415);
nand UO_265 (O_265,N_2672,N_2645);
nor UO_266 (O_266,N_2655,N_2822);
and UO_267 (O_267,N_2668,N_2711);
nand UO_268 (O_268,N_2434,N_2794);
nand UO_269 (O_269,N_2466,N_2878);
nand UO_270 (O_270,N_2912,N_2629);
and UO_271 (O_271,N_2530,N_2760);
nand UO_272 (O_272,N_2999,N_2752);
and UO_273 (O_273,N_2900,N_2501);
and UO_274 (O_274,N_2523,N_2855);
or UO_275 (O_275,N_2400,N_2557);
and UO_276 (O_276,N_2943,N_2583);
and UO_277 (O_277,N_2930,N_2887);
nand UO_278 (O_278,N_2554,N_2426);
or UO_279 (O_279,N_2962,N_2477);
and UO_280 (O_280,N_2525,N_2506);
or UO_281 (O_281,N_2705,N_2531);
nor UO_282 (O_282,N_2909,N_2404);
and UO_283 (O_283,N_2491,N_2737);
xnor UO_284 (O_284,N_2981,N_2926);
nor UO_285 (O_285,N_2667,N_2594);
or UO_286 (O_286,N_2726,N_2658);
and UO_287 (O_287,N_2748,N_2653);
xor UO_288 (O_288,N_2732,N_2897);
nand UO_289 (O_289,N_2839,N_2815);
nor UO_290 (O_290,N_2766,N_2991);
nor UO_291 (O_291,N_2785,N_2889);
xor UO_292 (O_292,N_2528,N_2700);
or UO_293 (O_293,N_2472,N_2623);
nor UO_294 (O_294,N_2819,N_2548);
nand UO_295 (O_295,N_2971,N_2529);
and UO_296 (O_296,N_2867,N_2901);
xnor UO_297 (O_297,N_2443,N_2457);
nor UO_298 (O_298,N_2908,N_2555);
xor UO_299 (O_299,N_2797,N_2513);
nand UO_300 (O_300,N_2580,N_2968);
nand UO_301 (O_301,N_2749,N_2879);
nor UO_302 (O_302,N_2541,N_2986);
nor UO_303 (O_303,N_2520,N_2905);
nand UO_304 (O_304,N_2474,N_2902);
nand UO_305 (O_305,N_2619,N_2648);
and UO_306 (O_306,N_2964,N_2698);
nand UO_307 (O_307,N_2794,N_2431);
xnor UO_308 (O_308,N_2461,N_2852);
xnor UO_309 (O_309,N_2432,N_2656);
nor UO_310 (O_310,N_2688,N_2885);
and UO_311 (O_311,N_2675,N_2709);
nand UO_312 (O_312,N_2795,N_2484);
and UO_313 (O_313,N_2901,N_2940);
nor UO_314 (O_314,N_2522,N_2675);
xnor UO_315 (O_315,N_2540,N_2861);
nor UO_316 (O_316,N_2618,N_2647);
nor UO_317 (O_317,N_2766,N_2666);
and UO_318 (O_318,N_2474,N_2668);
or UO_319 (O_319,N_2847,N_2973);
xor UO_320 (O_320,N_2762,N_2658);
and UO_321 (O_321,N_2425,N_2821);
nand UO_322 (O_322,N_2533,N_2880);
or UO_323 (O_323,N_2800,N_2991);
nor UO_324 (O_324,N_2710,N_2453);
nand UO_325 (O_325,N_2685,N_2717);
nand UO_326 (O_326,N_2900,N_2819);
nor UO_327 (O_327,N_2544,N_2966);
or UO_328 (O_328,N_2736,N_2699);
nor UO_329 (O_329,N_2945,N_2743);
and UO_330 (O_330,N_2854,N_2602);
nor UO_331 (O_331,N_2496,N_2656);
nand UO_332 (O_332,N_2501,N_2464);
xnor UO_333 (O_333,N_2484,N_2736);
or UO_334 (O_334,N_2519,N_2932);
and UO_335 (O_335,N_2705,N_2971);
and UO_336 (O_336,N_2665,N_2424);
and UO_337 (O_337,N_2615,N_2777);
or UO_338 (O_338,N_2876,N_2802);
or UO_339 (O_339,N_2902,N_2461);
nand UO_340 (O_340,N_2666,N_2679);
or UO_341 (O_341,N_2890,N_2433);
or UO_342 (O_342,N_2659,N_2861);
and UO_343 (O_343,N_2560,N_2929);
and UO_344 (O_344,N_2771,N_2855);
xnor UO_345 (O_345,N_2402,N_2478);
and UO_346 (O_346,N_2875,N_2815);
nand UO_347 (O_347,N_2531,N_2875);
nor UO_348 (O_348,N_2748,N_2695);
xor UO_349 (O_349,N_2934,N_2997);
or UO_350 (O_350,N_2537,N_2552);
and UO_351 (O_351,N_2685,N_2785);
and UO_352 (O_352,N_2446,N_2736);
or UO_353 (O_353,N_2685,N_2743);
nor UO_354 (O_354,N_2945,N_2456);
nor UO_355 (O_355,N_2851,N_2961);
and UO_356 (O_356,N_2699,N_2903);
nand UO_357 (O_357,N_2418,N_2708);
and UO_358 (O_358,N_2662,N_2492);
and UO_359 (O_359,N_2840,N_2464);
and UO_360 (O_360,N_2553,N_2712);
nand UO_361 (O_361,N_2774,N_2891);
and UO_362 (O_362,N_2435,N_2878);
and UO_363 (O_363,N_2912,N_2413);
nand UO_364 (O_364,N_2479,N_2631);
xnor UO_365 (O_365,N_2508,N_2723);
or UO_366 (O_366,N_2879,N_2892);
xnor UO_367 (O_367,N_2691,N_2791);
nand UO_368 (O_368,N_2617,N_2641);
nand UO_369 (O_369,N_2754,N_2516);
and UO_370 (O_370,N_2436,N_2697);
or UO_371 (O_371,N_2618,N_2807);
nand UO_372 (O_372,N_2946,N_2718);
nor UO_373 (O_373,N_2905,N_2961);
xor UO_374 (O_374,N_2556,N_2737);
nor UO_375 (O_375,N_2563,N_2591);
and UO_376 (O_376,N_2862,N_2764);
and UO_377 (O_377,N_2634,N_2414);
nor UO_378 (O_378,N_2483,N_2982);
nand UO_379 (O_379,N_2684,N_2559);
nor UO_380 (O_380,N_2945,N_2498);
nand UO_381 (O_381,N_2986,N_2969);
and UO_382 (O_382,N_2489,N_2967);
nor UO_383 (O_383,N_2510,N_2943);
nand UO_384 (O_384,N_2416,N_2582);
and UO_385 (O_385,N_2682,N_2889);
nor UO_386 (O_386,N_2705,N_2688);
nand UO_387 (O_387,N_2468,N_2548);
and UO_388 (O_388,N_2722,N_2886);
or UO_389 (O_389,N_2452,N_2779);
or UO_390 (O_390,N_2500,N_2745);
nor UO_391 (O_391,N_2946,N_2963);
nand UO_392 (O_392,N_2974,N_2608);
and UO_393 (O_393,N_2891,N_2995);
and UO_394 (O_394,N_2605,N_2825);
nor UO_395 (O_395,N_2460,N_2944);
nand UO_396 (O_396,N_2594,N_2963);
or UO_397 (O_397,N_2974,N_2805);
nand UO_398 (O_398,N_2400,N_2948);
and UO_399 (O_399,N_2530,N_2516);
nor UO_400 (O_400,N_2751,N_2647);
or UO_401 (O_401,N_2413,N_2469);
nor UO_402 (O_402,N_2537,N_2621);
xor UO_403 (O_403,N_2855,N_2693);
nand UO_404 (O_404,N_2612,N_2561);
or UO_405 (O_405,N_2788,N_2748);
or UO_406 (O_406,N_2784,N_2816);
xor UO_407 (O_407,N_2667,N_2468);
or UO_408 (O_408,N_2709,N_2499);
xor UO_409 (O_409,N_2509,N_2762);
and UO_410 (O_410,N_2414,N_2517);
nand UO_411 (O_411,N_2927,N_2922);
nor UO_412 (O_412,N_2434,N_2960);
and UO_413 (O_413,N_2669,N_2579);
nor UO_414 (O_414,N_2712,N_2492);
and UO_415 (O_415,N_2627,N_2742);
and UO_416 (O_416,N_2423,N_2921);
nor UO_417 (O_417,N_2716,N_2864);
nor UO_418 (O_418,N_2939,N_2523);
or UO_419 (O_419,N_2728,N_2761);
nand UO_420 (O_420,N_2713,N_2807);
nor UO_421 (O_421,N_2843,N_2672);
xnor UO_422 (O_422,N_2459,N_2918);
nor UO_423 (O_423,N_2763,N_2895);
and UO_424 (O_424,N_2974,N_2890);
xnor UO_425 (O_425,N_2914,N_2723);
nor UO_426 (O_426,N_2844,N_2752);
nand UO_427 (O_427,N_2423,N_2837);
nand UO_428 (O_428,N_2796,N_2851);
xnor UO_429 (O_429,N_2772,N_2478);
nand UO_430 (O_430,N_2554,N_2684);
nand UO_431 (O_431,N_2600,N_2927);
and UO_432 (O_432,N_2449,N_2473);
nor UO_433 (O_433,N_2643,N_2576);
and UO_434 (O_434,N_2989,N_2635);
or UO_435 (O_435,N_2769,N_2423);
and UO_436 (O_436,N_2849,N_2845);
or UO_437 (O_437,N_2602,N_2472);
and UO_438 (O_438,N_2889,N_2758);
nand UO_439 (O_439,N_2932,N_2776);
nor UO_440 (O_440,N_2818,N_2442);
nor UO_441 (O_441,N_2738,N_2441);
nor UO_442 (O_442,N_2669,N_2794);
and UO_443 (O_443,N_2970,N_2665);
nand UO_444 (O_444,N_2770,N_2858);
and UO_445 (O_445,N_2881,N_2916);
or UO_446 (O_446,N_2718,N_2852);
nand UO_447 (O_447,N_2872,N_2556);
or UO_448 (O_448,N_2572,N_2581);
or UO_449 (O_449,N_2611,N_2880);
or UO_450 (O_450,N_2663,N_2852);
nand UO_451 (O_451,N_2529,N_2564);
nor UO_452 (O_452,N_2819,N_2834);
and UO_453 (O_453,N_2578,N_2677);
nor UO_454 (O_454,N_2852,N_2987);
nor UO_455 (O_455,N_2891,N_2968);
nand UO_456 (O_456,N_2678,N_2901);
nor UO_457 (O_457,N_2679,N_2774);
or UO_458 (O_458,N_2617,N_2760);
and UO_459 (O_459,N_2706,N_2494);
nand UO_460 (O_460,N_2485,N_2468);
and UO_461 (O_461,N_2945,N_2536);
xor UO_462 (O_462,N_2881,N_2480);
nor UO_463 (O_463,N_2735,N_2982);
or UO_464 (O_464,N_2886,N_2433);
or UO_465 (O_465,N_2637,N_2965);
or UO_466 (O_466,N_2882,N_2921);
nor UO_467 (O_467,N_2912,N_2535);
and UO_468 (O_468,N_2599,N_2400);
nor UO_469 (O_469,N_2847,N_2637);
xor UO_470 (O_470,N_2899,N_2646);
or UO_471 (O_471,N_2465,N_2587);
nand UO_472 (O_472,N_2856,N_2831);
and UO_473 (O_473,N_2659,N_2833);
nand UO_474 (O_474,N_2498,N_2521);
nor UO_475 (O_475,N_2731,N_2440);
or UO_476 (O_476,N_2988,N_2499);
nand UO_477 (O_477,N_2708,N_2817);
nand UO_478 (O_478,N_2562,N_2756);
nand UO_479 (O_479,N_2905,N_2901);
nand UO_480 (O_480,N_2946,N_2904);
and UO_481 (O_481,N_2521,N_2491);
and UO_482 (O_482,N_2451,N_2977);
nor UO_483 (O_483,N_2927,N_2725);
or UO_484 (O_484,N_2437,N_2579);
nand UO_485 (O_485,N_2652,N_2664);
nor UO_486 (O_486,N_2745,N_2498);
nor UO_487 (O_487,N_2494,N_2606);
or UO_488 (O_488,N_2936,N_2524);
nand UO_489 (O_489,N_2619,N_2476);
nand UO_490 (O_490,N_2897,N_2563);
and UO_491 (O_491,N_2763,N_2525);
xnor UO_492 (O_492,N_2511,N_2848);
or UO_493 (O_493,N_2802,N_2566);
and UO_494 (O_494,N_2872,N_2420);
or UO_495 (O_495,N_2842,N_2401);
or UO_496 (O_496,N_2673,N_2818);
or UO_497 (O_497,N_2971,N_2942);
and UO_498 (O_498,N_2609,N_2884);
or UO_499 (O_499,N_2850,N_2700);
endmodule