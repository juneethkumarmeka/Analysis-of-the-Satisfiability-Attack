module basic_500_3000_500_50_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_417,In_362);
nand U1 (N_1,In_328,In_70);
nand U2 (N_2,In_146,In_42);
or U3 (N_3,In_389,In_221);
nand U4 (N_4,In_404,In_354);
and U5 (N_5,In_304,In_229);
and U6 (N_6,In_485,In_147);
and U7 (N_7,In_211,In_444);
or U8 (N_8,In_111,In_63);
and U9 (N_9,In_468,In_240);
and U10 (N_10,In_39,In_38);
nor U11 (N_11,In_258,In_290);
and U12 (N_12,In_381,In_357);
or U13 (N_13,In_453,In_225);
nand U14 (N_14,In_432,In_117);
or U15 (N_15,In_7,In_277);
and U16 (N_16,In_448,In_65);
nand U17 (N_17,In_334,In_185);
nand U18 (N_18,In_497,In_455);
nand U19 (N_19,In_450,In_219);
and U20 (N_20,In_251,In_447);
and U21 (N_21,In_152,In_297);
nor U22 (N_22,In_479,In_28);
nand U23 (N_23,In_246,In_391);
nor U24 (N_24,In_10,In_428);
nor U25 (N_25,In_406,In_437);
and U26 (N_26,In_414,In_93);
and U27 (N_27,In_215,In_168);
nor U28 (N_28,In_60,In_238);
or U29 (N_29,In_136,In_114);
or U30 (N_30,In_139,In_281);
nand U31 (N_31,In_143,In_69);
or U32 (N_32,In_127,In_314);
or U33 (N_33,In_423,In_312);
or U34 (N_34,In_376,In_426);
nor U35 (N_35,In_394,In_399);
and U36 (N_36,In_199,In_403);
and U37 (N_37,In_237,In_87);
nand U38 (N_38,In_31,In_411);
nor U39 (N_39,In_96,In_1);
or U40 (N_40,In_440,In_125);
nor U41 (N_41,In_164,In_186);
and U42 (N_42,In_295,In_167);
and U43 (N_43,In_388,In_310);
nand U44 (N_44,In_492,In_44);
or U45 (N_45,In_126,In_313);
nand U46 (N_46,In_467,In_35);
and U47 (N_47,In_308,In_192);
or U48 (N_48,In_375,In_332);
and U49 (N_49,In_436,In_74);
or U50 (N_50,In_18,In_371);
or U51 (N_51,In_5,In_190);
and U52 (N_52,In_330,In_161);
and U53 (N_53,In_269,In_148);
nor U54 (N_54,In_487,In_9);
or U55 (N_55,In_283,In_400);
xnor U56 (N_56,In_110,In_155);
nand U57 (N_57,In_288,In_317);
and U58 (N_58,In_265,In_178);
and U59 (N_59,In_272,In_208);
nor U60 (N_60,In_442,In_408);
nand U61 (N_61,In_395,In_257);
nand U62 (N_62,In_141,N_13);
or U63 (N_63,In_260,In_239);
and U64 (N_64,In_153,In_254);
and U65 (N_65,In_478,N_50);
and U66 (N_66,In_476,In_441);
nand U67 (N_67,In_438,In_392);
nor U68 (N_68,In_378,In_390);
and U69 (N_69,In_159,In_105);
xnor U70 (N_70,In_475,N_52);
and U71 (N_71,In_232,In_81);
or U72 (N_72,In_279,In_171);
nand U73 (N_73,In_103,N_9);
nand U74 (N_74,In_494,N_8);
nor U75 (N_75,In_355,In_116);
or U76 (N_76,N_21,In_274);
and U77 (N_77,In_309,In_256);
nand U78 (N_78,N_17,In_224);
nand U79 (N_79,N_18,In_489);
nand U80 (N_80,In_36,In_303);
and U81 (N_81,In_307,In_195);
or U82 (N_82,N_20,In_348);
and U83 (N_83,In_306,In_337);
nor U84 (N_84,In_109,In_369);
or U85 (N_85,In_121,In_300);
nand U86 (N_86,In_416,In_15);
or U87 (N_87,In_112,In_187);
nand U88 (N_88,In_212,In_429);
and U89 (N_89,In_459,In_298);
and U90 (N_90,In_104,In_361);
and U91 (N_91,In_14,In_101);
nor U92 (N_92,In_252,N_14);
nor U93 (N_93,In_352,In_207);
or U94 (N_94,In_51,In_245);
nand U95 (N_95,In_446,In_387);
or U96 (N_96,N_27,In_234);
nor U97 (N_97,In_79,In_318);
nor U98 (N_98,In_53,In_386);
nand U99 (N_99,In_94,In_316);
nor U100 (N_100,In_276,N_53);
or U101 (N_101,In_471,In_89);
xor U102 (N_102,In_78,In_130);
nand U103 (N_103,In_202,In_353);
nor U104 (N_104,In_261,In_336);
nand U105 (N_105,N_40,In_449);
or U106 (N_106,In_48,In_135);
nand U107 (N_107,In_499,In_255);
and U108 (N_108,N_37,In_21);
or U109 (N_109,N_55,In_80);
or U110 (N_110,In_131,N_51);
xnor U111 (N_111,In_299,N_30);
nand U112 (N_112,In_339,In_24);
and U113 (N_113,In_173,In_323);
or U114 (N_114,In_289,In_333);
nor U115 (N_115,In_372,In_204);
and U116 (N_116,In_359,In_62);
nand U117 (N_117,In_140,In_122);
nor U118 (N_118,In_193,In_345);
or U119 (N_119,In_123,In_356);
or U120 (N_120,In_346,In_377);
and U121 (N_121,In_54,In_341);
nand U122 (N_122,In_157,In_250);
or U123 (N_123,N_109,N_63);
and U124 (N_124,In_55,In_226);
or U125 (N_125,In_460,In_464);
or U126 (N_126,In_12,N_54);
nand U127 (N_127,In_291,N_0);
nor U128 (N_128,In_249,In_85);
nor U129 (N_129,In_64,In_160);
nor U130 (N_130,In_443,In_118);
nor U131 (N_131,In_165,In_335);
or U132 (N_132,In_40,N_32);
nor U133 (N_133,N_26,N_95);
nor U134 (N_134,In_99,In_498);
or U135 (N_135,N_111,In_458);
or U136 (N_136,In_86,In_68);
and U137 (N_137,In_194,N_67);
nor U138 (N_138,In_231,N_103);
and U139 (N_139,In_113,In_469);
nand U140 (N_140,In_177,In_418);
and U141 (N_141,In_46,In_129);
and U142 (N_142,In_247,In_268);
or U143 (N_143,N_118,In_91);
or U144 (N_144,N_85,In_350);
nand U145 (N_145,In_197,N_107);
and U146 (N_146,In_236,In_427);
or U147 (N_147,N_56,In_120);
or U148 (N_148,In_223,In_128);
nor U149 (N_149,In_4,In_174);
and U150 (N_150,In_67,In_439);
and U151 (N_151,N_84,In_434);
and U152 (N_152,In_66,In_379);
nand U153 (N_153,N_7,N_115);
and U154 (N_154,In_366,N_70);
and U155 (N_155,In_17,In_34);
nor U156 (N_156,In_301,N_22);
nor U157 (N_157,In_92,In_214);
nor U158 (N_158,N_48,N_46);
xnor U159 (N_159,In_196,In_338);
or U160 (N_160,In_456,In_61);
nand U161 (N_161,In_222,In_16);
or U162 (N_162,In_25,In_396);
nand U163 (N_163,In_321,In_27);
nand U164 (N_164,N_29,N_69);
and U165 (N_165,In_270,In_220);
nor U166 (N_166,In_209,In_3);
nor U167 (N_167,In_480,In_235);
nor U168 (N_168,N_75,N_66);
nor U169 (N_169,N_59,In_115);
or U170 (N_170,N_76,In_430);
or U171 (N_171,In_20,N_62);
or U172 (N_172,N_105,In_98);
and U173 (N_173,In_45,N_41);
or U174 (N_174,In_151,N_114);
nand U175 (N_175,N_44,In_156);
xnor U176 (N_176,N_42,N_43);
and U177 (N_177,In_95,N_49);
or U178 (N_178,In_97,N_119);
nor U179 (N_179,N_87,In_189);
and U180 (N_180,In_287,N_128);
nor U181 (N_181,In_82,N_164);
and U182 (N_182,N_170,N_140);
and U183 (N_183,N_45,N_175);
nor U184 (N_184,N_141,In_280);
nor U185 (N_185,N_168,N_162);
nand U186 (N_186,In_43,In_420);
or U187 (N_187,In_433,N_161);
nand U188 (N_188,N_112,In_198);
nor U189 (N_189,In_2,In_302);
or U190 (N_190,In_474,In_343);
or U191 (N_191,N_10,In_319);
nand U192 (N_192,N_15,In_180);
nor U193 (N_193,N_139,In_138);
nand U194 (N_194,In_71,N_92);
or U195 (N_195,In_324,In_266);
nor U196 (N_196,In_495,In_382);
xnor U197 (N_197,N_172,In_384);
nand U198 (N_198,In_326,N_68);
nand U199 (N_199,N_5,N_178);
xor U200 (N_200,In_76,N_125);
nor U201 (N_201,In_452,In_37);
or U202 (N_202,N_149,N_3);
xor U203 (N_203,In_367,In_150);
nand U204 (N_204,N_131,In_169);
nor U205 (N_205,N_93,N_88);
nand U206 (N_206,In_216,In_413);
and U207 (N_207,In_210,In_241);
nor U208 (N_208,In_175,In_132);
nor U209 (N_209,In_26,In_472);
nand U210 (N_210,In_496,In_370);
and U211 (N_211,In_0,N_110);
or U212 (N_212,In_285,In_412);
nand U213 (N_213,In_205,In_107);
nand U214 (N_214,In_203,In_405);
nand U215 (N_215,N_177,N_90);
nor U216 (N_216,In_166,N_136);
and U217 (N_217,In_47,In_410);
nor U218 (N_218,In_422,In_30);
nor U219 (N_219,N_91,In_286);
and U220 (N_220,In_402,In_267);
nand U221 (N_221,In_293,In_72);
nor U222 (N_222,N_104,N_165);
and U223 (N_223,In_347,N_2);
nand U224 (N_224,N_143,N_1);
nand U225 (N_225,In_142,In_275);
nor U226 (N_226,In_415,In_483);
nand U227 (N_227,In_200,N_135);
xnor U228 (N_228,N_113,N_151);
nand U229 (N_229,N_72,N_160);
and U230 (N_230,N_6,N_83);
and U231 (N_231,In_213,N_38);
nor U232 (N_232,In_228,In_477);
nand U233 (N_233,In_393,In_6);
or U234 (N_234,N_153,N_133);
and U235 (N_235,In_425,In_119);
nand U236 (N_236,In_243,N_159);
nand U237 (N_237,N_122,In_457);
and U238 (N_238,In_259,N_16);
or U239 (N_239,In_325,N_134);
nor U240 (N_240,N_34,In_358);
and U241 (N_241,In_52,N_237);
or U242 (N_242,N_203,In_217);
or U243 (N_243,In_88,N_152);
and U244 (N_244,In_145,N_171);
nor U245 (N_245,N_200,N_25);
nand U246 (N_246,N_138,N_193);
nor U247 (N_247,N_82,In_84);
and U248 (N_248,In_470,N_197);
xor U249 (N_249,In_351,In_363);
nor U250 (N_250,In_263,In_163);
nand U251 (N_251,In_264,N_96);
nand U252 (N_252,N_214,N_201);
nand U253 (N_253,In_364,In_29);
or U254 (N_254,In_397,In_75);
and U255 (N_255,N_130,In_108);
xor U256 (N_256,In_305,In_385);
nand U257 (N_257,N_205,N_132);
nor U258 (N_258,In_248,In_253);
and U259 (N_259,N_146,N_229);
or U260 (N_260,N_31,In_431);
nand U261 (N_261,N_217,N_23);
and U262 (N_262,In_419,N_230);
nor U263 (N_263,N_126,In_179);
or U264 (N_264,In_398,N_81);
nor U265 (N_265,N_79,In_329);
or U266 (N_266,In_365,N_225);
or U267 (N_267,In_73,N_236);
or U268 (N_268,N_117,N_142);
or U269 (N_269,N_167,N_204);
nor U270 (N_270,In_463,N_222);
or U271 (N_271,N_231,N_194);
and U272 (N_272,In_11,N_12);
nand U273 (N_273,In_294,In_124);
and U274 (N_274,N_184,In_59);
and U275 (N_275,In_83,In_134);
nor U276 (N_276,In_172,In_311);
nor U277 (N_277,N_206,In_176);
nand U278 (N_278,In_466,In_284);
nand U279 (N_279,N_124,In_486);
and U280 (N_280,N_145,In_57);
nand U281 (N_281,In_106,N_180);
xor U282 (N_282,N_209,In_407);
nand U283 (N_283,N_183,N_78);
and U284 (N_284,N_58,In_102);
or U285 (N_285,In_462,In_373);
or U286 (N_286,In_58,N_181);
nor U287 (N_287,In_191,N_227);
nor U288 (N_288,In_374,In_144);
nor U289 (N_289,In_383,In_445);
nand U290 (N_290,N_39,In_23);
nand U291 (N_291,In_162,In_33);
or U292 (N_292,N_156,N_198);
nand U293 (N_293,N_235,In_368);
and U294 (N_294,In_154,In_41);
nor U295 (N_295,N_4,N_157);
and U296 (N_296,N_35,N_108);
nand U297 (N_297,In_184,N_187);
nor U298 (N_298,N_221,N_101);
or U299 (N_299,N_97,In_218);
or U300 (N_300,N_99,In_181);
and U301 (N_301,In_230,In_242);
or U302 (N_302,In_233,In_149);
or U303 (N_303,In_182,N_247);
and U304 (N_304,N_28,N_188);
nand U305 (N_305,N_278,N_176);
and U306 (N_306,N_223,N_275);
nand U307 (N_307,N_120,N_89);
nor U308 (N_308,N_182,N_174);
nand U309 (N_309,In_262,N_190);
or U310 (N_310,N_218,In_435);
and U311 (N_311,N_249,In_409);
and U312 (N_312,N_240,N_77);
nor U313 (N_313,N_226,N_215);
or U314 (N_314,N_179,In_454);
nor U315 (N_315,N_94,In_273);
nand U316 (N_316,In_49,N_191);
and U317 (N_317,In_100,N_253);
and U318 (N_318,N_292,N_158);
and U319 (N_319,In_188,N_129);
and U320 (N_320,In_278,In_461);
nand U321 (N_321,N_279,N_144);
nor U322 (N_322,N_224,N_286);
and U323 (N_323,In_331,In_90);
nand U324 (N_324,N_147,In_158);
and U325 (N_325,N_290,N_74);
and U326 (N_326,N_155,In_282);
xnor U327 (N_327,N_271,In_22);
or U328 (N_328,N_220,N_258);
or U329 (N_329,N_267,In_473);
nor U330 (N_330,In_133,In_206);
and U331 (N_331,N_297,N_294);
or U332 (N_332,N_192,N_216);
or U333 (N_333,N_261,N_123);
or U334 (N_334,N_33,N_64);
nand U335 (N_335,In_170,N_127);
or U336 (N_336,N_211,N_264);
nor U337 (N_337,In_296,N_61);
nor U338 (N_338,N_246,N_251);
and U339 (N_339,N_277,In_380);
nor U340 (N_340,N_163,N_173);
and U341 (N_341,N_287,N_47);
nand U342 (N_342,In_327,N_116);
nor U343 (N_343,In_227,In_401);
or U344 (N_344,N_24,N_102);
nand U345 (N_345,N_268,In_32);
nor U346 (N_346,In_322,N_166);
and U347 (N_347,N_270,N_71);
and U348 (N_348,In_424,N_273);
nand U349 (N_349,N_291,In_77);
nand U350 (N_350,N_255,N_289);
and U351 (N_351,N_248,In_50);
xnor U352 (N_352,N_276,N_189);
or U353 (N_353,N_282,N_207);
nor U354 (N_354,N_288,In_183);
and U355 (N_355,N_254,N_259);
nand U356 (N_356,N_266,In_491);
or U357 (N_357,In_340,N_196);
nand U358 (N_358,N_244,In_349);
nor U359 (N_359,N_100,N_281);
nor U360 (N_360,In_344,N_313);
or U361 (N_361,N_260,N_293);
or U362 (N_362,N_339,N_345);
nor U363 (N_363,N_338,N_121);
nor U364 (N_364,N_269,N_219);
and U365 (N_365,In_451,N_274);
or U366 (N_366,In_244,N_280);
nor U367 (N_367,In_421,N_80);
nand U368 (N_368,N_239,In_481);
or U369 (N_369,N_298,In_465);
nand U370 (N_370,N_320,N_137);
nor U371 (N_371,N_300,N_213);
nor U372 (N_372,N_238,N_343);
nor U373 (N_373,N_317,N_232);
or U374 (N_374,N_195,N_252);
or U375 (N_375,N_319,N_307);
or U376 (N_376,N_250,N_323);
or U377 (N_377,N_256,N_243);
nand U378 (N_378,N_312,N_334);
or U379 (N_379,N_318,N_228);
and U380 (N_380,N_305,N_272);
or U381 (N_381,N_210,N_283);
nand U382 (N_382,N_233,In_490);
or U383 (N_383,In_292,N_358);
nand U384 (N_384,N_303,N_311);
nor U385 (N_385,N_354,N_357);
or U386 (N_386,N_310,N_314);
and U387 (N_387,N_349,N_208);
and U388 (N_388,N_315,In_493);
nand U389 (N_389,N_350,N_65);
and U390 (N_390,In_8,N_352);
and U391 (N_391,N_324,In_201);
nand U392 (N_392,N_199,N_326);
nor U393 (N_393,N_185,N_341);
nor U394 (N_394,In_342,N_328);
nand U395 (N_395,N_308,N_257);
and U396 (N_396,N_19,N_304);
and U397 (N_397,N_11,N_241);
or U398 (N_398,N_333,N_359);
and U399 (N_399,N_265,N_295);
nand U400 (N_400,N_337,N_356);
or U401 (N_401,N_242,N_336);
xnor U402 (N_402,N_60,N_322);
or U403 (N_403,In_484,N_284);
nor U404 (N_404,N_154,N_86);
nor U405 (N_405,In_488,N_332);
nor U406 (N_406,In_19,In_137);
and U407 (N_407,N_36,N_285);
nand U408 (N_408,N_329,In_482);
nand U409 (N_409,N_245,N_344);
or U410 (N_410,N_299,N_106);
nand U411 (N_411,N_186,N_347);
nor U412 (N_412,N_351,N_98);
nand U413 (N_413,N_330,N_321);
nor U414 (N_414,N_340,In_315);
and U415 (N_415,N_355,N_342);
or U416 (N_416,N_73,N_353);
nand U417 (N_417,In_320,N_309);
nor U418 (N_418,N_263,N_148);
and U419 (N_419,N_169,N_212);
and U420 (N_420,N_306,N_363);
nand U421 (N_421,N_406,N_381);
and U422 (N_422,N_389,N_384);
and U423 (N_423,N_302,N_234);
or U424 (N_424,N_369,N_400);
or U425 (N_425,N_373,N_395);
nand U426 (N_426,In_13,N_403);
nor U427 (N_427,N_404,N_412);
nand U428 (N_428,N_374,N_301);
and U429 (N_429,N_408,N_390);
nand U430 (N_430,N_410,In_56);
and U431 (N_431,N_386,N_202);
nand U432 (N_432,N_399,N_417);
nand U433 (N_433,N_396,N_335);
nand U434 (N_434,N_57,N_376);
and U435 (N_435,N_370,N_366);
nor U436 (N_436,N_377,N_393);
or U437 (N_437,N_397,N_385);
nand U438 (N_438,N_348,N_150);
and U439 (N_439,N_391,N_367);
nand U440 (N_440,N_316,N_379);
nand U441 (N_441,N_380,N_361);
nand U442 (N_442,N_411,N_368);
or U443 (N_443,N_402,N_364);
nand U444 (N_444,N_415,N_365);
or U445 (N_445,N_372,N_383);
nor U446 (N_446,N_409,N_388);
nor U447 (N_447,In_271,N_405);
nor U448 (N_448,N_414,N_362);
nor U449 (N_449,N_346,N_296);
and U450 (N_450,N_413,N_382);
nand U451 (N_451,N_407,N_392);
and U452 (N_452,N_371,N_331);
or U453 (N_453,N_394,N_360);
and U454 (N_454,N_418,N_387);
and U455 (N_455,N_401,N_375);
or U456 (N_456,N_398,N_262);
nand U457 (N_457,N_416,N_327);
nand U458 (N_458,N_325,In_360);
nand U459 (N_459,N_378,N_419);
nor U460 (N_460,N_391,N_361);
and U461 (N_461,N_386,N_393);
and U462 (N_462,In_13,N_391);
or U463 (N_463,N_361,In_56);
and U464 (N_464,N_388,N_368);
nor U465 (N_465,N_413,N_394);
nor U466 (N_466,N_296,N_394);
xnor U467 (N_467,N_409,N_335);
nor U468 (N_468,N_301,N_378);
or U469 (N_469,N_367,N_57);
nand U470 (N_470,N_388,N_413);
xnor U471 (N_471,N_372,N_404);
nor U472 (N_472,N_405,N_380);
and U473 (N_473,N_379,N_366);
nand U474 (N_474,N_301,N_150);
and U475 (N_475,N_397,N_365);
or U476 (N_476,N_382,N_415);
and U477 (N_477,N_380,N_296);
or U478 (N_478,N_365,N_374);
nand U479 (N_479,N_408,N_398);
nor U480 (N_480,N_452,N_474);
nor U481 (N_481,N_445,N_470);
nand U482 (N_482,N_427,N_478);
nor U483 (N_483,N_421,N_424);
or U484 (N_484,N_430,N_447);
nor U485 (N_485,N_435,N_476);
and U486 (N_486,N_439,N_455);
or U487 (N_487,N_461,N_477);
or U488 (N_488,N_479,N_472);
or U489 (N_489,N_426,N_425);
or U490 (N_490,N_464,N_453);
nand U491 (N_491,N_457,N_444);
and U492 (N_492,N_443,N_441);
nor U493 (N_493,N_454,N_465);
nor U494 (N_494,N_423,N_463);
and U495 (N_495,N_433,N_466);
or U496 (N_496,N_460,N_420);
nor U497 (N_497,N_429,N_434);
and U498 (N_498,N_422,N_442);
and U499 (N_499,N_451,N_440);
nand U500 (N_500,N_446,N_437);
and U501 (N_501,N_448,N_449);
nor U502 (N_502,N_458,N_462);
and U503 (N_503,N_436,N_456);
or U504 (N_504,N_467,N_428);
and U505 (N_505,N_469,N_473);
nand U506 (N_506,N_468,N_431);
or U507 (N_507,N_475,N_450);
and U508 (N_508,N_471,N_459);
or U509 (N_509,N_432,N_438);
or U510 (N_510,N_429,N_432);
nor U511 (N_511,N_471,N_424);
nor U512 (N_512,N_469,N_465);
nor U513 (N_513,N_456,N_458);
nor U514 (N_514,N_429,N_475);
nor U515 (N_515,N_458,N_452);
nand U516 (N_516,N_440,N_441);
or U517 (N_517,N_426,N_432);
and U518 (N_518,N_429,N_444);
or U519 (N_519,N_455,N_430);
and U520 (N_520,N_448,N_475);
nand U521 (N_521,N_477,N_473);
nand U522 (N_522,N_442,N_468);
and U523 (N_523,N_470,N_447);
nand U524 (N_524,N_453,N_466);
and U525 (N_525,N_438,N_479);
nand U526 (N_526,N_456,N_477);
or U527 (N_527,N_457,N_474);
xnor U528 (N_528,N_438,N_441);
nor U529 (N_529,N_458,N_453);
nor U530 (N_530,N_478,N_458);
and U531 (N_531,N_422,N_455);
nand U532 (N_532,N_421,N_464);
or U533 (N_533,N_420,N_474);
or U534 (N_534,N_428,N_468);
or U535 (N_535,N_441,N_469);
nand U536 (N_536,N_466,N_469);
xnor U537 (N_537,N_455,N_429);
or U538 (N_538,N_462,N_460);
nand U539 (N_539,N_422,N_433);
and U540 (N_540,N_486,N_512);
nand U541 (N_541,N_484,N_503);
nand U542 (N_542,N_532,N_504);
and U543 (N_543,N_489,N_536);
nand U544 (N_544,N_531,N_507);
nand U545 (N_545,N_538,N_527);
nand U546 (N_546,N_521,N_525);
nor U547 (N_547,N_523,N_533);
and U548 (N_548,N_539,N_491);
nor U549 (N_549,N_519,N_499);
and U550 (N_550,N_487,N_511);
nand U551 (N_551,N_520,N_490);
nor U552 (N_552,N_505,N_517);
nand U553 (N_553,N_500,N_494);
and U554 (N_554,N_495,N_530);
or U555 (N_555,N_518,N_496);
nand U556 (N_556,N_485,N_537);
nand U557 (N_557,N_502,N_510);
nand U558 (N_558,N_493,N_522);
nor U559 (N_559,N_482,N_488);
and U560 (N_560,N_498,N_497);
and U561 (N_561,N_524,N_481);
xor U562 (N_562,N_526,N_508);
or U563 (N_563,N_516,N_501);
nand U564 (N_564,N_515,N_514);
nor U565 (N_565,N_529,N_480);
nand U566 (N_566,N_509,N_535);
and U567 (N_567,N_513,N_534);
nor U568 (N_568,N_483,N_528);
nand U569 (N_569,N_506,N_492);
nor U570 (N_570,N_537,N_508);
nand U571 (N_571,N_536,N_510);
nor U572 (N_572,N_500,N_528);
nand U573 (N_573,N_514,N_485);
and U574 (N_574,N_534,N_499);
and U575 (N_575,N_503,N_519);
nor U576 (N_576,N_507,N_486);
nand U577 (N_577,N_514,N_492);
nand U578 (N_578,N_523,N_499);
or U579 (N_579,N_527,N_528);
or U580 (N_580,N_497,N_480);
or U581 (N_581,N_526,N_496);
and U582 (N_582,N_509,N_496);
nand U583 (N_583,N_515,N_481);
nor U584 (N_584,N_503,N_487);
or U585 (N_585,N_512,N_506);
nor U586 (N_586,N_493,N_510);
and U587 (N_587,N_484,N_513);
nor U588 (N_588,N_516,N_521);
and U589 (N_589,N_520,N_483);
and U590 (N_590,N_489,N_510);
xor U591 (N_591,N_488,N_500);
or U592 (N_592,N_524,N_523);
nand U593 (N_593,N_486,N_506);
or U594 (N_594,N_480,N_493);
nor U595 (N_595,N_534,N_500);
nor U596 (N_596,N_503,N_486);
nand U597 (N_597,N_504,N_537);
nor U598 (N_598,N_487,N_526);
xor U599 (N_599,N_521,N_504);
nand U600 (N_600,N_590,N_546);
or U601 (N_601,N_560,N_598);
nor U602 (N_602,N_585,N_545);
and U603 (N_603,N_574,N_594);
nand U604 (N_604,N_561,N_552);
or U605 (N_605,N_556,N_568);
xor U606 (N_606,N_558,N_548);
nor U607 (N_607,N_588,N_599);
and U608 (N_608,N_597,N_550);
or U609 (N_609,N_572,N_596);
nor U610 (N_610,N_549,N_551);
nand U611 (N_611,N_595,N_554);
or U612 (N_612,N_565,N_570);
and U613 (N_613,N_584,N_544);
xnor U614 (N_614,N_592,N_540);
nor U615 (N_615,N_573,N_567);
or U616 (N_616,N_566,N_589);
or U617 (N_617,N_591,N_547);
or U618 (N_618,N_541,N_583);
nand U619 (N_619,N_553,N_593);
or U620 (N_620,N_559,N_580);
nor U621 (N_621,N_579,N_577);
or U622 (N_622,N_575,N_586);
nor U623 (N_623,N_563,N_562);
and U624 (N_624,N_557,N_576);
nand U625 (N_625,N_578,N_581);
or U626 (N_626,N_569,N_555);
nor U627 (N_627,N_543,N_571);
nand U628 (N_628,N_564,N_542);
and U629 (N_629,N_582,N_587);
nand U630 (N_630,N_542,N_553);
nor U631 (N_631,N_551,N_569);
nand U632 (N_632,N_555,N_577);
and U633 (N_633,N_540,N_543);
nor U634 (N_634,N_559,N_593);
and U635 (N_635,N_582,N_565);
and U636 (N_636,N_544,N_546);
nor U637 (N_637,N_541,N_540);
nand U638 (N_638,N_576,N_556);
and U639 (N_639,N_555,N_561);
and U640 (N_640,N_580,N_561);
nand U641 (N_641,N_554,N_589);
and U642 (N_642,N_562,N_599);
nor U643 (N_643,N_564,N_554);
nor U644 (N_644,N_576,N_596);
or U645 (N_645,N_578,N_562);
or U646 (N_646,N_559,N_594);
nor U647 (N_647,N_591,N_567);
or U648 (N_648,N_597,N_572);
or U649 (N_649,N_562,N_571);
nand U650 (N_650,N_598,N_553);
nor U651 (N_651,N_567,N_565);
nor U652 (N_652,N_583,N_547);
nor U653 (N_653,N_590,N_545);
nor U654 (N_654,N_568,N_599);
nand U655 (N_655,N_570,N_566);
or U656 (N_656,N_581,N_590);
nand U657 (N_657,N_541,N_581);
and U658 (N_658,N_594,N_566);
and U659 (N_659,N_558,N_570);
or U660 (N_660,N_601,N_647);
and U661 (N_661,N_641,N_619);
nand U662 (N_662,N_638,N_612);
nand U663 (N_663,N_649,N_628);
and U664 (N_664,N_650,N_615);
or U665 (N_665,N_657,N_602);
or U666 (N_666,N_603,N_613);
or U667 (N_667,N_604,N_652);
nand U668 (N_668,N_624,N_631);
or U669 (N_669,N_639,N_616);
and U670 (N_670,N_634,N_622);
nor U671 (N_671,N_623,N_609);
nor U672 (N_672,N_600,N_644);
nor U673 (N_673,N_605,N_635);
and U674 (N_674,N_643,N_645);
and U675 (N_675,N_659,N_627);
and U676 (N_676,N_629,N_608);
nor U677 (N_677,N_621,N_617);
and U678 (N_678,N_636,N_620);
nor U679 (N_679,N_606,N_646);
nand U680 (N_680,N_611,N_651);
nor U681 (N_681,N_633,N_655);
nand U682 (N_682,N_640,N_653);
nand U683 (N_683,N_656,N_630);
nor U684 (N_684,N_607,N_610);
and U685 (N_685,N_625,N_648);
nor U686 (N_686,N_618,N_632);
nand U687 (N_687,N_626,N_642);
nor U688 (N_688,N_658,N_654);
or U689 (N_689,N_614,N_637);
nand U690 (N_690,N_635,N_655);
nand U691 (N_691,N_616,N_606);
xnor U692 (N_692,N_638,N_654);
or U693 (N_693,N_607,N_623);
and U694 (N_694,N_635,N_634);
nor U695 (N_695,N_610,N_648);
nand U696 (N_696,N_658,N_623);
and U697 (N_697,N_617,N_624);
and U698 (N_698,N_642,N_649);
or U699 (N_699,N_656,N_613);
nand U700 (N_700,N_638,N_602);
and U701 (N_701,N_647,N_659);
and U702 (N_702,N_607,N_647);
and U703 (N_703,N_615,N_611);
nand U704 (N_704,N_601,N_627);
nand U705 (N_705,N_648,N_630);
nand U706 (N_706,N_639,N_631);
and U707 (N_707,N_643,N_622);
and U708 (N_708,N_634,N_632);
nand U709 (N_709,N_623,N_612);
or U710 (N_710,N_611,N_659);
nand U711 (N_711,N_639,N_651);
nor U712 (N_712,N_647,N_645);
or U713 (N_713,N_612,N_620);
or U714 (N_714,N_611,N_608);
and U715 (N_715,N_624,N_647);
nand U716 (N_716,N_657,N_620);
nor U717 (N_717,N_634,N_631);
or U718 (N_718,N_613,N_651);
nand U719 (N_719,N_650,N_655);
or U720 (N_720,N_719,N_701);
nand U721 (N_721,N_678,N_673);
nor U722 (N_722,N_697,N_672);
nor U723 (N_723,N_677,N_669);
nor U724 (N_724,N_692,N_703);
xnor U725 (N_725,N_693,N_688);
nand U726 (N_726,N_670,N_702);
nor U727 (N_727,N_665,N_684);
and U728 (N_728,N_714,N_695);
nor U729 (N_729,N_675,N_664);
nor U730 (N_730,N_662,N_667);
nand U731 (N_731,N_707,N_713);
and U732 (N_732,N_680,N_710);
nand U733 (N_733,N_705,N_694);
nand U734 (N_734,N_716,N_685);
nor U735 (N_735,N_715,N_682);
or U736 (N_736,N_712,N_708);
or U737 (N_737,N_704,N_674);
nand U738 (N_738,N_699,N_666);
and U739 (N_739,N_676,N_687);
or U740 (N_740,N_709,N_717);
nand U741 (N_741,N_671,N_690);
and U742 (N_742,N_679,N_681);
or U743 (N_743,N_661,N_718);
and U744 (N_744,N_696,N_686);
nand U745 (N_745,N_668,N_689);
nor U746 (N_746,N_683,N_698);
or U747 (N_747,N_663,N_691);
or U748 (N_748,N_706,N_700);
xnor U749 (N_749,N_711,N_660);
nor U750 (N_750,N_671,N_706);
or U751 (N_751,N_700,N_703);
nand U752 (N_752,N_679,N_704);
or U753 (N_753,N_682,N_687);
or U754 (N_754,N_681,N_700);
nand U755 (N_755,N_701,N_690);
or U756 (N_756,N_679,N_715);
nor U757 (N_757,N_661,N_668);
nand U758 (N_758,N_697,N_719);
nand U759 (N_759,N_706,N_705);
or U760 (N_760,N_661,N_690);
and U761 (N_761,N_700,N_680);
and U762 (N_762,N_664,N_685);
nand U763 (N_763,N_717,N_675);
nor U764 (N_764,N_696,N_718);
nand U765 (N_765,N_699,N_684);
or U766 (N_766,N_668,N_662);
and U767 (N_767,N_687,N_711);
or U768 (N_768,N_707,N_689);
nand U769 (N_769,N_660,N_709);
and U770 (N_770,N_710,N_699);
and U771 (N_771,N_698,N_687);
xor U772 (N_772,N_662,N_713);
nor U773 (N_773,N_673,N_714);
and U774 (N_774,N_674,N_695);
or U775 (N_775,N_707,N_712);
nand U776 (N_776,N_707,N_665);
nor U777 (N_777,N_704,N_678);
or U778 (N_778,N_717,N_676);
nand U779 (N_779,N_660,N_700);
and U780 (N_780,N_745,N_763);
nand U781 (N_781,N_729,N_750);
xor U782 (N_782,N_762,N_721);
nor U783 (N_783,N_722,N_735);
and U784 (N_784,N_754,N_737);
nand U785 (N_785,N_760,N_736);
nand U786 (N_786,N_724,N_767);
and U787 (N_787,N_738,N_775);
nor U788 (N_788,N_730,N_756);
or U789 (N_789,N_774,N_761);
or U790 (N_790,N_725,N_776);
nor U791 (N_791,N_749,N_771);
nor U792 (N_792,N_743,N_741);
nand U793 (N_793,N_769,N_759);
xnor U794 (N_794,N_772,N_765);
nor U795 (N_795,N_748,N_744);
nor U796 (N_796,N_720,N_757);
or U797 (N_797,N_770,N_742);
nand U798 (N_798,N_758,N_731);
and U799 (N_799,N_733,N_779);
or U800 (N_800,N_752,N_728);
or U801 (N_801,N_755,N_739);
nand U802 (N_802,N_740,N_747);
and U803 (N_803,N_773,N_726);
nor U804 (N_804,N_732,N_777);
or U805 (N_805,N_751,N_778);
xor U806 (N_806,N_766,N_746);
nor U807 (N_807,N_727,N_734);
or U808 (N_808,N_753,N_768);
or U809 (N_809,N_723,N_764);
nand U810 (N_810,N_761,N_771);
nand U811 (N_811,N_755,N_767);
nor U812 (N_812,N_725,N_720);
nor U813 (N_813,N_769,N_724);
and U814 (N_814,N_733,N_742);
or U815 (N_815,N_764,N_744);
and U816 (N_816,N_768,N_732);
nor U817 (N_817,N_745,N_733);
or U818 (N_818,N_738,N_759);
or U819 (N_819,N_756,N_722);
or U820 (N_820,N_744,N_749);
nand U821 (N_821,N_721,N_737);
nand U822 (N_822,N_743,N_744);
and U823 (N_823,N_773,N_751);
nor U824 (N_824,N_763,N_754);
and U825 (N_825,N_769,N_749);
nand U826 (N_826,N_736,N_750);
or U827 (N_827,N_767,N_744);
nor U828 (N_828,N_737,N_730);
nor U829 (N_829,N_730,N_720);
and U830 (N_830,N_772,N_778);
nand U831 (N_831,N_779,N_774);
nor U832 (N_832,N_737,N_777);
or U833 (N_833,N_738,N_772);
and U834 (N_834,N_730,N_757);
or U835 (N_835,N_776,N_770);
nand U836 (N_836,N_727,N_728);
nor U837 (N_837,N_764,N_738);
nand U838 (N_838,N_731,N_761);
or U839 (N_839,N_740,N_776);
or U840 (N_840,N_793,N_815);
and U841 (N_841,N_825,N_811);
and U842 (N_842,N_783,N_803);
nand U843 (N_843,N_795,N_801);
nor U844 (N_844,N_812,N_785);
and U845 (N_845,N_806,N_830);
or U846 (N_846,N_833,N_839);
nor U847 (N_847,N_820,N_813);
nor U848 (N_848,N_827,N_837);
or U849 (N_849,N_826,N_786);
or U850 (N_850,N_796,N_788);
nor U851 (N_851,N_821,N_805);
and U852 (N_852,N_807,N_836);
nor U853 (N_853,N_808,N_800);
and U854 (N_854,N_784,N_818);
or U855 (N_855,N_835,N_814);
or U856 (N_856,N_838,N_829);
or U857 (N_857,N_802,N_816);
nand U858 (N_858,N_791,N_797);
or U859 (N_859,N_828,N_798);
or U860 (N_860,N_834,N_790);
or U861 (N_861,N_787,N_817);
and U862 (N_862,N_810,N_780);
xor U863 (N_863,N_832,N_781);
nand U864 (N_864,N_782,N_804);
and U865 (N_865,N_794,N_799);
nand U866 (N_866,N_789,N_824);
or U867 (N_867,N_792,N_819);
nor U868 (N_868,N_831,N_809);
and U869 (N_869,N_822,N_823);
nor U870 (N_870,N_782,N_818);
and U871 (N_871,N_784,N_838);
nand U872 (N_872,N_816,N_803);
nor U873 (N_873,N_808,N_784);
nor U874 (N_874,N_838,N_830);
nor U875 (N_875,N_802,N_823);
and U876 (N_876,N_829,N_796);
and U877 (N_877,N_821,N_788);
or U878 (N_878,N_786,N_830);
nand U879 (N_879,N_806,N_788);
and U880 (N_880,N_825,N_808);
or U881 (N_881,N_791,N_785);
nor U882 (N_882,N_782,N_825);
nor U883 (N_883,N_808,N_837);
and U884 (N_884,N_793,N_836);
or U885 (N_885,N_831,N_814);
or U886 (N_886,N_802,N_833);
and U887 (N_887,N_837,N_824);
and U888 (N_888,N_831,N_782);
or U889 (N_889,N_838,N_828);
and U890 (N_890,N_785,N_799);
nor U891 (N_891,N_786,N_815);
nor U892 (N_892,N_795,N_812);
or U893 (N_893,N_800,N_833);
nand U894 (N_894,N_783,N_801);
and U895 (N_895,N_837,N_832);
and U896 (N_896,N_801,N_790);
nand U897 (N_897,N_799,N_807);
nor U898 (N_898,N_831,N_794);
or U899 (N_899,N_782,N_827);
nand U900 (N_900,N_888,N_841);
and U901 (N_901,N_855,N_897);
and U902 (N_902,N_866,N_850);
nor U903 (N_903,N_886,N_842);
or U904 (N_904,N_843,N_880);
and U905 (N_905,N_868,N_858);
nand U906 (N_906,N_857,N_859);
nor U907 (N_907,N_863,N_899);
nand U908 (N_908,N_860,N_882);
and U909 (N_909,N_867,N_878);
nand U910 (N_910,N_851,N_847);
and U911 (N_911,N_890,N_877);
or U912 (N_912,N_865,N_876);
and U913 (N_913,N_854,N_870);
and U914 (N_914,N_889,N_864);
and U915 (N_915,N_856,N_892);
or U916 (N_916,N_884,N_873);
nand U917 (N_917,N_872,N_879);
or U918 (N_918,N_893,N_848);
nor U919 (N_919,N_845,N_883);
nand U920 (N_920,N_891,N_894);
or U921 (N_921,N_896,N_869);
nor U922 (N_922,N_887,N_875);
nor U923 (N_923,N_874,N_895);
and U924 (N_924,N_853,N_840);
nand U925 (N_925,N_844,N_871);
and U926 (N_926,N_849,N_885);
and U927 (N_927,N_862,N_846);
xnor U928 (N_928,N_881,N_861);
nand U929 (N_929,N_852,N_898);
and U930 (N_930,N_853,N_848);
nor U931 (N_931,N_883,N_886);
nand U932 (N_932,N_878,N_850);
nor U933 (N_933,N_867,N_880);
nand U934 (N_934,N_860,N_867);
and U935 (N_935,N_883,N_856);
nor U936 (N_936,N_873,N_850);
nor U937 (N_937,N_879,N_883);
nor U938 (N_938,N_869,N_844);
or U939 (N_939,N_883,N_887);
or U940 (N_940,N_887,N_873);
nand U941 (N_941,N_857,N_853);
xnor U942 (N_942,N_861,N_898);
nor U943 (N_943,N_891,N_867);
nor U944 (N_944,N_867,N_881);
nand U945 (N_945,N_862,N_882);
nor U946 (N_946,N_850,N_879);
nand U947 (N_947,N_847,N_870);
nand U948 (N_948,N_885,N_865);
and U949 (N_949,N_864,N_859);
nor U950 (N_950,N_878,N_887);
or U951 (N_951,N_869,N_852);
and U952 (N_952,N_860,N_864);
nand U953 (N_953,N_871,N_854);
nor U954 (N_954,N_890,N_843);
nand U955 (N_955,N_897,N_841);
and U956 (N_956,N_847,N_886);
nand U957 (N_957,N_853,N_897);
nand U958 (N_958,N_899,N_874);
nor U959 (N_959,N_883,N_858);
and U960 (N_960,N_956,N_915);
nor U961 (N_961,N_906,N_942);
and U962 (N_962,N_924,N_918);
or U963 (N_963,N_957,N_903);
nand U964 (N_964,N_921,N_949);
or U965 (N_965,N_940,N_913);
nand U966 (N_966,N_948,N_955);
nor U967 (N_967,N_925,N_900);
nor U968 (N_968,N_926,N_919);
xor U969 (N_969,N_945,N_954);
nor U970 (N_970,N_930,N_905);
nor U971 (N_971,N_941,N_908);
or U972 (N_972,N_909,N_914);
nand U973 (N_973,N_953,N_904);
nand U974 (N_974,N_950,N_936);
nor U975 (N_975,N_928,N_920);
and U976 (N_976,N_927,N_951);
or U977 (N_977,N_933,N_937);
or U978 (N_978,N_917,N_902);
and U979 (N_979,N_944,N_938);
and U980 (N_980,N_910,N_907);
or U981 (N_981,N_923,N_934);
or U982 (N_982,N_959,N_935);
nor U983 (N_983,N_931,N_911);
and U984 (N_984,N_922,N_952);
nor U985 (N_985,N_943,N_901);
and U986 (N_986,N_958,N_912);
and U987 (N_987,N_947,N_939);
and U988 (N_988,N_929,N_946);
or U989 (N_989,N_916,N_932);
or U990 (N_990,N_919,N_933);
and U991 (N_991,N_907,N_905);
or U992 (N_992,N_956,N_937);
or U993 (N_993,N_907,N_927);
xnor U994 (N_994,N_914,N_923);
or U995 (N_995,N_936,N_955);
or U996 (N_996,N_930,N_912);
and U997 (N_997,N_903,N_958);
or U998 (N_998,N_907,N_912);
nand U999 (N_999,N_942,N_941);
and U1000 (N_1000,N_957,N_947);
and U1001 (N_1001,N_922,N_932);
or U1002 (N_1002,N_903,N_944);
nand U1003 (N_1003,N_942,N_937);
nor U1004 (N_1004,N_926,N_942);
nand U1005 (N_1005,N_924,N_957);
and U1006 (N_1006,N_900,N_915);
nand U1007 (N_1007,N_956,N_959);
nor U1008 (N_1008,N_915,N_919);
and U1009 (N_1009,N_903,N_919);
nor U1010 (N_1010,N_928,N_935);
or U1011 (N_1011,N_917,N_910);
or U1012 (N_1012,N_939,N_932);
nor U1013 (N_1013,N_953,N_941);
nand U1014 (N_1014,N_935,N_912);
nand U1015 (N_1015,N_928,N_958);
nand U1016 (N_1016,N_934,N_938);
nor U1017 (N_1017,N_941,N_948);
and U1018 (N_1018,N_926,N_921);
nor U1019 (N_1019,N_911,N_953);
and U1020 (N_1020,N_985,N_1004);
and U1021 (N_1021,N_1014,N_1015);
and U1022 (N_1022,N_1008,N_1002);
nor U1023 (N_1023,N_988,N_995);
nor U1024 (N_1024,N_983,N_981);
or U1025 (N_1025,N_1013,N_1010);
and U1026 (N_1026,N_979,N_976);
nor U1027 (N_1027,N_964,N_1003);
or U1028 (N_1028,N_998,N_960);
and U1029 (N_1029,N_963,N_962);
and U1030 (N_1030,N_1009,N_975);
or U1031 (N_1031,N_980,N_994);
or U1032 (N_1032,N_987,N_1000);
or U1033 (N_1033,N_961,N_1018);
nor U1034 (N_1034,N_973,N_1019);
and U1035 (N_1035,N_990,N_966);
nor U1036 (N_1036,N_986,N_1011);
nand U1037 (N_1037,N_1006,N_974);
or U1038 (N_1038,N_997,N_971);
and U1039 (N_1039,N_968,N_991);
nand U1040 (N_1040,N_1017,N_982);
nand U1041 (N_1041,N_967,N_1012);
nand U1042 (N_1042,N_978,N_1005);
or U1043 (N_1043,N_969,N_999);
xnor U1044 (N_1044,N_992,N_1016);
or U1045 (N_1045,N_996,N_965);
or U1046 (N_1046,N_989,N_984);
and U1047 (N_1047,N_972,N_993);
nand U1048 (N_1048,N_970,N_1001);
nor U1049 (N_1049,N_977,N_1007);
nand U1050 (N_1050,N_983,N_1013);
nor U1051 (N_1051,N_975,N_1011);
and U1052 (N_1052,N_967,N_979);
nand U1053 (N_1053,N_991,N_975);
nand U1054 (N_1054,N_997,N_1012);
nand U1055 (N_1055,N_979,N_1019);
and U1056 (N_1056,N_994,N_1008);
nor U1057 (N_1057,N_992,N_994);
or U1058 (N_1058,N_960,N_966);
and U1059 (N_1059,N_1005,N_995);
or U1060 (N_1060,N_1013,N_985);
nor U1061 (N_1061,N_984,N_1003);
nand U1062 (N_1062,N_990,N_1004);
or U1063 (N_1063,N_963,N_1018);
nor U1064 (N_1064,N_1016,N_977);
or U1065 (N_1065,N_973,N_994);
or U1066 (N_1066,N_1019,N_997);
and U1067 (N_1067,N_1018,N_1015);
or U1068 (N_1068,N_961,N_982);
nor U1069 (N_1069,N_1013,N_992);
or U1070 (N_1070,N_1015,N_996);
or U1071 (N_1071,N_990,N_993);
nor U1072 (N_1072,N_990,N_1016);
or U1073 (N_1073,N_993,N_962);
nand U1074 (N_1074,N_989,N_985);
or U1075 (N_1075,N_973,N_981);
and U1076 (N_1076,N_964,N_1005);
nor U1077 (N_1077,N_990,N_960);
nor U1078 (N_1078,N_961,N_991);
nand U1079 (N_1079,N_962,N_1003);
nand U1080 (N_1080,N_1026,N_1049);
or U1081 (N_1081,N_1028,N_1052);
xor U1082 (N_1082,N_1065,N_1033);
nor U1083 (N_1083,N_1050,N_1072);
nor U1084 (N_1084,N_1022,N_1066);
or U1085 (N_1085,N_1043,N_1035);
or U1086 (N_1086,N_1039,N_1031);
and U1087 (N_1087,N_1056,N_1078);
nand U1088 (N_1088,N_1063,N_1038);
or U1089 (N_1089,N_1070,N_1057);
nand U1090 (N_1090,N_1047,N_1067);
xor U1091 (N_1091,N_1046,N_1079);
or U1092 (N_1092,N_1069,N_1025);
nand U1093 (N_1093,N_1045,N_1062);
or U1094 (N_1094,N_1053,N_1020);
nor U1095 (N_1095,N_1023,N_1029);
nand U1096 (N_1096,N_1034,N_1077);
nand U1097 (N_1097,N_1073,N_1061);
nand U1098 (N_1098,N_1048,N_1051);
nand U1099 (N_1099,N_1054,N_1071);
nor U1100 (N_1100,N_1068,N_1074);
nor U1101 (N_1101,N_1060,N_1032);
nand U1102 (N_1102,N_1042,N_1024);
or U1103 (N_1103,N_1021,N_1075);
nand U1104 (N_1104,N_1064,N_1040);
and U1105 (N_1105,N_1030,N_1058);
or U1106 (N_1106,N_1036,N_1076);
nor U1107 (N_1107,N_1027,N_1041);
nand U1108 (N_1108,N_1037,N_1059);
nor U1109 (N_1109,N_1044,N_1055);
nor U1110 (N_1110,N_1069,N_1056);
nand U1111 (N_1111,N_1040,N_1045);
or U1112 (N_1112,N_1025,N_1071);
or U1113 (N_1113,N_1069,N_1043);
nand U1114 (N_1114,N_1022,N_1068);
and U1115 (N_1115,N_1074,N_1056);
nand U1116 (N_1116,N_1074,N_1070);
and U1117 (N_1117,N_1035,N_1037);
xor U1118 (N_1118,N_1060,N_1059);
or U1119 (N_1119,N_1032,N_1061);
nand U1120 (N_1120,N_1056,N_1031);
and U1121 (N_1121,N_1034,N_1037);
nor U1122 (N_1122,N_1068,N_1041);
nand U1123 (N_1123,N_1064,N_1028);
or U1124 (N_1124,N_1057,N_1024);
nand U1125 (N_1125,N_1044,N_1051);
and U1126 (N_1126,N_1066,N_1078);
nand U1127 (N_1127,N_1023,N_1041);
nand U1128 (N_1128,N_1055,N_1035);
xor U1129 (N_1129,N_1050,N_1078);
nor U1130 (N_1130,N_1076,N_1024);
nor U1131 (N_1131,N_1037,N_1048);
and U1132 (N_1132,N_1075,N_1061);
and U1133 (N_1133,N_1071,N_1026);
xnor U1134 (N_1134,N_1055,N_1020);
nand U1135 (N_1135,N_1020,N_1070);
nor U1136 (N_1136,N_1027,N_1070);
nand U1137 (N_1137,N_1056,N_1043);
or U1138 (N_1138,N_1075,N_1066);
nand U1139 (N_1139,N_1061,N_1040);
or U1140 (N_1140,N_1137,N_1085);
or U1141 (N_1141,N_1098,N_1122);
nand U1142 (N_1142,N_1103,N_1101);
nor U1143 (N_1143,N_1084,N_1081);
nand U1144 (N_1144,N_1131,N_1086);
and U1145 (N_1145,N_1132,N_1094);
nor U1146 (N_1146,N_1092,N_1129);
and U1147 (N_1147,N_1093,N_1100);
nand U1148 (N_1148,N_1134,N_1126);
or U1149 (N_1149,N_1138,N_1091);
or U1150 (N_1150,N_1120,N_1115);
nand U1151 (N_1151,N_1121,N_1107);
nor U1152 (N_1152,N_1112,N_1125);
nand U1153 (N_1153,N_1109,N_1108);
and U1154 (N_1154,N_1139,N_1136);
nand U1155 (N_1155,N_1135,N_1111);
nor U1156 (N_1156,N_1114,N_1097);
or U1157 (N_1157,N_1095,N_1105);
and U1158 (N_1158,N_1102,N_1128);
or U1159 (N_1159,N_1089,N_1123);
or U1160 (N_1160,N_1082,N_1116);
or U1161 (N_1161,N_1106,N_1117);
nor U1162 (N_1162,N_1080,N_1088);
nand U1163 (N_1163,N_1130,N_1090);
nand U1164 (N_1164,N_1133,N_1104);
and U1165 (N_1165,N_1110,N_1118);
nor U1166 (N_1166,N_1124,N_1127);
and U1167 (N_1167,N_1119,N_1083);
and U1168 (N_1168,N_1099,N_1113);
and U1169 (N_1169,N_1087,N_1096);
and U1170 (N_1170,N_1133,N_1103);
nand U1171 (N_1171,N_1087,N_1126);
and U1172 (N_1172,N_1082,N_1137);
or U1173 (N_1173,N_1093,N_1119);
or U1174 (N_1174,N_1106,N_1136);
and U1175 (N_1175,N_1111,N_1102);
or U1176 (N_1176,N_1134,N_1100);
and U1177 (N_1177,N_1109,N_1131);
nand U1178 (N_1178,N_1095,N_1127);
nand U1179 (N_1179,N_1127,N_1122);
and U1180 (N_1180,N_1101,N_1095);
nand U1181 (N_1181,N_1101,N_1127);
nor U1182 (N_1182,N_1124,N_1082);
nor U1183 (N_1183,N_1083,N_1114);
nor U1184 (N_1184,N_1111,N_1112);
and U1185 (N_1185,N_1138,N_1094);
and U1186 (N_1186,N_1084,N_1116);
nand U1187 (N_1187,N_1080,N_1082);
nor U1188 (N_1188,N_1115,N_1099);
xnor U1189 (N_1189,N_1104,N_1121);
nor U1190 (N_1190,N_1092,N_1100);
and U1191 (N_1191,N_1122,N_1138);
nand U1192 (N_1192,N_1082,N_1139);
nor U1193 (N_1193,N_1110,N_1098);
and U1194 (N_1194,N_1131,N_1125);
or U1195 (N_1195,N_1107,N_1129);
nor U1196 (N_1196,N_1098,N_1119);
or U1197 (N_1197,N_1117,N_1088);
or U1198 (N_1198,N_1086,N_1094);
nand U1199 (N_1199,N_1121,N_1099);
xor U1200 (N_1200,N_1198,N_1189);
nand U1201 (N_1201,N_1163,N_1181);
nor U1202 (N_1202,N_1162,N_1141);
nand U1203 (N_1203,N_1153,N_1157);
and U1204 (N_1204,N_1151,N_1185);
and U1205 (N_1205,N_1146,N_1197);
nor U1206 (N_1206,N_1168,N_1186);
nor U1207 (N_1207,N_1193,N_1194);
and U1208 (N_1208,N_1145,N_1173);
nor U1209 (N_1209,N_1158,N_1142);
nor U1210 (N_1210,N_1192,N_1161);
nand U1211 (N_1211,N_1195,N_1171);
and U1212 (N_1212,N_1179,N_1172);
nand U1213 (N_1213,N_1174,N_1150);
or U1214 (N_1214,N_1159,N_1154);
or U1215 (N_1215,N_1143,N_1188);
nand U1216 (N_1216,N_1175,N_1182);
nand U1217 (N_1217,N_1155,N_1183);
nand U1218 (N_1218,N_1140,N_1170);
nand U1219 (N_1219,N_1191,N_1187);
nor U1220 (N_1220,N_1180,N_1166);
nand U1221 (N_1221,N_1169,N_1144);
nor U1222 (N_1222,N_1149,N_1178);
nand U1223 (N_1223,N_1176,N_1152);
nand U1224 (N_1224,N_1184,N_1148);
nor U1225 (N_1225,N_1165,N_1199);
nor U1226 (N_1226,N_1164,N_1160);
nand U1227 (N_1227,N_1156,N_1177);
xor U1228 (N_1228,N_1167,N_1196);
or U1229 (N_1229,N_1190,N_1147);
nor U1230 (N_1230,N_1180,N_1175);
nand U1231 (N_1231,N_1157,N_1181);
or U1232 (N_1232,N_1183,N_1161);
nor U1233 (N_1233,N_1185,N_1148);
nand U1234 (N_1234,N_1177,N_1166);
nand U1235 (N_1235,N_1150,N_1143);
nor U1236 (N_1236,N_1140,N_1167);
xor U1237 (N_1237,N_1195,N_1142);
or U1238 (N_1238,N_1168,N_1145);
nand U1239 (N_1239,N_1188,N_1168);
nand U1240 (N_1240,N_1140,N_1166);
nand U1241 (N_1241,N_1156,N_1168);
nand U1242 (N_1242,N_1150,N_1167);
or U1243 (N_1243,N_1148,N_1162);
nand U1244 (N_1244,N_1166,N_1157);
nor U1245 (N_1245,N_1195,N_1176);
or U1246 (N_1246,N_1172,N_1141);
and U1247 (N_1247,N_1193,N_1183);
nand U1248 (N_1248,N_1144,N_1152);
and U1249 (N_1249,N_1190,N_1143);
nand U1250 (N_1250,N_1174,N_1167);
nand U1251 (N_1251,N_1195,N_1198);
nor U1252 (N_1252,N_1165,N_1198);
nand U1253 (N_1253,N_1183,N_1176);
nor U1254 (N_1254,N_1197,N_1182);
or U1255 (N_1255,N_1161,N_1151);
and U1256 (N_1256,N_1140,N_1175);
nor U1257 (N_1257,N_1190,N_1163);
or U1258 (N_1258,N_1177,N_1155);
nor U1259 (N_1259,N_1155,N_1141);
or U1260 (N_1260,N_1217,N_1240);
nor U1261 (N_1261,N_1225,N_1242);
and U1262 (N_1262,N_1241,N_1235);
nand U1263 (N_1263,N_1256,N_1222);
nand U1264 (N_1264,N_1245,N_1216);
nor U1265 (N_1265,N_1213,N_1239);
nand U1266 (N_1266,N_1211,N_1218);
nand U1267 (N_1267,N_1253,N_1250);
or U1268 (N_1268,N_1238,N_1246);
nand U1269 (N_1269,N_1227,N_1206);
or U1270 (N_1270,N_1237,N_1223);
nor U1271 (N_1271,N_1259,N_1204);
nor U1272 (N_1272,N_1201,N_1251);
or U1273 (N_1273,N_1202,N_1248);
nor U1274 (N_1274,N_1209,N_1249);
nor U1275 (N_1275,N_1255,N_1215);
nor U1276 (N_1276,N_1229,N_1214);
or U1277 (N_1277,N_1212,N_1228);
nor U1278 (N_1278,N_1200,N_1224);
and U1279 (N_1279,N_1226,N_1244);
nand U1280 (N_1280,N_1219,N_1208);
xor U1281 (N_1281,N_1220,N_1203);
nand U1282 (N_1282,N_1236,N_1257);
and U1283 (N_1283,N_1231,N_1254);
and U1284 (N_1284,N_1247,N_1234);
or U1285 (N_1285,N_1230,N_1221);
nand U1286 (N_1286,N_1210,N_1258);
nand U1287 (N_1287,N_1205,N_1207);
and U1288 (N_1288,N_1243,N_1232);
nand U1289 (N_1289,N_1233,N_1252);
and U1290 (N_1290,N_1207,N_1237);
or U1291 (N_1291,N_1255,N_1200);
nand U1292 (N_1292,N_1221,N_1223);
or U1293 (N_1293,N_1228,N_1247);
or U1294 (N_1294,N_1217,N_1242);
or U1295 (N_1295,N_1205,N_1214);
nand U1296 (N_1296,N_1207,N_1256);
nor U1297 (N_1297,N_1234,N_1208);
or U1298 (N_1298,N_1235,N_1239);
nor U1299 (N_1299,N_1258,N_1243);
and U1300 (N_1300,N_1258,N_1225);
nand U1301 (N_1301,N_1237,N_1256);
nor U1302 (N_1302,N_1227,N_1220);
or U1303 (N_1303,N_1206,N_1221);
nand U1304 (N_1304,N_1250,N_1255);
and U1305 (N_1305,N_1226,N_1253);
and U1306 (N_1306,N_1216,N_1252);
or U1307 (N_1307,N_1244,N_1227);
or U1308 (N_1308,N_1239,N_1205);
or U1309 (N_1309,N_1241,N_1212);
and U1310 (N_1310,N_1212,N_1220);
nor U1311 (N_1311,N_1244,N_1245);
and U1312 (N_1312,N_1222,N_1215);
or U1313 (N_1313,N_1213,N_1257);
and U1314 (N_1314,N_1205,N_1248);
nor U1315 (N_1315,N_1246,N_1249);
nand U1316 (N_1316,N_1223,N_1203);
nand U1317 (N_1317,N_1217,N_1215);
nand U1318 (N_1318,N_1215,N_1230);
nor U1319 (N_1319,N_1222,N_1211);
nand U1320 (N_1320,N_1312,N_1292);
nor U1321 (N_1321,N_1293,N_1283);
and U1322 (N_1322,N_1310,N_1260);
and U1323 (N_1323,N_1279,N_1304);
or U1324 (N_1324,N_1269,N_1274);
nor U1325 (N_1325,N_1290,N_1285);
and U1326 (N_1326,N_1300,N_1282);
nand U1327 (N_1327,N_1307,N_1319);
and U1328 (N_1328,N_1275,N_1303);
nor U1329 (N_1329,N_1273,N_1267);
or U1330 (N_1330,N_1264,N_1316);
or U1331 (N_1331,N_1305,N_1296);
and U1332 (N_1332,N_1314,N_1288);
nand U1333 (N_1333,N_1278,N_1263);
nor U1334 (N_1334,N_1271,N_1299);
nand U1335 (N_1335,N_1286,N_1272);
or U1336 (N_1336,N_1281,N_1268);
and U1337 (N_1337,N_1262,N_1291);
or U1338 (N_1338,N_1315,N_1295);
and U1339 (N_1339,N_1302,N_1289);
nor U1340 (N_1340,N_1306,N_1301);
nor U1341 (N_1341,N_1284,N_1308);
nand U1342 (N_1342,N_1270,N_1265);
nand U1343 (N_1343,N_1311,N_1298);
nand U1344 (N_1344,N_1276,N_1297);
xor U1345 (N_1345,N_1309,N_1294);
and U1346 (N_1346,N_1280,N_1277);
nor U1347 (N_1347,N_1287,N_1317);
and U1348 (N_1348,N_1266,N_1313);
and U1349 (N_1349,N_1261,N_1318);
nor U1350 (N_1350,N_1282,N_1315);
nor U1351 (N_1351,N_1312,N_1261);
or U1352 (N_1352,N_1290,N_1295);
or U1353 (N_1353,N_1293,N_1285);
and U1354 (N_1354,N_1305,N_1269);
or U1355 (N_1355,N_1299,N_1287);
nor U1356 (N_1356,N_1307,N_1305);
nor U1357 (N_1357,N_1295,N_1303);
nand U1358 (N_1358,N_1262,N_1310);
and U1359 (N_1359,N_1292,N_1270);
and U1360 (N_1360,N_1263,N_1282);
nor U1361 (N_1361,N_1265,N_1281);
or U1362 (N_1362,N_1295,N_1297);
or U1363 (N_1363,N_1308,N_1314);
or U1364 (N_1364,N_1286,N_1319);
nand U1365 (N_1365,N_1307,N_1302);
or U1366 (N_1366,N_1279,N_1290);
and U1367 (N_1367,N_1274,N_1262);
and U1368 (N_1368,N_1309,N_1301);
or U1369 (N_1369,N_1264,N_1295);
and U1370 (N_1370,N_1261,N_1264);
and U1371 (N_1371,N_1304,N_1299);
nand U1372 (N_1372,N_1267,N_1270);
nand U1373 (N_1373,N_1315,N_1273);
and U1374 (N_1374,N_1281,N_1273);
nor U1375 (N_1375,N_1303,N_1306);
nand U1376 (N_1376,N_1265,N_1286);
or U1377 (N_1377,N_1305,N_1314);
nor U1378 (N_1378,N_1313,N_1278);
or U1379 (N_1379,N_1294,N_1276);
nor U1380 (N_1380,N_1321,N_1329);
nand U1381 (N_1381,N_1326,N_1343);
and U1382 (N_1382,N_1327,N_1324);
and U1383 (N_1383,N_1328,N_1372);
nand U1384 (N_1384,N_1377,N_1338);
and U1385 (N_1385,N_1344,N_1355);
and U1386 (N_1386,N_1369,N_1352);
nand U1387 (N_1387,N_1360,N_1356);
nand U1388 (N_1388,N_1346,N_1363);
and U1389 (N_1389,N_1368,N_1322);
and U1390 (N_1390,N_1374,N_1339);
or U1391 (N_1391,N_1379,N_1337);
nor U1392 (N_1392,N_1342,N_1365);
and U1393 (N_1393,N_1348,N_1323);
nor U1394 (N_1394,N_1341,N_1347);
or U1395 (N_1395,N_1340,N_1345);
and U1396 (N_1396,N_1333,N_1354);
or U1397 (N_1397,N_1362,N_1335);
nor U1398 (N_1398,N_1332,N_1320);
nand U1399 (N_1399,N_1330,N_1361);
nand U1400 (N_1400,N_1366,N_1325);
nor U1401 (N_1401,N_1376,N_1334);
or U1402 (N_1402,N_1367,N_1331);
nor U1403 (N_1403,N_1353,N_1364);
and U1404 (N_1404,N_1371,N_1370);
or U1405 (N_1405,N_1378,N_1375);
or U1406 (N_1406,N_1350,N_1351);
nand U1407 (N_1407,N_1358,N_1349);
and U1408 (N_1408,N_1336,N_1373);
nand U1409 (N_1409,N_1359,N_1357);
nor U1410 (N_1410,N_1349,N_1333);
nor U1411 (N_1411,N_1336,N_1349);
nor U1412 (N_1412,N_1353,N_1322);
and U1413 (N_1413,N_1360,N_1364);
nor U1414 (N_1414,N_1322,N_1347);
nand U1415 (N_1415,N_1331,N_1350);
and U1416 (N_1416,N_1378,N_1358);
or U1417 (N_1417,N_1373,N_1339);
and U1418 (N_1418,N_1376,N_1326);
and U1419 (N_1419,N_1332,N_1340);
nand U1420 (N_1420,N_1372,N_1357);
and U1421 (N_1421,N_1368,N_1328);
nor U1422 (N_1422,N_1343,N_1320);
nand U1423 (N_1423,N_1367,N_1349);
or U1424 (N_1424,N_1373,N_1347);
nor U1425 (N_1425,N_1321,N_1334);
or U1426 (N_1426,N_1354,N_1361);
nand U1427 (N_1427,N_1353,N_1336);
or U1428 (N_1428,N_1336,N_1344);
or U1429 (N_1429,N_1362,N_1357);
nor U1430 (N_1430,N_1322,N_1356);
and U1431 (N_1431,N_1328,N_1337);
and U1432 (N_1432,N_1350,N_1337);
nor U1433 (N_1433,N_1345,N_1338);
or U1434 (N_1434,N_1376,N_1333);
xnor U1435 (N_1435,N_1371,N_1363);
or U1436 (N_1436,N_1320,N_1328);
nand U1437 (N_1437,N_1368,N_1352);
xor U1438 (N_1438,N_1367,N_1355);
or U1439 (N_1439,N_1320,N_1379);
and U1440 (N_1440,N_1385,N_1419);
and U1441 (N_1441,N_1437,N_1427);
and U1442 (N_1442,N_1383,N_1438);
nor U1443 (N_1443,N_1398,N_1411);
nor U1444 (N_1444,N_1414,N_1380);
nand U1445 (N_1445,N_1388,N_1410);
nor U1446 (N_1446,N_1391,N_1404);
nand U1447 (N_1447,N_1409,N_1393);
and U1448 (N_1448,N_1416,N_1406);
and U1449 (N_1449,N_1382,N_1387);
nor U1450 (N_1450,N_1389,N_1426);
nor U1451 (N_1451,N_1407,N_1432);
nor U1452 (N_1452,N_1425,N_1436);
or U1453 (N_1453,N_1433,N_1395);
and U1454 (N_1454,N_1430,N_1423);
xor U1455 (N_1455,N_1421,N_1386);
nor U1456 (N_1456,N_1396,N_1428);
nand U1457 (N_1457,N_1418,N_1399);
or U1458 (N_1458,N_1400,N_1403);
and U1459 (N_1459,N_1381,N_1405);
or U1460 (N_1460,N_1415,N_1408);
nand U1461 (N_1461,N_1435,N_1390);
or U1462 (N_1462,N_1434,N_1439);
and U1463 (N_1463,N_1394,N_1412);
nor U1464 (N_1464,N_1413,N_1420);
and U1465 (N_1465,N_1417,N_1422);
nor U1466 (N_1466,N_1384,N_1431);
nor U1467 (N_1467,N_1402,N_1424);
or U1468 (N_1468,N_1401,N_1429);
and U1469 (N_1469,N_1392,N_1397);
and U1470 (N_1470,N_1434,N_1408);
and U1471 (N_1471,N_1409,N_1433);
nor U1472 (N_1472,N_1420,N_1428);
or U1473 (N_1473,N_1418,N_1413);
nor U1474 (N_1474,N_1405,N_1426);
or U1475 (N_1475,N_1391,N_1398);
nor U1476 (N_1476,N_1395,N_1390);
nor U1477 (N_1477,N_1383,N_1433);
and U1478 (N_1478,N_1407,N_1396);
nor U1479 (N_1479,N_1392,N_1429);
nor U1480 (N_1480,N_1439,N_1389);
nor U1481 (N_1481,N_1403,N_1430);
nand U1482 (N_1482,N_1425,N_1402);
or U1483 (N_1483,N_1427,N_1411);
nor U1484 (N_1484,N_1423,N_1408);
nor U1485 (N_1485,N_1425,N_1411);
or U1486 (N_1486,N_1409,N_1383);
and U1487 (N_1487,N_1436,N_1424);
xor U1488 (N_1488,N_1414,N_1400);
or U1489 (N_1489,N_1400,N_1382);
or U1490 (N_1490,N_1394,N_1433);
and U1491 (N_1491,N_1392,N_1418);
or U1492 (N_1492,N_1397,N_1438);
nand U1493 (N_1493,N_1421,N_1388);
and U1494 (N_1494,N_1436,N_1389);
and U1495 (N_1495,N_1439,N_1401);
and U1496 (N_1496,N_1425,N_1393);
or U1497 (N_1497,N_1400,N_1397);
nor U1498 (N_1498,N_1384,N_1382);
nor U1499 (N_1499,N_1382,N_1437);
or U1500 (N_1500,N_1498,N_1480);
nor U1501 (N_1501,N_1476,N_1453);
or U1502 (N_1502,N_1458,N_1462);
and U1503 (N_1503,N_1471,N_1444);
nand U1504 (N_1504,N_1446,N_1455);
nand U1505 (N_1505,N_1489,N_1443);
and U1506 (N_1506,N_1497,N_1452);
and U1507 (N_1507,N_1495,N_1461);
nor U1508 (N_1508,N_1445,N_1459);
and U1509 (N_1509,N_1457,N_1463);
nand U1510 (N_1510,N_1491,N_1440);
or U1511 (N_1511,N_1487,N_1468);
nand U1512 (N_1512,N_1451,N_1466);
or U1513 (N_1513,N_1470,N_1441);
or U1514 (N_1514,N_1479,N_1493);
nor U1515 (N_1515,N_1464,N_1472);
and U1516 (N_1516,N_1499,N_1469);
or U1517 (N_1517,N_1454,N_1465);
and U1518 (N_1518,N_1484,N_1478);
or U1519 (N_1519,N_1473,N_1442);
or U1520 (N_1520,N_1482,N_1475);
nand U1521 (N_1521,N_1481,N_1456);
xnor U1522 (N_1522,N_1494,N_1488);
nand U1523 (N_1523,N_1492,N_1449);
and U1524 (N_1524,N_1496,N_1448);
and U1525 (N_1525,N_1477,N_1474);
and U1526 (N_1526,N_1483,N_1486);
or U1527 (N_1527,N_1447,N_1450);
nor U1528 (N_1528,N_1485,N_1467);
and U1529 (N_1529,N_1460,N_1490);
and U1530 (N_1530,N_1468,N_1477);
or U1531 (N_1531,N_1460,N_1497);
and U1532 (N_1532,N_1499,N_1470);
nor U1533 (N_1533,N_1493,N_1459);
nand U1534 (N_1534,N_1474,N_1471);
or U1535 (N_1535,N_1490,N_1467);
nand U1536 (N_1536,N_1487,N_1481);
nand U1537 (N_1537,N_1480,N_1449);
and U1538 (N_1538,N_1491,N_1495);
nor U1539 (N_1539,N_1488,N_1466);
nor U1540 (N_1540,N_1451,N_1481);
or U1541 (N_1541,N_1484,N_1477);
nor U1542 (N_1542,N_1496,N_1445);
and U1543 (N_1543,N_1442,N_1468);
or U1544 (N_1544,N_1463,N_1454);
nor U1545 (N_1545,N_1482,N_1483);
and U1546 (N_1546,N_1467,N_1471);
nor U1547 (N_1547,N_1481,N_1440);
or U1548 (N_1548,N_1491,N_1443);
nand U1549 (N_1549,N_1487,N_1459);
or U1550 (N_1550,N_1480,N_1445);
and U1551 (N_1551,N_1480,N_1490);
nand U1552 (N_1552,N_1475,N_1486);
xnor U1553 (N_1553,N_1446,N_1440);
and U1554 (N_1554,N_1482,N_1457);
and U1555 (N_1555,N_1450,N_1440);
or U1556 (N_1556,N_1462,N_1440);
nand U1557 (N_1557,N_1485,N_1488);
nand U1558 (N_1558,N_1453,N_1471);
or U1559 (N_1559,N_1486,N_1474);
and U1560 (N_1560,N_1532,N_1554);
nor U1561 (N_1561,N_1521,N_1550);
nand U1562 (N_1562,N_1553,N_1530);
nand U1563 (N_1563,N_1557,N_1534);
and U1564 (N_1564,N_1549,N_1515);
nor U1565 (N_1565,N_1537,N_1503);
or U1566 (N_1566,N_1502,N_1551);
and U1567 (N_1567,N_1512,N_1509);
or U1568 (N_1568,N_1559,N_1522);
nor U1569 (N_1569,N_1505,N_1533);
nor U1570 (N_1570,N_1519,N_1548);
and U1571 (N_1571,N_1523,N_1542);
and U1572 (N_1572,N_1501,N_1544);
or U1573 (N_1573,N_1508,N_1526);
nand U1574 (N_1574,N_1524,N_1514);
or U1575 (N_1575,N_1535,N_1536);
or U1576 (N_1576,N_1507,N_1500);
or U1577 (N_1577,N_1541,N_1506);
nand U1578 (N_1578,N_1552,N_1527);
xnor U1579 (N_1579,N_1520,N_1518);
xor U1580 (N_1580,N_1517,N_1529);
nand U1581 (N_1581,N_1525,N_1510);
nand U1582 (N_1582,N_1555,N_1558);
or U1583 (N_1583,N_1531,N_1538);
or U1584 (N_1584,N_1556,N_1543);
or U1585 (N_1585,N_1511,N_1545);
or U1586 (N_1586,N_1539,N_1513);
nand U1587 (N_1587,N_1547,N_1528);
and U1588 (N_1588,N_1540,N_1546);
nor U1589 (N_1589,N_1516,N_1504);
nor U1590 (N_1590,N_1547,N_1537);
nor U1591 (N_1591,N_1542,N_1551);
or U1592 (N_1592,N_1512,N_1501);
nor U1593 (N_1593,N_1513,N_1507);
or U1594 (N_1594,N_1513,N_1524);
or U1595 (N_1595,N_1540,N_1550);
or U1596 (N_1596,N_1509,N_1534);
and U1597 (N_1597,N_1534,N_1537);
and U1598 (N_1598,N_1509,N_1520);
and U1599 (N_1599,N_1524,N_1516);
or U1600 (N_1600,N_1516,N_1525);
nand U1601 (N_1601,N_1544,N_1555);
and U1602 (N_1602,N_1524,N_1543);
nor U1603 (N_1603,N_1559,N_1557);
nand U1604 (N_1604,N_1541,N_1527);
or U1605 (N_1605,N_1528,N_1537);
or U1606 (N_1606,N_1505,N_1542);
or U1607 (N_1607,N_1535,N_1546);
and U1608 (N_1608,N_1549,N_1520);
nor U1609 (N_1609,N_1530,N_1532);
nand U1610 (N_1610,N_1512,N_1542);
or U1611 (N_1611,N_1538,N_1534);
nand U1612 (N_1612,N_1515,N_1533);
nor U1613 (N_1613,N_1555,N_1522);
and U1614 (N_1614,N_1538,N_1541);
nand U1615 (N_1615,N_1504,N_1515);
nor U1616 (N_1616,N_1550,N_1541);
nor U1617 (N_1617,N_1519,N_1533);
or U1618 (N_1618,N_1500,N_1514);
or U1619 (N_1619,N_1517,N_1536);
or U1620 (N_1620,N_1573,N_1568);
and U1621 (N_1621,N_1561,N_1564);
nor U1622 (N_1622,N_1604,N_1563);
nor U1623 (N_1623,N_1565,N_1574);
nand U1624 (N_1624,N_1577,N_1562);
and U1625 (N_1625,N_1617,N_1609);
or U1626 (N_1626,N_1606,N_1592);
nor U1627 (N_1627,N_1612,N_1608);
xor U1628 (N_1628,N_1580,N_1581);
nand U1629 (N_1629,N_1582,N_1570);
and U1630 (N_1630,N_1616,N_1590);
or U1631 (N_1631,N_1560,N_1584);
or U1632 (N_1632,N_1578,N_1615);
nand U1633 (N_1633,N_1589,N_1610);
nand U1634 (N_1634,N_1593,N_1607);
and U1635 (N_1635,N_1569,N_1600);
nand U1636 (N_1636,N_1619,N_1572);
or U1637 (N_1637,N_1603,N_1583);
nor U1638 (N_1638,N_1614,N_1576);
or U1639 (N_1639,N_1596,N_1585);
and U1640 (N_1640,N_1611,N_1571);
and U1641 (N_1641,N_1588,N_1598);
and U1642 (N_1642,N_1567,N_1605);
nor U1643 (N_1643,N_1594,N_1613);
nor U1644 (N_1644,N_1575,N_1587);
nor U1645 (N_1645,N_1601,N_1599);
or U1646 (N_1646,N_1579,N_1618);
nor U1647 (N_1647,N_1591,N_1602);
nand U1648 (N_1648,N_1586,N_1597);
nand U1649 (N_1649,N_1595,N_1566);
nand U1650 (N_1650,N_1580,N_1577);
or U1651 (N_1651,N_1569,N_1606);
or U1652 (N_1652,N_1608,N_1602);
nand U1653 (N_1653,N_1604,N_1608);
or U1654 (N_1654,N_1613,N_1607);
and U1655 (N_1655,N_1615,N_1619);
or U1656 (N_1656,N_1608,N_1598);
nor U1657 (N_1657,N_1572,N_1586);
nand U1658 (N_1658,N_1618,N_1596);
nand U1659 (N_1659,N_1590,N_1611);
and U1660 (N_1660,N_1617,N_1598);
nand U1661 (N_1661,N_1606,N_1567);
xor U1662 (N_1662,N_1587,N_1608);
or U1663 (N_1663,N_1603,N_1582);
nor U1664 (N_1664,N_1564,N_1574);
nor U1665 (N_1665,N_1585,N_1562);
and U1666 (N_1666,N_1614,N_1570);
nand U1667 (N_1667,N_1575,N_1617);
nand U1668 (N_1668,N_1582,N_1566);
nand U1669 (N_1669,N_1591,N_1612);
nor U1670 (N_1670,N_1613,N_1574);
nor U1671 (N_1671,N_1605,N_1584);
nand U1672 (N_1672,N_1560,N_1606);
and U1673 (N_1673,N_1594,N_1595);
or U1674 (N_1674,N_1573,N_1601);
nor U1675 (N_1675,N_1573,N_1572);
nand U1676 (N_1676,N_1609,N_1577);
nand U1677 (N_1677,N_1585,N_1593);
or U1678 (N_1678,N_1568,N_1570);
nor U1679 (N_1679,N_1594,N_1602);
nand U1680 (N_1680,N_1642,N_1641);
or U1681 (N_1681,N_1652,N_1629);
and U1682 (N_1682,N_1644,N_1670);
nand U1683 (N_1683,N_1653,N_1655);
and U1684 (N_1684,N_1654,N_1672);
or U1685 (N_1685,N_1669,N_1668);
or U1686 (N_1686,N_1648,N_1678);
or U1687 (N_1687,N_1664,N_1646);
and U1688 (N_1688,N_1650,N_1625);
nand U1689 (N_1689,N_1639,N_1626);
or U1690 (N_1690,N_1636,N_1647);
and U1691 (N_1691,N_1643,N_1675);
and U1692 (N_1692,N_1631,N_1656);
nand U1693 (N_1693,N_1637,N_1661);
nor U1694 (N_1694,N_1640,N_1665);
nand U1695 (N_1695,N_1658,N_1624);
and U1696 (N_1696,N_1679,N_1621);
and U1697 (N_1697,N_1666,N_1663);
nand U1698 (N_1698,N_1676,N_1635);
nor U1699 (N_1699,N_1638,N_1627);
nor U1700 (N_1700,N_1628,N_1671);
nor U1701 (N_1701,N_1657,N_1662);
nand U1702 (N_1702,N_1677,N_1651);
nand U1703 (N_1703,N_1630,N_1667);
nor U1704 (N_1704,N_1623,N_1674);
nor U1705 (N_1705,N_1659,N_1649);
nand U1706 (N_1706,N_1632,N_1622);
or U1707 (N_1707,N_1620,N_1634);
or U1708 (N_1708,N_1633,N_1673);
nand U1709 (N_1709,N_1660,N_1645);
or U1710 (N_1710,N_1652,N_1654);
or U1711 (N_1711,N_1621,N_1649);
and U1712 (N_1712,N_1621,N_1677);
nand U1713 (N_1713,N_1666,N_1650);
nor U1714 (N_1714,N_1648,N_1650);
and U1715 (N_1715,N_1638,N_1634);
or U1716 (N_1716,N_1664,N_1653);
and U1717 (N_1717,N_1642,N_1649);
or U1718 (N_1718,N_1652,N_1647);
and U1719 (N_1719,N_1660,N_1634);
and U1720 (N_1720,N_1647,N_1640);
or U1721 (N_1721,N_1640,N_1622);
nor U1722 (N_1722,N_1645,N_1666);
and U1723 (N_1723,N_1646,N_1677);
or U1724 (N_1724,N_1645,N_1642);
nand U1725 (N_1725,N_1620,N_1671);
nor U1726 (N_1726,N_1635,N_1638);
and U1727 (N_1727,N_1677,N_1673);
nor U1728 (N_1728,N_1673,N_1639);
nor U1729 (N_1729,N_1629,N_1648);
or U1730 (N_1730,N_1630,N_1620);
and U1731 (N_1731,N_1626,N_1656);
nor U1732 (N_1732,N_1652,N_1648);
or U1733 (N_1733,N_1661,N_1657);
and U1734 (N_1734,N_1660,N_1676);
nor U1735 (N_1735,N_1650,N_1645);
or U1736 (N_1736,N_1658,N_1636);
and U1737 (N_1737,N_1622,N_1676);
or U1738 (N_1738,N_1667,N_1623);
or U1739 (N_1739,N_1633,N_1664);
nor U1740 (N_1740,N_1736,N_1686);
or U1741 (N_1741,N_1726,N_1734);
and U1742 (N_1742,N_1709,N_1728);
nor U1743 (N_1743,N_1720,N_1702);
and U1744 (N_1744,N_1713,N_1699);
or U1745 (N_1745,N_1717,N_1681);
nor U1746 (N_1746,N_1682,N_1691);
or U1747 (N_1747,N_1707,N_1706);
and U1748 (N_1748,N_1724,N_1733);
or U1749 (N_1749,N_1687,N_1695);
nor U1750 (N_1750,N_1730,N_1737);
or U1751 (N_1751,N_1732,N_1692);
nor U1752 (N_1752,N_1708,N_1731);
nor U1753 (N_1753,N_1716,N_1684);
nor U1754 (N_1754,N_1738,N_1722);
or U1755 (N_1755,N_1711,N_1694);
or U1756 (N_1756,N_1685,N_1700);
or U1757 (N_1757,N_1683,N_1698);
nand U1758 (N_1758,N_1727,N_1721);
or U1759 (N_1759,N_1725,N_1719);
xnor U1760 (N_1760,N_1715,N_1735);
or U1761 (N_1761,N_1701,N_1697);
and U1762 (N_1762,N_1718,N_1712);
or U1763 (N_1763,N_1703,N_1688);
and U1764 (N_1764,N_1710,N_1739);
or U1765 (N_1765,N_1680,N_1689);
and U1766 (N_1766,N_1696,N_1723);
and U1767 (N_1767,N_1690,N_1704);
nand U1768 (N_1768,N_1729,N_1705);
nand U1769 (N_1769,N_1714,N_1693);
xnor U1770 (N_1770,N_1690,N_1705);
or U1771 (N_1771,N_1723,N_1694);
nor U1772 (N_1772,N_1716,N_1714);
or U1773 (N_1773,N_1702,N_1693);
nor U1774 (N_1774,N_1733,N_1680);
and U1775 (N_1775,N_1683,N_1729);
and U1776 (N_1776,N_1717,N_1720);
and U1777 (N_1777,N_1680,N_1724);
or U1778 (N_1778,N_1738,N_1719);
and U1779 (N_1779,N_1712,N_1723);
nand U1780 (N_1780,N_1709,N_1731);
nand U1781 (N_1781,N_1709,N_1714);
nor U1782 (N_1782,N_1709,N_1716);
nand U1783 (N_1783,N_1684,N_1715);
nor U1784 (N_1784,N_1705,N_1698);
and U1785 (N_1785,N_1724,N_1732);
nor U1786 (N_1786,N_1738,N_1696);
or U1787 (N_1787,N_1735,N_1734);
nand U1788 (N_1788,N_1696,N_1718);
nand U1789 (N_1789,N_1688,N_1717);
and U1790 (N_1790,N_1732,N_1731);
nand U1791 (N_1791,N_1728,N_1694);
or U1792 (N_1792,N_1680,N_1716);
nor U1793 (N_1793,N_1721,N_1695);
xnor U1794 (N_1794,N_1716,N_1733);
or U1795 (N_1795,N_1720,N_1727);
and U1796 (N_1796,N_1698,N_1716);
and U1797 (N_1797,N_1688,N_1683);
nor U1798 (N_1798,N_1687,N_1688);
nor U1799 (N_1799,N_1727,N_1703);
xnor U1800 (N_1800,N_1788,N_1774);
nor U1801 (N_1801,N_1741,N_1752);
and U1802 (N_1802,N_1775,N_1765);
nor U1803 (N_1803,N_1777,N_1763);
or U1804 (N_1804,N_1780,N_1785);
nor U1805 (N_1805,N_1745,N_1767);
nor U1806 (N_1806,N_1772,N_1766);
nor U1807 (N_1807,N_1764,N_1793);
nand U1808 (N_1808,N_1799,N_1757);
and U1809 (N_1809,N_1753,N_1787);
nand U1810 (N_1810,N_1798,N_1743);
xor U1811 (N_1811,N_1778,N_1789);
nor U1812 (N_1812,N_1794,N_1756);
nor U1813 (N_1813,N_1759,N_1791);
or U1814 (N_1814,N_1790,N_1744);
nand U1815 (N_1815,N_1748,N_1746);
and U1816 (N_1816,N_1773,N_1755);
nor U1817 (N_1817,N_1771,N_1740);
nand U1818 (N_1818,N_1769,N_1768);
or U1819 (N_1819,N_1776,N_1797);
nand U1820 (N_1820,N_1796,N_1770);
nand U1821 (N_1821,N_1760,N_1782);
or U1822 (N_1822,N_1762,N_1761);
or U1823 (N_1823,N_1754,N_1758);
or U1824 (N_1824,N_1742,N_1795);
or U1825 (N_1825,N_1751,N_1747);
nor U1826 (N_1826,N_1779,N_1792);
nand U1827 (N_1827,N_1784,N_1749);
or U1828 (N_1828,N_1786,N_1783);
nor U1829 (N_1829,N_1750,N_1781);
nor U1830 (N_1830,N_1754,N_1793);
and U1831 (N_1831,N_1786,N_1788);
nand U1832 (N_1832,N_1781,N_1786);
nor U1833 (N_1833,N_1749,N_1772);
or U1834 (N_1834,N_1765,N_1780);
or U1835 (N_1835,N_1742,N_1782);
nor U1836 (N_1836,N_1756,N_1780);
nand U1837 (N_1837,N_1760,N_1783);
nand U1838 (N_1838,N_1769,N_1755);
nand U1839 (N_1839,N_1770,N_1764);
nor U1840 (N_1840,N_1773,N_1789);
and U1841 (N_1841,N_1782,N_1764);
nand U1842 (N_1842,N_1771,N_1778);
nand U1843 (N_1843,N_1774,N_1773);
nand U1844 (N_1844,N_1766,N_1784);
nor U1845 (N_1845,N_1761,N_1750);
or U1846 (N_1846,N_1787,N_1767);
or U1847 (N_1847,N_1779,N_1755);
or U1848 (N_1848,N_1793,N_1783);
and U1849 (N_1849,N_1753,N_1747);
and U1850 (N_1850,N_1778,N_1781);
and U1851 (N_1851,N_1741,N_1753);
nand U1852 (N_1852,N_1755,N_1799);
and U1853 (N_1853,N_1794,N_1771);
and U1854 (N_1854,N_1772,N_1755);
nor U1855 (N_1855,N_1760,N_1754);
nor U1856 (N_1856,N_1745,N_1740);
nand U1857 (N_1857,N_1768,N_1756);
nand U1858 (N_1858,N_1778,N_1747);
and U1859 (N_1859,N_1755,N_1749);
nor U1860 (N_1860,N_1851,N_1804);
and U1861 (N_1861,N_1826,N_1848);
nand U1862 (N_1862,N_1815,N_1813);
or U1863 (N_1863,N_1811,N_1806);
or U1864 (N_1864,N_1819,N_1821);
and U1865 (N_1865,N_1810,N_1853);
and U1866 (N_1866,N_1831,N_1837);
nand U1867 (N_1867,N_1800,N_1818);
nor U1868 (N_1868,N_1805,N_1825);
or U1869 (N_1869,N_1802,N_1830);
or U1870 (N_1870,N_1841,N_1842);
nor U1871 (N_1871,N_1820,N_1839);
and U1872 (N_1872,N_1854,N_1801);
and U1873 (N_1873,N_1844,N_1838);
nor U1874 (N_1874,N_1840,N_1814);
or U1875 (N_1875,N_1836,N_1843);
and U1876 (N_1876,N_1850,N_1833);
nand U1877 (N_1877,N_1849,N_1855);
nand U1878 (N_1878,N_1832,N_1845);
nand U1879 (N_1879,N_1809,N_1847);
nor U1880 (N_1880,N_1812,N_1827);
nand U1881 (N_1881,N_1829,N_1856);
or U1882 (N_1882,N_1816,N_1807);
or U1883 (N_1883,N_1803,N_1817);
nor U1884 (N_1884,N_1846,N_1852);
nand U1885 (N_1885,N_1857,N_1828);
or U1886 (N_1886,N_1858,N_1834);
nor U1887 (N_1887,N_1823,N_1824);
or U1888 (N_1888,N_1808,N_1822);
nor U1889 (N_1889,N_1835,N_1859);
nor U1890 (N_1890,N_1833,N_1836);
nor U1891 (N_1891,N_1850,N_1856);
and U1892 (N_1892,N_1854,N_1804);
nor U1893 (N_1893,N_1846,N_1855);
nor U1894 (N_1894,N_1834,N_1817);
nor U1895 (N_1895,N_1824,N_1851);
or U1896 (N_1896,N_1810,N_1858);
nand U1897 (N_1897,N_1818,N_1851);
and U1898 (N_1898,N_1851,N_1829);
nor U1899 (N_1899,N_1844,N_1800);
and U1900 (N_1900,N_1834,N_1821);
nor U1901 (N_1901,N_1823,N_1837);
or U1902 (N_1902,N_1843,N_1826);
nor U1903 (N_1903,N_1823,N_1822);
and U1904 (N_1904,N_1823,N_1816);
and U1905 (N_1905,N_1836,N_1827);
nor U1906 (N_1906,N_1857,N_1834);
nand U1907 (N_1907,N_1859,N_1830);
nor U1908 (N_1908,N_1811,N_1840);
nor U1909 (N_1909,N_1835,N_1840);
nor U1910 (N_1910,N_1850,N_1812);
nor U1911 (N_1911,N_1846,N_1812);
nand U1912 (N_1912,N_1857,N_1811);
or U1913 (N_1913,N_1816,N_1859);
or U1914 (N_1914,N_1805,N_1852);
or U1915 (N_1915,N_1807,N_1811);
nand U1916 (N_1916,N_1818,N_1806);
and U1917 (N_1917,N_1813,N_1828);
nor U1918 (N_1918,N_1845,N_1808);
nor U1919 (N_1919,N_1808,N_1821);
nand U1920 (N_1920,N_1876,N_1908);
and U1921 (N_1921,N_1871,N_1870);
nand U1922 (N_1922,N_1911,N_1893);
or U1923 (N_1923,N_1879,N_1886);
or U1924 (N_1924,N_1895,N_1902);
and U1925 (N_1925,N_1878,N_1863);
nand U1926 (N_1926,N_1888,N_1882);
or U1927 (N_1927,N_1885,N_1907);
nor U1928 (N_1928,N_1881,N_1873);
or U1929 (N_1929,N_1869,N_1898);
or U1930 (N_1930,N_1903,N_1915);
nor U1931 (N_1931,N_1896,N_1877);
and U1932 (N_1932,N_1919,N_1865);
nor U1933 (N_1933,N_1872,N_1899);
nand U1934 (N_1934,N_1862,N_1900);
nand U1935 (N_1935,N_1904,N_1894);
nand U1936 (N_1936,N_1916,N_1913);
or U1937 (N_1937,N_1867,N_1891);
or U1938 (N_1938,N_1875,N_1905);
nor U1939 (N_1939,N_1912,N_1866);
and U1940 (N_1940,N_1892,N_1887);
nand U1941 (N_1941,N_1864,N_1917);
xnor U1942 (N_1942,N_1868,N_1860);
nand U1943 (N_1943,N_1880,N_1906);
and U1944 (N_1944,N_1897,N_1883);
and U1945 (N_1945,N_1889,N_1884);
or U1946 (N_1946,N_1918,N_1910);
nand U1947 (N_1947,N_1914,N_1890);
nand U1948 (N_1948,N_1861,N_1909);
xnor U1949 (N_1949,N_1874,N_1901);
nor U1950 (N_1950,N_1886,N_1896);
nand U1951 (N_1951,N_1883,N_1862);
nand U1952 (N_1952,N_1908,N_1888);
nor U1953 (N_1953,N_1889,N_1909);
or U1954 (N_1954,N_1875,N_1860);
nand U1955 (N_1955,N_1866,N_1914);
nor U1956 (N_1956,N_1909,N_1914);
and U1957 (N_1957,N_1866,N_1889);
or U1958 (N_1958,N_1919,N_1884);
nor U1959 (N_1959,N_1897,N_1876);
nand U1960 (N_1960,N_1917,N_1881);
nand U1961 (N_1961,N_1899,N_1907);
nor U1962 (N_1962,N_1862,N_1897);
nand U1963 (N_1963,N_1901,N_1876);
and U1964 (N_1964,N_1864,N_1881);
nor U1965 (N_1965,N_1875,N_1894);
nor U1966 (N_1966,N_1911,N_1913);
nor U1967 (N_1967,N_1869,N_1895);
xnor U1968 (N_1968,N_1901,N_1866);
nand U1969 (N_1969,N_1892,N_1875);
nor U1970 (N_1970,N_1903,N_1904);
nand U1971 (N_1971,N_1912,N_1898);
nor U1972 (N_1972,N_1881,N_1912);
nor U1973 (N_1973,N_1889,N_1875);
nor U1974 (N_1974,N_1909,N_1863);
or U1975 (N_1975,N_1903,N_1896);
nand U1976 (N_1976,N_1868,N_1869);
nand U1977 (N_1977,N_1873,N_1899);
nand U1978 (N_1978,N_1919,N_1867);
nand U1979 (N_1979,N_1913,N_1892);
or U1980 (N_1980,N_1978,N_1948);
or U1981 (N_1981,N_1971,N_1977);
and U1982 (N_1982,N_1941,N_1949);
nor U1983 (N_1983,N_1979,N_1974);
or U1984 (N_1984,N_1935,N_1923);
nand U1985 (N_1985,N_1958,N_1942);
and U1986 (N_1986,N_1951,N_1933);
nand U1987 (N_1987,N_1924,N_1946);
nor U1988 (N_1988,N_1963,N_1936);
or U1989 (N_1989,N_1954,N_1925);
nand U1990 (N_1990,N_1937,N_1944);
nand U1991 (N_1991,N_1960,N_1973);
nand U1992 (N_1992,N_1931,N_1970);
nand U1993 (N_1993,N_1934,N_1929);
or U1994 (N_1994,N_1961,N_1938);
or U1995 (N_1995,N_1965,N_1930);
nor U1996 (N_1996,N_1926,N_1920);
and U1997 (N_1997,N_1972,N_1955);
and U1998 (N_1998,N_1959,N_1957);
nand U1999 (N_1999,N_1966,N_1939);
or U2000 (N_2000,N_1950,N_1962);
or U2001 (N_2001,N_1969,N_1945);
nor U2002 (N_2002,N_1967,N_1964);
nand U2003 (N_2003,N_1953,N_1943);
or U2004 (N_2004,N_1975,N_1932);
nor U2005 (N_2005,N_1952,N_1940);
or U2006 (N_2006,N_1921,N_1956);
xor U2007 (N_2007,N_1947,N_1922);
or U2008 (N_2008,N_1927,N_1928);
nor U2009 (N_2009,N_1976,N_1968);
or U2010 (N_2010,N_1926,N_1960);
and U2011 (N_2011,N_1924,N_1939);
nor U2012 (N_2012,N_1927,N_1952);
or U2013 (N_2013,N_1944,N_1977);
and U2014 (N_2014,N_1969,N_1920);
nor U2015 (N_2015,N_1958,N_1962);
nand U2016 (N_2016,N_1936,N_1926);
nand U2017 (N_2017,N_1937,N_1934);
nor U2018 (N_2018,N_1975,N_1926);
and U2019 (N_2019,N_1970,N_1935);
or U2020 (N_2020,N_1976,N_1951);
and U2021 (N_2021,N_1934,N_1960);
or U2022 (N_2022,N_1923,N_1966);
nand U2023 (N_2023,N_1928,N_1954);
and U2024 (N_2024,N_1932,N_1965);
nor U2025 (N_2025,N_1962,N_1976);
nor U2026 (N_2026,N_1924,N_1957);
or U2027 (N_2027,N_1935,N_1950);
or U2028 (N_2028,N_1957,N_1952);
nand U2029 (N_2029,N_1953,N_1942);
or U2030 (N_2030,N_1933,N_1956);
and U2031 (N_2031,N_1936,N_1952);
and U2032 (N_2032,N_1931,N_1960);
nand U2033 (N_2033,N_1927,N_1960);
and U2034 (N_2034,N_1951,N_1957);
nand U2035 (N_2035,N_1956,N_1954);
nor U2036 (N_2036,N_1956,N_1969);
nand U2037 (N_2037,N_1934,N_1977);
nand U2038 (N_2038,N_1946,N_1932);
nor U2039 (N_2039,N_1922,N_1969);
xnor U2040 (N_2040,N_2014,N_2025);
nand U2041 (N_2041,N_1996,N_2009);
nand U2042 (N_2042,N_2010,N_2012);
and U2043 (N_2043,N_1989,N_2034);
nor U2044 (N_2044,N_2038,N_1993);
and U2045 (N_2045,N_1988,N_2033);
and U2046 (N_2046,N_2001,N_2024);
nor U2047 (N_2047,N_1999,N_2037);
or U2048 (N_2048,N_2029,N_2027);
nand U2049 (N_2049,N_1997,N_2008);
or U2050 (N_2050,N_1986,N_2022);
nor U2051 (N_2051,N_1995,N_2036);
and U2052 (N_2052,N_2007,N_2026);
and U2053 (N_2053,N_1982,N_1992);
and U2054 (N_2054,N_2023,N_1983);
nor U2055 (N_2055,N_2006,N_1994);
nand U2056 (N_2056,N_2013,N_2020);
and U2057 (N_2057,N_2039,N_2028);
nand U2058 (N_2058,N_2031,N_1998);
or U2059 (N_2059,N_2015,N_2000);
or U2060 (N_2060,N_1985,N_2030);
or U2061 (N_2061,N_2016,N_1980);
and U2062 (N_2062,N_2035,N_2019);
xor U2063 (N_2063,N_2017,N_2003);
or U2064 (N_2064,N_1991,N_2011);
nand U2065 (N_2065,N_2002,N_1990);
nand U2066 (N_2066,N_2032,N_1984);
and U2067 (N_2067,N_1987,N_2005);
and U2068 (N_2068,N_1981,N_2021);
nand U2069 (N_2069,N_2004,N_2018);
and U2070 (N_2070,N_1987,N_2037);
nor U2071 (N_2071,N_2018,N_2032);
nand U2072 (N_2072,N_2030,N_2032);
or U2073 (N_2073,N_1994,N_1982);
nor U2074 (N_2074,N_2024,N_2011);
or U2075 (N_2075,N_2036,N_1988);
and U2076 (N_2076,N_2019,N_2018);
nand U2077 (N_2077,N_2016,N_1990);
and U2078 (N_2078,N_2000,N_1986);
nor U2079 (N_2079,N_2022,N_2038);
xnor U2080 (N_2080,N_1991,N_2032);
xor U2081 (N_2081,N_1990,N_1987);
or U2082 (N_2082,N_2016,N_2008);
nand U2083 (N_2083,N_2036,N_2023);
and U2084 (N_2084,N_2023,N_2027);
nor U2085 (N_2085,N_1992,N_2021);
and U2086 (N_2086,N_2000,N_2039);
or U2087 (N_2087,N_2019,N_1981);
or U2088 (N_2088,N_1985,N_2007);
nor U2089 (N_2089,N_2039,N_2003);
or U2090 (N_2090,N_2013,N_2001);
and U2091 (N_2091,N_2021,N_1989);
or U2092 (N_2092,N_2038,N_1995);
nor U2093 (N_2093,N_1993,N_1987);
nor U2094 (N_2094,N_2027,N_2028);
or U2095 (N_2095,N_2000,N_1987);
or U2096 (N_2096,N_2010,N_2011);
xor U2097 (N_2097,N_2019,N_2031);
nand U2098 (N_2098,N_2016,N_2020);
nand U2099 (N_2099,N_2003,N_1996);
nand U2100 (N_2100,N_2071,N_2057);
and U2101 (N_2101,N_2091,N_2099);
nand U2102 (N_2102,N_2070,N_2067);
nor U2103 (N_2103,N_2056,N_2051);
and U2104 (N_2104,N_2076,N_2072);
and U2105 (N_2105,N_2080,N_2083);
and U2106 (N_2106,N_2045,N_2085);
nand U2107 (N_2107,N_2073,N_2078);
nand U2108 (N_2108,N_2064,N_2053);
nand U2109 (N_2109,N_2066,N_2044);
nand U2110 (N_2110,N_2097,N_2069);
nand U2111 (N_2111,N_2094,N_2062);
or U2112 (N_2112,N_2059,N_2084);
or U2113 (N_2113,N_2079,N_2074);
nand U2114 (N_2114,N_2060,N_2095);
and U2115 (N_2115,N_2049,N_2058);
and U2116 (N_2116,N_2096,N_2043);
nor U2117 (N_2117,N_2075,N_2077);
nor U2118 (N_2118,N_2052,N_2050);
and U2119 (N_2119,N_2093,N_2098);
xnor U2120 (N_2120,N_2041,N_2089);
or U2121 (N_2121,N_2063,N_2087);
and U2122 (N_2122,N_2055,N_2065);
and U2123 (N_2123,N_2090,N_2068);
and U2124 (N_2124,N_2086,N_2054);
and U2125 (N_2125,N_2061,N_2081);
nor U2126 (N_2126,N_2048,N_2046);
nand U2127 (N_2127,N_2047,N_2092);
or U2128 (N_2128,N_2042,N_2040);
nor U2129 (N_2129,N_2088,N_2082);
nand U2130 (N_2130,N_2081,N_2079);
nand U2131 (N_2131,N_2094,N_2049);
and U2132 (N_2132,N_2040,N_2089);
or U2133 (N_2133,N_2094,N_2059);
and U2134 (N_2134,N_2051,N_2067);
nand U2135 (N_2135,N_2092,N_2094);
or U2136 (N_2136,N_2094,N_2047);
or U2137 (N_2137,N_2077,N_2044);
or U2138 (N_2138,N_2066,N_2076);
and U2139 (N_2139,N_2056,N_2098);
xor U2140 (N_2140,N_2090,N_2098);
nand U2141 (N_2141,N_2086,N_2055);
nor U2142 (N_2142,N_2072,N_2092);
and U2143 (N_2143,N_2090,N_2089);
nor U2144 (N_2144,N_2059,N_2043);
nor U2145 (N_2145,N_2051,N_2064);
nor U2146 (N_2146,N_2056,N_2040);
or U2147 (N_2147,N_2095,N_2088);
and U2148 (N_2148,N_2072,N_2081);
or U2149 (N_2149,N_2079,N_2096);
nor U2150 (N_2150,N_2048,N_2067);
and U2151 (N_2151,N_2042,N_2051);
and U2152 (N_2152,N_2086,N_2063);
or U2153 (N_2153,N_2044,N_2071);
nand U2154 (N_2154,N_2056,N_2059);
or U2155 (N_2155,N_2069,N_2056);
and U2156 (N_2156,N_2093,N_2055);
and U2157 (N_2157,N_2098,N_2088);
and U2158 (N_2158,N_2070,N_2043);
or U2159 (N_2159,N_2044,N_2045);
or U2160 (N_2160,N_2122,N_2129);
and U2161 (N_2161,N_2131,N_2149);
and U2162 (N_2162,N_2151,N_2150);
nand U2163 (N_2163,N_2108,N_2133);
nor U2164 (N_2164,N_2155,N_2140);
nand U2165 (N_2165,N_2143,N_2141);
nand U2166 (N_2166,N_2124,N_2119);
and U2167 (N_2167,N_2138,N_2102);
nand U2168 (N_2168,N_2130,N_2159);
or U2169 (N_2169,N_2121,N_2146);
and U2170 (N_2170,N_2123,N_2116);
or U2171 (N_2171,N_2101,N_2132);
and U2172 (N_2172,N_2114,N_2139);
nor U2173 (N_2173,N_2111,N_2126);
nor U2174 (N_2174,N_2113,N_2105);
nor U2175 (N_2175,N_2142,N_2156);
and U2176 (N_2176,N_2152,N_2118);
nor U2177 (N_2177,N_2134,N_2154);
and U2178 (N_2178,N_2128,N_2157);
nand U2179 (N_2179,N_2107,N_2106);
nand U2180 (N_2180,N_2144,N_2103);
nor U2181 (N_2181,N_2136,N_2110);
nor U2182 (N_2182,N_2100,N_2127);
nand U2183 (N_2183,N_2115,N_2148);
nor U2184 (N_2184,N_2112,N_2117);
nand U2185 (N_2185,N_2109,N_2120);
nand U2186 (N_2186,N_2104,N_2125);
and U2187 (N_2187,N_2145,N_2147);
xnor U2188 (N_2188,N_2137,N_2158);
xnor U2189 (N_2189,N_2153,N_2135);
nor U2190 (N_2190,N_2109,N_2110);
nand U2191 (N_2191,N_2147,N_2140);
or U2192 (N_2192,N_2157,N_2119);
nor U2193 (N_2193,N_2154,N_2131);
nor U2194 (N_2194,N_2110,N_2122);
nor U2195 (N_2195,N_2144,N_2135);
or U2196 (N_2196,N_2117,N_2135);
nand U2197 (N_2197,N_2132,N_2103);
nand U2198 (N_2198,N_2102,N_2104);
nor U2199 (N_2199,N_2148,N_2111);
nand U2200 (N_2200,N_2138,N_2103);
and U2201 (N_2201,N_2116,N_2121);
or U2202 (N_2202,N_2139,N_2158);
nor U2203 (N_2203,N_2145,N_2138);
nor U2204 (N_2204,N_2155,N_2144);
nand U2205 (N_2205,N_2151,N_2145);
or U2206 (N_2206,N_2115,N_2108);
nor U2207 (N_2207,N_2114,N_2146);
or U2208 (N_2208,N_2100,N_2156);
and U2209 (N_2209,N_2119,N_2139);
and U2210 (N_2210,N_2141,N_2126);
xor U2211 (N_2211,N_2102,N_2100);
nand U2212 (N_2212,N_2111,N_2155);
or U2213 (N_2213,N_2144,N_2113);
nor U2214 (N_2214,N_2159,N_2123);
nor U2215 (N_2215,N_2132,N_2113);
and U2216 (N_2216,N_2121,N_2119);
xor U2217 (N_2217,N_2136,N_2130);
or U2218 (N_2218,N_2110,N_2153);
nand U2219 (N_2219,N_2134,N_2120);
nor U2220 (N_2220,N_2204,N_2168);
nor U2221 (N_2221,N_2196,N_2173);
and U2222 (N_2222,N_2164,N_2184);
nand U2223 (N_2223,N_2186,N_2194);
and U2224 (N_2224,N_2187,N_2193);
nor U2225 (N_2225,N_2161,N_2216);
and U2226 (N_2226,N_2201,N_2213);
and U2227 (N_2227,N_2211,N_2214);
nor U2228 (N_2228,N_2212,N_2218);
and U2229 (N_2229,N_2189,N_2165);
or U2230 (N_2230,N_2171,N_2183);
nand U2231 (N_2231,N_2215,N_2192);
or U2232 (N_2232,N_2185,N_2207);
or U2233 (N_2233,N_2198,N_2197);
and U2234 (N_2234,N_2182,N_2162);
and U2235 (N_2235,N_2178,N_2160);
nor U2236 (N_2236,N_2191,N_2206);
and U2237 (N_2237,N_2208,N_2202);
nor U2238 (N_2238,N_2163,N_2210);
or U2239 (N_2239,N_2179,N_2172);
nor U2240 (N_2240,N_2175,N_2169);
nor U2241 (N_2241,N_2205,N_2167);
and U2242 (N_2242,N_2166,N_2176);
or U2243 (N_2243,N_2219,N_2203);
xnor U2244 (N_2244,N_2209,N_2188);
nor U2245 (N_2245,N_2200,N_2181);
nor U2246 (N_2246,N_2174,N_2195);
nand U2247 (N_2247,N_2180,N_2199);
nor U2248 (N_2248,N_2170,N_2217);
and U2249 (N_2249,N_2177,N_2190);
and U2250 (N_2250,N_2189,N_2162);
and U2251 (N_2251,N_2182,N_2190);
and U2252 (N_2252,N_2174,N_2164);
and U2253 (N_2253,N_2192,N_2190);
nand U2254 (N_2254,N_2183,N_2197);
and U2255 (N_2255,N_2166,N_2185);
nand U2256 (N_2256,N_2200,N_2172);
or U2257 (N_2257,N_2191,N_2170);
or U2258 (N_2258,N_2194,N_2201);
or U2259 (N_2259,N_2162,N_2164);
nor U2260 (N_2260,N_2179,N_2212);
or U2261 (N_2261,N_2182,N_2183);
or U2262 (N_2262,N_2194,N_2202);
nor U2263 (N_2263,N_2191,N_2200);
nor U2264 (N_2264,N_2162,N_2205);
or U2265 (N_2265,N_2162,N_2166);
or U2266 (N_2266,N_2191,N_2160);
and U2267 (N_2267,N_2174,N_2206);
nor U2268 (N_2268,N_2198,N_2183);
and U2269 (N_2269,N_2192,N_2183);
nand U2270 (N_2270,N_2169,N_2216);
and U2271 (N_2271,N_2182,N_2202);
or U2272 (N_2272,N_2219,N_2217);
or U2273 (N_2273,N_2209,N_2216);
nor U2274 (N_2274,N_2171,N_2178);
nor U2275 (N_2275,N_2206,N_2208);
nor U2276 (N_2276,N_2162,N_2204);
or U2277 (N_2277,N_2218,N_2194);
nor U2278 (N_2278,N_2218,N_2219);
or U2279 (N_2279,N_2170,N_2207);
and U2280 (N_2280,N_2243,N_2247);
xor U2281 (N_2281,N_2263,N_2239);
and U2282 (N_2282,N_2237,N_2233);
xnor U2283 (N_2283,N_2258,N_2273);
or U2284 (N_2284,N_2234,N_2220);
nor U2285 (N_2285,N_2277,N_2221);
xnor U2286 (N_2286,N_2236,N_2232);
nand U2287 (N_2287,N_2249,N_2265);
or U2288 (N_2288,N_2272,N_2256);
and U2289 (N_2289,N_2257,N_2223);
or U2290 (N_2290,N_2266,N_2261);
nand U2291 (N_2291,N_2267,N_2252);
or U2292 (N_2292,N_2279,N_2245);
or U2293 (N_2293,N_2248,N_2251);
nor U2294 (N_2294,N_2242,N_2255);
nor U2295 (N_2295,N_2260,N_2246);
nand U2296 (N_2296,N_2270,N_2238);
nand U2297 (N_2297,N_2254,N_2222);
nand U2298 (N_2298,N_2262,N_2224);
nor U2299 (N_2299,N_2241,N_2231);
nor U2300 (N_2300,N_2228,N_2259);
nor U2301 (N_2301,N_2253,N_2275);
or U2302 (N_2302,N_2269,N_2274);
and U2303 (N_2303,N_2229,N_2235);
nand U2304 (N_2304,N_2278,N_2244);
or U2305 (N_2305,N_2226,N_2268);
nor U2306 (N_2306,N_2250,N_2225);
and U2307 (N_2307,N_2264,N_2240);
or U2308 (N_2308,N_2230,N_2227);
nor U2309 (N_2309,N_2276,N_2271);
nand U2310 (N_2310,N_2230,N_2253);
and U2311 (N_2311,N_2220,N_2222);
or U2312 (N_2312,N_2239,N_2268);
nand U2313 (N_2313,N_2244,N_2270);
and U2314 (N_2314,N_2244,N_2277);
and U2315 (N_2315,N_2246,N_2264);
nand U2316 (N_2316,N_2238,N_2235);
or U2317 (N_2317,N_2225,N_2251);
nor U2318 (N_2318,N_2251,N_2245);
and U2319 (N_2319,N_2235,N_2271);
or U2320 (N_2320,N_2220,N_2257);
and U2321 (N_2321,N_2257,N_2272);
nand U2322 (N_2322,N_2229,N_2250);
nand U2323 (N_2323,N_2252,N_2266);
nand U2324 (N_2324,N_2228,N_2270);
nand U2325 (N_2325,N_2251,N_2279);
or U2326 (N_2326,N_2277,N_2228);
or U2327 (N_2327,N_2275,N_2257);
and U2328 (N_2328,N_2233,N_2228);
and U2329 (N_2329,N_2243,N_2234);
or U2330 (N_2330,N_2236,N_2254);
and U2331 (N_2331,N_2261,N_2238);
nand U2332 (N_2332,N_2270,N_2232);
nand U2333 (N_2333,N_2244,N_2249);
nand U2334 (N_2334,N_2240,N_2229);
nand U2335 (N_2335,N_2228,N_2247);
and U2336 (N_2336,N_2267,N_2273);
or U2337 (N_2337,N_2220,N_2235);
or U2338 (N_2338,N_2259,N_2277);
and U2339 (N_2339,N_2242,N_2265);
and U2340 (N_2340,N_2322,N_2316);
or U2341 (N_2341,N_2335,N_2306);
nor U2342 (N_2342,N_2339,N_2281);
or U2343 (N_2343,N_2331,N_2313);
or U2344 (N_2344,N_2291,N_2312);
nand U2345 (N_2345,N_2326,N_2320);
and U2346 (N_2346,N_2299,N_2310);
or U2347 (N_2347,N_2294,N_2332);
or U2348 (N_2348,N_2307,N_2317);
and U2349 (N_2349,N_2297,N_2300);
xor U2350 (N_2350,N_2286,N_2314);
or U2351 (N_2351,N_2318,N_2315);
or U2352 (N_2352,N_2324,N_2305);
and U2353 (N_2353,N_2330,N_2336);
nor U2354 (N_2354,N_2282,N_2333);
or U2355 (N_2355,N_2327,N_2285);
nor U2356 (N_2356,N_2311,N_2292);
and U2357 (N_2357,N_2319,N_2301);
or U2358 (N_2358,N_2321,N_2283);
or U2359 (N_2359,N_2302,N_2287);
nor U2360 (N_2360,N_2309,N_2289);
nor U2361 (N_2361,N_2296,N_2337);
or U2362 (N_2362,N_2325,N_2338);
nand U2363 (N_2363,N_2308,N_2288);
and U2364 (N_2364,N_2323,N_2303);
nor U2365 (N_2365,N_2293,N_2295);
and U2366 (N_2366,N_2298,N_2290);
nor U2367 (N_2367,N_2280,N_2329);
nor U2368 (N_2368,N_2334,N_2304);
xor U2369 (N_2369,N_2284,N_2328);
nor U2370 (N_2370,N_2338,N_2329);
and U2371 (N_2371,N_2335,N_2329);
nand U2372 (N_2372,N_2324,N_2319);
nand U2373 (N_2373,N_2305,N_2287);
nor U2374 (N_2374,N_2308,N_2313);
and U2375 (N_2375,N_2312,N_2323);
nor U2376 (N_2376,N_2300,N_2323);
nand U2377 (N_2377,N_2299,N_2339);
nor U2378 (N_2378,N_2335,N_2324);
nor U2379 (N_2379,N_2328,N_2304);
or U2380 (N_2380,N_2295,N_2298);
xnor U2381 (N_2381,N_2339,N_2291);
nand U2382 (N_2382,N_2282,N_2290);
nor U2383 (N_2383,N_2321,N_2337);
nor U2384 (N_2384,N_2293,N_2285);
or U2385 (N_2385,N_2284,N_2337);
or U2386 (N_2386,N_2334,N_2333);
nand U2387 (N_2387,N_2339,N_2336);
nor U2388 (N_2388,N_2306,N_2339);
or U2389 (N_2389,N_2313,N_2311);
or U2390 (N_2390,N_2299,N_2327);
nand U2391 (N_2391,N_2285,N_2287);
nor U2392 (N_2392,N_2329,N_2327);
and U2393 (N_2393,N_2296,N_2331);
or U2394 (N_2394,N_2321,N_2336);
nor U2395 (N_2395,N_2292,N_2281);
nor U2396 (N_2396,N_2300,N_2310);
and U2397 (N_2397,N_2321,N_2305);
and U2398 (N_2398,N_2286,N_2306);
and U2399 (N_2399,N_2305,N_2312);
nor U2400 (N_2400,N_2375,N_2350);
nand U2401 (N_2401,N_2368,N_2359);
or U2402 (N_2402,N_2342,N_2351);
and U2403 (N_2403,N_2347,N_2346);
nor U2404 (N_2404,N_2353,N_2385);
nor U2405 (N_2405,N_2394,N_2376);
nor U2406 (N_2406,N_2356,N_2392);
and U2407 (N_2407,N_2352,N_2390);
or U2408 (N_2408,N_2388,N_2358);
nor U2409 (N_2409,N_2397,N_2382);
nor U2410 (N_2410,N_2354,N_2378);
nor U2411 (N_2411,N_2395,N_2391);
and U2412 (N_2412,N_2344,N_2367);
or U2413 (N_2413,N_2363,N_2383);
nand U2414 (N_2414,N_2380,N_2343);
nand U2415 (N_2415,N_2364,N_2357);
nand U2416 (N_2416,N_2398,N_2370);
and U2417 (N_2417,N_2348,N_2386);
and U2418 (N_2418,N_2396,N_2384);
nand U2419 (N_2419,N_2369,N_2355);
nand U2420 (N_2420,N_2381,N_2374);
nand U2421 (N_2421,N_2377,N_2373);
nor U2422 (N_2422,N_2372,N_2371);
nor U2423 (N_2423,N_2341,N_2340);
or U2424 (N_2424,N_2345,N_2360);
nor U2425 (N_2425,N_2399,N_2389);
xnor U2426 (N_2426,N_2362,N_2366);
and U2427 (N_2427,N_2365,N_2379);
and U2428 (N_2428,N_2361,N_2393);
nand U2429 (N_2429,N_2349,N_2387);
and U2430 (N_2430,N_2393,N_2380);
nand U2431 (N_2431,N_2377,N_2360);
or U2432 (N_2432,N_2374,N_2361);
and U2433 (N_2433,N_2394,N_2369);
or U2434 (N_2434,N_2396,N_2341);
or U2435 (N_2435,N_2366,N_2389);
nor U2436 (N_2436,N_2368,N_2379);
nand U2437 (N_2437,N_2349,N_2378);
nand U2438 (N_2438,N_2368,N_2362);
and U2439 (N_2439,N_2351,N_2397);
nand U2440 (N_2440,N_2371,N_2382);
or U2441 (N_2441,N_2392,N_2370);
nand U2442 (N_2442,N_2354,N_2359);
nor U2443 (N_2443,N_2399,N_2356);
or U2444 (N_2444,N_2353,N_2397);
nand U2445 (N_2445,N_2375,N_2381);
nand U2446 (N_2446,N_2383,N_2378);
nor U2447 (N_2447,N_2340,N_2374);
and U2448 (N_2448,N_2359,N_2348);
and U2449 (N_2449,N_2379,N_2374);
or U2450 (N_2450,N_2346,N_2354);
or U2451 (N_2451,N_2341,N_2381);
nor U2452 (N_2452,N_2371,N_2396);
nor U2453 (N_2453,N_2354,N_2393);
nor U2454 (N_2454,N_2359,N_2355);
nor U2455 (N_2455,N_2394,N_2358);
xor U2456 (N_2456,N_2360,N_2353);
or U2457 (N_2457,N_2379,N_2376);
and U2458 (N_2458,N_2361,N_2355);
or U2459 (N_2459,N_2342,N_2343);
nand U2460 (N_2460,N_2406,N_2408);
and U2461 (N_2461,N_2439,N_2434);
nand U2462 (N_2462,N_2411,N_2416);
nand U2463 (N_2463,N_2457,N_2415);
and U2464 (N_2464,N_2407,N_2446);
nor U2465 (N_2465,N_2435,N_2403);
or U2466 (N_2466,N_2440,N_2402);
and U2467 (N_2467,N_2414,N_2421);
xnor U2468 (N_2468,N_2427,N_2404);
or U2469 (N_2469,N_2455,N_2444);
or U2470 (N_2470,N_2412,N_2458);
nand U2471 (N_2471,N_2436,N_2425);
nand U2472 (N_2472,N_2424,N_2423);
nor U2473 (N_2473,N_2445,N_2454);
nand U2474 (N_2474,N_2400,N_2419);
and U2475 (N_2475,N_2449,N_2428);
nand U2476 (N_2476,N_2433,N_2432);
nand U2477 (N_2477,N_2418,N_2422);
or U2478 (N_2478,N_2448,N_2409);
or U2479 (N_2479,N_2441,N_2430);
and U2480 (N_2480,N_2456,N_2452);
or U2481 (N_2481,N_2431,N_2442);
or U2482 (N_2482,N_2459,N_2401);
nor U2483 (N_2483,N_2429,N_2451);
nor U2484 (N_2484,N_2410,N_2443);
or U2485 (N_2485,N_2437,N_2417);
nand U2486 (N_2486,N_2450,N_2426);
or U2487 (N_2487,N_2447,N_2420);
or U2488 (N_2488,N_2453,N_2413);
nand U2489 (N_2489,N_2405,N_2438);
and U2490 (N_2490,N_2420,N_2400);
nor U2491 (N_2491,N_2414,N_2458);
and U2492 (N_2492,N_2401,N_2447);
nand U2493 (N_2493,N_2444,N_2426);
nand U2494 (N_2494,N_2400,N_2417);
nand U2495 (N_2495,N_2426,N_2403);
nand U2496 (N_2496,N_2459,N_2453);
and U2497 (N_2497,N_2453,N_2428);
nor U2498 (N_2498,N_2440,N_2452);
or U2499 (N_2499,N_2406,N_2455);
and U2500 (N_2500,N_2414,N_2433);
or U2501 (N_2501,N_2404,N_2424);
and U2502 (N_2502,N_2412,N_2457);
and U2503 (N_2503,N_2436,N_2403);
or U2504 (N_2504,N_2421,N_2437);
and U2505 (N_2505,N_2429,N_2444);
nand U2506 (N_2506,N_2429,N_2415);
and U2507 (N_2507,N_2443,N_2424);
or U2508 (N_2508,N_2400,N_2412);
nor U2509 (N_2509,N_2408,N_2407);
nand U2510 (N_2510,N_2447,N_2448);
nand U2511 (N_2511,N_2426,N_2445);
and U2512 (N_2512,N_2422,N_2417);
nor U2513 (N_2513,N_2446,N_2419);
and U2514 (N_2514,N_2411,N_2419);
nand U2515 (N_2515,N_2404,N_2458);
nand U2516 (N_2516,N_2406,N_2436);
nand U2517 (N_2517,N_2445,N_2419);
nand U2518 (N_2518,N_2427,N_2456);
nor U2519 (N_2519,N_2444,N_2458);
nand U2520 (N_2520,N_2515,N_2483);
and U2521 (N_2521,N_2511,N_2495);
or U2522 (N_2522,N_2517,N_2508);
nor U2523 (N_2523,N_2505,N_2518);
or U2524 (N_2524,N_2476,N_2490);
or U2525 (N_2525,N_2497,N_2493);
and U2526 (N_2526,N_2478,N_2510);
and U2527 (N_2527,N_2463,N_2509);
and U2528 (N_2528,N_2471,N_2501);
or U2529 (N_2529,N_2477,N_2482);
and U2530 (N_2530,N_2506,N_2492);
and U2531 (N_2531,N_2519,N_2516);
nor U2532 (N_2532,N_2466,N_2472);
nor U2533 (N_2533,N_2480,N_2461);
nand U2534 (N_2534,N_2464,N_2498);
or U2535 (N_2535,N_2475,N_2462);
nand U2536 (N_2536,N_2486,N_2503);
or U2537 (N_2537,N_2474,N_2465);
nand U2538 (N_2538,N_2470,N_2502);
and U2539 (N_2539,N_2473,N_2467);
and U2540 (N_2540,N_2514,N_2504);
nor U2541 (N_2541,N_2491,N_2469);
or U2542 (N_2542,N_2513,N_2496);
nand U2543 (N_2543,N_2487,N_2500);
nand U2544 (N_2544,N_2507,N_2489);
and U2545 (N_2545,N_2479,N_2494);
and U2546 (N_2546,N_2481,N_2484);
nor U2547 (N_2547,N_2488,N_2468);
nand U2548 (N_2548,N_2499,N_2460);
nand U2549 (N_2549,N_2512,N_2485);
and U2550 (N_2550,N_2514,N_2483);
and U2551 (N_2551,N_2506,N_2474);
and U2552 (N_2552,N_2511,N_2461);
nor U2553 (N_2553,N_2492,N_2519);
or U2554 (N_2554,N_2479,N_2485);
or U2555 (N_2555,N_2486,N_2508);
and U2556 (N_2556,N_2482,N_2473);
nor U2557 (N_2557,N_2460,N_2477);
nand U2558 (N_2558,N_2462,N_2516);
or U2559 (N_2559,N_2461,N_2516);
xor U2560 (N_2560,N_2490,N_2492);
and U2561 (N_2561,N_2510,N_2468);
nor U2562 (N_2562,N_2512,N_2505);
or U2563 (N_2563,N_2465,N_2480);
or U2564 (N_2564,N_2481,N_2470);
nor U2565 (N_2565,N_2501,N_2496);
or U2566 (N_2566,N_2477,N_2502);
nand U2567 (N_2567,N_2508,N_2465);
and U2568 (N_2568,N_2478,N_2492);
nand U2569 (N_2569,N_2487,N_2515);
or U2570 (N_2570,N_2464,N_2502);
nand U2571 (N_2571,N_2506,N_2464);
and U2572 (N_2572,N_2495,N_2514);
nor U2573 (N_2573,N_2484,N_2485);
nor U2574 (N_2574,N_2476,N_2503);
nand U2575 (N_2575,N_2487,N_2506);
and U2576 (N_2576,N_2501,N_2489);
nor U2577 (N_2577,N_2504,N_2461);
nand U2578 (N_2578,N_2515,N_2504);
nor U2579 (N_2579,N_2485,N_2464);
nand U2580 (N_2580,N_2547,N_2570);
and U2581 (N_2581,N_2548,N_2575);
nor U2582 (N_2582,N_2527,N_2564);
and U2583 (N_2583,N_2534,N_2558);
nand U2584 (N_2584,N_2540,N_2553);
nand U2585 (N_2585,N_2526,N_2533);
and U2586 (N_2586,N_2573,N_2552);
and U2587 (N_2587,N_2559,N_2550);
or U2588 (N_2588,N_2565,N_2560);
nand U2589 (N_2589,N_2566,N_2557);
and U2590 (N_2590,N_2562,N_2579);
and U2591 (N_2591,N_2535,N_2536);
nand U2592 (N_2592,N_2567,N_2555);
nor U2593 (N_2593,N_2578,N_2556);
or U2594 (N_2594,N_2537,N_2543);
or U2595 (N_2595,N_2554,N_2561);
nand U2596 (N_2596,N_2528,N_2546);
nor U2597 (N_2597,N_2525,N_2542);
nand U2598 (N_2598,N_2544,N_2521);
nand U2599 (N_2599,N_2577,N_2532);
nor U2600 (N_2600,N_2563,N_2574);
and U2601 (N_2601,N_2522,N_2529);
or U2602 (N_2602,N_2520,N_2568);
and U2603 (N_2603,N_2530,N_2539);
and U2604 (N_2604,N_2571,N_2549);
nor U2605 (N_2605,N_2541,N_2576);
nand U2606 (N_2606,N_2524,N_2545);
nor U2607 (N_2607,N_2569,N_2551);
or U2608 (N_2608,N_2531,N_2538);
nor U2609 (N_2609,N_2523,N_2572);
or U2610 (N_2610,N_2546,N_2537);
nand U2611 (N_2611,N_2525,N_2560);
nand U2612 (N_2612,N_2550,N_2534);
nor U2613 (N_2613,N_2532,N_2547);
nand U2614 (N_2614,N_2522,N_2541);
nor U2615 (N_2615,N_2553,N_2547);
nand U2616 (N_2616,N_2578,N_2550);
or U2617 (N_2617,N_2563,N_2535);
and U2618 (N_2618,N_2530,N_2524);
nor U2619 (N_2619,N_2553,N_2536);
xnor U2620 (N_2620,N_2554,N_2564);
nor U2621 (N_2621,N_2560,N_2531);
nand U2622 (N_2622,N_2530,N_2576);
or U2623 (N_2623,N_2574,N_2566);
nor U2624 (N_2624,N_2531,N_2539);
nand U2625 (N_2625,N_2550,N_2548);
nand U2626 (N_2626,N_2559,N_2551);
or U2627 (N_2627,N_2536,N_2575);
nor U2628 (N_2628,N_2540,N_2536);
nand U2629 (N_2629,N_2524,N_2565);
and U2630 (N_2630,N_2525,N_2570);
or U2631 (N_2631,N_2528,N_2520);
nor U2632 (N_2632,N_2553,N_2566);
or U2633 (N_2633,N_2537,N_2523);
nor U2634 (N_2634,N_2559,N_2572);
or U2635 (N_2635,N_2578,N_2567);
nor U2636 (N_2636,N_2536,N_2546);
nor U2637 (N_2637,N_2577,N_2567);
nor U2638 (N_2638,N_2533,N_2555);
or U2639 (N_2639,N_2520,N_2569);
or U2640 (N_2640,N_2606,N_2581);
nor U2641 (N_2641,N_2612,N_2620);
xnor U2642 (N_2642,N_2592,N_2604);
or U2643 (N_2643,N_2584,N_2601);
or U2644 (N_2644,N_2583,N_2605);
and U2645 (N_2645,N_2627,N_2621);
and U2646 (N_2646,N_2610,N_2624);
nand U2647 (N_2647,N_2586,N_2628);
or U2648 (N_2648,N_2611,N_2619);
nand U2649 (N_2649,N_2591,N_2613);
nand U2650 (N_2650,N_2602,N_2588);
or U2651 (N_2651,N_2622,N_2595);
xnor U2652 (N_2652,N_2632,N_2607);
and U2653 (N_2653,N_2609,N_2598);
nor U2654 (N_2654,N_2608,N_2603);
or U2655 (N_2655,N_2599,N_2615);
or U2656 (N_2656,N_2616,N_2585);
or U2657 (N_2657,N_2617,N_2637);
and U2658 (N_2658,N_2630,N_2633);
nor U2659 (N_2659,N_2629,N_2594);
and U2660 (N_2660,N_2636,N_2600);
and U2661 (N_2661,N_2639,N_2635);
or U2662 (N_2662,N_2587,N_2582);
and U2663 (N_2663,N_2631,N_2597);
and U2664 (N_2664,N_2634,N_2580);
xnor U2665 (N_2665,N_2590,N_2623);
nand U2666 (N_2666,N_2614,N_2596);
or U2667 (N_2667,N_2626,N_2625);
or U2668 (N_2668,N_2618,N_2638);
and U2669 (N_2669,N_2589,N_2593);
or U2670 (N_2670,N_2591,N_2608);
or U2671 (N_2671,N_2611,N_2620);
and U2672 (N_2672,N_2615,N_2619);
or U2673 (N_2673,N_2625,N_2635);
nand U2674 (N_2674,N_2635,N_2626);
and U2675 (N_2675,N_2632,N_2636);
or U2676 (N_2676,N_2596,N_2583);
nor U2677 (N_2677,N_2636,N_2637);
or U2678 (N_2678,N_2603,N_2623);
and U2679 (N_2679,N_2581,N_2608);
nand U2680 (N_2680,N_2619,N_2605);
nand U2681 (N_2681,N_2617,N_2605);
and U2682 (N_2682,N_2619,N_2628);
nand U2683 (N_2683,N_2626,N_2611);
or U2684 (N_2684,N_2590,N_2625);
and U2685 (N_2685,N_2621,N_2624);
or U2686 (N_2686,N_2592,N_2587);
or U2687 (N_2687,N_2601,N_2608);
nand U2688 (N_2688,N_2625,N_2581);
and U2689 (N_2689,N_2629,N_2625);
or U2690 (N_2690,N_2632,N_2585);
nor U2691 (N_2691,N_2637,N_2635);
or U2692 (N_2692,N_2630,N_2614);
nand U2693 (N_2693,N_2593,N_2618);
nor U2694 (N_2694,N_2611,N_2591);
nand U2695 (N_2695,N_2626,N_2627);
or U2696 (N_2696,N_2598,N_2624);
nand U2697 (N_2697,N_2600,N_2592);
or U2698 (N_2698,N_2615,N_2636);
and U2699 (N_2699,N_2627,N_2595);
and U2700 (N_2700,N_2679,N_2655);
or U2701 (N_2701,N_2663,N_2693);
or U2702 (N_2702,N_2683,N_2657);
or U2703 (N_2703,N_2695,N_2678);
or U2704 (N_2704,N_2659,N_2686);
nand U2705 (N_2705,N_2652,N_2661);
nand U2706 (N_2706,N_2680,N_2696);
nor U2707 (N_2707,N_2681,N_2674);
and U2708 (N_2708,N_2665,N_2648);
nand U2709 (N_2709,N_2656,N_2698);
and U2710 (N_2710,N_2662,N_2682);
nand U2711 (N_2711,N_2692,N_2697);
nand U2712 (N_2712,N_2660,N_2669);
nand U2713 (N_2713,N_2649,N_2690);
xnor U2714 (N_2714,N_2670,N_2640);
or U2715 (N_2715,N_2664,N_2688);
or U2716 (N_2716,N_2651,N_2676);
nand U2717 (N_2717,N_2685,N_2689);
nor U2718 (N_2718,N_2645,N_2647);
or U2719 (N_2719,N_2667,N_2687);
and U2720 (N_2720,N_2684,N_2677);
xnor U2721 (N_2721,N_2691,N_2653);
and U2722 (N_2722,N_2666,N_2672);
or U2723 (N_2723,N_2646,N_2654);
nand U2724 (N_2724,N_2650,N_2641);
and U2725 (N_2725,N_2694,N_2673);
xor U2726 (N_2726,N_2644,N_2699);
or U2727 (N_2727,N_2671,N_2668);
nor U2728 (N_2728,N_2642,N_2675);
nor U2729 (N_2729,N_2643,N_2658);
or U2730 (N_2730,N_2660,N_2678);
and U2731 (N_2731,N_2662,N_2649);
nor U2732 (N_2732,N_2690,N_2670);
nand U2733 (N_2733,N_2650,N_2693);
nand U2734 (N_2734,N_2662,N_2672);
nor U2735 (N_2735,N_2669,N_2655);
nor U2736 (N_2736,N_2698,N_2662);
nand U2737 (N_2737,N_2673,N_2676);
nor U2738 (N_2738,N_2665,N_2653);
nand U2739 (N_2739,N_2668,N_2689);
or U2740 (N_2740,N_2683,N_2691);
and U2741 (N_2741,N_2685,N_2645);
or U2742 (N_2742,N_2642,N_2647);
nor U2743 (N_2743,N_2643,N_2642);
and U2744 (N_2744,N_2652,N_2688);
or U2745 (N_2745,N_2653,N_2680);
or U2746 (N_2746,N_2685,N_2661);
nor U2747 (N_2747,N_2643,N_2693);
or U2748 (N_2748,N_2665,N_2688);
and U2749 (N_2749,N_2690,N_2677);
nor U2750 (N_2750,N_2659,N_2684);
and U2751 (N_2751,N_2691,N_2663);
and U2752 (N_2752,N_2687,N_2644);
or U2753 (N_2753,N_2678,N_2643);
nand U2754 (N_2754,N_2676,N_2661);
nand U2755 (N_2755,N_2648,N_2683);
or U2756 (N_2756,N_2673,N_2686);
or U2757 (N_2757,N_2696,N_2655);
nand U2758 (N_2758,N_2645,N_2649);
nand U2759 (N_2759,N_2681,N_2665);
or U2760 (N_2760,N_2733,N_2710);
and U2761 (N_2761,N_2724,N_2737);
nor U2762 (N_2762,N_2756,N_2714);
nand U2763 (N_2763,N_2736,N_2731);
or U2764 (N_2764,N_2757,N_2708);
nand U2765 (N_2765,N_2706,N_2721);
xnor U2766 (N_2766,N_2741,N_2744);
or U2767 (N_2767,N_2726,N_2720);
nor U2768 (N_2768,N_2700,N_2742);
nor U2769 (N_2769,N_2723,N_2743);
and U2770 (N_2770,N_2717,N_2747);
nand U2771 (N_2771,N_2718,N_2754);
or U2772 (N_2772,N_2725,N_2701);
nand U2773 (N_2773,N_2729,N_2752);
and U2774 (N_2774,N_2722,N_2746);
or U2775 (N_2775,N_2728,N_2707);
nand U2776 (N_2776,N_2759,N_2703);
nor U2777 (N_2777,N_2758,N_2713);
or U2778 (N_2778,N_2732,N_2745);
nor U2779 (N_2779,N_2734,N_2711);
and U2780 (N_2780,N_2727,N_2702);
nor U2781 (N_2781,N_2751,N_2705);
xnor U2782 (N_2782,N_2750,N_2715);
or U2783 (N_2783,N_2730,N_2712);
or U2784 (N_2784,N_2740,N_2753);
nand U2785 (N_2785,N_2719,N_2709);
nor U2786 (N_2786,N_2738,N_2755);
or U2787 (N_2787,N_2704,N_2739);
and U2788 (N_2788,N_2716,N_2749);
or U2789 (N_2789,N_2748,N_2735);
nor U2790 (N_2790,N_2748,N_2711);
and U2791 (N_2791,N_2710,N_2738);
nand U2792 (N_2792,N_2742,N_2736);
nand U2793 (N_2793,N_2731,N_2725);
nand U2794 (N_2794,N_2754,N_2710);
nor U2795 (N_2795,N_2717,N_2702);
and U2796 (N_2796,N_2742,N_2729);
or U2797 (N_2797,N_2705,N_2753);
or U2798 (N_2798,N_2733,N_2735);
nor U2799 (N_2799,N_2710,N_2740);
or U2800 (N_2800,N_2751,N_2728);
nand U2801 (N_2801,N_2719,N_2701);
or U2802 (N_2802,N_2713,N_2716);
nor U2803 (N_2803,N_2736,N_2737);
nand U2804 (N_2804,N_2742,N_2706);
nand U2805 (N_2805,N_2712,N_2738);
nor U2806 (N_2806,N_2738,N_2734);
and U2807 (N_2807,N_2759,N_2712);
and U2808 (N_2808,N_2753,N_2717);
and U2809 (N_2809,N_2752,N_2727);
nand U2810 (N_2810,N_2714,N_2701);
and U2811 (N_2811,N_2759,N_2707);
nand U2812 (N_2812,N_2754,N_2731);
and U2813 (N_2813,N_2709,N_2701);
or U2814 (N_2814,N_2736,N_2724);
nand U2815 (N_2815,N_2739,N_2752);
nor U2816 (N_2816,N_2717,N_2712);
xnor U2817 (N_2817,N_2722,N_2749);
nor U2818 (N_2818,N_2710,N_2737);
or U2819 (N_2819,N_2742,N_2741);
and U2820 (N_2820,N_2791,N_2775);
nor U2821 (N_2821,N_2804,N_2762);
nor U2822 (N_2822,N_2763,N_2803);
or U2823 (N_2823,N_2784,N_2767);
nor U2824 (N_2824,N_2764,N_2806);
nand U2825 (N_2825,N_2812,N_2807);
or U2826 (N_2826,N_2818,N_2815);
and U2827 (N_2827,N_2785,N_2805);
nand U2828 (N_2828,N_2776,N_2814);
and U2829 (N_2829,N_2801,N_2810);
nand U2830 (N_2830,N_2813,N_2819);
nor U2831 (N_2831,N_2798,N_2772);
and U2832 (N_2832,N_2792,N_2760);
nand U2833 (N_2833,N_2777,N_2808);
and U2834 (N_2834,N_2797,N_2794);
and U2835 (N_2835,N_2817,N_2788);
or U2836 (N_2836,N_2789,N_2766);
or U2837 (N_2837,N_2770,N_2786);
nand U2838 (N_2838,N_2761,N_2799);
and U2839 (N_2839,N_2795,N_2768);
or U2840 (N_2840,N_2793,N_2790);
or U2841 (N_2841,N_2778,N_2787);
or U2842 (N_2842,N_2769,N_2811);
or U2843 (N_2843,N_2802,N_2780);
nor U2844 (N_2844,N_2800,N_2816);
xor U2845 (N_2845,N_2782,N_2779);
nand U2846 (N_2846,N_2783,N_2773);
and U2847 (N_2847,N_2774,N_2781);
nand U2848 (N_2848,N_2771,N_2809);
or U2849 (N_2849,N_2765,N_2796);
and U2850 (N_2850,N_2764,N_2787);
and U2851 (N_2851,N_2806,N_2773);
nor U2852 (N_2852,N_2818,N_2809);
and U2853 (N_2853,N_2814,N_2787);
or U2854 (N_2854,N_2793,N_2775);
and U2855 (N_2855,N_2768,N_2796);
and U2856 (N_2856,N_2772,N_2789);
nor U2857 (N_2857,N_2794,N_2781);
nand U2858 (N_2858,N_2790,N_2768);
and U2859 (N_2859,N_2806,N_2781);
and U2860 (N_2860,N_2812,N_2817);
nand U2861 (N_2861,N_2814,N_2798);
or U2862 (N_2862,N_2773,N_2777);
nand U2863 (N_2863,N_2788,N_2794);
nor U2864 (N_2864,N_2763,N_2775);
nand U2865 (N_2865,N_2798,N_2761);
nor U2866 (N_2866,N_2763,N_2808);
or U2867 (N_2867,N_2798,N_2776);
nor U2868 (N_2868,N_2769,N_2809);
or U2869 (N_2869,N_2773,N_2782);
and U2870 (N_2870,N_2813,N_2774);
and U2871 (N_2871,N_2777,N_2763);
nand U2872 (N_2872,N_2794,N_2767);
nor U2873 (N_2873,N_2802,N_2764);
and U2874 (N_2874,N_2779,N_2796);
nor U2875 (N_2875,N_2798,N_2782);
or U2876 (N_2876,N_2807,N_2808);
and U2877 (N_2877,N_2799,N_2774);
or U2878 (N_2878,N_2783,N_2813);
nand U2879 (N_2879,N_2768,N_2816);
and U2880 (N_2880,N_2855,N_2840);
nand U2881 (N_2881,N_2847,N_2843);
and U2882 (N_2882,N_2873,N_2828);
or U2883 (N_2883,N_2820,N_2878);
and U2884 (N_2884,N_2858,N_2846);
xor U2885 (N_2885,N_2879,N_2845);
nor U2886 (N_2886,N_2838,N_2822);
nand U2887 (N_2887,N_2848,N_2837);
xor U2888 (N_2888,N_2844,N_2870);
nor U2889 (N_2889,N_2859,N_2824);
xnor U2890 (N_2890,N_2875,N_2866);
and U2891 (N_2891,N_2821,N_2854);
nor U2892 (N_2892,N_2852,N_2874);
xor U2893 (N_2893,N_2856,N_2860);
and U2894 (N_2894,N_2867,N_2872);
nand U2895 (N_2895,N_2829,N_2850);
nand U2896 (N_2896,N_2861,N_2827);
nor U2897 (N_2897,N_2834,N_2841);
nand U2898 (N_2898,N_2830,N_2836);
nand U2899 (N_2899,N_2823,N_2853);
nand U2900 (N_2900,N_2862,N_2857);
nor U2901 (N_2901,N_2877,N_2868);
and U2902 (N_2902,N_2865,N_2826);
nand U2903 (N_2903,N_2851,N_2849);
nand U2904 (N_2904,N_2871,N_2835);
and U2905 (N_2905,N_2869,N_2839);
nand U2906 (N_2906,N_2864,N_2832);
nand U2907 (N_2907,N_2876,N_2831);
xnor U2908 (N_2908,N_2825,N_2863);
xnor U2909 (N_2909,N_2833,N_2842);
and U2910 (N_2910,N_2851,N_2835);
nor U2911 (N_2911,N_2843,N_2844);
nand U2912 (N_2912,N_2872,N_2845);
nand U2913 (N_2913,N_2834,N_2870);
and U2914 (N_2914,N_2859,N_2872);
nand U2915 (N_2915,N_2846,N_2854);
or U2916 (N_2916,N_2829,N_2865);
or U2917 (N_2917,N_2824,N_2855);
and U2918 (N_2918,N_2832,N_2870);
nand U2919 (N_2919,N_2868,N_2848);
and U2920 (N_2920,N_2824,N_2853);
nor U2921 (N_2921,N_2839,N_2858);
or U2922 (N_2922,N_2875,N_2842);
and U2923 (N_2923,N_2866,N_2827);
nand U2924 (N_2924,N_2836,N_2820);
or U2925 (N_2925,N_2830,N_2853);
xnor U2926 (N_2926,N_2840,N_2848);
and U2927 (N_2927,N_2832,N_2837);
and U2928 (N_2928,N_2849,N_2827);
nor U2929 (N_2929,N_2850,N_2862);
nand U2930 (N_2930,N_2848,N_2867);
nor U2931 (N_2931,N_2827,N_2864);
or U2932 (N_2932,N_2852,N_2873);
nor U2933 (N_2933,N_2869,N_2860);
nand U2934 (N_2934,N_2846,N_2875);
or U2935 (N_2935,N_2826,N_2856);
or U2936 (N_2936,N_2861,N_2864);
nand U2937 (N_2937,N_2828,N_2852);
nor U2938 (N_2938,N_2860,N_2826);
xnor U2939 (N_2939,N_2828,N_2835);
nand U2940 (N_2940,N_2904,N_2888);
and U2941 (N_2941,N_2912,N_2884);
and U2942 (N_2942,N_2935,N_2903);
or U2943 (N_2943,N_2899,N_2898);
or U2944 (N_2944,N_2891,N_2909);
nor U2945 (N_2945,N_2924,N_2881);
and U2946 (N_2946,N_2893,N_2892);
and U2947 (N_2947,N_2927,N_2897);
nor U2948 (N_2948,N_2933,N_2887);
and U2949 (N_2949,N_2905,N_2907);
or U2950 (N_2950,N_2908,N_2900);
nor U2951 (N_2951,N_2917,N_2915);
nor U2952 (N_2952,N_2921,N_2931);
and U2953 (N_2953,N_2882,N_2902);
nand U2954 (N_2954,N_2913,N_2929);
xor U2955 (N_2955,N_2886,N_2937);
nor U2956 (N_2956,N_2920,N_2883);
and U2957 (N_2957,N_2910,N_2932);
and U2958 (N_2958,N_2926,N_2885);
nor U2959 (N_2959,N_2925,N_2914);
and U2960 (N_2960,N_2906,N_2916);
and U2961 (N_2961,N_2895,N_2928);
and U2962 (N_2962,N_2939,N_2930);
nand U2963 (N_2963,N_2880,N_2923);
nand U2964 (N_2964,N_2894,N_2890);
nand U2965 (N_2965,N_2889,N_2919);
or U2966 (N_2966,N_2896,N_2911);
nor U2967 (N_2967,N_2938,N_2922);
nand U2968 (N_2968,N_2934,N_2901);
nor U2969 (N_2969,N_2918,N_2936);
and U2970 (N_2970,N_2911,N_2887);
xor U2971 (N_2971,N_2896,N_2891);
or U2972 (N_2972,N_2912,N_2894);
nor U2973 (N_2973,N_2890,N_2923);
nand U2974 (N_2974,N_2883,N_2928);
nand U2975 (N_2975,N_2895,N_2899);
and U2976 (N_2976,N_2884,N_2917);
and U2977 (N_2977,N_2903,N_2893);
or U2978 (N_2978,N_2912,N_2932);
or U2979 (N_2979,N_2937,N_2903);
and U2980 (N_2980,N_2935,N_2906);
and U2981 (N_2981,N_2922,N_2917);
nor U2982 (N_2982,N_2889,N_2902);
and U2983 (N_2983,N_2901,N_2891);
or U2984 (N_2984,N_2883,N_2904);
or U2985 (N_2985,N_2883,N_2933);
nand U2986 (N_2986,N_2899,N_2883);
nand U2987 (N_2987,N_2897,N_2911);
nand U2988 (N_2988,N_2893,N_2930);
nor U2989 (N_2989,N_2885,N_2902);
and U2990 (N_2990,N_2920,N_2928);
or U2991 (N_2991,N_2906,N_2904);
nand U2992 (N_2992,N_2884,N_2939);
nor U2993 (N_2993,N_2919,N_2917);
nor U2994 (N_2994,N_2924,N_2901);
or U2995 (N_2995,N_2918,N_2906);
nand U2996 (N_2996,N_2916,N_2929);
nor U2997 (N_2997,N_2920,N_2901);
or U2998 (N_2998,N_2930,N_2902);
nand U2999 (N_2999,N_2937,N_2894);
nand UO_0 (O_0,N_2994,N_2948);
nand UO_1 (O_1,N_2964,N_2956);
and UO_2 (O_2,N_2979,N_2947);
or UO_3 (O_3,N_2953,N_2959);
and UO_4 (O_4,N_2992,N_2972);
nor UO_5 (O_5,N_2984,N_2970);
nor UO_6 (O_6,N_2975,N_2997);
nand UO_7 (O_7,N_2941,N_2976);
nor UO_8 (O_8,N_2955,N_2962);
or UO_9 (O_9,N_2973,N_2977);
and UO_10 (O_10,N_2993,N_2985);
and UO_11 (O_11,N_2991,N_2988);
or UO_12 (O_12,N_2946,N_2942);
or UO_13 (O_13,N_2978,N_2967);
nand UO_14 (O_14,N_2957,N_2961);
and UO_15 (O_15,N_2983,N_2980);
nor UO_16 (O_16,N_2969,N_2952);
and UO_17 (O_17,N_2954,N_2944);
or UO_18 (O_18,N_2963,N_2989);
and UO_19 (O_19,N_2958,N_2950);
and UO_20 (O_20,N_2949,N_2968);
nor UO_21 (O_21,N_2995,N_2981);
nand UO_22 (O_22,N_2974,N_2951);
or UO_23 (O_23,N_2982,N_2999);
nand UO_24 (O_24,N_2966,N_2996);
or UO_25 (O_25,N_2971,N_2990);
nor UO_26 (O_26,N_2998,N_2940);
or UO_27 (O_27,N_2986,N_2945);
or UO_28 (O_28,N_2965,N_2960);
or UO_29 (O_29,N_2987,N_2943);
and UO_30 (O_30,N_2961,N_2944);
nor UO_31 (O_31,N_2976,N_2954);
nor UO_32 (O_32,N_2950,N_2970);
and UO_33 (O_33,N_2986,N_2941);
and UO_34 (O_34,N_2981,N_2942);
nand UO_35 (O_35,N_2961,N_2974);
and UO_36 (O_36,N_2971,N_2977);
and UO_37 (O_37,N_2996,N_2975);
and UO_38 (O_38,N_2983,N_2986);
nand UO_39 (O_39,N_2981,N_2970);
nor UO_40 (O_40,N_2970,N_2946);
and UO_41 (O_41,N_2940,N_2975);
and UO_42 (O_42,N_2966,N_2964);
and UO_43 (O_43,N_2995,N_2991);
nor UO_44 (O_44,N_2989,N_2961);
and UO_45 (O_45,N_2945,N_2961);
and UO_46 (O_46,N_2959,N_2981);
and UO_47 (O_47,N_2994,N_2965);
nor UO_48 (O_48,N_2951,N_2965);
or UO_49 (O_49,N_2960,N_2957);
or UO_50 (O_50,N_2952,N_2947);
and UO_51 (O_51,N_2979,N_2996);
or UO_52 (O_52,N_2961,N_2941);
nand UO_53 (O_53,N_2940,N_2955);
or UO_54 (O_54,N_2943,N_2954);
nor UO_55 (O_55,N_2967,N_2973);
or UO_56 (O_56,N_2990,N_2943);
or UO_57 (O_57,N_2950,N_2994);
or UO_58 (O_58,N_2985,N_2964);
nor UO_59 (O_59,N_2941,N_2960);
nand UO_60 (O_60,N_2942,N_2954);
xor UO_61 (O_61,N_2957,N_2959);
nand UO_62 (O_62,N_2971,N_2945);
nand UO_63 (O_63,N_2971,N_2959);
or UO_64 (O_64,N_2953,N_2957);
or UO_65 (O_65,N_2978,N_2965);
and UO_66 (O_66,N_2964,N_2994);
nor UO_67 (O_67,N_2996,N_2963);
nand UO_68 (O_68,N_2959,N_2952);
nand UO_69 (O_69,N_2993,N_2998);
or UO_70 (O_70,N_2985,N_2981);
and UO_71 (O_71,N_2949,N_2997);
or UO_72 (O_72,N_2956,N_2974);
and UO_73 (O_73,N_2957,N_2944);
or UO_74 (O_74,N_2942,N_2959);
nand UO_75 (O_75,N_2940,N_2984);
and UO_76 (O_76,N_2995,N_2967);
or UO_77 (O_77,N_2957,N_2991);
nand UO_78 (O_78,N_2993,N_2976);
or UO_79 (O_79,N_2941,N_2962);
xnor UO_80 (O_80,N_2959,N_2946);
nor UO_81 (O_81,N_2991,N_2975);
and UO_82 (O_82,N_2993,N_2942);
or UO_83 (O_83,N_2943,N_2984);
nand UO_84 (O_84,N_2982,N_2943);
or UO_85 (O_85,N_2956,N_2962);
or UO_86 (O_86,N_2994,N_2990);
or UO_87 (O_87,N_2989,N_2977);
and UO_88 (O_88,N_2973,N_2952);
or UO_89 (O_89,N_2963,N_2977);
nand UO_90 (O_90,N_2973,N_2998);
or UO_91 (O_91,N_2997,N_2955);
nand UO_92 (O_92,N_2995,N_2962);
and UO_93 (O_93,N_2958,N_2947);
or UO_94 (O_94,N_2981,N_2994);
xor UO_95 (O_95,N_2954,N_2940);
nor UO_96 (O_96,N_2975,N_2976);
and UO_97 (O_97,N_2962,N_2989);
or UO_98 (O_98,N_2987,N_2975);
and UO_99 (O_99,N_2987,N_2948);
xor UO_100 (O_100,N_2940,N_2983);
nor UO_101 (O_101,N_2996,N_2956);
nand UO_102 (O_102,N_2947,N_2973);
nor UO_103 (O_103,N_2995,N_2999);
and UO_104 (O_104,N_2951,N_2980);
or UO_105 (O_105,N_2949,N_2988);
and UO_106 (O_106,N_2970,N_2969);
or UO_107 (O_107,N_2987,N_2997);
or UO_108 (O_108,N_2975,N_2949);
nand UO_109 (O_109,N_2994,N_2978);
nand UO_110 (O_110,N_2977,N_2978);
nand UO_111 (O_111,N_2978,N_2957);
nor UO_112 (O_112,N_2963,N_2950);
or UO_113 (O_113,N_2946,N_2992);
nand UO_114 (O_114,N_2987,N_2974);
and UO_115 (O_115,N_2990,N_2953);
or UO_116 (O_116,N_2952,N_2967);
and UO_117 (O_117,N_2996,N_2969);
nor UO_118 (O_118,N_2992,N_2980);
nor UO_119 (O_119,N_2986,N_2940);
or UO_120 (O_120,N_2947,N_2957);
nand UO_121 (O_121,N_2999,N_2963);
and UO_122 (O_122,N_2940,N_2946);
or UO_123 (O_123,N_2998,N_2981);
and UO_124 (O_124,N_2982,N_2970);
nand UO_125 (O_125,N_2975,N_2953);
nand UO_126 (O_126,N_2969,N_2986);
nand UO_127 (O_127,N_2983,N_2977);
xnor UO_128 (O_128,N_2995,N_2990);
nand UO_129 (O_129,N_2953,N_2999);
nand UO_130 (O_130,N_2951,N_2959);
or UO_131 (O_131,N_2965,N_2950);
nand UO_132 (O_132,N_2996,N_2978);
or UO_133 (O_133,N_2991,N_2992);
xor UO_134 (O_134,N_2972,N_2953);
nand UO_135 (O_135,N_2996,N_2993);
or UO_136 (O_136,N_2979,N_2966);
nor UO_137 (O_137,N_2983,N_2987);
nor UO_138 (O_138,N_2956,N_2943);
and UO_139 (O_139,N_2940,N_2964);
nor UO_140 (O_140,N_2957,N_2988);
and UO_141 (O_141,N_2954,N_2957);
and UO_142 (O_142,N_2971,N_2994);
or UO_143 (O_143,N_2957,N_2949);
or UO_144 (O_144,N_2966,N_2987);
and UO_145 (O_145,N_2981,N_2979);
nor UO_146 (O_146,N_2997,N_2974);
nor UO_147 (O_147,N_2941,N_2966);
or UO_148 (O_148,N_2988,N_2968);
or UO_149 (O_149,N_2991,N_2985);
xnor UO_150 (O_150,N_2994,N_2974);
or UO_151 (O_151,N_2953,N_2997);
and UO_152 (O_152,N_2956,N_2967);
or UO_153 (O_153,N_2987,N_2946);
or UO_154 (O_154,N_2941,N_2948);
xnor UO_155 (O_155,N_2958,N_2988);
and UO_156 (O_156,N_2993,N_2997);
nand UO_157 (O_157,N_2942,N_2945);
nor UO_158 (O_158,N_2996,N_2944);
nor UO_159 (O_159,N_2982,N_2958);
nand UO_160 (O_160,N_2988,N_2963);
nor UO_161 (O_161,N_2960,N_2975);
or UO_162 (O_162,N_2968,N_2971);
nor UO_163 (O_163,N_2980,N_2993);
nor UO_164 (O_164,N_2961,N_2946);
nor UO_165 (O_165,N_2960,N_2983);
xnor UO_166 (O_166,N_2948,N_2966);
and UO_167 (O_167,N_2943,N_2953);
and UO_168 (O_168,N_2950,N_2968);
or UO_169 (O_169,N_2989,N_2983);
xor UO_170 (O_170,N_2980,N_2945);
and UO_171 (O_171,N_2996,N_2965);
or UO_172 (O_172,N_2994,N_2988);
or UO_173 (O_173,N_2948,N_2943);
or UO_174 (O_174,N_2994,N_2996);
xnor UO_175 (O_175,N_2946,N_2991);
or UO_176 (O_176,N_2948,N_2940);
nand UO_177 (O_177,N_2957,N_2951);
nor UO_178 (O_178,N_2954,N_2946);
and UO_179 (O_179,N_2997,N_2940);
and UO_180 (O_180,N_2953,N_2951);
or UO_181 (O_181,N_2941,N_2993);
and UO_182 (O_182,N_2942,N_2986);
nor UO_183 (O_183,N_2972,N_2955);
or UO_184 (O_184,N_2977,N_2953);
or UO_185 (O_185,N_2943,N_2955);
nand UO_186 (O_186,N_2947,N_2985);
xnor UO_187 (O_187,N_2994,N_2980);
nand UO_188 (O_188,N_2970,N_2954);
nor UO_189 (O_189,N_2966,N_2940);
or UO_190 (O_190,N_2977,N_2994);
nor UO_191 (O_191,N_2980,N_2997);
nand UO_192 (O_192,N_2978,N_2995);
nand UO_193 (O_193,N_2998,N_2992);
nor UO_194 (O_194,N_2956,N_2941);
nor UO_195 (O_195,N_2971,N_2943);
nand UO_196 (O_196,N_2972,N_2999);
or UO_197 (O_197,N_2949,N_2984);
nor UO_198 (O_198,N_2965,N_2986);
nor UO_199 (O_199,N_2999,N_2967);
nand UO_200 (O_200,N_2959,N_2961);
and UO_201 (O_201,N_2991,N_2987);
nor UO_202 (O_202,N_2965,N_2999);
and UO_203 (O_203,N_2968,N_2997);
and UO_204 (O_204,N_2953,N_2993);
and UO_205 (O_205,N_2974,N_2960);
nand UO_206 (O_206,N_2947,N_2943);
or UO_207 (O_207,N_2958,N_2998);
or UO_208 (O_208,N_2956,N_2973);
and UO_209 (O_209,N_2941,N_2972);
and UO_210 (O_210,N_2951,N_2994);
and UO_211 (O_211,N_2983,N_2997);
nand UO_212 (O_212,N_2999,N_2956);
nor UO_213 (O_213,N_2990,N_2970);
nand UO_214 (O_214,N_2951,N_2975);
nor UO_215 (O_215,N_2967,N_2955);
and UO_216 (O_216,N_2979,N_2982);
or UO_217 (O_217,N_2966,N_2957);
or UO_218 (O_218,N_2966,N_2944);
nand UO_219 (O_219,N_2953,N_2946);
or UO_220 (O_220,N_2996,N_2989);
nor UO_221 (O_221,N_2995,N_2969);
nor UO_222 (O_222,N_2964,N_2996);
nor UO_223 (O_223,N_2978,N_2956);
nor UO_224 (O_224,N_2974,N_2943);
or UO_225 (O_225,N_2956,N_2987);
and UO_226 (O_226,N_2995,N_2949);
nand UO_227 (O_227,N_2998,N_2950);
or UO_228 (O_228,N_2968,N_2995);
and UO_229 (O_229,N_2990,N_2991);
and UO_230 (O_230,N_2944,N_2985);
nand UO_231 (O_231,N_2974,N_2945);
and UO_232 (O_232,N_2955,N_2995);
or UO_233 (O_233,N_2949,N_2991);
nand UO_234 (O_234,N_2949,N_2945);
or UO_235 (O_235,N_2941,N_2951);
or UO_236 (O_236,N_2955,N_2998);
nand UO_237 (O_237,N_2952,N_2988);
nor UO_238 (O_238,N_2972,N_2978);
and UO_239 (O_239,N_2993,N_2967);
or UO_240 (O_240,N_2961,N_2963);
or UO_241 (O_241,N_2984,N_2953);
nand UO_242 (O_242,N_2967,N_2970);
xor UO_243 (O_243,N_2955,N_2976);
xnor UO_244 (O_244,N_2958,N_2942);
nor UO_245 (O_245,N_2999,N_2986);
nand UO_246 (O_246,N_2996,N_2972);
or UO_247 (O_247,N_2971,N_2965);
nor UO_248 (O_248,N_2964,N_2970);
nand UO_249 (O_249,N_2960,N_2943);
or UO_250 (O_250,N_2994,N_2940);
or UO_251 (O_251,N_2968,N_2977);
nand UO_252 (O_252,N_2959,N_2982);
nand UO_253 (O_253,N_2999,N_2945);
nor UO_254 (O_254,N_2967,N_2979);
and UO_255 (O_255,N_2968,N_2951);
nand UO_256 (O_256,N_2945,N_2948);
or UO_257 (O_257,N_2971,N_2962);
nand UO_258 (O_258,N_2989,N_2988);
and UO_259 (O_259,N_2994,N_2966);
nor UO_260 (O_260,N_2959,N_2949);
nand UO_261 (O_261,N_2972,N_2989);
nand UO_262 (O_262,N_2971,N_2952);
or UO_263 (O_263,N_2956,N_2988);
xnor UO_264 (O_264,N_2985,N_2949);
nand UO_265 (O_265,N_2983,N_2970);
and UO_266 (O_266,N_2973,N_2996);
and UO_267 (O_267,N_2952,N_2993);
and UO_268 (O_268,N_2968,N_2947);
nand UO_269 (O_269,N_2945,N_2975);
nor UO_270 (O_270,N_2947,N_2988);
nor UO_271 (O_271,N_2950,N_2985);
or UO_272 (O_272,N_2989,N_2945);
nor UO_273 (O_273,N_2951,N_2973);
nor UO_274 (O_274,N_2941,N_2965);
or UO_275 (O_275,N_2950,N_2960);
nor UO_276 (O_276,N_2966,N_2977);
and UO_277 (O_277,N_2965,N_2972);
nor UO_278 (O_278,N_2999,N_2957);
nand UO_279 (O_279,N_2946,N_2963);
nand UO_280 (O_280,N_2968,N_2994);
nand UO_281 (O_281,N_2954,N_2941);
or UO_282 (O_282,N_2940,N_2988);
nand UO_283 (O_283,N_2993,N_2956);
or UO_284 (O_284,N_2962,N_2946);
nor UO_285 (O_285,N_2960,N_2979);
nand UO_286 (O_286,N_2977,N_2997);
or UO_287 (O_287,N_2963,N_2997);
and UO_288 (O_288,N_2953,N_2952);
and UO_289 (O_289,N_2958,N_2985);
nand UO_290 (O_290,N_2982,N_2946);
nand UO_291 (O_291,N_2947,N_2940);
or UO_292 (O_292,N_2950,N_2952);
nor UO_293 (O_293,N_2962,N_2979);
xor UO_294 (O_294,N_2971,N_2988);
or UO_295 (O_295,N_2992,N_2967);
or UO_296 (O_296,N_2952,N_2974);
nand UO_297 (O_297,N_2999,N_2968);
and UO_298 (O_298,N_2988,N_2974);
nor UO_299 (O_299,N_2953,N_2948);
and UO_300 (O_300,N_2985,N_2999);
and UO_301 (O_301,N_2975,N_2971);
and UO_302 (O_302,N_2967,N_2953);
and UO_303 (O_303,N_2961,N_2954);
and UO_304 (O_304,N_2988,N_2966);
nand UO_305 (O_305,N_2987,N_2950);
or UO_306 (O_306,N_2965,N_2947);
or UO_307 (O_307,N_2954,N_2995);
nand UO_308 (O_308,N_2957,N_2992);
nand UO_309 (O_309,N_2968,N_2989);
and UO_310 (O_310,N_2992,N_2968);
nor UO_311 (O_311,N_2989,N_2998);
and UO_312 (O_312,N_2963,N_2982);
nand UO_313 (O_313,N_2980,N_2940);
or UO_314 (O_314,N_2996,N_2982);
and UO_315 (O_315,N_2944,N_2949);
nand UO_316 (O_316,N_2982,N_2984);
nor UO_317 (O_317,N_2967,N_2977);
or UO_318 (O_318,N_2973,N_2988);
nor UO_319 (O_319,N_2967,N_2941);
nor UO_320 (O_320,N_2947,N_2969);
nand UO_321 (O_321,N_2955,N_2963);
nor UO_322 (O_322,N_2952,N_2941);
nor UO_323 (O_323,N_2955,N_2981);
or UO_324 (O_324,N_2989,N_2975);
or UO_325 (O_325,N_2987,N_2981);
nand UO_326 (O_326,N_2982,N_2954);
and UO_327 (O_327,N_2956,N_2955);
and UO_328 (O_328,N_2955,N_2942);
and UO_329 (O_329,N_2995,N_2971);
or UO_330 (O_330,N_2958,N_2956);
or UO_331 (O_331,N_2942,N_2948);
and UO_332 (O_332,N_2947,N_2970);
nand UO_333 (O_333,N_2998,N_2965);
nor UO_334 (O_334,N_2947,N_2994);
nor UO_335 (O_335,N_2995,N_2997);
and UO_336 (O_336,N_2966,N_2995);
or UO_337 (O_337,N_2985,N_2998);
or UO_338 (O_338,N_2951,N_2962);
or UO_339 (O_339,N_2985,N_2955);
and UO_340 (O_340,N_2970,N_2962);
and UO_341 (O_341,N_2979,N_2984);
nor UO_342 (O_342,N_2991,N_2956);
or UO_343 (O_343,N_2993,N_2964);
nand UO_344 (O_344,N_2968,N_2980);
and UO_345 (O_345,N_2973,N_2981);
or UO_346 (O_346,N_2974,N_2946);
and UO_347 (O_347,N_2961,N_2992);
nand UO_348 (O_348,N_2977,N_2940);
nor UO_349 (O_349,N_2964,N_2995);
nand UO_350 (O_350,N_2998,N_2999);
and UO_351 (O_351,N_2954,N_2991);
and UO_352 (O_352,N_2945,N_2969);
nor UO_353 (O_353,N_2971,N_2991);
nand UO_354 (O_354,N_2943,N_2967);
nand UO_355 (O_355,N_2959,N_2999);
nor UO_356 (O_356,N_2995,N_2974);
nand UO_357 (O_357,N_2973,N_2984);
or UO_358 (O_358,N_2986,N_2966);
nor UO_359 (O_359,N_2996,N_2984);
nor UO_360 (O_360,N_2983,N_2992);
nor UO_361 (O_361,N_2943,N_2998);
and UO_362 (O_362,N_2971,N_2967);
nor UO_363 (O_363,N_2990,N_2974);
nand UO_364 (O_364,N_2964,N_2990);
nor UO_365 (O_365,N_2968,N_2958);
and UO_366 (O_366,N_2956,N_2952);
or UO_367 (O_367,N_2940,N_2945);
nor UO_368 (O_368,N_2956,N_2946);
and UO_369 (O_369,N_2950,N_2991);
or UO_370 (O_370,N_2986,N_2953);
nor UO_371 (O_371,N_2983,N_2991);
nand UO_372 (O_372,N_2953,N_2965);
and UO_373 (O_373,N_2974,N_2977);
and UO_374 (O_374,N_2972,N_2966);
nand UO_375 (O_375,N_2999,N_2966);
and UO_376 (O_376,N_2942,N_2983);
and UO_377 (O_377,N_2989,N_2964);
nor UO_378 (O_378,N_2984,N_2942);
nor UO_379 (O_379,N_2990,N_2940);
or UO_380 (O_380,N_2976,N_2995);
or UO_381 (O_381,N_2959,N_2940);
nor UO_382 (O_382,N_2963,N_2959);
nor UO_383 (O_383,N_2959,N_2976);
or UO_384 (O_384,N_2946,N_2985);
and UO_385 (O_385,N_2975,N_2998);
or UO_386 (O_386,N_2978,N_2960);
and UO_387 (O_387,N_2979,N_2983);
or UO_388 (O_388,N_2970,N_2966);
or UO_389 (O_389,N_2973,N_2971);
nor UO_390 (O_390,N_2942,N_2989);
nand UO_391 (O_391,N_2985,N_2967);
nand UO_392 (O_392,N_2961,N_2975);
nand UO_393 (O_393,N_2970,N_2973);
nand UO_394 (O_394,N_2940,N_2979);
nor UO_395 (O_395,N_2995,N_2983);
or UO_396 (O_396,N_2954,N_2987);
and UO_397 (O_397,N_2978,N_2985);
nand UO_398 (O_398,N_2996,N_2948);
nor UO_399 (O_399,N_2942,N_2971);
and UO_400 (O_400,N_2957,N_2948);
nand UO_401 (O_401,N_2975,N_2948);
and UO_402 (O_402,N_2998,N_2967);
or UO_403 (O_403,N_2956,N_2954);
or UO_404 (O_404,N_2975,N_2995);
or UO_405 (O_405,N_2977,N_2962);
xnor UO_406 (O_406,N_2964,N_2988);
and UO_407 (O_407,N_2981,N_2974);
or UO_408 (O_408,N_2951,N_2996);
and UO_409 (O_409,N_2986,N_2972);
and UO_410 (O_410,N_2984,N_2963);
or UO_411 (O_411,N_2981,N_2954);
nand UO_412 (O_412,N_2993,N_2981);
and UO_413 (O_413,N_2987,N_2960);
nand UO_414 (O_414,N_2964,N_2952);
or UO_415 (O_415,N_2973,N_2995);
nand UO_416 (O_416,N_2996,N_2968);
nand UO_417 (O_417,N_2992,N_2943);
or UO_418 (O_418,N_2997,N_2990);
nor UO_419 (O_419,N_2991,N_2953);
nand UO_420 (O_420,N_2963,N_2998);
and UO_421 (O_421,N_2978,N_2986);
or UO_422 (O_422,N_2992,N_2963);
nor UO_423 (O_423,N_2978,N_2971);
and UO_424 (O_424,N_2948,N_2993);
nor UO_425 (O_425,N_2985,N_2948);
nor UO_426 (O_426,N_2941,N_2999);
and UO_427 (O_427,N_2959,N_2965);
nand UO_428 (O_428,N_2947,N_2975);
nor UO_429 (O_429,N_2974,N_2953);
nor UO_430 (O_430,N_2990,N_2999);
nand UO_431 (O_431,N_2964,N_2997);
or UO_432 (O_432,N_2970,N_2960);
xor UO_433 (O_433,N_2971,N_2958);
xnor UO_434 (O_434,N_2991,N_2970);
or UO_435 (O_435,N_2951,N_2948);
nor UO_436 (O_436,N_2975,N_2973);
nor UO_437 (O_437,N_2979,N_2941);
or UO_438 (O_438,N_2988,N_2969);
or UO_439 (O_439,N_2978,N_2941);
and UO_440 (O_440,N_2990,N_2947);
or UO_441 (O_441,N_2985,N_2963);
nand UO_442 (O_442,N_2967,N_2983);
and UO_443 (O_443,N_2973,N_2992);
nor UO_444 (O_444,N_2998,N_2944);
nand UO_445 (O_445,N_2994,N_2976);
xor UO_446 (O_446,N_2944,N_2983);
nand UO_447 (O_447,N_2982,N_2975);
or UO_448 (O_448,N_2954,N_2959);
nor UO_449 (O_449,N_2978,N_2959);
nand UO_450 (O_450,N_2972,N_2954);
or UO_451 (O_451,N_2951,N_2956);
nor UO_452 (O_452,N_2956,N_2986);
nor UO_453 (O_453,N_2945,N_2957);
nor UO_454 (O_454,N_2968,N_2981);
xnor UO_455 (O_455,N_2968,N_2985);
nor UO_456 (O_456,N_2956,N_2995);
nor UO_457 (O_457,N_2970,N_2997);
nor UO_458 (O_458,N_2995,N_2944);
and UO_459 (O_459,N_2992,N_2944);
or UO_460 (O_460,N_2975,N_2977);
nand UO_461 (O_461,N_2953,N_2971);
and UO_462 (O_462,N_2944,N_2960);
or UO_463 (O_463,N_2983,N_2976);
nor UO_464 (O_464,N_2948,N_2992);
nand UO_465 (O_465,N_2956,N_2969);
and UO_466 (O_466,N_2986,N_2950);
nand UO_467 (O_467,N_2962,N_2961);
and UO_468 (O_468,N_2977,N_2988);
and UO_469 (O_469,N_2985,N_2956);
nand UO_470 (O_470,N_2960,N_2989);
and UO_471 (O_471,N_2953,N_2958);
or UO_472 (O_472,N_2993,N_2982);
nand UO_473 (O_473,N_2964,N_2948);
and UO_474 (O_474,N_2966,N_2993);
nand UO_475 (O_475,N_2947,N_2983);
nand UO_476 (O_476,N_2987,N_2959);
or UO_477 (O_477,N_2973,N_2964);
and UO_478 (O_478,N_2962,N_2986);
nor UO_479 (O_479,N_2960,N_2981);
nor UO_480 (O_480,N_2951,N_2972);
nand UO_481 (O_481,N_2980,N_2964);
nand UO_482 (O_482,N_2945,N_2997);
nand UO_483 (O_483,N_2945,N_2995);
or UO_484 (O_484,N_2954,N_2978);
nand UO_485 (O_485,N_2951,N_2947);
and UO_486 (O_486,N_2977,N_2976);
nand UO_487 (O_487,N_2953,N_2940);
and UO_488 (O_488,N_2980,N_2962);
nor UO_489 (O_489,N_2971,N_2941);
nand UO_490 (O_490,N_2991,N_2984);
and UO_491 (O_491,N_2954,N_2977);
and UO_492 (O_492,N_2955,N_2986);
nor UO_493 (O_493,N_2989,N_2976);
xor UO_494 (O_494,N_2948,N_2971);
and UO_495 (O_495,N_2973,N_2978);
or UO_496 (O_496,N_2955,N_2988);
nand UO_497 (O_497,N_2950,N_2999);
nor UO_498 (O_498,N_2991,N_2981);
xnor UO_499 (O_499,N_2993,N_2990);
endmodule