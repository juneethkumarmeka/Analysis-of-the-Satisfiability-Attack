module basic_2000_20000_2500_40_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_1643,In_910);
and U1 (N_1,In_1070,In_929);
xor U2 (N_2,In_774,In_972);
or U3 (N_3,In_730,In_1360);
xnor U4 (N_4,In_1109,In_1671);
xnor U5 (N_5,In_47,In_917);
and U6 (N_6,In_679,In_79);
or U7 (N_7,In_537,In_1475);
nand U8 (N_8,In_347,In_513);
and U9 (N_9,In_299,In_1670);
xnor U10 (N_10,In_403,In_603);
and U11 (N_11,In_446,In_578);
and U12 (N_12,In_853,In_646);
nand U13 (N_13,In_765,In_726);
xnor U14 (N_14,In_698,In_1444);
nor U15 (N_15,In_1861,In_949);
nand U16 (N_16,In_1378,In_850);
nand U17 (N_17,In_536,In_1214);
and U18 (N_18,In_636,In_964);
nor U19 (N_19,In_1417,In_1341);
nand U20 (N_20,In_715,In_761);
nor U21 (N_21,In_1930,In_1950);
and U22 (N_22,In_1128,In_633);
nand U23 (N_23,In_1408,In_1542);
nand U24 (N_24,In_716,In_404);
or U25 (N_25,In_281,In_952);
xnor U26 (N_26,In_463,In_189);
nand U27 (N_27,In_1072,In_992);
or U28 (N_28,In_305,In_789);
and U29 (N_29,In_363,In_1168);
or U30 (N_30,In_1712,In_583);
nor U31 (N_31,In_1743,In_1543);
xor U32 (N_32,In_443,In_1493);
xnor U33 (N_33,In_33,In_1393);
and U34 (N_34,In_1218,In_1365);
nor U35 (N_35,In_232,In_360);
nand U36 (N_36,In_1802,In_563);
nand U37 (N_37,In_811,In_128);
and U38 (N_38,In_1352,In_709);
xor U39 (N_39,In_1222,In_1915);
nand U40 (N_40,In_282,In_1235);
or U41 (N_41,In_1040,In_1100);
nor U42 (N_42,In_263,In_139);
nor U43 (N_43,In_847,In_1011);
xnor U44 (N_44,In_450,In_1063);
and U45 (N_45,In_1526,In_311);
nand U46 (N_46,In_212,In_1812);
and U47 (N_47,In_1064,In_205);
xnor U48 (N_48,In_652,In_792);
nor U49 (N_49,In_1017,In_1344);
xnor U50 (N_50,In_406,In_108);
nor U51 (N_51,In_921,In_1702);
or U52 (N_52,In_1596,In_832);
nand U53 (N_53,In_621,In_110);
and U54 (N_54,In_876,In_401);
or U55 (N_55,In_1441,In_800);
or U56 (N_56,In_1061,In_948);
nand U57 (N_57,In_173,In_1056);
xnor U58 (N_58,In_916,In_1962);
nor U59 (N_59,In_148,In_398);
nand U60 (N_60,In_1217,In_678);
or U61 (N_61,In_1704,In_346);
and U62 (N_62,In_237,In_1661);
xor U63 (N_63,In_32,In_1528);
nand U64 (N_64,In_162,In_1136);
and U65 (N_65,In_1446,In_1923);
xnor U66 (N_66,In_512,In_806);
nor U67 (N_67,In_1955,In_292);
or U68 (N_68,In_1464,In_223);
or U69 (N_69,In_1937,In_1374);
xor U70 (N_70,In_1589,In_1669);
nand U71 (N_71,In_649,In_1953);
or U72 (N_72,In_931,In_1357);
nand U73 (N_73,In_228,In_1964);
xor U74 (N_74,In_1716,In_596);
and U75 (N_75,In_760,In_741);
xnor U76 (N_76,In_994,In_751);
xor U77 (N_77,In_624,In_54);
nor U78 (N_78,In_67,In_1648);
xor U79 (N_79,In_440,In_451);
and U80 (N_80,In_1085,In_70);
or U81 (N_81,In_1871,In_1166);
nor U82 (N_82,In_1460,In_490);
xor U83 (N_83,In_975,In_638);
nand U84 (N_84,In_1328,In_985);
nor U85 (N_85,In_1368,In_225);
xor U86 (N_86,In_1199,In_834);
or U87 (N_87,In_1143,In_270);
and U88 (N_88,In_1466,In_1709);
or U89 (N_89,In_1111,In_1794);
and U90 (N_90,In_872,In_623);
xor U91 (N_91,In_1603,In_1399);
xor U92 (N_92,In_1630,In_1244);
nand U93 (N_93,In_7,In_1867);
nor U94 (N_94,In_631,In_1711);
or U95 (N_95,In_435,In_177);
or U96 (N_96,In_412,In_267);
nor U97 (N_97,In_1032,In_941);
and U98 (N_98,In_1397,In_224);
and U99 (N_99,In_573,In_906);
nor U100 (N_100,In_1878,In_312);
and U101 (N_101,In_1785,In_1008);
or U102 (N_102,In_1811,In_154);
and U103 (N_103,In_1834,In_1824);
or U104 (N_104,In_1349,In_456);
and U105 (N_105,In_693,In_1197);
nor U106 (N_106,In_1180,In_1749);
nor U107 (N_107,In_265,In_1133);
nor U108 (N_108,In_1209,In_1550);
xor U109 (N_109,In_327,In_820);
nand U110 (N_110,In_1488,In_199);
or U111 (N_111,In_1185,In_220);
xor U112 (N_112,In_40,In_1383);
or U113 (N_113,In_339,In_1877);
nor U114 (N_114,In_241,In_589);
and U115 (N_115,In_1337,In_1348);
nor U116 (N_116,In_179,In_970);
nor U117 (N_117,In_1595,In_691);
xor U118 (N_118,In_15,In_695);
xor U119 (N_119,In_1855,In_1590);
or U120 (N_120,In_1092,In_1120);
nand U121 (N_121,In_688,In_1534);
nand U122 (N_122,In_1260,In_169);
or U123 (N_123,In_534,In_1333);
nand U124 (N_124,In_1114,In_1073);
nor U125 (N_125,In_1625,In_28);
xor U126 (N_126,In_620,In_1082);
or U127 (N_127,In_81,In_76);
and U128 (N_128,In_1579,In_1585);
and U129 (N_129,In_597,In_1065);
xnor U130 (N_130,In_1409,In_1351);
xor U131 (N_131,In_1554,In_616);
nor U132 (N_132,In_1416,In_1993);
or U133 (N_133,In_1918,In_797);
or U134 (N_134,In_12,In_1617);
xnor U135 (N_135,In_190,In_1573);
and U136 (N_136,In_1266,In_752);
and U137 (N_137,In_1949,In_988);
nand U138 (N_138,In_905,In_1448);
nand U139 (N_139,In_144,In_1880);
xor U140 (N_140,In_999,In_995);
nand U141 (N_141,In_1339,In_1018);
nand U142 (N_142,In_1162,In_1765);
nor U143 (N_143,In_1924,In_318);
and U144 (N_144,In_1129,In_685);
and U145 (N_145,In_255,In_1605);
or U146 (N_146,In_1471,In_1771);
xnor U147 (N_147,In_737,In_644);
nand U148 (N_148,In_348,In_565);
nand U149 (N_149,In_1265,In_960);
or U150 (N_150,In_122,In_997);
or U151 (N_151,In_1006,In_1283);
and U152 (N_152,In_1631,In_478);
xnor U153 (N_153,In_1453,In_1445);
or U154 (N_154,In_236,In_475);
nand U155 (N_155,In_1175,In_1538);
and U156 (N_156,In_78,In_533);
and U157 (N_157,In_1483,In_1735);
and U158 (N_158,In_576,In_1287);
or U159 (N_159,In_1694,In_1828);
nor U160 (N_160,In_734,In_1705);
nand U161 (N_161,In_1776,In_1621);
xnor U162 (N_162,In_1899,In_1698);
or U163 (N_163,In_803,In_1676);
nand U164 (N_164,In_702,In_138);
xnor U165 (N_165,In_743,In_21);
or U166 (N_166,In_399,In_98);
xor U167 (N_167,In_1280,In_609);
nand U168 (N_168,In_468,In_1570);
nand U169 (N_169,In_219,In_1667);
or U170 (N_170,In_1844,In_1227);
or U171 (N_171,In_870,In_1340);
and U172 (N_172,In_1968,In_1234);
xnor U173 (N_173,In_521,In_1839);
and U174 (N_174,In_1872,In_405);
and U175 (N_175,In_817,In_180);
xor U176 (N_176,In_804,In_843);
nand U177 (N_177,In_202,In_1931);
nand U178 (N_178,In_1503,In_1591);
nand U179 (N_179,In_1809,In_1746);
and U180 (N_180,In_193,In_654);
xnor U181 (N_181,In_1237,In_1662);
xor U182 (N_182,In_1833,In_873);
and U183 (N_183,In_883,In_1467);
or U184 (N_184,In_250,In_126);
nand U185 (N_185,In_480,In_1299);
or U186 (N_186,In_1826,In_674);
or U187 (N_187,In_936,In_1938);
xor U188 (N_188,In_846,In_395);
and U189 (N_189,In_352,In_851);
nand U190 (N_190,In_1347,In_1284);
xor U191 (N_191,In_274,In_1051);
xnor U192 (N_192,In_1911,In_822);
and U193 (N_193,In_1097,In_1412);
or U194 (N_194,In_340,In_1219);
or U195 (N_195,In_1606,In_1979);
nand U196 (N_196,In_1273,In_791);
or U197 (N_197,In_591,In_1523);
or U198 (N_198,In_1515,In_1174);
nor U199 (N_199,In_1939,In_507);
and U200 (N_200,In_925,In_1960);
nand U201 (N_201,In_1866,In_801);
nand U202 (N_202,In_542,In_82);
nor U203 (N_203,In_1414,In_742);
or U204 (N_204,In_93,In_694);
or U205 (N_205,In_174,In_825);
nor U206 (N_206,In_37,In_291);
xor U207 (N_207,In_1679,In_768);
xnor U208 (N_208,In_1131,In_141);
nor U209 (N_209,In_1382,In_1186);
or U210 (N_210,In_1449,In_1994);
xor U211 (N_211,In_49,In_345);
nand U212 (N_212,In_123,In_508);
nor U213 (N_213,In_1058,In_158);
nand U214 (N_214,In_1014,In_90);
or U215 (N_215,In_1117,In_1303);
nand U216 (N_216,In_1015,In_408);
nand U217 (N_217,In_1741,In_1564);
or U218 (N_218,In_764,In_73);
xnor U219 (N_219,In_1646,In_1577);
and U220 (N_220,In_370,In_657);
nand U221 (N_221,In_1026,In_1118);
nand U222 (N_222,In_1571,In_955);
and U223 (N_223,In_1122,In_708);
and U224 (N_224,In_1108,In_1619);
nand U225 (N_225,In_486,In_1271);
nor U226 (N_226,In_868,In_529);
or U227 (N_227,In_354,In_1054);
and U228 (N_228,In_759,In_895);
xor U229 (N_229,In_1933,In_417);
nor U230 (N_230,In_1583,In_1020);
or U231 (N_231,In_664,In_1838);
xor U232 (N_232,In_581,In_261);
nand U233 (N_233,In_983,In_1936);
nor U234 (N_234,In_1353,In_506);
and U235 (N_235,In_890,In_1587);
and U236 (N_236,In_1469,In_1759);
xnor U237 (N_237,In_1030,In_1691);
nand U238 (N_238,In_1304,In_247);
and U239 (N_239,In_472,In_1487);
nand U240 (N_240,In_671,In_1519);
nor U241 (N_241,In_87,In_1821);
xnor U242 (N_242,In_243,In_1841);
or U243 (N_243,In_300,In_1150);
nand U244 (N_244,In_1588,In_821);
nand U245 (N_245,In_1774,In_254);
nand U246 (N_246,In_328,In_326);
nor U247 (N_247,In_1484,In_781);
and U248 (N_248,In_1644,In_510);
or U249 (N_249,In_209,In_1411);
nor U250 (N_250,In_1195,In_125);
xnor U251 (N_251,In_771,In_441);
nand U252 (N_252,In_928,In_829);
xnor U253 (N_253,In_1456,In_191);
nand U254 (N_254,In_1849,In_454);
xor U255 (N_255,In_1048,In_314);
or U256 (N_256,In_1492,In_732);
and U257 (N_257,In_962,In_1744);
nand U258 (N_258,In_1091,In_296);
nand U259 (N_259,In_545,In_1112);
nand U260 (N_260,In_1203,In_1736);
or U261 (N_261,In_1103,In_1325);
nand U262 (N_262,In_747,In_725);
xnor U263 (N_263,In_0,In_455);
nand U264 (N_264,In_31,In_1315);
or U265 (N_265,In_877,In_91);
and U266 (N_266,In_1173,In_387);
xnor U267 (N_267,In_1433,In_64);
and U268 (N_268,In_1971,In_499);
nand U269 (N_269,In_1514,In_1213);
or U270 (N_270,In_1426,In_1804);
nand U271 (N_271,In_377,In_1666);
nor U272 (N_272,In_810,In_535);
and U273 (N_273,In_1864,In_944);
or U274 (N_274,In_1236,In_268);
nand U275 (N_275,In_1405,In_104);
xor U276 (N_276,In_900,In_656);
and U277 (N_277,In_239,In_1154);
xnor U278 (N_278,In_231,In_1345);
or U279 (N_279,In_1327,In_1178);
xor U280 (N_280,In_1293,In_1555);
and U281 (N_281,In_251,In_903);
or U282 (N_282,In_206,In_1813);
and U283 (N_283,In_1309,In_1229);
nor U284 (N_284,In_517,In_1586);
xor U285 (N_285,In_1132,In_1733);
xnor U286 (N_286,In_1820,In_1815);
xnor U287 (N_287,In_385,In_1773);
xnor U288 (N_288,In_201,In_538);
or U289 (N_289,In_1990,In_750);
or U290 (N_290,In_1485,In_469);
and U291 (N_291,In_216,In_1027);
nand U292 (N_292,In_107,In_1852);
or U293 (N_293,In_1163,In_518);
nor U294 (N_294,In_1096,In_1262);
or U295 (N_295,In_755,In_1893);
and U296 (N_296,In_786,In_302);
and U297 (N_297,In_974,In_495);
and U298 (N_298,In_618,In_968);
or U299 (N_299,In_252,In_458);
nor U300 (N_300,In_1208,In_266);
nand U301 (N_301,In_710,In_1090);
nand U302 (N_302,In_1738,In_1113);
nor U303 (N_303,In_198,In_57);
nand U304 (N_304,In_1707,In_95);
and U305 (N_305,In_1093,In_1259);
nor U306 (N_306,In_432,In_349);
or U307 (N_307,In_445,In_1474);
or U308 (N_308,In_1655,In_749);
or U309 (N_309,In_993,In_956);
xor U310 (N_310,In_1689,In_324);
nor U311 (N_311,In_316,In_1221);
nor U312 (N_312,In_1380,In_610);
nand U313 (N_313,In_1465,In_996);
and U314 (N_314,In_1330,In_1101);
or U315 (N_315,In_1270,In_1810);
xnor U316 (N_316,In_544,In_1170);
xnor U317 (N_317,In_1859,In_1976);
or U318 (N_318,In_612,In_132);
xor U319 (N_319,In_1710,In_1319);
or U320 (N_320,In_200,In_775);
or U321 (N_321,In_1566,In_1317);
nor U322 (N_322,In_1517,In_845);
and U323 (N_323,In_22,In_1533);
nor U324 (N_324,In_1608,In_1322);
xor U325 (N_325,In_1803,In_355);
or U326 (N_326,In_1246,In_1521);
xor U327 (N_327,In_1879,In_86);
nand U328 (N_328,In_1121,In_1278);
and U329 (N_329,In_69,In_394);
nand U330 (N_330,In_1198,In_320);
xor U331 (N_331,In_1391,In_1231);
and U332 (N_332,In_1697,In_24);
and U333 (N_333,In_717,In_1398);
nand U334 (N_334,In_1305,In_598);
nand U335 (N_335,In_579,In_594);
xor U336 (N_336,In_782,In_1754);
nand U337 (N_337,In_491,In_111);
xnor U338 (N_338,In_1761,In_176);
and U339 (N_339,In_161,In_1628);
and U340 (N_340,In_1629,In_539);
or U341 (N_341,In_1370,In_343);
nand U342 (N_342,In_559,In_1201);
nor U343 (N_343,In_1258,In_285);
nor U344 (N_344,In_724,In_1281);
nor U345 (N_345,In_748,In_476);
nor U346 (N_346,In_639,In_319);
or U347 (N_347,In_1215,In_1454);
nand U348 (N_348,In_117,In_953);
xor U349 (N_349,In_332,In_1302);
nand U350 (N_350,In_625,In_430);
xnor U351 (N_351,In_1530,In_1323);
xor U352 (N_352,In_635,In_807);
nor U353 (N_353,In_208,In_361);
nand U354 (N_354,In_338,In_1623);
nor U355 (N_355,In_20,In_359);
nor U356 (N_356,In_697,In_1329);
or U357 (N_357,In_439,In_1141);
nor U358 (N_358,In_1137,In_256);
nand U359 (N_359,In_74,In_182);
xnor U360 (N_360,In_234,In_1377);
nand U361 (N_361,In_298,In_1518);
nor U362 (N_362,In_1511,In_699);
nand U363 (N_363,In_235,In_647);
and U364 (N_364,In_1567,In_951);
or U365 (N_365,In_783,In_264);
xnor U366 (N_366,In_892,In_1164);
nor U367 (N_367,In_546,In_1184);
nor U368 (N_368,In_1297,In_823);
or U369 (N_369,In_959,In_1076);
or U370 (N_370,In_950,In_871);
nor U371 (N_371,In_736,In_1343);
or U372 (N_372,In_1913,In_1581);
or U373 (N_373,In_286,In_912);
nand U374 (N_374,In_283,In_1983);
and U375 (N_375,In_146,In_1756);
or U376 (N_376,In_1793,In_400);
or U377 (N_377,In_494,In_164);
or U378 (N_378,In_1052,In_1848);
nand U379 (N_379,In_1240,In_1827);
and U380 (N_380,In_1560,In_1984);
or U381 (N_381,In_1706,In_1592);
nand U382 (N_382,In_1985,In_907);
nor U383 (N_383,In_773,In_374);
and U384 (N_384,In_1665,In_1437);
nand U385 (N_385,In_181,In_665);
nand U386 (N_386,In_1727,In_46);
or U387 (N_387,In_1598,In_1798);
nor U388 (N_388,In_244,In_1300);
xnor U389 (N_389,In_1039,In_805);
and U390 (N_390,In_1860,In_1135);
or U391 (N_391,In_1350,In_1144);
nand U392 (N_392,In_333,In_1775);
nor U393 (N_393,In_1479,In_568);
nand U394 (N_394,In_758,In_1068);
and U395 (N_395,In_965,In_707);
and U396 (N_396,In_818,In_1612);
and U397 (N_397,In_686,In_1025);
or U398 (N_398,In_745,In_1675);
or U399 (N_399,In_1638,In_362);
or U400 (N_400,In_1886,In_878);
nor U401 (N_401,In_1896,In_1537);
or U402 (N_402,In_1415,In_498);
or U403 (N_403,In_924,In_1788);
nor U404 (N_404,In_168,In_365);
nor U405 (N_405,In_1395,In_1151);
and U406 (N_406,In_946,In_1683);
nand U407 (N_407,In_1696,In_943);
xor U408 (N_408,In_967,In_1256);
nor U409 (N_409,In_1171,In_932);
nand U410 (N_410,In_1814,In_1932);
nor U411 (N_411,In_1272,In_1681);
xnor U412 (N_412,In_142,In_259);
or U413 (N_413,In_1882,In_1998);
or U414 (N_414,In_1037,In_1336);
nand U415 (N_415,In_273,In_1726);
or U416 (N_416,In_1012,In_392);
and U417 (N_417,In_438,In_72);
or U418 (N_418,In_611,In_1038);
or U419 (N_419,In_1193,In_1961);
nand U420 (N_420,In_1948,In_839);
xor U421 (N_421,In_276,In_1862);
xor U422 (N_422,In_1753,In_1447);
nand U423 (N_423,In_1326,In_911);
or U424 (N_424,In_1870,In_1049);
nand U425 (N_425,In_453,In_1752);
nor U426 (N_426,In_1582,In_230);
and U427 (N_427,In_841,In_1463);
xor U428 (N_428,In_1313,In_421);
nand U429 (N_429,In_894,In_858);
and U430 (N_430,In_77,In_1685);
and U431 (N_431,In_942,In_481);
and U432 (N_432,In_1640,In_1687);
nand U433 (N_433,In_1970,In_1495);
xor U434 (N_434,In_1242,In_1633);
and U435 (N_435,In_893,In_680);
and U436 (N_436,In_315,In_971);
xnor U437 (N_437,In_1895,In_402);
xor U438 (N_438,In_1869,In_229);
nor U439 (N_439,In_935,In_712);
nor U440 (N_440,In_1247,In_836);
nand U441 (N_441,In_880,In_1723);
xor U442 (N_442,In_278,In_1884);
xor U443 (N_443,In_706,In_1921);
or U444 (N_444,In_1611,In_1830);
nand U445 (N_445,In_1574,In_431);
or U446 (N_446,In_1430,In_1807);
nand U447 (N_447,In_1883,In_214);
nand U448 (N_448,In_1652,In_473);
or U449 (N_449,In_1760,In_1552);
nor U450 (N_450,In_1190,In_1682);
nand U451 (N_451,In_526,In_1062);
nor U452 (N_452,In_186,In_1396);
nand U453 (N_453,In_1693,In_192);
or U454 (N_454,In_1005,In_1013);
nor U455 (N_455,In_1386,In_272);
and U456 (N_456,In_1786,In_92);
nor U457 (N_457,In_1684,In_1138);
nor U458 (N_458,In_114,In_1451);
or U459 (N_459,In_1668,In_1034);
nand U460 (N_460,In_898,In_336);
and U461 (N_461,In_555,In_407);
and U462 (N_462,In_143,In_548);
xnor U463 (N_463,In_682,In_1212);
and U464 (N_464,In_378,In_713);
xnor U465 (N_465,In_442,In_1480);
and U466 (N_466,In_1192,In_727);
nor U467 (N_467,In_1853,In_62);
or U468 (N_468,In_414,In_136);
or U469 (N_469,In_550,In_661);
nor U470 (N_470,In_700,In_1799);
or U471 (N_471,In_1461,In_1413);
nor U472 (N_472,In_663,In_99);
and U473 (N_473,In_1455,In_587);
xnor U474 (N_474,In_641,In_1900);
xnor U475 (N_475,In_1531,In_1914);
xnor U476 (N_476,In_165,In_844);
nand U477 (N_477,In_586,In_784);
and U478 (N_478,In_634,In_500);
and U479 (N_479,In_1945,In_248);
nand U480 (N_480,In_1257,In_980);
xor U481 (N_481,In_188,In_178);
xor U482 (N_482,In_643,In_577);
or U483 (N_483,In_1419,In_570);
nand U484 (N_484,In_1028,In_1110);
and U485 (N_485,In_1400,In_1187);
and U486 (N_486,In_482,In_253);
or U487 (N_487,In_1232,In_34);
xor U488 (N_488,In_1818,In_1817);
xor U489 (N_489,In_703,In_1338);
and U490 (N_490,In_1713,In_36);
or U491 (N_491,In_233,In_614);
and U492 (N_492,In_1009,In_1715);
nor U493 (N_493,In_1699,In_14);
or U494 (N_494,In_1053,In_1780);
xnor U495 (N_495,In_1181,In_1610);
nand U496 (N_496,In_1083,In_240);
nand U497 (N_497,In_1954,In_1719);
and U498 (N_498,In_1854,In_1840);
xor U499 (N_499,In_1657,In_1403);
nor U500 (N_500,In_840,In_650);
nand U501 (N_501,In_1783,N_496);
or U502 (N_502,In_89,In_1285);
or U503 (N_503,In_434,In_1751);
nor U504 (N_504,In_1614,In_1010);
or U505 (N_505,In_561,N_402);
xnor U506 (N_506,In_582,N_391);
nand U507 (N_507,N_124,In_1874);
or U508 (N_508,N_485,In_819);
and U509 (N_509,N_36,N_185);
or U510 (N_510,N_403,N_469);
or U511 (N_511,In_1226,In_723);
xnor U512 (N_512,N_237,In_1275);
or U513 (N_513,In_295,In_1388);
nor U514 (N_514,In_1077,N_273);
xor U515 (N_515,N_307,In_1764);
and U516 (N_516,In_195,In_303);
nor U517 (N_517,N_151,In_350);
xor U518 (N_518,N_375,In_828);
and U519 (N_519,In_1369,In_1541);
xor U520 (N_520,In_1512,In_121);
nor U521 (N_521,N_90,N_8);
nand U522 (N_522,In_1019,In_831);
nor U523 (N_523,In_1251,In_393);
and U524 (N_524,N_406,In_528);
nor U525 (N_525,In_799,N_134);
or U526 (N_526,N_251,In_1354);
xnor U527 (N_527,In_1334,In_1672);
nand U528 (N_528,N_247,N_325);
xnor U529 (N_529,In_1384,N_131);
or U530 (N_530,In_1873,In_884);
nand U531 (N_531,N_230,N_302);
nor U532 (N_532,N_317,In_1500);
and U533 (N_533,In_145,In_600);
xnor U534 (N_534,N_184,In_1410);
nand U535 (N_535,In_1887,In_540);
nand U536 (N_536,In_857,In_655);
nor U537 (N_537,In_852,In_762);
xor U538 (N_538,N_97,In_1940);
nor U539 (N_539,In_739,In_464);
nor U540 (N_540,In_1045,In_670);
and U541 (N_541,In_304,N_371);
xnor U542 (N_542,In_886,In_60);
xor U543 (N_543,In_1134,In_1087);
and U544 (N_544,In_1604,N_288);
or U545 (N_545,N_27,N_217);
and U546 (N_546,In_1837,In_1762);
xor U547 (N_547,N_299,In_599);
and U548 (N_548,In_1903,In_1740);
and U549 (N_549,In_1593,In_584);
nor U550 (N_550,In_1730,In_814);
and U551 (N_551,In_1372,In_909);
or U552 (N_552,N_386,In_1792);
nand U553 (N_553,In_1777,N_88);
nand U554 (N_554,In_1597,In_284);
or U555 (N_555,In_1664,In_1972);
or U556 (N_556,N_56,N_270);
and U557 (N_557,In_184,N_225);
or U558 (N_558,In_1650,In_622);
nand U559 (N_559,In_48,In_1926);
or U560 (N_560,In_590,In_1578);
nand U561 (N_561,In_918,In_849);
nor U562 (N_562,In_1157,In_301);
nand U563 (N_563,N_204,In_1607);
xor U564 (N_564,N_130,N_339);
or U565 (N_565,In_331,In_809);
xor U566 (N_566,In_1060,In_1865);
and U567 (N_567,N_279,N_259);
or U568 (N_568,N_303,In_1975);
and U569 (N_569,In_966,In_731);
nand U570 (N_570,In_1245,N_39);
nor U571 (N_571,In_1289,In_602);
xor U572 (N_572,In_1739,N_311);
and U573 (N_573,In_919,N_12);
nand U574 (N_574,In_1701,In_945);
or U575 (N_575,In_592,N_78);
and U576 (N_576,In_368,N_84);
nand U577 (N_577,In_1796,N_242);
or U578 (N_578,In_1194,In_2);
or U579 (N_579,In_1497,In_1656);
or U580 (N_580,In_289,In_1228);
or U581 (N_581,N_119,In_720);
or U582 (N_582,N_285,In_1172);
xnor U583 (N_583,In_915,In_501);
nand U584 (N_584,N_30,In_1980);
nand U585 (N_585,In_530,In_1066);
nor U586 (N_586,In_551,In_1594);
xnor U587 (N_587,N_383,In_1321);
or U588 (N_588,In_862,In_879);
xnor U589 (N_589,In_1489,In_1836);
and U590 (N_590,In_1080,In_1563);
or U591 (N_591,N_440,In_1308);
and U592 (N_592,N_149,N_385);
and U593 (N_593,In_1905,N_221);
and U594 (N_594,In_838,N_319);
or U595 (N_595,In_1458,N_349);
nor U596 (N_596,In_675,In_991);
xnor U597 (N_597,In_1146,In_1361);
or U598 (N_598,N_269,In_279);
xnor U599 (N_599,In_1119,In_601);
nor U600 (N_600,N_16,N_65);
or U601 (N_601,N_494,N_467);
and U602 (N_602,In_604,In_129);
nand U603 (N_603,In_901,In_1651);
or U604 (N_604,In_353,N_414);
and U605 (N_605,N_104,In_1919);
xnor U606 (N_606,In_777,N_176);
and U607 (N_607,N_68,In_667);
and U608 (N_608,In_425,In_1856);
or U609 (N_609,In_1767,N_328);
xnor U610 (N_610,N_355,N_60);
nand U611 (N_611,In_58,In_683);
or U612 (N_612,In_1216,N_47);
xnor U613 (N_613,N_369,In_1513);
nor U614 (N_614,In_1888,In_1708);
or U615 (N_615,In_492,In_105);
xor U616 (N_616,In_1379,In_221);
or U617 (N_617,In_1301,In_1999);
or U618 (N_618,N_474,N_263);
or U619 (N_619,N_11,In_1569);
nand U620 (N_620,In_585,In_543);
or U621 (N_621,In_989,In_669);
nand U622 (N_622,In_637,In_887);
nor U623 (N_623,In_334,In_424);
nor U624 (N_624,In_619,N_266);
and U625 (N_625,N_441,N_71);
and U626 (N_626,In_124,In_1094);
nor U627 (N_627,In_1238,In_1390);
nand U628 (N_628,In_1912,In_640);
xor U629 (N_629,N_89,In_371);
nand U630 (N_630,N_277,N_350);
nor U631 (N_631,N_75,In_1654);
xor U632 (N_632,In_383,N_108);
or U633 (N_633,N_459,In_1452);
and U634 (N_634,In_793,N_278);
or U635 (N_635,In_1126,In_1050);
and U636 (N_636,N_378,N_495);
xnor U637 (N_637,In_1967,In_1402);
xnor U638 (N_638,In_1929,In_1335);
xnor U639 (N_639,In_1429,In_1770);
nand U640 (N_640,In_1191,In_1358);
nor U641 (N_641,In_558,In_519);
or U642 (N_642,N_362,In_567);
nand U643 (N_643,In_416,In_1645);
nor U644 (N_644,In_808,In_1635);
nor U645 (N_645,In_294,In_575);
xnor U646 (N_646,In_899,In_1288);
nor U647 (N_647,In_1700,In_1261);
nor U648 (N_648,In_1997,N_458);
or U649 (N_649,In_1572,In_779);
nand U650 (N_650,In_217,In_1059);
and U651 (N_651,N_227,In_554);
nor U652 (N_652,In_606,N_427);
nor U653 (N_653,In_55,N_499);
or U654 (N_654,In_1145,In_835);
nand U655 (N_655,In_692,In_153);
xor U656 (N_656,N_374,In_444);
nor U657 (N_657,In_628,N_418);
nor U658 (N_658,In_864,In_1580);
or U659 (N_659,In_812,N_31);
nor U660 (N_660,N_192,N_122);
and U661 (N_661,In_389,In_1996);
xnor U662 (N_662,N_377,In_84);
nor U663 (N_663,In_1613,N_486);
xnor U664 (N_664,In_766,In_1407);
nor U665 (N_665,N_413,In_1428);
nor U666 (N_666,N_51,In_630);
nor U667 (N_667,In_1568,In_1626);
and U668 (N_668,N_73,N_468);
or U669 (N_669,In_379,N_208);
nand U670 (N_670,N_234,In_1023);
and U671 (N_671,In_902,N_255);
nand U672 (N_672,N_305,N_276);
nor U673 (N_673,N_140,N_198);
and U674 (N_674,In_1421,N_111);
and U675 (N_675,In_388,In_1387);
and U676 (N_676,N_443,N_26);
and U677 (N_677,In_672,In_1772);
nand U678 (N_678,In_238,In_1107);
and U679 (N_679,N_62,In_1024);
xor U680 (N_680,In_778,N_155);
xnor U681 (N_681,N_38,In_547);
nand U682 (N_682,N_390,N_314);
and U683 (N_683,In_1624,N_40);
xnor U684 (N_684,N_82,In_1001);
nor U685 (N_685,In_183,N_271);
nor U686 (N_686,In_888,In_51);
or U687 (N_687,In_325,N_59);
or U688 (N_688,In_1659,N_207);
xor U689 (N_689,In_1946,In_1978);
xor U690 (N_690,In_1167,In_1432);
and U691 (N_691,In_1910,In_290);
nand U692 (N_692,N_129,In_1084);
nor U693 (N_693,In_437,In_467);
nand U694 (N_694,In_795,N_457);
nand U695 (N_695,N_246,In_1747);
nor U696 (N_696,In_1714,In_396);
or U697 (N_697,In_1158,In_1422);
and U698 (N_698,N_6,In_171);
or U699 (N_699,In_172,In_1196);
and U700 (N_700,In_1498,N_239);
or U701 (N_701,In_275,In_262);
nor U702 (N_702,In_1536,In_1800);
nand U703 (N_703,N_28,In_1248);
nand U704 (N_704,In_1703,In_1724);
or U705 (N_705,N_439,In_1095);
xor U706 (N_706,In_1891,N_409);
nand U707 (N_707,In_372,In_1941);
xnor U708 (N_708,In_1373,In_287);
or U709 (N_709,In_1440,In_1647);
nor U710 (N_710,In_1692,In_798);
xor U711 (N_711,In_1179,In_1423);
nand U712 (N_712,N_240,In_1680);
xnor U713 (N_713,In_569,In_1989);
nand U714 (N_714,In_1420,In_1916);
and U715 (N_715,In_1717,N_431);
xor U716 (N_716,In_1296,In_787);
nor U717 (N_717,In_1142,In_882);
or U718 (N_718,In_1003,N_284);
nand U719 (N_719,In_1958,In_1205);
xor U720 (N_720,In_681,In_719);
or U721 (N_721,In_1876,In_608);
and U722 (N_722,In_520,N_373);
nor U723 (N_723,In_1041,N_98);
xnor U724 (N_724,In_1982,N_175);
nor U725 (N_725,In_1732,N_76);
nor U726 (N_726,In_1267,N_447);
nand U727 (N_727,N_256,In_18);
or U728 (N_728,N_103,N_133);
nor U729 (N_729,In_1858,In_1755);
and U730 (N_730,In_1310,In_1842);
or U731 (N_731,In_651,In_1992);
or U732 (N_732,In_856,In_908);
or U733 (N_733,N_281,N_381);
or U734 (N_734,In_337,In_101);
or U735 (N_735,N_479,N_370);
and U736 (N_736,In_187,In_1674);
nand U737 (N_737,N_52,In_185);
xor U738 (N_738,N_5,N_424);
xnor U739 (N_739,In_1637,In_155);
nor U740 (N_740,In_52,N_182);
and U741 (N_741,N_126,In_39);
nor U742 (N_742,In_1462,In_42);
nand U743 (N_743,In_213,In_629);
nor U744 (N_744,In_133,In_1481);
nand U745 (N_745,N_478,N_261);
or U746 (N_746,In_772,In_1532);
nand U747 (N_747,In_869,In_313);
nand U748 (N_748,N_372,N_15);
xor U749 (N_749,N_118,In_525);
nand U750 (N_750,In_1189,In_1729);
and U751 (N_751,In_427,In_1956);
and U752 (N_752,In_462,In_676);
nor U753 (N_753,N_352,In_785);
nand U754 (N_754,In_627,In_449);
nand U755 (N_755,In_1943,N_382);
xnor U756 (N_756,In_1332,In_341);
nand U757 (N_757,In_23,In_1071);
or U758 (N_758,In_826,In_1401);
xnor U759 (N_759,In_1649,N_470);
or U760 (N_760,In_896,In_1748);
nor U761 (N_761,N_331,In_1404);
or U762 (N_762,In_308,N_178);
nand U763 (N_763,N_357,N_34);
xor U764 (N_764,N_218,N_205);
nand U765 (N_765,In_1312,In_203);
nor U766 (N_766,In_96,In_134);
nand U767 (N_767,In_613,In_1966);
nand U768 (N_768,N_268,In_1890);
nor U769 (N_769,In_249,In_137);
nand U770 (N_770,N_477,N_61);
nand U771 (N_771,In_1295,In_118);
or U772 (N_772,In_35,In_891);
nor U773 (N_773,In_1324,N_298);
nand U774 (N_774,In_729,In_474);
xnor U775 (N_775,N_393,In_422);
nor U776 (N_776,N_2,In_1516);
xor U777 (N_777,In_260,In_753);
and U778 (N_778,In_733,N_146);
and U779 (N_779,In_429,In_307);
and U780 (N_780,In_1249,In_1863);
xnor U781 (N_781,N_451,In_1263);
or U782 (N_782,In_1385,In_460);
xor U783 (N_783,In_645,N_337);
and U784 (N_784,In_1556,In_1152);
and U785 (N_785,In_1366,In_1995);
and U786 (N_786,In_756,N_327);
xnor U787 (N_787,N_164,In_794);
and U788 (N_788,In_71,N_310);
and U789 (N_789,In_1482,In_1225);
and U790 (N_790,N_330,In_1069);
xnor U791 (N_791,N_145,In_1);
and U792 (N_792,N_18,In_1678);
and U793 (N_793,In_418,N_160);
or U794 (N_794,In_979,N_48);
or U795 (N_795,In_833,In_1959);
nor U796 (N_796,In_1722,In_30);
or U797 (N_797,N_329,N_13);
xor U798 (N_798,In_790,In_342);
nand U799 (N_799,N_180,In_1636);
nor U800 (N_800,N_387,N_77);
xnor U801 (N_801,In_210,In_1973);
nand U802 (N_802,In_1104,In_1161);
and U803 (N_803,In_1658,N_85);
or U804 (N_804,In_130,N_157);
or U805 (N_805,N_489,In_1545);
nor U806 (N_806,N_399,N_482);
nor U807 (N_807,N_45,N_228);
or U808 (N_808,In_1808,N_113);
nor U809 (N_809,N_304,In_100);
nor U810 (N_810,In_1089,In_68);
nor U811 (N_811,In_1686,N_177);
nand U812 (N_812,N_171,In_1632);
nand U813 (N_813,In_65,In_1639);
nand U814 (N_814,N_224,In_1906);
nor U815 (N_815,In_595,In_170);
nor U816 (N_816,In_1183,In_1904);
or U817 (N_817,In_470,N_95);
or U818 (N_818,In_1210,N_473);
nor U819 (N_819,N_161,N_222);
and U820 (N_820,N_14,In_549);
nand U821 (N_821,In_43,N_120);
or U822 (N_822,N_365,N_231);
and U823 (N_823,In_1436,N_324);
or U824 (N_824,In_1520,N_37);
xnor U825 (N_825,In_1031,In_1508);
xnor U826 (N_826,In_531,N_196);
nor U827 (N_827,N_419,In_3);
or U828 (N_828,N_170,N_142);
xnor U829 (N_829,In_1220,N_125);
or U830 (N_830,In_1105,In_13);
nor U831 (N_831,N_472,N_143);
and U832 (N_832,In_1806,In_1963);
xor U833 (N_833,In_1908,N_348);
xor U834 (N_834,In_493,In_1898);
and U835 (N_835,In_1147,N_466);
xor U836 (N_836,In_246,N_364);
xnor U837 (N_837,In_1832,In_1947);
nor U838 (N_838,In_1206,In_112);
or U839 (N_839,In_27,In_969);
nor U840 (N_840,N_361,In_1406);
nor U841 (N_841,In_323,N_159);
nand U842 (N_842,In_1478,In_45);
nor U843 (N_843,In_984,N_21);
and U844 (N_844,In_1721,N_455);
and U845 (N_845,In_1252,In_149);
nor U846 (N_846,N_267,In_1055);
nor U847 (N_847,N_487,In_1046);
xnor U848 (N_848,In_1544,In_373);
nand U849 (N_849,In_215,In_1047);
and U850 (N_850,In_1677,In_1443);
nand U851 (N_851,In_1074,N_359);
and U852 (N_852,In_1156,N_464);
or U853 (N_853,In_1922,In_973);
nor U854 (N_854,In_116,In_1502);
or U855 (N_855,In_1557,In_1033);
and U856 (N_856,In_147,In_1737);
xor U857 (N_857,N_289,N_127);
nor U858 (N_858,In_1991,In_1253);
xor U859 (N_859,In_881,In_211);
and U860 (N_860,N_292,N_367);
or U861 (N_861,N_435,In_1507);
nor U862 (N_862,N_454,N_282);
or U863 (N_863,N_42,In_1177);
nor U864 (N_864,In_1504,N_9);
xor U865 (N_865,In_977,N_232);
xor U866 (N_866,In_297,N_203);
nand U867 (N_867,N_188,N_165);
xor U868 (N_868,N_49,N_80);
or U869 (N_869,In_483,In_1254);
nor U870 (N_870,In_1016,N_395);
nor U871 (N_871,N_411,In_1546);
or U872 (N_872,N_115,N_450);
nor U873 (N_873,In_1561,In_522);
xor U874 (N_874,N_400,In_1894);
or U875 (N_875,N_405,In_1831);
and U876 (N_876,In_1468,N_318);
nor U877 (N_877,N_81,N_147);
or U878 (N_878,In_358,In_571);
and U879 (N_879,N_449,In_1660);
nand U880 (N_880,N_154,In_411);
xor U881 (N_881,In_127,In_25);
nand U882 (N_882,In_1529,In_1851);
xor U883 (N_883,N_462,N_483);
and U884 (N_884,N_10,In_1434);
or U885 (N_885,N_417,In_1363);
xnor U886 (N_886,In_436,In_1371);
xor U887 (N_887,N_183,N_235);
and U888 (N_888,In_1885,N_294);
nor U889 (N_889,In_1944,In_1286);
xor U890 (N_890,In_351,In_1067);
xor U891 (N_891,In_824,N_92);
xor U892 (N_892,N_41,N_64);
or U893 (N_893,N_3,In_718);
and U894 (N_894,In_802,In_939);
nand U895 (N_895,In_119,N_87);
nor U896 (N_896,N_444,In_1846);
nand U897 (N_897,In_976,N_189);
xnor U898 (N_898,In_958,N_214);
or U899 (N_899,In_11,In_1294);
xnor U900 (N_900,In_867,In_1086);
and U901 (N_901,In_848,In_1745);
nor U902 (N_902,In_150,In_1688);
and U903 (N_903,N_181,In_1927);
and U904 (N_904,In_668,N_241);
nor U905 (N_905,N_452,N_172);
nor U906 (N_906,In_1233,In_648);
and U907 (N_907,N_296,In_687);
and U908 (N_908,In_194,N_420);
nor U909 (N_909,N_322,N_168);
xor U910 (N_910,N_426,In_1320);
and U911 (N_911,N_94,N_315);
nand U912 (N_912,In_660,In_109);
or U913 (N_913,N_425,N_422);
nor U914 (N_914,In_309,In_156);
nor U915 (N_915,In_689,N_389);
and U916 (N_916,In_658,N_408);
and U917 (N_917,In_738,In_1381);
nand U918 (N_918,In_159,N_216);
or U919 (N_919,In_813,In_1160);
and U920 (N_920,In_367,In_855);
and U921 (N_921,N_309,In_1435);
and U922 (N_922,N_213,In_1169);
nand U923 (N_923,N_429,N_423);
nand U924 (N_924,N_138,In_1207);
and U925 (N_925,In_1277,In_1241);
or U926 (N_926,N_353,In_1892);
nand U927 (N_927,In_1472,In_1829);
nand U928 (N_928,In_157,In_1952);
nor U929 (N_929,In_1424,N_55);
xor U930 (N_930,In_166,In_356);
nor U931 (N_931,In_242,In_413);
nand U932 (N_932,In_1274,N_54);
or U933 (N_933,In_1551,In_1728);
and U934 (N_934,In_306,In_562);
nor U935 (N_935,In_1098,N_50);
or U936 (N_936,N_112,N_0);
nor U937 (N_937,In_1907,In_1527);
xnor U938 (N_938,In_1951,N_297);
nor U939 (N_939,In_937,In_375);
xnor U940 (N_940,N_23,In_1805);
or U941 (N_941,In_947,In_593);
xor U942 (N_942,N_481,N_74);
nor U943 (N_943,In_1139,N_167);
nand U944 (N_944,In_321,In_954);
xor U945 (N_945,In_1763,N_326);
nor U946 (N_946,In_553,In_1290);
or U947 (N_947,N_25,In_1510);
nand U948 (N_948,N_70,In_1004);
nand U949 (N_949,In_428,N_245);
nand U950 (N_950,In_1450,In_152);
nor U951 (N_951,In_1496,In_1125);
xor U952 (N_952,In_677,N_200);
and U953 (N_953,In_484,In_714);
nand U954 (N_954,In_1584,N_201);
xnor U955 (N_955,In_776,In_1316);
nand U956 (N_956,In_1742,In_1734);
nand U957 (N_957,N_215,In_860);
nor U958 (N_958,In_865,In_163);
or U959 (N_959,In_874,N_340);
nand U960 (N_960,In_364,N_173);
nand U961 (N_961,In_1148,In_990);
nand U962 (N_962,In_1268,N_174);
or U963 (N_963,N_301,N_44);
and U964 (N_964,N_407,N_295);
and U965 (N_965,N_430,In_922);
nand U966 (N_966,In_1364,In_487);
nor U967 (N_967,N_162,In_511);
nor U968 (N_968,N_158,In_1376);
nand U969 (N_969,N_7,In_704);
or U970 (N_970,In_17,In_1615);
nor U971 (N_971,In_701,N_244);
and U972 (N_972,In_1057,In_271);
nor U973 (N_973,N_338,In_981);
and U974 (N_974,N_415,N_114);
nand U975 (N_975,In_503,In_1801);
and U976 (N_976,In_502,N_316);
nand U977 (N_977,N_163,N_363);
xnor U978 (N_978,In_1720,In_527);
and U979 (N_979,In_830,In_1791);
nand U980 (N_980,N_199,In_763);
nor U981 (N_981,In_842,In_696);
nor U982 (N_982,In_1522,In_106);
or U983 (N_983,In_1291,In_1823);
or U984 (N_984,N_438,In_1477);
nor U985 (N_985,In_496,N_107);
nand U986 (N_986,N_347,In_1499);
or U987 (N_987,In_1889,In_914);
xnor U988 (N_988,N_153,In_1243);
nand U989 (N_989,In_423,In_1875);
xor U990 (N_990,In_930,In_933);
or U991 (N_991,In_1757,N_412);
nand U992 (N_992,In_1264,In_897);
and U993 (N_993,N_43,In_1766);
and U994 (N_994,N_498,In_515);
nor U995 (N_995,N_437,In_1981);
nor U996 (N_996,In_957,N_238);
or U997 (N_997,In_1494,In_938);
xnor U998 (N_998,In_1021,In_386);
and U999 (N_999,N_150,In_1306);
nor U1000 (N_1000,In_1149,In_1769);
nor U1001 (N_1001,In_1075,In_1601);
xnor U1002 (N_1002,N_4,In_1239);
nor U1003 (N_1003,N_582,N_780);
or U1004 (N_1004,N_1,N_562);
and U1005 (N_1005,N_642,N_674);
and U1006 (N_1006,N_719,In_788);
nor U1007 (N_1007,N_835,N_471);
xor U1008 (N_1008,In_135,N_717);
or U1009 (N_1009,N_747,N_380);
nand U1010 (N_1010,In_447,In_662);
or U1011 (N_1011,N_865,N_69);
nand U1012 (N_1012,N_646,N_714);
and U1013 (N_1013,N_961,In_767);
xnor U1014 (N_1014,In_1342,In_1620);
and U1015 (N_1015,N_860,N_777);
nor U1016 (N_1016,In_1986,In_1928);
or U1017 (N_1017,N_492,N_926);
and U1018 (N_1018,N_738,N_576);
and U1019 (N_1019,N_834,N_250);
or U1020 (N_1020,In_410,In_1079);
or U1021 (N_1021,N_287,N_607);
xnor U1022 (N_1022,In_1394,N_532);
and U1023 (N_1023,N_636,N_323);
or U1024 (N_1024,N_600,In_632);
or U1025 (N_1025,In_615,N_608);
nor U1026 (N_1026,N_594,N_293);
and U1027 (N_1027,N_982,N_779);
and U1028 (N_1028,In_381,N_515);
or U1029 (N_1029,N_506,N_771);
and U1030 (N_1030,In_257,In_1690);
or U1031 (N_1031,N_893,N_803);
and U1032 (N_1032,N_723,N_769);
and U1033 (N_1033,N_590,In_1124);
and U1034 (N_1034,In_556,N_644);
nand U1035 (N_1035,N_445,N_932);
nor U1036 (N_1036,N_592,In_102);
nor U1037 (N_1037,N_977,N_632);
nor U1038 (N_1038,In_986,N_758);
nor U1039 (N_1039,In_1115,N_935);
nand U1040 (N_1040,In_426,N_574);
nand U1041 (N_1041,N_598,In_120);
or U1042 (N_1042,N_650,In_605);
and U1043 (N_1043,N_565,N_897);
nor U1044 (N_1044,N_950,N_677);
or U1045 (N_1045,N_853,N_634);
nor U1046 (N_1046,N_306,N_566);
nand U1047 (N_1047,N_629,N_729);
or U1048 (N_1048,In_607,N_291);
nand U1049 (N_1049,In_1917,In_288);
nand U1050 (N_1050,N_404,In_1356);
xnor U1051 (N_1051,In_889,In_75);
nor U1052 (N_1052,In_245,In_509);
and U1053 (N_1053,N_658,In_277);
and U1054 (N_1054,In_1418,In_1868);
xnor U1055 (N_1055,N_857,N_610);
xnor U1056 (N_1056,In_258,N_748);
nor U1057 (N_1057,N_750,N_100);
xor U1058 (N_1058,N_917,N_807);
or U1059 (N_1059,N_567,In_711);
nand U1060 (N_1060,In_452,N_905);
nor U1061 (N_1061,N_991,N_531);
nand U1062 (N_1062,In_1476,N_583);
or U1063 (N_1063,In_1642,In_866);
nor U1064 (N_1064,N_595,N_283);
or U1065 (N_1065,In_1490,N_676);
nand U1066 (N_1066,N_211,In_465);
nor U1067 (N_1067,N_33,In_1000);
nand U1068 (N_1068,N_609,In_1965);
nand U1069 (N_1069,In_1822,N_722);
nor U1070 (N_1070,N_981,In_721);
and U1071 (N_1071,N_806,N_527);
and U1072 (N_1072,N_448,N_915);
nand U1073 (N_1073,N_432,N_702);
nand U1074 (N_1074,N_730,N_823);
nand U1075 (N_1075,N_797,N_586);
nor U1076 (N_1076,N_785,N_683);
xor U1077 (N_1077,In_982,N_446);
nor U1078 (N_1078,N_675,N_57);
xnor U1079 (N_1079,N_493,In_10);
nor U1080 (N_1080,N_772,N_637);
nor U1081 (N_1081,In_479,In_26);
nand U1082 (N_1082,N_460,N_840);
and U1083 (N_1083,N_17,N_930);
xnor U1084 (N_1084,N_770,N_541);
or U1085 (N_1085,N_596,N_698);
nand U1086 (N_1086,N_19,N_191);
nor U1087 (N_1087,N_999,In_466);
nor U1088 (N_1088,N_793,N_376);
nand U1089 (N_1089,N_396,N_265);
or U1090 (N_1090,N_505,N_392);
nand U1091 (N_1091,In_1224,N_808);
xnor U1092 (N_1092,In_204,N_667);
and U1093 (N_1093,In_115,N_951);
nor U1094 (N_1094,N_659,N_144);
and U1095 (N_1095,N_919,In_269);
nor U1096 (N_1096,N_573,In_735);
or U1097 (N_1097,In_1845,In_1725);
nor U1098 (N_1098,In_497,N_943);
and U1099 (N_1099,N_914,N_442);
nand U1100 (N_1100,N_249,N_508);
nand U1101 (N_1101,In_541,In_1359);
nand U1102 (N_1102,N_816,N_680);
and U1103 (N_1103,N_662,N_633);
xnor U1104 (N_1104,In_103,In_1565);
and U1105 (N_1105,In_566,N_742);
nand U1106 (N_1106,N_942,N_253);
xnor U1107 (N_1107,In_1787,N_997);
or U1108 (N_1108,N_954,In_390);
nor U1109 (N_1109,N_512,In_796);
and U1110 (N_1110,N_899,N_96);
nor U1111 (N_1111,N_944,In_113);
xor U1112 (N_1112,N_585,In_1768);
and U1113 (N_1113,N_229,N_931);
xnor U1114 (N_1114,In_59,N_628);
xnor U1115 (N_1115,N_649,N_751);
and U1116 (N_1116,N_351,N_720);
nand U1117 (N_1117,N_694,N_814);
or U1118 (N_1118,In_41,N_121);
nor U1119 (N_1119,N_274,N_643);
and U1120 (N_1120,N_980,In_1525);
nand U1121 (N_1121,In_1779,N_836);
xor U1122 (N_1122,N_976,In_1211);
and U1123 (N_1123,N_332,N_219);
or U1124 (N_1124,In_1539,N_819);
xor U1125 (N_1125,N_928,N_885);
and U1126 (N_1126,N_728,In_1641);
nor U1127 (N_1127,N_929,In_1438);
and U1128 (N_1128,In_1459,N_890);
nand U1129 (N_1129,N_190,N_463);
xnor U1130 (N_1130,N_907,N_883);
nand U1131 (N_1131,In_1784,N_781);
nor U1132 (N_1132,In_1202,N_762);
and U1133 (N_1133,N_978,In_1106);
nor U1134 (N_1134,In_1548,N_186);
xor U1135 (N_1135,N_837,N_992);
xor U1136 (N_1136,N_578,N_490);
xnor U1137 (N_1137,N_821,N_875);
xnor U1138 (N_1138,N_904,N_491);
xor U1139 (N_1139,In_653,N_734);
xor U1140 (N_1140,N_966,N_533);
and U1141 (N_1141,N_557,N_612);
and U1142 (N_1142,N_888,N_861);
and U1143 (N_1143,In_1988,In_19);
xor U1144 (N_1144,N_604,N_733);
xor U1145 (N_1145,In_580,N_560);
or U1146 (N_1146,N_356,In_1029);
or U1147 (N_1147,N_546,In_1653);
nand U1148 (N_1148,N_625,In_419);
and U1149 (N_1149,N_264,N_724);
nand U1150 (N_1150,N_358,N_630);
or U1151 (N_1151,In_557,In_1558);
nand U1152 (N_1152,In_1439,In_1602);
xnor U1153 (N_1153,In_1731,In_4);
nor U1154 (N_1154,N_872,In_44);
nor U1155 (N_1155,In_1427,N_563);
xor U1156 (N_1156,N_631,N_640);
or U1157 (N_1157,In_1695,N_623);
or U1158 (N_1158,In_488,N_827);
nor U1159 (N_1159,In_1116,N_156);
xor U1160 (N_1160,N_635,N_666);
or U1161 (N_1161,In_1897,In_448);
and U1162 (N_1162,N_193,N_817);
or U1163 (N_1163,In_1506,N_801);
xor U1164 (N_1164,In_861,N_735);
xnor U1165 (N_1165,N_336,In_1007);
or U1166 (N_1166,N_593,N_152);
and U1167 (N_1167,N_903,N_968);
or U1168 (N_1168,In_1781,In_1843);
and U1169 (N_1169,N_796,In_1942);
and U1170 (N_1170,In_722,N_555);
nand U1171 (N_1171,In_88,N_656);
nor U1172 (N_1172,In_1795,N_572);
or U1173 (N_1173,In_1609,N_985);
and U1174 (N_1174,N_715,In_1392);
and U1175 (N_1175,In_380,N_262);
xor U1176 (N_1176,In_1035,N_937);
and U1177 (N_1177,N_398,In_1600);
nor U1178 (N_1178,In_1974,In_998);
and U1179 (N_1179,N_681,N_461);
and U1180 (N_1180,N_870,In_1575);
xor U1181 (N_1181,N_761,In_1778);
or U1182 (N_1182,N_105,N_941);
nand U1183 (N_1183,N_707,In_1634);
and U1184 (N_1184,In_1346,N_916);
nand U1185 (N_1185,N_401,N_535);
nor U1186 (N_1186,In_1375,N_599);
xnor U1187 (N_1187,In_1123,N_434);
nand U1188 (N_1188,In_744,N_804);
xnor U1189 (N_1189,In_859,N_179);
nand U1190 (N_1190,N_994,In_1847);
or U1191 (N_1191,In_1987,N_476);
or U1192 (N_1192,N_550,N_767);
and U1193 (N_1193,N_530,N_959);
nand U1194 (N_1194,In_1797,In_1127);
or U1195 (N_1195,N_653,In_160);
or U1196 (N_1196,In_1431,N_669);
nand U1197 (N_1197,In_1599,N_502);
nor U1198 (N_1198,N_672,N_776);
nor U1199 (N_1199,N_838,In_85);
and U1200 (N_1200,N_212,N_805);
nand U1201 (N_1201,N_900,N_866);
nor U1202 (N_1202,N_744,N_782);
and U1203 (N_1203,N_745,In_197);
or U1204 (N_1204,N_290,In_167);
and U1205 (N_1205,N_575,In_63);
nor U1206 (N_1206,In_1909,N_272);
and U1207 (N_1207,N_257,N_972);
xor U1208 (N_1208,N_475,N_66);
nor U1209 (N_1209,N_679,In_1835);
and U1210 (N_1210,In_1627,N_248);
nor U1211 (N_1211,N_936,N_924);
and U1212 (N_1212,N_784,N_614);
or U1213 (N_1213,N_902,N_774);
nor U1214 (N_1214,N_741,N_202);
or U1215 (N_1215,N_209,N_989);
nor U1216 (N_1216,In_1044,N_712);
nand U1217 (N_1217,N_206,In_9);
nand U1218 (N_1218,N_588,In_280);
xor U1219 (N_1219,N_965,N_718);
nor U1220 (N_1220,N_116,N_690);
or U1221 (N_1221,In_1782,N_864);
or U1222 (N_1222,In_728,In_564);
or U1223 (N_1223,N_699,In_780);
and U1224 (N_1224,N_137,N_611);
or U1225 (N_1225,N_243,N_947);
or U1226 (N_1226,N_765,In_524);
xnor U1227 (N_1227,In_684,In_317);
and U1228 (N_1228,In_131,N_894);
nor U1229 (N_1229,N_135,In_83);
or U1230 (N_1230,N_537,In_815);
nor U1231 (N_1231,In_875,In_1540);
or U1232 (N_1232,In_1230,N_948);
and U1233 (N_1233,In_923,N_695);
xor U1234 (N_1234,N_660,N_746);
or U1235 (N_1235,N_661,N_436);
nor U1236 (N_1236,N_922,N_545);
nor U1237 (N_1237,N_394,N_911);
or U1238 (N_1238,N_945,N_645);
and U1239 (N_1239,N_67,N_549);
xnor U1240 (N_1240,N_547,N_881);
nand U1241 (N_1241,N_91,N_691);
nor U1242 (N_1242,N_987,In_1022);
or U1243 (N_1243,In_1043,In_1790);
and U1244 (N_1244,N_513,N_678);
or U1245 (N_1245,In_1819,N_616);
or U1246 (N_1246,N_320,In_335);
nor U1247 (N_1247,N_511,In_673);
xor U1248 (N_1248,In_1331,N_601);
and U1249 (N_1249,N_543,N_20);
and U1250 (N_1250,In_560,N_484);
or U1251 (N_1251,N_856,In_1935);
nand U1252 (N_1252,N_664,In_384);
nor U1253 (N_1253,N_850,N_521);
nor U1254 (N_1254,In_310,N_749);
nand U1255 (N_1255,In_1165,N_798);
and U1256 (N_1256,N_704,In_885);
nor U1257 (N_1257,N_613,N_556);
xor U1258 (N_1258,In_1553,N_974);
nand U1259 (N_1259,In_1491,N_397);
xnor U1260 (N_1260,In_572,N_846);
nor U1261 (N_1261,N_708,N_313);
xnor U1262 (N_1262,N_428,N_236);
and U1263 (N_1263,N_939,In_505);
nor U1264 (N_1264,N_148,N_688);
and U1265 (N_1265,N_848,N_570);
nand U1266 (N_1266,N_874,N_921);
or U1267 (N_1267,N_141,N_571);
and U1268 (N_1268,In_1130,N_844);
and U1269 (N_1269,N_971,N_668);
and U1270 (N_1270,In_391,In_1934);
nand U1271 (N_1271,In_1957,In_477);
nor U1272 (N_1272,N_132,N_842);
nand U1273 (N_1273,N_716,In_1457);
nor U1274 (N_1274,In_1099,N_920);
nand U1275 (N_1275,N_970,N_706);
or U1276 (N_1276,N_952,In_366);
nand U1277 (N_1277,N_584,N_953);
xnor U1278 (N_1278,N_624,N_106);
or U1279 (N_1279,In_1616,N_536);
xnor U1280 (N_1280,N_187,In_666);
and U1281 (N_1281,In_1176,N_869);
and U1282 (N_1282,In_1535,In_369);
and U1283 (N_1283,In_1318,N_892);
or U1284 (N_1284,N_354,N_260);
xnor U1285 (N_1285,In_1269,N_651);
nor U1286 (N_1286,N_757,N_652);
nand U1287 (N_1287,N_810,N_128);
xnor U1288 (N_1288,In_29,N_908);
nor U1289 (N_1289,N_433,N_587);
and U1290 (N_1290,N_568,N_453);
nor U1291 (N_1291,N_731,N_342);
xor U1292 (N_1292,In_1547,In_196);
and U1293 (N_1293,N_99,In_226);
xnor U1294 (N_1294,N_843,N_687);
or U1295 (N_1295,N_46,N_528);
or U1296 (N_1296,N_641,N_622);
and U1297 (N_1297,N_794,N_300);
and U1298 (N_1298,N_534,In_227);
and U1299 (N_1299,In_61,N_671);
and U1300 (N_1300,In_642,N_517);
nand U1301 (N_1301,In_415,N_783);
xnor U1302 (N_1302,N_852,N_194);
nor U1303 (N_1303,N_873,N_993);
xor U1304 (N_1304,N_841,In_140);
or U1305 (N_1305,N_795,In_754);
xor U1306 (N_1306,N_510,In_1036);
nor U1307 (N_1307,N_561,N_579);
nand U1308 (N_1308,In_1159,In_904);
nor U1309 (N_1309,N_83,N_544);
and U1310 (N_1310,N_488,N_32);
xnor U1311 (N_1311,In_854,N_755);
or U1312 (N_1312,In_175,N_863);
nor U1313 (N_1313,N_727,In_920);
and U1314 (N_1314,In_1501,N_829);
and U1315 (N_1315,N_809,In_1663);
nand U1316 (N_1316,N_851,N_696);
nor U1317 (N_1317,N_787,In_1901);
nand U1318 (N_1318,N_102,N_887);
nor U1319 (N_1319,N_345,In_552);
or U1320 (N_1320,In_6,In_97);
xor U1321 (N_1321,N_552,N_53);
or U1322 (N_1322,N_995,N_520);
or U1323 (N_1323,N_822,In_1367);
or U1324 (N_1324,N_686,N_768);
and U1325 (N_1325,N_591,N_346);
xnor U1326 (N_1326,N_665,In_1920);
xnor U1327 (N_1327,N_626,N_709);
or U1328 (N_1328,In_1140,N_605);
xnor U1329 (N_1329,N_621,In_376);
and U1330 (N_1330,N_539,N_960);
xnor U1331 (N_1331,N_826,N_480);
nand U1332 (N_1332,N_773,In_1857);
xor U1333 (N_1333,N_753,In_816);
nor U1334 (N_1334,In_489,N_136);
or U1335 (N_1335,In_978,N_701);
nor U1336 (N_1336,N_553,N_949);
nand U1337 (N_1337,In_1473,N_923);
or U1338 (N_1338,N_538,In_1102);
nor U1339 (N_1339,N_366,N_967);
or U1340 (N_1340,N_726,N_275);
nand U1341 (N_1341,In_56,N_388);
or U1342 (N_1342,In_1977,N_606);
or U1343 (N_1343,N_617,In_1850);
nor U1344 (N_1344,In_409,N_597);
and U1345 (N_1345,N_799,N_86);
xnor U1346 (N_1346,N_825,N_925);
or U1347 (N_1347,In_1622,In_1155);
or U1348 (N_1348,In_382,N_800);
nor U1349 (N_1349,N_811,N_333);
xnor U1350 (N_1350,In_433,In_16);
or U1351 (N_1351,N_559,In_626);
nand U1352 (N_1352,In_1505,N_760);
xor U1353 (N_1353,N_663,In_1902);
or U1354 (N_1354,N_500,N_254);
nand U1355 (N_1355,N_996,N_602);
nand U1356 (N_1356,In_1881,N_522);
and U1357 (N_1357,N_603,N_63);
nand U1358 (N_1358,N_858,In_485);
nor U1359 (N_1359,In_420,N_862);
nor U1360 (N_1360,In_1311,In_322);
or U1361 (N_1361,In_1355,In_740);
nor U1362 (N_1362,N_933,N_998);
nor U1363 (N_1363,In_863,In_1223);
nor U1364 (N_1364,N_72,In_1509);
or U1365 (N_1365,N_580,N_58);
and U1366 (N_1366,N_410,N_117);
and U1367 (N_1367,N_697,N_901);
xor U1368 (N_1368,In_1576,N_786);
nor U1369 (N_1369,N_940,N_898);
nand U1370 (N_1370,In_1188,In_514);
xnor U1371 (N_1371,N_828,In_293);
nor U1372 (N_1372,In_659,N_548);
nand U1373 (N_1373,N_754,In_1250);
and U1374 (N_1374,N_22,N_620);
nor U1375 (N_1375,In_1182,In_66);
xnor U1376 (N_1376,In_913,N_896);
and U1377 (N_1377,N_964,N_421);
xnor U1378 (N_1378,N_831,N_29);
nand U1379 (N_1379,In_1362,N_540);
nor U1380 (N_1380,In_1153,N_955);
and U1381 (N_1381,N_815,N_523);
and U1382 (N_1382,N_705,N_732);
nor U1383 (N_1383,In_1276,N_524);
nor U1384 (N_1384,In_1825,N_657);
nor U1385 (N_1385,N_223,N_518);
and U1386 (N_1386,N_169,N_344);
and U1387 (N_1387,In_837,N_895);
and U1388 (N_1388,N_984,N_884);
xnor U1389 (N_1389,N_820,In_963);
nor U1390 (N_1390,In_1078,In_80);
or U1391 (N_1391,In_1255,N_963);
nand U1392 (N_1392,N_618,N_736);
and U1393 (N_1393,In_1562,In_461);
nand U1394 (N_1394,N_764,N_910);
nand U1395 (N_1395,In_1718,N_957);
nand U1396 (N_1396,In_934,In_1088);
nand U1397 (N_1397,N_673,In_770);
xor U1398 (N_1398,N_689,N_654);
or U1399 (N_1399,In_927,N_682);
or U1400 (N_1400,N_867,N_465);
nand U1401 (N_1401,In_1002,In_588);
nor U1402 (N_1402,N_139,N_110);
or U1403 (N_1403,N_886,In_1292);
nand U1404 (N_1404,In_1200,N_876);
nand U1405 (N_1405,N_79,N_775);
or U1406 (N_1406,N_551,In_1758);
nor U1407 (N_1407,N_849,N_983);
or U1408 (N_1408,N_526,N_525);
or U1409 (N_1409,In_5,N_558);
nor U1410 (N_1410,N_507,N_839);
nand U1411 (N_1411,In_523,In_987);
nand U1412 (N_1412,In_617,N_35);
or U1413 (N_1413,N_564,N_946);
nand U1414 (N_1414,N_956,N_648);
and U1415 (N_1415,In_940,N_503);
and U1416 (N_1416,N_721,In_705);
nor U1417 (N_1417,N_589,N_627);
and U1418 (N_1418,N_684,In_516);
nor U1419 (N_1419,N_123,In_1969);
nor U1420 (N_1420,N_581,In_1750);
nor U1421 (N_1421,N_855,N_962);
nand U1422 (N_1422,N_824,In_746);
and U1423 (N_1423,N_912,N_788);
nor U1424 (N_1424,In_344,N_280);
xnor U1425 (N_1425,N_384,N_516);
xnor U1426 (N_1426,In_926,N_766);
xor U1427 (N_1427,N_233,N_252);
nor U1428 (N_1428,N_368,N_878);
xor U1429 (N_1429,N_334,N_847);
xnor U1430 (N_1430,N_791,N_286);
or U1431 (N_1431,N_655,N_416);
nor U1432 (N_1432,N_725,N_845);
and U1433 (N_1433,N_790,N_308);
and U1434 (N_1434,N_973,In_207);
and U1435 (N_1435,N_927,N_880);
and U1436 (N_1436,N_509,N_321);
and U1437 (N_1437,In_1081,In_1789);
nor U1438 (N_1438,N_988,N_700);
or U1439 (N_1439,In_1549,N_871);
nand U1440 (N_1440,In_1314,N_859);
nand U1441 (N_1441,In_397,N_830);
or U1442 (N_1442,N_685,In_218);
xor U1443 (N_1443,In_1298,N_906);
xnor U1444 (N_1444,N_24,N_868);
nand U1445 (N_1445,In_1559,N_693);
nor U1446 (N_1446,In_53,N_638);
xnor U1447 (N_1447,N_752,N_692);
and U1448 (N_1448,In_459,N_737);
nor U1449 (N_1449,N_918,In_8);
or U1450 (N_1450,In_94,N_101);
or U1451 (N_1451,N_529,N_166);
nand U1452 (N_1452,N_854,N_639);
xnor U1453 (N_1453,In_50,In_757);
nand U1454 (N_1454,N_109,N_360);
and U1455 (N_1455,In_222,In_769);
nor U1456 (N_1456,N_990,In_1425);
nor U1457 (N_1457,N_877,In_1389);
nor U1458 (N_1458,N_456,In_961);
nor U1459 (N_1459,N_909,In_1925);
nor U1460 (N_1460,N_740,In_1618);
and U1461 (N_1461,N_710,N_703);
nor U1462 (N_1462,N_519,N_833);
xnor U1463 (N_1463,N_619,In_827);
or U1464 (N_1464,N_743,In_457);
xnor U1465 (N_1465,In_1673,N_879);
nand U1466 (N_1466,N_504,N_759);
and U1467 (N_1467,In_1816,N_789);
xor U1468 (N_1468,N_312,N_93);
xnor U1469 (N_1469,In_330,N_969);
nor U1470 (N_1470,In_1524,N_501);
nor U1471 (N_1471,N_975,N_818);
nor U1472 (N_1472,In_574,N_891);
or U1473 (N_1473,N_813,N_195);
nand U1474 (N_1474,N_739,N_335);
nand U1475 (N_1475,In_690,N_379);
xnor U1476 (N_1476,N_756,N_913);
nor U1477 (N_1477,N_812,N_554);
nor U1478 (N_1478,In_504,N_514);
nand U1479 (N_1479,N_341,In_1470);
or U1480 (N_1480,N_934,N_220);
nand U1481 (N_1481,N_882,In_38);
and U1482 (N_1482,N_615,In_471);
or U1483 (N_1483,N_497,N_542);
and U1484 (N_1484,In_1442,N_713);
or U1485 (N_1485,N_343,In_1279);
nand U1486 (N_1486,In_532,In_329);
and U1487 (N_1487,N_577,In_1042);
or U1488 (N_1488,N_258,N_832);
nand U1489 (N_1489,N_197,In_1282);
nand U1490 (N_1490,N_958,In_357);
or U1491 (N_1491,In_1307,In_1486);
and U1492 (N_1492,N_711,N_763);
and U1493 (N_1493,N_802,N_979);
xnor U1494 (N_1494,N_986,In_151);
xnor U1495 (N_1495,In_1204,N_210);
or U1496 (N_1496,N_792,N_569);
nor U1497 (N_1497,N_938,N_226);
and U1498 (N_1498,N_647,N_670);
nand U1499 (N_1499,N_778,N_889);
nor U1500 (N_1500,N_1118,N_1063);
xnor U1501 (N_1501,N_1089,N_1369);
or U1502 (N_1502,N_1488,N_1188);
and U1503 (N_1503,N_1301,N_1231);
nand U1504 (N_1504,N_1236,N_1145);
nand U1505 (N_1505,N_1211,N_1430);
and U1506 (N_1506,N_1273,N_1179);
xnor U1507 (N_1507,N_1127,N_1128);
or U1508 (N_1508,N_1280,N_1096);
or U1509 (N_1509,N_1029,N_1472);
nor U1510 (N_1510,N_1135,N_1092);
xnor U1511 (N_1511,N_1348,N_1104);
nand U1512 (N_1512,N_1015,N_1186);
nand U1513 (N_1513,N_1033,N_1398);
and U1514 (N_1514,N_1454,N_1489);
nand U1515 (N_1515,N_1498,N_1125);
nor U1516 (N_1516,N_1252,N_1335);
nand U1517 (N_1517,N_1134,N_1260);
nand U1518 (N_1518,N_1368,N_1317);
or U1519 (N_1519,N_1378,N_1446);
and U1520 (N_1520,N_1081,N_1285);
or U1521 (N_1521,N_1164,N_1133);
and U1522 (N_1522,N_1026,N_1069);
and U1523 (N_1523,N_1414,N_1372);
xnor U1524 (N_1524,N_1396,N_1499);
and U1525 (N_1525,N_1198,N_1084);
nand U1526 (N_1526,N_1223,N_1204);
or U1527 (N_1527,N_1436,N_1074);
or U1528 (N_1528,N_1320,N_1143);
or U1529 (N_1529,N_1195,N_1115);
and U1530 (N_1530,N_1213,N_1381);
nor U1531 (N_1531,N_1497,N_1462);
and U1532 (N_1532,N_1422,N_1185);
or U1533 (N_1533,N_1177,N_1232);
nand U1534 (N_1534,N_1058,N_1064);
or U1535 (N_1535,N_1068,N_1352);
xor U1536 (N_1536,N_1022,N_1205);
and U1537 (N_1537,N_1391,N_1382);
nand U1538 (N_1538,N_1336,N_1221);
nand U1539 (N_1539,N_1228,N_1097);
nor U1540 (N_1540,N_1018,N_1102);
nand U1541 (N_1541,N_1075,N_1191);
nor U1542 (N_1542,N_1001,N_1056);
and U1543 (N_1543,N_1024,N_1288);
nand U1544 (N_1544,N_1019,N_1367);
nand U1545 (N_1545,N_1464,N_1250);
nor U1546 (N_1546,N_1337,N_1356);
nand U1547 (N_1547,N_1131,N_1152);
and U1548 (N_1548,N_1370,N_1385);
nand U1549 (N_1549,N_1375,N_1256);
xnor U1550 (N_1550,N_1100,N_1031);
nor U1551 (N_1551,N_1116,N_1387);
xnor U1552 (N_1552,N_1479,N_1261);
nor U1553 (N_1553,N_1267,N_1389);
and U1554 (N_1554,N_1163,N_1054);
and U1555 (N_1555,N_1230,N_1399);
or U1556 (N_1556,N_1027,N_1051);
nand U1557 (N_1557,N_1235,N_1078);
and U1558 (N_1558,N_1023,N_1340);
xor U1559 (N_1559,N_1264,N_1300);
nand U1560 (N_1560,N_1234,N_1277);
xnor U1561 (N_1561,N_1302,N_1392);
nand U1562 (N_1562,N_1207,N_1243);
and U1563 (N_1563,N_1443,N_1136);
or U1564 (N_1564,N_1435,N_1222);
or U1565 (N_1565,N_1376,N_1463);
nor U1566 (N_1566,N_1431,N_1365);
or U1567 (N_1567,N_1478,N_1047);
nand U1568 (N_1568,N_1475,N_1107);
or U1569 (N_1569,N_1296,N_1388);
xor U1570 (N_1570,N_1466,N_1150);
xnor U1571 (N_1571,N_1245,N_1407);
nor U1572 (N_1572,N_1065,N_1121);
or U1573 (N_1573,N_1404,N_1181);
or U1574 (N_1574,N_1247,N_1111);
and U1575 (N_1575,N_1386,N_1343);
nor U1576 (N_1576,N_1050,N_1468);
nor U1577 (N_1577,N_1339,N_1172);
and U1578 (N_1578,N_1455,N_1000);
and U1579 (N_1579,N_1345,N_1060);
xnor U1580 (N_1580,N_1306,N_1044);
or U1581 (N_1581,N_1105,N_1144);
nand U1582 (N_1582,N_1427,N_1461);
nand U1583 (N_1583,N_1088,N_1411);
nand U1584 (N_1584,N_1083,N_1091);
xor U1585 (N_1585,N_1483,N_1149);
and U1586 (N_1586,N_1076,N_1477);
nor U1587 (N_1587,N_1201,N_1450);
nor U1588 (N_1588,N_1009,N_1330);
xnor U1589 (N_1589,N_1259,N_1032);
or U1590 (N_1590,N_1106,N_1341);
xnor U1591 (N_1591,N_1216,N_1274);
nor U1592 (N_1592,N_1449,N_1405);
xnor U1593 (N_1593,N_1268,N_1408);
nor U1594 (N_1594,N_1094,N_1217);
or U1595 (N_1595,N_1049,N_1242);
xnor U1596 (N_1596,N_1007,N_1303);
xnor U1597 (N_1597,N_1086,N_1434);
nand U1598 (N_1598,N_1239,N_1157);
nor U1599 (N_1599,N_1020,N_1326);
nand U1600 (N_1600,N_1401,N_1146);
or U1601 (N_1601,N_1254,N_1495);
or U1602 (N_1602,N_1142,N_1406);
or U1603 (N_1603,N_1328,N_1278);
nor U1604 (N_1604,N_1439,N_1428);
and U1605 (N_1605,N_1041,N_1344);
nand U1606 (N_1606,N_1038,N_1469);
and U1607 (N_1607,N_1218,N_1057);
nand U1608 (N_1608,N_1453,N_1309);
nand U1609 (N_1609,N_1305,N_1079);
and U1610 (N_1610,N_1008,N_1117);
nor U1611 (N_1611,N_1113,N_1036);
nand U1612 (N_1612,N_1166,N_1156);
or U1613 (N_1613,N_1039,N_1310);
or U1614 (N_1614,N_1052,N_1290);
or U1615 (N_1615,N_1419,N_1071);
nor U1616 (N_1616,N_1161,N_1006);
nand U1617 (N_1617,N_1444,N_1109);
and U1618 (N_1618,N_1194,N_1284);
nand U1619 (N_1619,N_1410,N_1424);
nor U1620 (N_1620,N_1490,N_1394);
or U1621 (N_1621,N_1390,N_1361);
or U1622 (N_1622,N_1312,N_1458);
and U1623 (N_1623,N_1486,N_1255);
and U1624 (N_1624,N_1315,N_1126);
nor U1625 (N_1625,N_1360,N_1103);
nand U1626 (N_1626,N_1190,N_1002);
and U1627 (N_1627,N_1160,N_1313);
nand U1628 (N_1628,N_1433,N_1077);
nand U1629 (N_1629,N_1298,N_1383);
xnor U1630 (N_1630,N_1279,N_1429);
nand U1631 (N_1631,N_1214,N_1212);
xnor U1632 (N_1632,N_1307,N_1045);
or U1633 (N_1633,N_1493,N_1281);
nor U1634 (N_1634,N_1349,N_1293);
xnor U1635 (N_1635,N_1175,N_1187);
nor U1636 (N_1636,N_1403,N_1451);
and U1637 (N_1637,N_1353,N_1017);
nor U1638 (N_1638,N_1359,N_1229);
nand U1639 (N_1639,N_1035,N_1492);
or U1640 (N_1640,N_1496,N_1016);
and U1641 (N_1641,N_1093,N_1366);
or U1642 (N_1642,N_1206,N_1173);
nand U1643 (N_1643,N_1192,N_1225);
nand U1644 (N_1644,N_1141,N_1110);
or U1645 (N_1645,N_1059,N_1482);
nand U1646 (N_1646,N_1095,N_1416);
and U1647 (N_1647,N_1122,N_1354);
nand U1648 (N_1648,N_1154,N_1295);
or U1649 (N_1649,N_1400,N_1415);
and U1650 (N_1650,N_1271,N_1210);
xor U1651 (N_1651,N_1233,N_1108);
nor U1652 (N_1652,N_1459,N_1304);
xor U1653 (N_1653,N_1046,N_1474);
or U1654 (N_1654,N_1262,N_1276);
xnor U1655 (N_1655,N_1090,N_1413);
nand U1656 (N_1656,N_1248,N_1476);
nor U1657 (N_1657,N_1253,N_1323);
and U1658 (N_1658,N_1005,N_1409);
or U1659 (N_1659,N_1299,N_1358);
nor U1660 (N_1660,N_1004,N_1010);
and U1661 (N_1661,N_1123,N_1350);
or U1662 (N_1662,N_1316,N_1165);
nand U1663 (N_1663,N_1332,N_1291);
nor U1664 (N_1664,N_1119,N_1132);
and U1665 (N_1665,N_1030,N_1257);
nand U1666 (N_1666,N_1270,N_1470);
or U1667 (N_1667,N_1028,N_1275);
xor U1668 (N_1668,N_1003,N_1043);
and U1669 (N_1669,N_1140,N_1171);
nor U1670 (N_1670,N_1355,N_1178);
nand U1671 (N_1671,N_1485,N_1034);
nor U1672 (N_1672,N_1287,N_1491);
or U1673 (N_1673,N_1066,N_1139);
or U1674 (N_1674,N_1438,N_1246);
and U1675 (N_1675,N_1138,N_1114);
or U1676 (N_1676,N_1040,N_1471);
xnor U1677 (N_1677,N_1199,N_1425);
xnor U1678 (N_1678,N_1120,N_1319);
xor U1679 (N_1679,N_1189,N_1374);
and U1680 (N_1680,N_1238,N_1465);
or U1681 (N_1681,N_1447,N_1013);
and U1682 (N_1682,N_1318,N_1042);
and U1683 (N_1683,N_1011,N_1174);
or U1684 (N_1684,N_1266,N_1395);
and U1685 (N_1685,N_1265,N_1130);
nor U1686 (N_1686,N_1437,N_1329);
and U1687 (N_1687,N_1292,N_1258);
or U1688 (N_1688,N_1202,N_1460);
nand U1689 (N_1689,N_1012,N_1176);
nor U1690 (N_1690,N_1421,N_1321);
or U1691 (N_1691,N_1070,N_1209);
and U1692 (N_1692,N_1331,N_1347);
nor U1693 (N_1693,N_1220,N_1170);
or U1694 (N_1694,N_1197,N_1481);
nand U1695 (N_1695,N_1193,N_1112);
xor U1696 (N_1696,N_1333,N_1494);
xor U1697 (N_1697,N_1393,N_1062);
nor U1698 (N_1698,N_1241,N_1147);
and U1699 (N_1699,N_1053,N_1467);
and U1700 (N_1700,N_1371,N_1351);
or U1701 (N_1701,N_1240,N_1480);
or U1702 (N_1702,N_1440,N_1101);
nor U1703 (N_1703,N_1324,N_1373);
or U1704 (N_1704,N_1269,N_1338);
xor U1705 (N_1705,N_1021,N_1308);
or U1706 (N_1706,N_1037,N_1249);
nor U1707 (N_1707,N_1484,N_1162);
and U1708 (N_1708,N_1215,N_1473);
nor U1709 (N_1709,N_1168,N_1423);
or U1710 (N_1710,N_1448,N_1151);
nor U1711 (N_1711,N_1420,N_1283);
nor U1712 (N_1712,N_1418,N_1342);
nand U1713 (N_1713,N_1487,N_1073);
nor U1714 (N_1714,N_1124,N_1452);
nand U1715 (N_1715,N_1203,N_1048);
or U1716 (N_1716,N_1208,N_1182);
or U1717 (N_1717,N_1237,N_1379);
and U1718 (N_1718,N_1180,N_1227);
xor U1719 (N_1719,N_1155,N_1397);
nor U1720 (N_1720,N_1196,N_1224);
xor U1721 (N_1721,N_1098,N_1432);
or U1722 (N_1722,N_1325,N_1080);
nor U1723 (N_1723,N_1129,N_1363);
nor U1724 (N_1724,N_1169,N_1286);
nand U1725 (N_1725,N_1380,N_1314);
and U1726 (N_1726,N_1014,N_1384);
or U1727 (N_1727,N_1159,N_1426);
nand U1728 (N_1728,N_1377,N_1087);
nand U1729 (N_1729,N_1282,N_1025);
nor U1730 (N_1730,N_1226,N_1219);
nor U1731 (N_1731,N_1364,N_1417);
nand U1732 (N_1732,N_1334,N_1311);
nand U1733 (N_1733,N_1085,N_1456);
or U1734 (N_1734,N_1137,N_1072);
xnor U1735 (N_1735,N_1322,N_1402);
nand U1736 (N_1736,N_1184,N_1445);
nand U1737 (N_1737,N_1297,N_1357);
xor U1738 (N_1738,N_1099,N_1441);
and U1739 (N_1739,N_1148,N_1272);
nand U1740 (N_1740,N_1067,N_1082);
and U1741 (N_1741,N_1167,N_1327);
and U1742 (N_1742,N_1362,N_1200);
and U1743 (N_1743,N_1153,N_1263);
xnor U1744 (N_1744,N_1346,N_1251);
nor U1745 (N_1745,N_1158,N_1457);
or U1746 (N_1746,N_1183,N_1412);
nand U1747 (N_1747,N_1442,N_1294);
nor U1748 (N_1748,N_1289,N_1244);
xor U1749 (N_1749,N_1055,N_1061);
or U1750 (N_1750,N_1278,N_1178);
xnor U1751 (N_1751,N_1060,N_1333);
nand U1752 (N_1752,N_1187,N_1054);
nor U1753 (N_1753,N_1488,N_1476);
nor U1754 (N_1754,N_1310,N_1108);
and U1755 (N_1755,N_1110,N_1209);
and U1756 (N_1756,N_1376,N_1397);
or U1757 (N_1757,N_1197,N_1417);
nor U1758 (N_1758,N_1401,N_1012);
and U1759 (N_1759,N_1017,N_1290);
nand U1760 (N_1760,N_1044,N_1385);
or U1761 (N_1761,N_1372,N_1112);
nor U1762 (N_1762,N_1447,N_1146);
and U1763 (N_1763,N_1067,N_1268);
nand U1764 (N_1764,N_1191,N_1093);
nand U1765 (N_1765,N_1061,N_1050);
and U1766 (N_1766,N_1437,N_1462);
nor U1767 (N_1767,N_1317,N_1405);
nor U1768 (N_1768,N_1061,N_1330);
nand U1769 (N_1769,N_1063,N_1481);
and U1770 (N_1770,N_1367,N_1014);
xor U1771 (N_1771,N_1472,N_1243);
or U1772 (N_1772,N_1147,N_1234);
nand U1773 (N_1773,N_1153,N_1195);
and U1774 (N_1774,N_1254,N_1371);
nor U1775 (N_1775,N_1154,N_1045);
xor U1776 (N_1776,N_1093,N_1418);
or U1777 (N_1777,N_1390,N_1378);
and U1778 (N_1778,N_1181,N_1141);
xor U1779 (N_1779,N_1466,N_1266);
or U1780 (N_1780,N_1159,N_1168);
xor U1781 (N_1781,N_1074,N_1348);
nand U1782 (N_1782,N_1242,N_1180);
and U1783 (N_1783,N_1464,N_1014);
nor U1784 (N_1784,N_1251,N_1266);
or U1785 (N_1785,N_1410,N_1006);
xor U1786 (N_1786,N_1489,N_1081);
or U1787 (N_1787,N_1199,N_1029);
nor U1788 (N_1788,N_1499,N_1283);
nor U1789 (N_1789,N_1278,N_1067);
and U1790 (N_1790,N_1116,N_1268);
or U1791 (N_1791,N_1191,N_1038);
nand U1792 (N_1792,N_1427,N_1178);
nand U1793 (N_1793,N_1059,N_1370);
nand U1794 (N_1794,N_1164,N_1395);
xnor U1795 (N_1795,N_1274,N_1247);
nor U1796 (N_1796,N_1160,N_1449);
and U1797 (N_1797,N_1233,N_1429);
xnor U1798 (N_1798,N_1197,N_1103);
xor U1799 (N_1799,N_1457,N_1305);
xor U1800 (N_1800,N_1204,N_1483);
nand U1801 (N_1801,N_1225,N_1157);
and U1802 (N_1802,N_1157,N_1220);
xnor U1803 (N_1803,N_1395,N_1494);
nor U1804 (N_1804,N_1105,N_1313);
nand U1805 (N_1805,N_1429,N_1157);
and U1806 (N_1806,N_1040,N_1432);
and U1807 (N_1807,N_1402,N_1220);
nand U1808 (N_1808,N_1212,N_1341);
and U1809 (N_1809,N_1055,N_1377);
nand U1810 (N_1810,N_1263,N_1056);
and U1811 (N_1811,N_1386,N_1074);
or U1812 (N_1812,N_1448,N_1366);
and U1813 (N_1813,N_1401,N_1440);
nor U1814 (N_1814,N_1100,N_1092);
nand U1815 (N_1815,N_1297,N_1199);
nor U1816 (N_1816,N_1002,N_1206);
xor U1817 (N_1817,N_1191,N_1470);
nor U1818 (N_1818,N_1306,N_1094);
and U1819 (N_1819,N_1499,N_1193);
nor U1820 (N_1820,N_1146,N_1180);
xnor U1821 (N_1821,N_1061,N_1225);
nand U1822 (N_1822,N_1043,N_1265);
nor U1823 (N_1823,N_1125,N_1222);
nand U1824 (N_1824,N_1287,N_1160);
nor U1825 (N_1825,N_1490,N_1037);
xor U1826 (N_1826,N_1024,N_1068);
and U1827 (N_1827,N_1332,N_1444);
nand U1828 (N_1828,N_1368,N_1089);
xor U1829 (N_1829,N_1414,N_1249);
xnor U1830 (N_1830,N_1362,N_1257);
xnor U1831 (N_1831,N_1030,N_1227);
or U1832 (N_1832,N_1387,N_1024);
or U1833 (N_1833,N_1297,N_1065);
and U1834 (N_1834,N_1275,N_1279);
nand U1835 (N_1835,N_1285,N_1414);
or U1836 (N_1836,N_1406,N_1215);
and U1837 (N_1837,N_1423,N_1091);
nand U1838 (N_1838,N_1384,N_1307);
and U1839 (N_1839,N_1411,N_1121);
xnor U1840 (N_1840,N_1127,N_1135);
and U1841 (N_1841,N_1244,N_1031);
or U1842 (N_1842,N_1019,N_1412);
xnor U1843 (N_1843,N_1223,N_1332);
xor U1844 (N_1844,N_1110,N_1046);
nor U1845 (N_1845,N_1442,N_1114);
nand U1846 (N_1846,N_1015,N_1036);
nand U1847 (N_1847,N_1144,N_1404);
xor U1848 (N_1848,N_1429,N_1470);
or U1849 (N_1849,N_1425,N_1441);
and U1850 (N_1850,N_1126,N_1387);
nor U1851 (N_1851,N_1232,N_1418);
nor U1852 (N_1852,N_1339,N_1492);
nand U1853 (N_1853,N_1460,N_1100);
xnor U1854 (N_1854,N_1335,N_1458);
nor U1855 (N_1855,N_1080,N_1486);
or U1856 (N_1856,N_1023,N_1123);
nand U1857 (N_1857,N_1064,N_1076);
nor U1858 (N_1858,N_1004,N_1270);
and U1859 (N_1859,N_1158,N_1309);
or U1860 (N_1860,N_1368,N_1405);
xnor U1861 (N_1861,N_1215,N_1018);
xor U1862 (N_1862,N_1007,N_1080);
or U1863 (N_1863,N_1170,N_1312);
or U1864 (N_1864,N_1029,N_1270);
xor U1865 (N_1865,N_1406,N_1357);
xor U1866 (N_1866,N_1446,N_1437);
nand U1867 (N_1867,N_1256,N_1295);
and U1868 (N_1868,N_1390,N_1294);
xor U1869 (N_1869,N_1162,N_1485);
nand U1870 (N_1870,N_1381,N_1346);
nand U1871 (N_1871,N_1383,N_1438);
xnor U1872 (N_1872,N_1316,N_1140);
nand U1873 (N_1873,N_1263,N_1016);
or U1874 (N_1874,N_1132,N_1060);
or U1875 (N_1875,N_1034,N_1197);
nor U1876 (N_1876,N_1203,N_1042);
and U1877 (N_1877,N_1218,N_1422);
nand U1878 (N_1878,N_1208,N_1322);
nand U1879 (N_1879,N_1137,N_1011);
xor U1880 (N_1880,N_1107,N_1271);
or U1881 (N_1881,N_1092,N_1166);
nand U1882 (N_1882,N_1320,N_1307);
nand U1883 (N_1883,N_1181,N_1483);
and U1884 (N_1884,N_1484,N_1086);
nand U1885 (N_1885,N_1374,N_1141);
nand U1886 (N_1886,N_1230,N_1471);
nand U1887 (N_1887,N_1352,N_1320);
and U1888 (N_1888,N_1184,N_1186);
nor U1889 (N_1889,N_1034,N_1133);
nor U1890 (N_1890,N_1163,N_1321);
nand U1891 (N_1891,N_1267,N_1121);
nand U1892 (N_1892,N_1046,N_1327);
xnor U1893 (N_1893,N_1071,N_1219);
and U1894 (N_1894,N_1211,N_1215);
nand U1895 (N_1895,N_1488,N_1308);
nor U1896 (N_1896,N_1045,N_1323);
nand U1897 (N_1897,N_1118,N_1206);
nand U1898 (N_1898,N_1348,N_1030);
nand U1899 (N_1899,N_1479,N_1263);
or U1900 (N_1900,N_1396,N_1342);
or U1901 (N_1901,N_1224,N_1080);
or U1902 (N_1902,N_1345,N_1134);
and U1903 (N_1903,N_1360,N_1070);
xnor U1904 (N_1904,N_1109,N_1232);
nor U1905 (N_1905,N_1153,N_1428);
and U1906 (N_1906,N_1361,N_1157);
or U1907 (N_1907,N_1210,N_1280);
or U1908 (N_1908,N_1183,N_1045);
nor U1909 (N_1909,N_1143,N_1206);
nand U1910 (N_1910,N_1399,N_1246);
nand U1911 (N_1911,N_1215,N_1420);
and U1912 (N_1912,N_1413,N_1108);
nand U1913 (N_1913,N_1345,N_1138);
nor U1914 (N_1914,N_1463,N_1345);
xnor U1915 (N_1915,N_1054,N_1434);
or U1916 (N_1916,N_1190,N_1192);
and U1917 (N_1917,N_1142,N_1109);
nand U1918 (N_1918,N_1275,N_1119);
nor U1919 (N_1919,N_1216,N_1470);
and U1920 (N_1920,N_1191,N_1489);
nor U1921 (N_1921,N_1364,N_1095);
xnor U1922 (N_1922,N_1174,N_1466);
or U1923 (N_1923,N_1370,N_1465);
nand U1924 (N_1924,N_1100,N_1042);
nor U1925 (N_1925,N_1022,N_1117);
and U1926 (N_1926,N_1138,N_1488);
or U1927 (N_1927,N_1367,N_1011);
nor U1928 (N_1928,N_1293,N_1351);
nor U1929 (N_1929,N_1109,N_1318);
or U1930 (N_1930,N_1082,N_1102);
or U1931 (N_1931,N_1151,N_1378);
xnor U1932 (N_1932,N_1167,N_1437);
or U1933 (N_1933,N_1144,N_1038);
nor U1934 (N_1934,N_1144,N_1145);
or U1935 (N_1935,N_1059,N_1014);
and U1936 (N_1936,N_1215,N_1395);
nand U1937 (N_1937,N_1237,N_1246);
xnor U1938 (N_1938,N_1112,N_1077);
or U1939 (N_1939,N_1395,N_1129);
nor U1940 (N_1940,N_1280,N_1497);
nor U1941 (N_1941,N_1465,N_1058);
and U1942 (N_1942,N_1216,N_1317);
or U1943 (N_1943,N_1107,N_1106);
and U1944 (N_1944,N_1103,N_1145);
nor U1945 (N_1945,N_1323,N_1276);
nand U1946 (N_1946,N_1461,N_1496);
nand U1947 (N_1947,N_1409,N_1156);
or U1948 (N_1948,N_1055,N_1246);
nand U1949 (N_1949,N_1376,N_1264);
xnor U1950 (N_1950,N_1029,N_1356);
or U1951 (N_1951,N_1317,N_1342);
nand U1952 (N_1952,N_1101,N_1371);
nand U1953 (N_1953,N_1236,N_1400);
nor U1954 (N_1954,N_1250,N_1329);
and U1955 (N_1955,N_1250,N_1387);
or U1956 (N_1956,N_1367,N_1308);
xnor U1957 (N_1957,N_1305,N_1302);
and U1958 (N_1958,N_1139,N_1299);
xor U1959 (N_1959,N_1361,N_1256);
xnor U1960 (N_1960,N_1443,N_1056);
nand U1961 (N_1961,N_1193,N_1358);
xnor U1962 (N_1962,N_1220,N_1101);
nor U1963 (N_1963,N_1045,N_1189);
and U1964 (N_1964,N_1275,N_1262);
nand U1965 (N_1965,N_1086,N_1424);
nand U1966 (N_1966,N_1483,N_1275);
or U1967 (N_1967,N_1467,N_1138);
nand U1968 (N_1968,N_1007,N_1442);
and U1969 (N_1969,N_1075,N_1142);
nand U1970 (N_1970,N_1308,N_1136);
nor U1971 (N_1971,N_1465,N_1085);
or U1972 (N_1972,N_1069,N_1478);
xnor U1973 (N_1973,N_1296,N_1219);
nand U1974 (N_1974,N_1039,N_1452);
xor U1975 (N_1975,N_1325,N_1478);
nand U1976 (N_1976,N_1172,N_1246);
or U1977 (N_1977,N_1286,N_1170);
nor U1978 (N_1978,N_1363,N_1047);
or U1979 (N_1979,N_1049,N_1097);
xnor U1980 (N_1980,N_1134,N_1410);
or U1981 (N_1981,N_1198,N_1465);
and U1982 (N_1982,N_1052,N_1084);
xor U1983 (N_1983,N_1030,N_1098);
xor U1984 (N_1984,N_1264,N_1315);
and U1985 (N_1985,N_1462,N_1010);
or U1986 (N_1986,N_1090,N_1303);
or U1987 (N_1987,N_1408,N_1246);
nor U1988 (N_1988,N_1477,N_1494);
and U1989 (N_1989,N_1268,N_1125);
and U1990 (N_1990,N_1484,N_1077);
nor U1991 (N_1991,N_1382,N_1242);
nor U1992 (N_1992,N_1113,N_1148);
or U1993 (N_1993,N_1174,N_1190);
or U1994 (N_1994,N_1264,N_1295);
nand U1995 (N_1995,N_1191,N_1264);
xor U1996 (N_1996,N_1228,N_1198);
nand U1997 (N_1997,N_1342,N_1171);
or U1998 (N_1998,N_1337,N_1228);
or U1999 (N_1999,N_1103,N_1490);
or U2000 (N_2000,N_1728,N_1999);
nor U2001 (N_2001,N_1757,N_1841);
xnor U2002 (N_2002,N_1525,N_1900);
xor U2003 (N_2003,N_1897,N_1684);
xnor U2004 (N_2004,N_1520,N_1574);
and U2005 (N_2005,N_1537,N_1563);
nand U2006 (N_2006,N_1854,N_1699);
nor U2007 (N_2007,N_1805,N_1935);
xor U2008 (N_2008,N_1603,N_1503);
and U2009 (N_2009,N_1530,N_1814);
nand U2010 (N_2010,N_1949,N_1706);
nor U2011 (N_2011,N_1785,N_1670);
nand U2012 (N_2012,N_1830,N_1736);
or U2013 (N_2013,N_1746,N_1857);
and U2014 (N_2014,N_1501,N_1884);
nor U2015 (N_2015,N_1961,N_1981);
and U2016 (N_2016,N_1950,N_1808);
and U2017 (N_2017,N_1952,N_1708);
nand U2018 (N_2018,N_1716,N_1998);
nand U2019 (N_2019,N_1945,N_1681);
xnor U2020 (N_2020,N_1823,N_1820);
nand U2021 (N_2021,N_1564,N_1985);
or U2022 (N_2022,N_1738,N_1538);
nand U2023 (N_2023,N_1559,N_1722);
nand U2024 (N_2024,N_1558,N_1973);
xor U2025 (N_2025,N_1774,N_1509);
and U2026 (N_2026,N_1894,N_1575);
and U2027 (N_2027,N_1778,N_1694);
xor U2028 (N_2028,N_1861,N_1695);
nor U2029 (N_2029,N_1828,N_1636);
xor U2030 (N_2030,N_1697,N_1733);
or U2031 (N_2031,N_1764,N_1683);
xnor U2032 (N_2032,N_1522,N_1605);
nor U2033 (N_2033,N_1944,N_1580);
nand U2034 (N_2034,N_1989,N_1729);
nor U2035 (N_2035,N_1827,N_1844);
nand U2036 (N_2036,N_1565,N_1920);
and U2037 (N_2037,N_1658,N_1631);
nand U2038 (N_2038,N_1882,N_1782);
nor U2039 (N_2039,N_1514,N_1704);
or U2040 (N_2040,N_1506,N_1690);
nor U2041 (N_2041,N_1616,N_1640);
and U2042 (N_2042,N_1784,N_1671);
nand U2043 (N_2043,N_1531,N_1901);
nand U2044 (N_2044,N_1698,N_1758);
nand U2045 (N_2045,N_1578,N_1890);
nor U2046 (N_2046,N_1891,N_1995);
or U2047 (N_2047,N_1988,N_1980);
xor U2048 (N_2048,N_1510,N_1969);
or U2049 (N_2049,N_1773,N_1753);
or U2050 (N_2050,N_1652,N_1613);
nand U2051 (N_2051,N_1585,N_1789);
xor U2052 (N_2052,N_1769,N_1781);
and U2053 (N_2053,N_1889,N_1913);
nand U2054 (N_2054,N_1802,N_1860);
nor U2055 (N_2055,N_1731,N_1555);
and U2056 (N_2056,N_1819,N_1834);
and U2057 (N_2057,N_1798,N_1760);
and U2058 (N_2058,N_1502,N_1922);
or U2059 (N_2059,N_1957,N_1593);
nor U2060 (N_2060,N_1788,N_1546);
nand U2061 (N_2061,N_1919,N_1879);
and U2062 (N_2062,N_1902,N_1584);
xor U2063 (N_2063,N_1673,N_1598);
and U2064 (N_2064,N_1748,N_1526);
or U2065 (N_2065,N_1977,N_1549);
or U2066 (N_2066,N_1590,N_1840);
xor U2067 (N_2067,N_1835,N_1836);
and U2068 (N_2068,N_1553,N_1843);
and U2069 (N_2069,N_1818,N_1669);
or U2070 (N_2070,N_1915,N_1972);
or U2071 (N_2071,N_1982,N_1907);
and U2072 (N_2072,N_1679,N_1839);
nor U2073 (N_2073,N_1664,N_1693);
nor U2074 (N_2074,N_1606,N_1622);
xnor U2075 (N_2075,N_1872,N_1583);
nor U2076 (N_2076,N_1570,N_1617);
nor U2077 (N_2077,N_1682,N_1554);
xnor U2078 (N_2078,N_1749,N_1816);
xor U2079 (N_2079,N_1809,N_1858);
and U2080 (N_2080,N_1639,N_1633);
nand U2081 (N_2081,N_1507,N_1552);
nand U2082 (N_2082,N_1876,N_1523);
and U2083 (N_2083,N_1703,N_1938);
nor U2084 (N_2084,N_1667,N_1562);
and U2085 (N_2085,N_1833,N_1672);
nor U2086 (N_2086,N_1853,N_1511);
or U2087 (N_2087,N_1692,N_1568);
and U2088 (N_2088,N_1874,N_1971);
and U2089 (N_2089,N_1615,N_1655);
or U2090 (N_2090,N_1790,N_1638);
nand U2091 (N_2091,N_1586,N_1875);
nand U2092 (N_2092,N_1528,N_1625);
and U2093 (N_2093,N_1661,N_1926);
or U2094 (N_2094,N_1515,N_1817);
xnor U2095 (N_2095,N_1573,N_1850);
nor U2096 (N_2096,N_1536,N_1637);
or U2097 (N_2097,N_1803,N_1936);
and U2098 (N_2098,N_1963,N_1619);
and U2099 (N_2099,N_1842,N_1723);
nand U2100 (N_2100,N_1734,N_1826);
nor U2101 (N_2101,N_1984,N_1567);
nand U2102 (N_2102,N_1862,N_1621);
nor U2103 (N_2103,N_1801,N_1524);
xnor U2104 (N_2104,N_1966,N_1696);
nor U2105 (N_2105,N_1540,N_1591);
and U2106 (N_2106,N_1635,N_1620);
xnor U2107 (N_2107,N_1904,N_1737);
nand U2108 (N_2108,N_1940,N_1886);
or U2109 (N_2109,N_1707,N_1608);
and U2110 (N_2110,N_1800,N_1701);
nor U2111 (N_2111,N_1983,N_1687);
nor U2112 (N_2112,N_1856,N_1838);
and U2113 (N_2113,N_1614,N_1885);
xnor U2114 (N_2114,N_1965,N_1867);
and U2115 (N_2115,N_1676,N_1576);
and U2116 (N_2116,N_1776,N_1933);
and U2117 (N_2117,N_1718,N_1508);
and U2118 (N_2118,N_1715,N_1588);
nand U2119 (N_2119,N_1765,N_1986);
and U2120 (N_2120,N_1993,N_1812);
xnor U2121 (N_2121,N_1516,N_1551);
nor U2122 (N_2122,N_1914,N_1775);
nor U2123 (N_2123,N_1806,N_1767);
xor U2124 (N_2124,N_1651,N_1744);
and U2125 (N_2125,N_1990,N_1727);
nor U2126 (N_2126,N_1942,N_1877);
xor U2127 (N_2127,N_1941,N_1925);
and U2128 (N_2128,N_1864,N_1970);
nand U2129 (N_2129,N_1791,N_1632);
or U2130 (N_2130,N_1954,N_1712);
xnor U2131 (N_2131,N_1675,N_1871);
and U2132 (N_2132,N_1725,N_1500);
or U2133 (N_2133,N_1743,N_1624);
nor U2134 (N_2134,N_1618,N_1921);
nor U2135 (N_2135,N_1880,N_1717);
xor U2136 (N_2136,N_1866,N_1589);
and U2137 (N_2137,N_1943,N_1688);
or U2138 (N_2138,N_1710,N_1587);
xnor U2139 (N_2139,N_1566,N_1807);
or U2140 (N_2140,N_1815,N_1519);
nand U2141 (N_2141,N_1911,N_1822);
and U2142 (N_2142,N_1611,N_1918);
or U2143 (N_2143,N_1799,N_1931);
nand U2144 (N_2144,N_1662,N_1813);
xor U2145 (N_2145,N_1832,N_1974);
nand U2146 (N_2146,N_1689,N_1545);
nor U2147 (N_2147,N_1958,N_1997);
xnor U2148 (N_2148,N_1577,N_1724);
nand U2149 (N_2149,N_1649,N_1923);
and U2150 (N_2150,N_1992,N_1865);
nor U2151 (N_2151,N_1975,N_1711);
xnor U2152 (N_2152,N_1668,N_1595);
nor U2153 (N_2153,N_1794,N_1709);
xnor U2154 (N_2154,N_1740,N_1512);
xor U2155 (N_2155,N_1571,N_1592);
xor U2156 (N_2156,N_1561,N_1987);
xor U2157 (N_2157,N_1648,N_1582);
nor U2158 (N_2158,N_1599,N_1755);
or U2159 (N_2159,N_1930,N_1761);
nand U2160 (N_2160,N_1521,N_1542);
xnor U2161 (N_2161,N_1517,N_1581);
nor U2162 (N_2162,N_1654,N_1527);
or U2163 (N_2163,N_1906,N_1978);
nand U2164 (N_2164,N_1917,N_1887);
xor U2165 (N_2165,N_1825,N_1888);
or U2166 (N_2166,N_1653,N_1747);
or U2167 (N_2167,N_1645,N_1666);
and U2168 (N_2168,N_1869,N_1626);
and U2169 (N_2169,N_1529,N_1610);
and U2170 (N_2170,N_1903,N_1951);
xnor U2171 (N_2171,N_1873,N_1726);
xnor U2172 (N_2172,N_1685,N_1837);
nand U2173 (N_2173,N_1870,N_1910);
xor U2174 (N_2174,N_1787,N_1691);
or U2175 (N_2175,N_1560,N_1750);
xnor U2176 (N_2176,N_1678,N_1793);
xor U2177 (N_2177,N_1859,N_1629);
xnor U2178 (N_2178,N_1751,N_1602);
nor U2179 (N_2179,N_1770,N_1656);
xor U2180 (N_2180,N_1792,N_1532);
nand U2181 (N_2181,N_1641,N_1851);
or U2182 (N_2182,N_1612,N_1535);
or U2183 (N_2183,N_1766,N_1518);
nor U2184 (N_2184,N_1829,N_1948);
xnor U2185 (N_2185,N_1735,N_1924);
nor U2186 (N_2186,N_1821,N_1991);
or U2187 (N_2187,N_1883,N_1927);
nor U2188 (N_2188,N_1557,N_1643);
nand U2189 (N_2189,N_1804,N_1539);
and U2190 (N_2190,N_1634,N_1847);
nand U2191 (N_2191,N_1759,N_1763);
and U2192 (N_2192,N_1964,N_1863);
xnor U2193 (N_2193,N_1505,N_1541);
nor U2194 (N_2194,N_1777,N_1929);
or U2195 (N_2195,N_1786,N_1946);
nor U2196 (N_2196,N_1912,N_1579);
or U2197 (N_2197,N_1752,N_1601);
and U2198 (N_2198,N_1713,N_1721);
and U2199 (N_2199,N_1644,N_1534);
nand U2200 (N_2200,N_1953,N_1934);
nand U2201 (N_2201,N_1596,N_1979);
nand U2202 (N_2202,N_1771,N_1796);
or U2203 (N_2203,N_1650,N_1878);
or U2204 (N_2204,N_1756,N_1892);
nor U2205 (N_2205,N_1594,N_1881);
and U2206 (N_2206,N_1659,N_1895);
and U2207 (N_2207,N_1928,N_1848);
or U2208 (N_2208,N_1754,N_1810);
and U2209 (N_2209,N_1600,N_1623);
xor U2210 (N_2210,N_1959,N_1745);
or U2211 (N_2211,N_1908,N_1968);
xnor U2212 (N_2212,N_1607,N_1762);
or U2213 (N_2213,N_1896,N_1646);
nand U2214 (N_2214,N_1960,N_1956);
or U2215 (N_2215,N_1544,N_1939);
and U2216 (N_2216,N_1783,N_1852);
or U2217 (N_2217,N_1660,N_1994);
nor U2218 (N_2218,N_1811,N_1677);
or U2219 (N_2219,N_1720,N_1647);
nor U2220 (N_2220,N_1909,N_1597);
nor U2221 (N_2221,N_1665,N_1642);
nor U2222 (N_2222,N_1898,N_1609);
and U2223 (N_2223,N_1732,N_1947);
xnor U2224 (N_2224,N_1779,N_1996);
nor U2225 (N_2225,N_1627,N_1976);
and U2226 (N_2226,N_1937,N_1932);
nor U2227 (N_2227,N_1550,N_1849);
xor U2228 (N_2228,N_1702,N_1899);
and U2229 (N_2229,N_1780,N_1556);
nand U2230 (N_2230,N_1741,N_1705);
nor U2231 (N_2231,N_1797,N_1893);
or U2232 (N_2232,N_1962,N_1855);
and U2233 (N_2233,N_1768,N_1845);
nand U2234 (N_2234,N_1569,N_1739);
nor U2235 (N_2235,N_1868,N_1663);
nor U2236 (N_2236,N_1628,N_1742);
nand U2237 (N_2237,N_1846,N_1719);
and U2238 (N_2238,N_1916,N_1772);
and U2239 (N_2239,N_1831,N_1714);
nand U2240 (N_2240,N_1905,N_1630);
xor U2241 (N_2241,N_1657,N_1504);
and U2242 (N_2242,N_1700,N_1572);
and U2243 (N_2243,N_1513,N_1533);
or U2244 (N_2244,N_1955,N_1795);
nand U2245 (N_2245,N_1730,N_1824);
and U2246 (N_2246,N_1548,N_1967);
nand U2247 (N_2247,N_1674,N_1604);
xor U2248 (N_2248,N_1686,N_1543);
or U2249 (N_2249,N_1547,N_1680);
xnor U2250 (N_2250,N_1754,N_1680);
and U2251 (N_2251,N_1579,N_1776);
and U2252 (N_2252,N_1939,N_1597);
nor U2253 (N_2253,N_1501,N_1584);
nor U2254 (N_2254,N_1567,N_1568);
and U2255 (N_2255,N_1579,N_1622);
xor U2256 (N_2256,N_1932,N_1903);
nand U2257 (N_2257,N_1522,N_1988);
nor U2258 (N_2258,N_1778,N_1584);
and U2259 (N_2259,N_1763,N_1677);
xor U2260 (N_2260,N_1719,N_1643);
nor U2261 (N_2261,N_1629,N_1785);
nor U2262 (N_2262,N_1955,N_1680);
or U2263 (N_2263,N_1575,N_1756);
or U2264 (N_2264,N_1552,N_1930);
and U2265 (N_2265,N_1728,N_1526);
xor U2266 (N_2266,N_1566,N_1777);
or U2267 (N_2267,N_1527,N_1614);
or U2268 (N_2268,N_1979,N_1731);
nor U2269 (N_2269,N_1737,N_1990);
or U2270 (N_2270,N_1858,N_1950);
and U2271 (N_2271,N_1871,N_1714);
xnor U2272 (N_2272,N_1506,N_1607);
and U2273 (N_2273,N_1679,N_1700);
nand U2274 (N_2274,N_1564,N_1611);
xnor U2275 (N_2275,N_1932,N_1639);
and U2276 (N_2276,N_1777,N_1733);
nand U2277 (N_2277,N_1910,N_1715);
nor U2278 (N_2278,N_1643,N_1930);
nand U2279 (N_2279,N_1848,N_1996);
xnor U2280 (N_2280,N_1770,N_1505);
nand U2281 (N_2281,N_1947,N_1500);
or U2282 (N_2282,N_1921,N_1504);
or U2283 (N_2283,N_1968,N_1741);
and U2284 (N_2284,N_1988,N_1973);
nand U2285 (N_2285,N_1852,N_1741);
nor U2286 (N_2286,N_1515,N_1691);
nor U2287 (N_2287,N_1716,N_1973);
or U2288 (N_2288,N_1686,N_1983);
or U2289 (N_2289,N_1869,N_1786);
xor U2290 (N_2290,N_1533,N_1522);
xnor U2291 (N_2291,N_1843,N_1756);
and U2292 (N_2292,N_1870,N_1648);
and U2293 (N_2293,N_1895,N_1560);
or U2294 (N_2294,N_1888,N_1686);
nor U2295 (N_2295,N_1767,N_1651);
nor U2296 (N_2296,N_1625,N_1802);
xor U2297 (N_2297,N_1704,N_1981);
or U2298 (N_2298,N_1661,N_1899);
or U2299 (N_2299,N_1742,N_1656);
and U2300 (N_2300,N_1853,N_1860);
and U2301 (N_2301,N_1583,N_1864);
nand U2302 (N_2302,N_1795,N_1904);
xnor U2303 (N_2303,N_1981,N_1912);
xnor U2304 (N_2304,N_1585,N_1859);
or U2305 (N_2305,N_1740,N_1729);
nand U2306 (N_2306,N_1842,N_1548);
nor U2307 (N_2307,N_1866,N_1930);
or U2308 (N_2308,N_1755,N_1817);
xor U2309 (N_2309,N_1531,N_1601);
or U2310 (N_2310,N_1907,N_1714);
nor U2311 (N_2311,N_1895,N_1756);
or U2312 (N_2312,N_1858,N_1750);
or U2313 (N_2313,N_1872,N_1718);
and U2314 (N_2314,N_1590,N_1912);
xnor U2315 (N_2315,N_1567,N_1716);
and U2316 (N_2316,N_1982,N_1767);
or U2317 (N_2317,N_1578,N_1790);
nor U2318 (N_2318,N_1546,N_1784);
xnor U2319 (N_2319,N_1536,N_1772);
and U2320 (N_2320,N_1980,N_1627);
or U2321 (N_2321,N_1985,N_1683);
or U2322 (N_2322,N_1565,N_1720);
or U2323 (N_2323,N_1697,N_1833);
xor U2324 (N_2324,N_1884,N_1880);
nor U2325 (N_2325,N_1960,N_1852);
nand U2326 (N_2326,N_1904,N_1732);
nor U2327 (N_2327,N_1694,N_1709);
xor U2328 (N_2328,N_1922,N_1899);
nand U2329 (N_2329,N_1925,N_1898);
or U2330 (N_2330,N_1536,N_1845);
nor U2331 (N_2331,N_1810,N_1544);
nand U2332 (N_2332,N_1593,N_1533);
xor U2333 (N_2333,N_1785,N_1725);
or U2334 (N_2334,N_1832,N_1966);
and U2335 (N_2335,N_1868,N_1661);
xnor U2336 (N_2336,N_1860,N_1648);
xor U2337 (N_2337,N_1970,N_1687);
nor U2338 (N_2338,N_1877,N_1940);
nor U2339 (N_2339,N_1961,N_1953);
and U2340 (N_2340,N_1846,N_1835);
nand U2341 (N_2341,N_1613,N_1579);
nand U2342 (N_2342,N_1769,N_1941);
xnor U2343 (N_2343,N_1880,N_1941);
nand U2344 (N_2344,N_1690,N_1737);
nand U2345 (N_2345,N_1890,N_1723);
nand U2346 (N_2346,N_1678,N_1530);
and U2347 (N_2347,N_1514,N_1705);
xnor U2348 (N_2348,N_1689,N_1738);
nor U2349 (N_2349,N_1554,N_1795);
xor U2350 (N_2350,N_1649,N_1672);
or U2351 (N_2351,N_1772,N_1865);
nor U2352 (N_2352,N_1754,N_1830);
or U2353 (N_2353,N_1621,N_1596);
and U2354 (N_2354,N_1769,N_1816);
xor U2355 (N_2355,N_1992,N_1824);
and U2356 (N_2356,N_1522,N_1959);
and U2357 (N_2357,N_1829,N_1872);
xor U2358 (N_2358,N_1881,N_1812);
or U2359 (N_2359,N_1546,N_1753);
nand U2360 (N_2360,N_1880,N_1955);
nand U2361 (N_2361,N_1868,N_1697);
nand U2362 (N_2362,N_1643,N_1823);
and U2363 (N_2363,N_1751,N_1826);
xnor U2364 (N_2364,N_1649,N_1771);
or U2365 (N_2365,N_1504,N_1629);
and U2366 (N_2366,N_1746,N_1673);
nand U2367 (N_2367,N_1813,N_1748);
and U2368 (N_2368,N_1730,N_1650);
nor U2369 (N_2369,N_1966,N_1543);
or U2370 (N_2370,N_1602,N_1939);
or U2371 (N_2371,N_1596,N_1947);
or U2372 (N_2372,N_1846,N_1937);
and U2373 (N_2373,N_1596,N_1789);
and U2374 (N_2374,N_1913,N_1699);
or U2375 (N_2375,N_1861,N_1593);
xnor U2376 (N_2376,N_1571,N_1771);
and U2377 (N_2377,N_1850,N_1961);
xnor U2378 (N_2378,N_1982,N_1571);
nand U2379 (N_2379,N_1697,N_1713);
nand U2380 (N_2380,N_1942,N_1954);
xor U2381 (N_2381,N_1884,N_1608);
nor U2382 (N_2382,N_1741,N_1908);
or U2383 (N_2383,N_1862,N_1968);
or U2384 (N_2384,N_1703,N_1604);
xor U2385 (N_2385,N_1585,N_1793);
nand U2386 (N_2386,N_1819,N_1674);
or U2387 (N_2387,N_1512,N_1890);
nand U2388 (N_2388,N_1791,N_1569);
or U2389 (N_2389,N_1700,N_1640);
xor U2390 (N_2390,N_1628,N_1892);
nor U2391 (N_2391,N_1529,N_1917);
or U2392 (N_2392,N_1796,N_1533);
nand U2393 (N_2393,N_1843,N_1801);
nand U2394 (N_2394,N_1697,N_1968);
nor U2395 (N_2395,N_1665,N_1531);
and U2396 (N_2396,N_1978,N_1555);
nor U2397 (N_2397,N_1710,N_1849);
xnor U2398 (N_2398,N_1807,N_1837);
nor U2399 (N_2399,N_1842,N_1685);
or U2400 (N_2400,N_1690,N_1613);
or U2401 (N_2401,N_1633,N_1816);
xor U2402 (N_2402,N_1715,N_1973);
nor U2403 (N_2403,N_1803,N_1898);
nand U2404 (N_2404,N_1909,N_1973);
nand U2405 (N_2405,N_1542,N_1872);
nand U2406 (N_2406,N_1816,N_1664);
xor U2407 (N_2407,N_1869,N_1943);
nand U2408 (N_2408,N_1913,N_1798);
nor U2409 (N_2409,N_1765,N_1517);
nor U2410 (N_2410,N_1811,N_1854);
nor U2411 (N_2411,N_1502,N_1926);
and U2412 (N_2412,N_1920,N_1941);
nand U2413 (N_2413,N_1501,N_1676);
or U2414 (N_2414,N_1887,N_1650);
xor U2415 (N_2415,N_1583,N_1688);
xor U2416 (N_2416,N_1608,N_1940);
and U2417 (N_2417,N_1663,N_1884);
and U2418 (N_2418,N_1811,N_1809);
and U2419 (N_2419,N_1926,N_1653);
or U2420 (N_2420,N_1993,N_1910);
or U2421 (N_2421,N_1766,N_1529);
nand U2422 (N_2422,N_1612,N_1557);
nor U2423 (N_2423,N_1749,N_1809);
xor U2424 (N_2424,N_1864,N_1604);
and U2425 (N_2425,N_1918,N_1724);
xor U2426 (N_2426,N_1536,N_1551);
nand U2427 (N_2427,N_1697,N_1645);
or U2428 (N_2428,N_1965,N_1617);
xnor U2429 (N_2429,N_1587,N_1681);
or U2430 (N_2430,N_1554,N_1974);
and U2431 (N_2431,N_1731,N_1694);
xnor U2432 (N_2432,N_1659,N_1996);
xnor U2433 (N_2433,N_1983,N_1586);
or U2434 (N_2434,N_1888,N_1598);
nand U2435 (N_2435,N_1899,N_1926);
nand U2436 (N_2436,N_1717,N_1606);
and U2437 (N_2437,N_1823,N_1613);
or U2438 (N_2438,N_1715,N_1630);
nor U2439 (N_2439,N_1716,N_1590);
xnor U2440 (N_2440,N_1510,N_1585);
and U2441 (N_2441,N_1693,N_1537);
or U2442 (N_2442,N_1847,N_1671);
nor U2443 (N_2443,N_1505,N_1711);
xor U2444 (N_2444,N_1572,N_1826);
nor U2445 (N_2445,N_1581,N_1833);
or U2446 (N_2446,N_1632,N_1600);
nor U2447 (N_2447,N_1748,N_1945);
or U2448 (N_2448,N_1716,N_1723);
nor U2449 (N_2449,N_1925,N_1829);
nand U2450 (N_2450,N_1848,N_1807);
or U2451 (N_2451,N_1721,N_1623);
nand U2452 (N_2452,N_1755,N_1678);
nor U2453 (N_2453,N_1640,N_1631);
or U2454 (N_2454,N_1578,N_1767);
nor U2455 (N_2455,N_1759,N_1975);
nand U2456 (N_2456,N_1655,N_1694);
and U2457 (N_2457,N_1932,N_1606);
nor U2458 (N_2458,N_1709,N_1668);
or U2459 (N_2459,N_1903,N_1700);
nor U2460 (N_2460,N_1561,N_1796);
and U2461 (N_2461,N_1703,N_1747);
and U2462 (N_2462,N_1718,N_1779);
or U2463 (N_2463,N_1981,N_1893);
nand U2464 (N_2464,N_1794,N_1998);
and U2465 (N_2465,N_1836,N_1984);
and U2466 (N_2466,N_1772,N_1797);
nor U2467 (N_2467,N_1950,N_1619);
nor U2468 (N_2468,N_1635,N_1600);
nand U2469 (N_2469,N_1900,N_1664);
nand U2470 (N_2470,N_1657,N_1739);
xor U2471 (N_2471,N_1928,N_1573);
or U2472 (N_2472,N_1510,N_1927);
xor U2473 (N_2473,N_1994,N_1584);
or U2474 (N_2474,N_1802,N_1832);
nand U2475 (N_2475,N_1789,N_1600);
or U2476 (N_2476,N_1910,N_1685);
nand U2477 (N_2477,N_1590,N_1577);
and U2478 (N_2478,N_1576,N_1563);
or U2479 (N_2479,N_1631,N_1572);
or U2480 (N_2480,N_1849,N_1529);
and U2481 (N_2481,N_1525,N_1694);
and U2482 (N_2482,N_1576,N_1599);
nor U2483 (N_2483,N_1572,N_1607);
and U2484 (N_2484,N_1684,N_1537);
nor U2485 (N_2485,N_1794,N_1512);
and U2486 (N_2486,N_1873,N_1680);
nand U2487 (N_2487,N_1764,N_1675);
nor U2488 (N_2488,N_1947,N_1670);
xor U2489 (N_2489,N_1781,N_1812);
and U2490 (N_2490,N_1934,N_1595);
nor U2491 (N_2491,N_1566,N_1993);
nand U2492 (N_2492,N_1817,N_1797);
xor U2493 (N_2493,N_1938,N_1965);
and U2494 (N_2494,N_1610,N_1554);
xnor U2495 (N_2495,N_1718,N_1513);
nand U2496 (N_2496,N_1549,N_1969);
xnor U2497 (N_2497,N_1868,N_1557);
or U2498 (N_2498,N_1571,N_1621);
or U2499 (N_2499,N_1999,N_1925);
xnor U2500 (N_2500,N_2084,N_2319);
nor U2501 (N_2501,N_2348,N_2230);
or U2502 (N_2502,N_2106,N_2269);
nor U2503 (N_2503,N_2085,N_2119);
nand U2504 (N_2504,N_2429,N_2261);
xor U2505 (N_2505,N_2360,N_2449);
nand U2506 (N_2506,N_2292,N_2015);
or U2507 (N_2507,N_2477,N_2344);
and U2508 (N_2508,N_2253,N_2001);
nor U2509 (N_2509,N_2010,N_2441);
xnor U2510 (N_2510,N_2420,N_2494);
nand U2511 (N_2511,N_2112,N_2418);
and U2512 (N_2512,N_2213,N_2342);
or U2513 (N_2513,N_2279,N_2442);
or U2514 (N_2514,N_2147,N_2021);
and U2515 (N_2515,N_2254,N_2060);
nor U2516 (N_2516,N_2366,N_2309);
nand U2517 (N_2517,N_2465,N_2390);
xnor U2518 (N_2518,N_2093,N_2271);
and U2519 (N_2519,N_2053,N_2218);
and U2520 (N_2520,N_2296,N_2411);
and U2521 (N_2521,N_2485,N_2167);
nand U2522 (N_2522,N_2463,N_2351);
nand U2523 (N_2523,N_2159,N_2208);
xnor U2524 (N_2524,N_2235,N_2490);
nand U2525 (N_2525,N_2154,N_2438);
xor U2526 (N_2526,N_2312,N_2122);
nand U2527 (N_2527,N_2150,N_2410);
xnor U2528 (N_2528,N_2155,N_2008);
nor U2529 (N_2529,N_2302,N_2231);
or U2530 (N_2530,N_2337,N_2370);
nand U2531 (N_2531,N_2019,N_2346);
and U2532 (N_2532,N_2263,N_2229);
nand U2533 (N_2533,N_2216,N_2111);
or U2534 (N_2534,N_2482,N_2041);
or U2535 (N_2535,N_2156,N_2046);
nand U2536 (N_2536,N_2475,N_2075);
and U2537 (N_2537,N_2455,N_2334);
nor U2538 (N_2538,N_2489,N_2035);
xnor U2539 (N_2539,N_2116,N_2029);
xnor U2540 (N_2540,N_2343,N_2373);
or U2541 (N_2541,N_2293,N_2368);
xnor U2542 (N_2542,N_2182,N_2070);
xor U2543 (N_2543,N_2201,N_2083);
and U2544 (N_2544,N_2120,N_2300);
nand U2545 (N_2545,N_2097,N_2059);
xnor U2546 (N_2546,N_2163,N_2139);
nand U2547 (N_2547,N_2023,N_2425);
xor U2548 (N_2548,N_2495,N_2382);
xor U2549 (N_2549,N_2138,N_2247);
and U2550 (N_2550,N_2311,N_2326);
nor U2551 (N_2551,N_2320,N_2028);
or U2552 (N_2552,N_2426,N_2087);
nand U2553 (N_2553,N_2401,N_2081);
and U2554 (N_2554,N_2499,N_2051);
or U2555 (N_2555,N_2427,N_2259);
xnor U2556 (N_2556,N_2117,N_2157);
nand U2557 (N_2557,N_2166,N_2203);
nor U2558 (N_2558,N_2004,N_2340);
nand U2559 (N_2559,N_2137,N_2228);
xnor U2560 (N_2560,N_2472,N_2409);
xnor U2561 (N_2561,N_2371,N_2386);
or U2562 (N_2562,N_2406,N_2484);
or U2563 (N_2563,N_2240,N_2092);
or U2564 (N_2564,N_2392,N_2007);
or U2565 (N_2565,N_2314,N_2473);
nand U2566 (N_2566,N_2322,N_2483);
and U2567 (N_2567,N_2445,N_2324);
nor U2568 (N_2568,N_2339,N_2058);
or U2569 (N_2569,N_2383,N_2474);
nand U2570 (N_2570,N_2408,N_2113);
xor U2571 (N_2571,N_2009,N_2428);
or U2572 (N_2572,N_2124,N_2185);
or U2573 (N_2573,N_2435,N_2416);
xor U2574 (N_2574,N_2189,N_2123);
nand U2575 (N_2575,N_2486,N_2452);
or U2576 (N_2576,N_2252,N_2195);
or U2577 (N_2577,N_2135,N_2376);
nor U2578 (N_2578,N_2275,N_2361);
nor U2579 (N_2579,N_2196,N_2205);
xnor U2580 (N_2580,N_2437,N_2413);
xor U2581 (N_2581,N_2100,N_2128);
xnor U2582 (N_2582,N_2470,N_2064);
xnor U2583 (N_2583,N_2133,N_2394);
nand U2584 (N_2584,N_2049,N_2467);
or U2585 (N_2585,N_2448,N_2170);
or U2586 (N_2586,N_2315,N_2352);
or U2587 (N_2587,N_2024,N_2013);
nand U2588 (N_2588,N_2329,N_2379);
xor U2589 (N_2589,N_2063,N_2262);
or U2590 (N_2590,N_2082,N_2105);
xor U2591 (N_2591,N_2219,N_2462);
and U2592 (N_2592,N_2375,N_2333);
nor U2593 (N_2593,N_2129,N_2266);
xor U2594 (N_2594,N_2039,N_2108);
nor U2595 (N_2595,N_2264,N_2397);
nand U2596 (N_2596,N_2493,N_2062);
or U2597 (N_2597,N_2460,N_2215);
nor U2598 (N_2598,N_2297,N_2214);
nand U2599 (N_2599,N_2236,N_2212);
xnor U2600 (N_2600,N_2384,N_2047);
and U2601 (N_2601,N_2142,N_2178);
nor U2602 (N_2602,N_2057,N_2273);
nand U2603 (N_2603,N_2464,N_2202);
and U2604 (N_2604,N_2402,N_2144);
and U2605 (N_2605,N_2140,N_2487);
xnor U2606 (N_2606,N_2480,N_2466);
and U2607 (N_2607,N_2316,N_2032);
nor U2608 (N_2608,N_2358,N_2451);
and U2609 (N_2609,N_2169,N_2220);
nand U2610 (N_2610,N_2069,N_2130);
or U2611 (N_2611,N_2476,N_2094);
xor U2612 (N_2612,N_2389,N_2206);
and U2613 (N_2613,N_2412,N_2443);
nor U2614 (N_2614,N_2439,N_2488);
xnor U2615 (N_2615,N_2318,N_2200);
or U2616 (N_2616,N_2176,N_2423);
nor U2617 (N_2617,N_2125,N_2055);
and U2618 (N_2618,N_2282,N_2497);
nand U2619 (N_2619,N_2350,N_2199);
or U2620 (N_2620,N_2241,N_2450);
nand U2621 (N_2621,N_2440,N_2298);
or U2622 (N_2622,N_2018,N_2191);
nand U2623 (N_2623,N_2098,N_2288);
and U2624 (N_2624,N_2414,N_2323);
nand U2625 (N_2625,N_2468,N_2299);
xor U2626 (N_2626,N_2034,N_2459);
xor U2627 (N_2627,N_2050,N_2492);
or U2628 (N_2628,N_2255,N_2365);
nand U2629 (N_2629,N_2305,N_2152);
nand U2630 (N_2630,N_2385,N_2148);
nor U2631 (N_2631,N_2168,N_2265);
and U2632 (N_2632,N_2251,N_2457);
nor U2633 (N_2633,N_2149,N_2095);
or U2634 (N_2634,N_2325,N_2404);
nor U2635 (N_2635,N_2221,N_2204);
nand U2636 (N_2636,N_2011,N_2104);
nor U2637 (N_2637,N_2006,N_2031);
or U2638 (N_2638,N_2446,N_2458);
nor U2639 (N_2639,N_2183,N_2380);
nor U2640 (N_2640,N_2481,N_2190);
xor U2641 (N_2641,N_2303,N_2290);
xnor U2642 (N_2642,N_2160,N_2444);
xor U2643 (N_2643,N_2349,N_2061);
or U2644 (N_2644,N_2295,N_2395);
and U2645 (N_2645,N_2321,N_2301);
nor U2646 (N_2646,N_2091,N_2284);
nand U2647 (N_2647,N_2355,N_2249);
and U2648 (N_2648,N_2327,N_2399);
and U2649 (N_2649,N_2294,N_2136);
or U2650 (N_2650,N_2089,N_2192);
nand U2651 (N_2651,N_2407,N_2403);
or U2652 (N_2652,N_2012,N_2143);
or U2653 (N_2653,N_2158,N_2153);
and U2654 (N_2654,N_2074,N_2338);
or U2655 (N_2655,N_2478,N_2076);
and U2656 (N_2656,N_2210,N_2310);
xor U2657 (N_2657,N_2405,N_2456);
nand U2658 (N_2658,N_2020,N_2030);
and U2659 (N_2659,N_2042,N_2436);
nand U2660 (N_2660,N_2036,N_2026);
xnor U2661 (N_2661,N_2079,N_2281);
nor U2662 (N_2662,N_2179,N_2134);
xnor U2663 (N_2663,N_2391,N_2080);
xnor U2664 (N_2664,N_2177,N_2222);
xnor U2665 (N_2665,N_2194,N_2033);
nor U2666 (N_2666,N_2347,N_2172);
nor U2667 (N_2667,N_2161,N_2335);
nor U2668 (N_2668,N_2396,N_2072);
nand U2669 (N_2669,N_2367,N_2419);
or U2670 (N_2670,N_2077,N_2238);
and U2671 (N_2671,N_2118,N_2260);
and U2672 (N_2672,N_2126,N_2393);
xnor U2673 (N_2673,N_2422,N_2066);
nor U2674 (N_2674,N_2398,N_2005);
nand U2675 (N_2675,N_2431,N_2223);
nand U2676 (N_2676,N_2272,N_2071);
nor U2677 (N_2677,N_2328,N_2433);
nor U2678 (N_2678,N_2043,N_2308);
xnor U2679 (N_2679,N_2496,N_2025);
or U2680 (N_2680,N_2430,N_2022);
nor U2681 (N_2681,N_2217,N_2132);
and U2682 (N_2682,N_2357,N_2421);
nor U2683 (N_2683,N_2471,N_2491);
or U2684 (N_2684,N_2432,N_2479);
or U2685 (N_2685,N_2054,N_2381);
or U2686 (N_2686,N_2234,N_2274);
xnor U2687 (N_2687,N_2103,N_2131);
nor U2688 (N_2688,N_2186,N_2286);
nor U2689 (N_2689,N_2378,N_2174);
and U2690 (N_2690,N_2447,N_2267);
or U2691 (N_2691,N_2387,N_2362);
or U2692 (N_2692,N_2115,N_2304);
or U2693 (N_2693,N_2233,N_2313);
xnor U2694 (N_2694,N_2285,N_2354);
and U2695 (N_2695,N_2250,N_2345);
or U2696 (N_2696,N_2246,N_2027);
nand U2697 (N_2697,N_2096,N_2173);
xor U2698 (N_2698,N_2068,N_2151);
nand U2699 (N_2699,N_2341,N_2145);
xor U2700 (N_2700,N_2014,N_2270);
nand U2701 (N_2701,N_2044,N_2017);
xor U2702 (N_2702,N_2336,N_2127);
xnor U2703 (N_2703,N_2002,N_2289);
and U2704 (N_2704,N_2003,N_2107);
or U2705 (N_2705,N_2184,N_2086);
nand U2706 (N_2706,N_2283,N_2193);
nand U2707 (N_2707,N_2198,N_2278);
and U2708 (N_2708,N_2287,N_2141);
xor U2709 (N_2709,N_2171,N_2078);
and U2710 (N_2710,N_2038,N_2461);
or U2711 (N_2711,N_2369,N_2257);
or U2712 (N_2712,N_2258,N_2317);
nand U2713 (N_2713,N_2016,N_2239);
xnor U2714 (N_2714,N_2245,N_2237);
and U2715 (N_2715,N_2048,N_2052);
xnor U2716 (N_2716,N_2164,N_2065);
and U2717 (N_2717,N_2101,N_2146);
or U2718 (N_2718,N_2330,N_2331);
or U2719 (N_2719,N_2498,N_2332);
and U2720 (N_2720,N_2291,N_2377);
or U2721 (N_2721,N_2180,N_2102);
xor U2722 (N_2722,N_2248,N_2280);
and U2723 (N_2723,N_2037,N_2224);
or U2724 (N_2724,N_2090,N_2400);
nand U2725 (N_2725,N_2187,N_2109);
nand U2726 (N_2726,N_2256,N_2040);
or U2727 (N_2727,N_2088,N_2073);
and U2728 (N_2728,N_2211,N_2188);
and U2729 (N_2729,N_2469,N_2276);
nor U2730 (N_2730,N_2306,N_2067);
nand U2731 (N_2731,N_2165,N_2417);
or U2732 (N_2732,N_2353,N_2374);
xnor U2733 (N_2733,N_2232,N_2356);
xor U2734 (N_2734,N_2197,N_2207);
nand U2735 (N_2735,N_2000,N_2364);
and U2736 (N_2736,N_2359,N_2056);
nor U2737 (N_2737,N_2243,N_2045);
xor U2738 (N_2738,N_2114,N_2209);
xor U2739 (N_2739,N_2226,N_2162);
nor U2740 (N_2740,N_2099,N_2227);
nand U2741 (N_2741,N_2121,N_2242);
and U2742 (N_2742,N_2277,N_2363);
or U2743 (N_2743,N_2415,N_2175);
or U2744 (N_2744,N_2268,N_2454);
nand U2745 (N_2745,N_2181,N_2225);
and U2746 (N_2746,N_2453,N_2244);
nor U2747 (N_2747,N_2388,N_2424);
or U2748 (N_2748,N_2110,N_2372);
and U2749 (N_2749,N_2434,N_2307);
xnor U2750 (N_2750,N_2068,N_2134);
nand U2751 (N_2751,N_2456,N_2374);
and U2752 (N_2752,N_2007,N_2094);
nand U2753 (N_2753,N_2233,N_2090);
xnor U2754 (N_2754,N_2401,N_2133);
nor U2755 (N_2755,N_2421,N_2040);
nand U2756 (N_2756,N_2174,N_2484);
and U2757 (N_2757,N_2411,N_2079);
nand U2758 (N_2758,N_2055,N_2204);
or U2759 (N_2759,N_2113,N_2317);
nand U2760 (N_2760,N_2067,N_2115);
or U2761 (N_2761,N_2291,N_2197);
nand U2762 (N_2762,N_2085,N_2397);
nand U2763 (N_2763,N_2100,N_2230);
or U2764 (N_2764,N_2202,N_2497);
nor U2765 (N_2765,N_2163,N_2084);
nand U2766 (N_2766,N_2129,N_2383);
nor U2767 (N_2767,N_2021,N_2447);
nor U2768 (N_2768,N_2461,N_2094);
or U2769 (N_2769,N_2403,N_2269);
and U2770 (N_2770,N_2086,N_2347);
xor U2771 (N_2771,N_2038,N_2066);
nand U2772 (N_2772,N_2168,N_2474);
xor U2773 (N_2773,N_2315,N_2094);
or U2774 (N_2774,N_2157,N_2449);
nand U2775 (N_2775,N_2436,N_2118);
xnor U2776 (N_2776,N_2431,N_2308);
nand U2777 (N_2777,N_2293,N_2404);
xor U2778 (N_2778,N_2322,N_2370);
nand U2779 (N_2779,N_2065,N_2436);
xnor U2780 (N_2780,N_2353,N_2318);
xnor U2781 (N_2781,N_2302,N_2252);
xor U2782 (N_2782,N_2020,N_2161);
nand U2783 (N_2783,N_2241,N_2250);
nand U2784 (N_2784,N_2066,N_2394);
and U2785 (N_2785,N_2323,N_2306);
nor U2786 (N_2786,N_2214,N_2262);
xor U2787 (N_2787,N_2044,N_2447);
and U2788 (N_2788,N_2438,N_2486);
and U2789 (N_2789,N_2164,N_2324);
xnor U2790 (N_2790,N_2328,N_2287);
xor U2791 (N_2791,N_2129,N_2271);
nand U2792 (N_2792,N_2103,N_2149);
nor U2793 (N_2793,N_2022,N_2201);
nor U2794 (N_2794,N_2305,N_2296);
or U2795 (N_2795,N_2227,N_2326);
nor U2796 (N_2796,N_2115,N_2460);
and U2797 (N_2797,N_2331,N_2364);
and U2798 (N_2798,N_2194,N_2370);
xor U2799 (N_2799,N_2091,N_2082);
xnor U2800 (N_2800,N_2342,N_2256);
xor U2801 (N_2801,N_2319,N_2433);
xor U2802 (N_2802,N_2161,N_2155);
and U2803 (N_2803,N_2084,N_2447);
nor U2804 (N_2804,N_2339,N_2280);
nand U2805 (N_2805,N_2395,N_2289);
nand U2806 (N_2806,N_2070,N_2422);
and U2807 (N_2807,N_2203,N_2407);
nand U2808 (N_2808,N_2291,N_2261);
nand U2809 (N_2809,N_2265,N_2477);
and U2810 (N_2810,N_2351,N_2119);
nand U2811 (N_2811,N_2380,N_2240);
nor U2812 (N_2812,N_2143,N_2016);
nand U2813 (N_2813,N_2120,N_2206);
nand U2814 (N_2814,N_2239,N_2316);
nor U2815 (N_2815,N_2200,N_2237);
or U2816 (N_2816,N_2472,N_2297);
and U2817 (N_2817,N_2245,N_2044);
nand U2818 (N_2818,N_2373,N_2271);
nand U2819 (N_2819,N_2072,N_2134);
and U2820 (N_2820,N_2153,N_2258);
nand U2821 (N_2821,N_2237,N_2124);
nand U2822 (N_2822,N_2184,N_2023);
and U2823 (N_2823,N_2067,N_2310);
and U2824 (N_2824,N_2241,N_2110);
xnor U2825 (N_2825,N_2170,N_2013);
nor U2826 (N_2826,N_2350,N_2191);
or U2827 (N_2827,N_2085,N_2250);
nand U2828 (N_2828,N_2286,N_2398);
or U2829 (N_2829,N_2033,N_2299);
nand U2830 (N_2830,N_2451,N_2364);
xnor U2831 (N_2831,N_2315,N_2019);
nor U2832 (N_2832,N_2379,N_2453);
or U2833 (N_2833,N_2436,N_2426);
nand U2834 (N_2834,N_2122,N_2465);
xnor U2835 (N_2835,N_2445,N_2476);
or U2836 (N_2836,N_2023,N_2442);
nor U2837 (N_2837,N_2275,N_2116);
nor U2838 (N_2838,N_2379,N_2484);
and U2839 (N_2839,N_2221,N_2167);
nor U2840 (N_2840,N_2118,N_2475);
or U2841 (N_2841,N_2266,N_2451);
and U2842 (N_2842,N_2282,N_2103);
nand U2843 (N_2843,N_2269,N_2194);
or U2844 (N_2844,N_2418,N_2317);
xor U2845 (N_2845,N_2170,N_2436);
nor U2846 (N_2846,N_2169,N_2306);
xnor U2847 (N_2847,N_2439,N_2081);
and U2848 (N_2848,N_2414,N_2320);
nand U2849 (N_2849,N_2262,N_2109);
xor U2850 (N_2850,N_2127,N_2129);
or U2851 (N_2851,N_2135,N_2081);
nor U2852 (N_2852,N_2332,N_2446);
and U2853 (N_2853,N_2388,N_2100);
and U2854 (N_2854,N_2106,N_2031);
nand U2855 (N_2855,N_2296,N_2459);
nor U2856 (N_2856,N_2498,N_2380);
nand U2857 (N_2857,N_2005,N_2143);
nor U2858 (N_2858,N_2178,N_2230);
nand U2859 (N_2859,N_2372,N_2191);
and U2860 (N_2860,N_2015,N_2336);
or U2861 (N_2861,N_2133,N_2247);
xnor U2862 (N_2862,N_2065,N_2361);
nor U2863 (N_2863,N_2259,N_2207);
and U2864 (N_2864,N_2431,N_2028);
or U2865 (N_2865,N_2286,N_2281);
and U2866 (N_2866,N_2285,N_2061);
and U2867 (N_2867,N_2050,N_2188);
xnor U2868 (N_2868,N_2199,N_2454);
nor U2869 (N_2869,N_2305,N_2229);
or U2870 (N_2870,N_2208,N_2494);
xnor U2871 (N_2871,N_2388,N_2455);
or U2872 (N_2872,N_2016,N_2459);
nor U2873 (N_2873,N_2185,N_2048);
or U2874 (N_2874,N_2179,N_2180);
nand U2875 (N_2875,N_2070,N_2191);
nor U2876 (N_2876,N_2392,N_2055);
nand U2877 (N_2877,N_2150,N_2395);
nand U2878 (N_2878,N_2015,N_2374);
or U2879 (N_2879,N_2014,N_2141);
nand U2880 (N_2880,N_2486,N_2091);
and U2881 (N_2881,N_2052,N_2129);
nor U2882 (N_2882,N_2435,N_2399);
nand U2883 (N_2883,N_2197,N_2031);
nor U2884 (N_2884,N_2157,N_2247);
or U2885 (N_2885,N_2022,N_2398);
xor U2886 (N_2886,N_2294,N_2112);
or U2887 (N_2887,N_2359,N_2031);
or U2888 (N_2888,N_2366,N_2487);
and U2889 (N_2889,N_2324,N_2318);
or U2890 (N_2890,N_2439,N_2401);
xor U2891 (N_2891,N_2264,N_2346);
or U2892 (N_2892,N_2195,N_2181);
nor U2893 (N_2893,N_2224,N_2245);
or U2894 (N_2894,N_2199,N_2297);
and U2895 (N_2895,N_2443,N_2345);
nand U2896 (N_2896,N_2497,N_2268);
nor U2897 (N_2897,N_2451,N_2159);
and U2898 (N_2898,N_2246,N_2410);
or U2899 (N_2899,N_2068,N_2216);
xnor U2900 (N_2900,N_2052,N_2261);
nor U2901 (N_2901,N_2302,N_2374);
xor U2902 (N_2902,N_2325,N_2407);
and U2903 (N_2903,N_2496,N_2074);
xor U2904 (N_2904,N_2112,N_2278);
xnor U2905 (N_2905,N_2475,N_2015);
nor U2906 (N_2906,N_2482,N_2132);
xor U2907 (N_2907,N_2007,N_2059);
or U2908 (N_2908,N_2282,N_2384);
nand U2909 (N_2909,N_2431,N_2253);
and U2910 (N_2910,N_2309,N_2097);
xnor U2911 (N_2911,N_2477,N_2112);
and U2912 (N_2912,N_2440,N_2157);
nor U2913 (N_2913,N_2491,N_2126);
xnor U2914 (N_2914,N_2085,N_2404);
and U2915 (N_2915,N_2455,N_2055);
and U2916 (N_2916,N_2374,N_2117);
nand U2917 (N_2917,N_2020,N_2134);
nand U2918 (N_2918,N_2266,N_2112);
and U2919 (N_2919,N_2432,N_2203);
xor U2920 (N_2920,N_2327,N_2324);
and U2921 (N_2921,N_2253,N_2132);
nor U2922 (N_2922,N_2101,N_2244);
nor U2923 (N_2923,N_2046,N_2459);
nand U2924 (N_2924,N_2070,N_2281);
nor U2925 (N_2925,N_2477,N_2187);
and U2926 (N_2926,N_2328,N_2067);
and U2927 (N_2927,N_2252,N_2303);
or U2928 (N_2928,N_2296,N_2493);
or U2929 (N_2929,N_2167,N_2148);
and U2930 (N_2930,N_2292,N_2183);
nor U2931 (N_2931,N_2190,N_2312);
nor U2932 (N_2932,N_2149,N_2138);
nand U2933 (N_2933,N_2264,N_2471);
and U2934 (N_2934,N_2162,N_2155);
or U2935 (N_2935,N_2012,N_2254);
nand U2936 (N_2936,N_2461,N_2413);
xnor U2937 (N_2937,N_2260,N_2345);
or U2938 (N_2938,N_2490,N_2459);
nor U2939 (N_2939,N_2010,N_2238);
nand U2940 (N_2940,N_2063,N_2191);
or U2941 (N_2941,N_2184,N_2405);
and U2942 (N_2942,N_2116,N_2009);
nor U2943 (N_2943,N_2093,N_2440);
nand U2944 (N_2944,N_2215,N_2254);
or U2945 (N_2945,N_2404,N_2115);
or U2946 (N_2946,N_2246,N_2273);
or U2947 (N_2947,N_2200,N_2397);
and U2948 (N_2948,N_2486,N_2015);
nand U2949 (N_2949,N_2351,N_2291);
nand U2950 (N_2950,N_2210,N_2112);
and U2951 (N_2951,N_2037,N_2128);
xnor U2952 (N_2952,N_2290,N_2420);
or U2953 (N_2953,N_2031,N_2014);
nor U2954 (N_2954,N_2167,N_2375);
nor U2955 (N_2955,N_2184,N_2149);
xnor U2956 (N_2956,N_2318,N_2335);
and U2957 (N_2957,N_2137,N_2161);
and U2958 (N_2958,N_2317,N_2195);
nand U2959 (N_2959,N_2413,N_2089);
nor U2960 (N_2960,N_2461,N_2098);
nor U2961 (N_2961,N_2317,N_2260);
xor U2962 (N_2962,N_2492,N_2399);
nor U2963 (N_2963,N_2031,N_2079);
nor U2964 (N_2964,N_2417,N_2457);
nand U2965 (N_2965,N_2302,N_2472);
xor U2966 (N_2966,N_2112,N_2111);
or U2967 (N_2967,N_2008,N_2252);
and U2968 (N_2968,N_2340,N_2245);
nor U2969 (N_2969,N_2324,N_2158);
nor U2970 (N_2970,N_2094,N_2377);
nand U2971 (N_2971,N_2030,N_2222);
or U2972 (N_2972,N_2385,N_2040);
xor U2973 (N_2973,N_2170,N_2260);
or U2974 (N_2974,N_2008,N_2403);
nand U2975 (N_2975,N_2042,N_2325);
or U2976 (N_2976,N_2472,N_2355);
and U2977 (N_2977,N_2376,N_2437);
nand U2978 (N_2978,N_2171,N_2239);
and U2979 (N_2979,N_2405,N_2057);
and U2980 (N_2980,N_2414,N_2039);
and U2981 (N_2981,N_2477,N_2402);
and U2982 (N_2982,N_2256,N_2070);
and U2983 (N_2983,N_2093,N_2340);
or U2984 (N_2984,N_2258,N_2143);
xor U2985 (N_2985,N_2040,N_2139);
or U2986 (N_2986,N_2200,N_2166);
nand U2987 (N_2987,N_2440,N_2108);
and U2988 (N_2988,N_2062,N_2010);
or U2989 (N_2989,N_2338,N_2424);
and U2990 (N_2990,N_2040,N_2076);
or U2991 (N_2991,N_2496,N_2225);
and U2992 (N_2992,N_2271,N_2019);
nor U2993 (N_2993,N_2018,N_2249);
xnor U2994 (N_2994,N_2034,N_2444);
nand U2995 (N_2995,N_2047,N_2097);
or U2996 (N_2996,N_2195,N_2273);
nand U2997 (N_2997,N_2271,N_2127);
xnor U2998 (N_2998,N_2121,N_2199);
xor U2999 (N_2999,N_2285,N_2391);
nand U3000 (N_3000,N_2744,N_2876);
or U3001 (N_3001,N_2762,N_2793);
xor U3002 (N_3002,N_2860,N_2677);
or U3003 (N_3003,N_2808,N_2656);
and U3004 (N_3004,N_2942,N_2739);
xor U3005 (N_3005,N_2642,N_2814);
nor U3006 (N_3006,N_2584,N_2756);
or U3007 (N_3007,N_2888,N_2967);
nand U3008 (N_3008,N_2825,N_2631);
nand U3009 (N_3009,N_2775,N_2786);
or U3010 (N_3010,N_2985,N_2897);
nand U3011 (N_3011,N_2805,N_2921);
or U3012 (N_3012,N_2898,N_2521);
nand U3013 (N_3013,N_2634,N_2502);
or U3014 (N_3014,N_2993,N_2659);
and U3015 (N_3015,N_2872,N_2648);
and U3016 (N_3016,N_2563,N_2980);
nor U3017 (N_3017,N_2698,N_2787);
xor U3018 (N_3018,N_2530,N_2614);
xnor U3019 (N_3019,N_2730,N_2666);
and U3020 (N_3020,N_2514,N_2886);
nor U3021 (N_3021,N_2607,N_2588);
or U3022 (N_3022,N_2678,N_2819);
nor U3023 (N_3023,N_2834,N_2560);
xor U3024 (N_3024,N_2599,N_2968);
or U3025 (N_3025,N_2753,N_2806);
or U3026 (N_3026,N_2529,N_2957);
xor U3027 (N_3027,N_2875,N_2958);
nand U3028 (N_3028,N_2881,N_2571);
and U3029 (N_3029,N_2894,N_2721);
nand U3030 (N_3030,N_2674,N_2517);
and U3031 (N_3031,N_2840,N_2541);
nand U3032 (N_3032,N_2619,N_2785);
nor U3033 (N_3033,N_2914,N_2690);
and U3034 (N_3034,N_2685,N_2777);
nand U3035 (N_3035,N_2551,N_2526);
and U3036 (N_3036,N_2791,N_2542);
or U3037 (N_3037,N_2846,N_2663);
or U3038 (N_3038,N_2751,N_2635);
or U3039 (N_3039,N_2692,N_2844);
or U3040 (N_3040,N_2593,N_2760);
and U3041 (N_3041,N_2861,N_2802);
xnor U3042 (N_3042,N_2525,N_2550);
and U3043 (N_3043,N_2912,N_2729);
xor U3044 (N_3044,N_2585,N_2901);
or U3045 (N_3045,N_2507,N_2658);
nor U3046 (N_3046,N_2591,N_2889);
nor U3047 (N_3047,N_2969,N_2625);
nand U3048 (N_3048,N_2766,N_2655);
or U3049 (N_3049,N_2577,N_2649);
xor U3050 (N_3050,N_2722,N_2850);
xor U3051 (N_3051,N_2854,N_2772);
and U3052 (N_3052,N_2885,N_2682);
nor U3053 (N_3053,N_2691,N_2500);
or U3054 (N_3054,N_2841,N_2837);
xor U3055 (N_3055,N_2963,N_2546);
or U3056 (N_3056,N_2800,N_2624);
xor U3057 (N_3057,N_2725,N_2554);
and U3058 (N_3058,N_2618,N_2549);
nor U3059 (N_3059,N_2974,N_2538);
or U3060 (N_3060,N_2600,N_2911);
and U3061 (N_3061,N_2829,N_2810);
or U3062 (N_3062,N_2695,N_2984);
nand U3063 (N_3063,N_2966,N_2557);
or U3064 (N_3064,N_2741,N_2660);
xnor U3065 (N_3065,N_2759,N_2731);
or U3066 (N_3066,N_2848,N_2509);
and U3067 (N_3067,N_2713,N_2539);
nor U3068 (N_3068,N_2855,N_2617);
nand U3069 (N_3069,N_2555,N_2795);
and U3070 (N_3070,N_2605,N_2693);
or U3071 (N_3071,N_2516,N_2629);
and U3072 (N_3072,N_2831,N_2804);
and U3073 (N_3073,N_2639,N_2896);
and U3074 (N_3074,N_2638,N_2643);
nand U3075 (N_3075,N_2944,N_2827);
or U3076 (N_3076,N_2824,N_2511);
and U3077 (N_3077,N_2781,N_2803);
or U3078 (N_3078,N_2922,N_2671);
nand U3079 (N_3079,N_2651,N_2975);
xor U3080 (N_3080,N_2564,N_2681);
nand U3081 (N_3081,N_2851,N_2765);
or U3082 (N_3082,N_2790,N_2990);
and U3083 (N_3083,N_2612,N_2627);
or U3084 (N_3084,N_2843,N_2964);
xnor U3085 (N_3085,N_2512,N_2580);
nand U3086 (N_3086,N_2689,N_2783);
nand U3087 (N_3087,N_2566,N_2891);
xnor U3088 (N_3088,N_2796,N_2794);
xor U3089 (N_3089,N_2826,N_2675);
or U3090 (N_3090,N_2702,N_2913);
xnor U3091 (N_3091,N_2799,N_2879);
nand U3092 (N_3092,N_2972,N_2609);
nor U3093 (N_3093,N_2815,N_2915);
and U3094 (N_3094,N_2933,N_2833);
xor U3095 (N_3095,N_2616,N_2534);
nor U3096 (N_3096,N_2955,N_2823);
xor U3097 (N_3097,N_2628,N_2548);
nand U3098 (N_3098,N_2950,N_2845);
xor U3099 (N_3099,N_2665,N_2903);
nand U3100 (N_3100,N_2757,N_2746);
nand U3101 (N_3101,N_2636,N_2576);
and U3102 (N_3102,N_2701,N_2565);
or U3103 (N_3103,N_2962,N_2773);
nor U3104 (N_3104,N_2910,N_2847);
nor U3105 (N_3105,N_2904,N_2749);
xor U3106 (N_3106,N_2531,N_2884);
or U3107 (N_3107,N_2608,N_2996);
or U3108 (N_3108,N_2709,N_2988);
xor U3109 (N_3109,N_2707,N_2735);
xor U3110 (N_3110,N_2719,N_2532);
nor U3111 (N_3111,N_2991,N_2740);
xor U3112 (N_3112,N_2953,N_2982);
nor U3113 (N_3113,N_2943,N_2732);
xor U3114 (N_3114,N_2570,N_2973);
nand U3115 (N_3115,N_2644,N_2664);
nand U3116 (N_3116,N_2873,N_2925);
nor U3117 (N_3117,N_2956,N_2870);
and U3118 (N_3118,N_2838,N_2971);
and U3119 (N_3119,N_2835,N_2755);
or U3120 (N_3120,N_2641,N_2528);
or U3121 (N_3121,N_2750,N_2820);
nand U3122 (N_3122,N_2866,N_2553);
nand U3123 (N_3123,N_2779,N_2633);
nor U3124 (N_3124,N_2706,N_2523);
or U3125 (N_3125,N_2776,N_2640);
or U3126 (N_3126,N_2997,N_2763);
xor U3127 (N_3127,N_2717,N_2899);
xor U3128 (N_3128,N_2579,N_2994);
and U3129 (N_3129,N_2868,N_2874);
and U3130 (N_3130,N_2645,N_2699);
nor U3131 (N_3131,N_2935,N_2508);
and U3132 (N_3132,N_2998,N_2864);
xnor U3133 (N_3133,N_2780,N_2734);
or U3134 (N_3134,N_2515,N_2959);
nor U3135 (N_3135,N_2927,N_2518);
nand U3136 (N_3136,N_2992,N_2657);
nand U3137 (N_3137,N_2989,N_2726);
nand U3138 (N_3138,N_2856,N_2813);
and U3139 (N_3139,N_2503,N_2597);
and U3140 (N_3140,N_2907,N_2924);
or U3141 (N_3141,N_2880,N_2667);
nand U3142 (N_3142,N_2951,N_2737);
xnor U3143 (N_3143,N_2945,N_2598);
nor U3144 (N_3144,N_2604,N_2669);
and U3145 (N_3145,N_2696,N_2801);
and U3146 (N_3146,N_2582,N_2917);
nor U3147 (N_3147,N_2905,N_2939);
nor U3148 (N_3148,N_2710,N_2694);
nor U3149 (N_3149,N_2540,N_2736);
xor U3150 (N_3150,N_2738,N_2575);
nand U3151 (N_3151,N_2987,N_2620);
and U3152 (N_3152,N_2983,N_2680);
nand U3153 (N_3153,N_2932,N_2887);
and U3154 (N_3154,N_2583,N_2784);
xor U3155 (N_3155,N_2742,N_2811);
nor U3156 (N_3156,N_2919,N_2697);
or U3157 (N_3157,N_2857,N_2970);
nand U3158 (N_3158,N_2764,N_2906);
xnor U3159 (N_3159,N_2720,N_2832);
or U3160 (N_3160,N_2979,N_2807);
and U3161 (N_3161,N_2714,N_2798);
or U3162 (N_3162,N_2895,N_2908);
nand U3163 (N_3163,N_2504,N_2818);
xor U3164 (N_3164,N_2572,N_2778);
or U3165 (N_3165,N_2774,N_2587);
xnor U3166 (N_3166,N_2890,N_2916);
nand U3167 (N_3167,N_2849,N_2812);
and U3168 (N_3168,N_2859,N_2684);
xor U3169 (N_3169,N_2797,N_2603);
and U3170 (N_3170,N_2654,N_2703);
nor U3171 (N_3171,N_2952,N_2606);
or U3172 (N_3172,N_2688,N_2590);
or U3173 (N_3173,N_2977,N_2594);
nand U3174 (N_3174,N_2770,N_2830);
xnor U3175 (N_3175,N_2920,N_2533);
or U3176 (N_3176,N_2892,N_2562);
nand U3177 (N_3177,N_2581,N_2676);
nor U3178 (N_3178,N_2623,N_2986);
nor U3179 (N_3179,N_2862,N_2621);
nor U3180 (N_3180,N_2747,N_2661);
nor U3181 (N_3181,N_2728,N_2652);
and U3182 (N_3182,N_2981,N_2976);
and U3183 (N_3183,N_2946,N_2723);
and U3184 (N_3184,N_2941,N_2556);
or U3185 (N_3185,N_2936,N_2999);
and U3186 (N_3186,N_2960,N_2543);
xnor U3187 (N_3187,N_2817,N_2978);
or U3188 (N_3188,N_2668,N_2615);
or U3189 (N_3189,N_2711,N_2558);
nand U3190 (N_3190,N_2883,N_2506);
and U3191 (N_3191,N_2519,N_2877);
xor U3192 (N_3192,N_2573,N_2611);
xor U3193 (N_3193,N_2535,N_2524);
nand U3194 (N_3194,N_2718,N_2574);
nor U3195 (N_3195,N_2505,N_2909);
nor U3196 (N_3196,N_2949,N_2561);
and U3197 (N_3197,N_2947,N_2782);
or U3198 (N_3198,N_2601,N_2995);
xor U3199 (N_3199,N_2547,N_2761);
and U3200 (N_3200,N_2768,N_2544);
nand U3201 (N_3201,N_2863,N_2653);
or U3202 (N_3202,N_2926,N_2632);
nor U3203 (N_3203,N_2748,N_2792);
nor U3204 (N_3204,N_2940,N_2602);
and U3205 (N_3205,N_2771,N_2716);
xnor U3206 (N_3206,N_2626,N_2865);
nor U3207 (N_3207,N_2672,N_2867);
nor U3208 (N_3208,N_2769,N_2501);
xor U3209 (N_3209,N_2552,N_2630);
or U3210 (N_3210,N_2961,N_2536);
xor U3211 (N_3211,N_2537,N_2586);
or U3212 (N_3212,N_2646,N_2842);
or U3213 (N_3213,N_2828,N_2900);
nor U3214 (N_3214,N_2954,N_2923);
xor U3215 (N_3215,N_2705,N_2858);
nor U3216 (N_3216,N_2568,N_2758);
or U3217 (N_3217,N_2679,N_2520);
nand U3218 (N_3218,N_2902,N_2948);
xnor U3219 (N_3219,N_2893,N_2622);
nand U3220 (N_3220,N_2704,N_2662);
or U3221 (N_3221,N_2589,N_2569);
xnor U3222 (N_3222,N_2715,N_2821);
or U3223 (N_3223,N_2686,N_2647);
nor U3224 (N_3224,N_2712,N_2578);
nor U3225 (N_3225,N_2788,N_2727);
or U3226 (N_3226,N_2613,N_2595);
nand U3227 (N_3227,N_2610,N_2650);
nor U3228 (N_3228,N_2918,N_2687);
nand U3229 (N_3229,N_2700,N_2839);
or U3230 (N_3230,N_2670,N_2878);
nand U3231 (N_3231,N_2527,N_2708);
nor U3232 (N_3232,N_2567,N_2637);
xor U3233 (N_3233,N_2596,N_2931);
xnor U3234 (N_3234,N_2683,N_2928);
nor U3235 (N_3235,N_2673,N_2929);
nand U3236 (N_3236,N_2522,N_2816);
nor U3237 (N_3237,N_2513,N_2853);
or U3238 (N_3238,N_2930,N_2745);
nand U3239 (N_3239,N_2965,N_2822);
and U3240 (N_3240,N_2559,N_2869);
xnor U3241 (N_3241,N_2743,N_2767);
nor U3242 (N_3242,N_2510,N_2724);
xnor U3243 (N_3243,N_2852,N_2871);
nor U3244 (N_3244,N_2752,N_2733);
and U3245 (N_3245,N_2592,N_2754);
or U3246 (N_3246,N_2934,N_2937);
nor U3247 (N_3247,N_2836,N_2789);
xnor U3248 (N_3248,N_2938,N_2545);
nand U3249 (N_3249,N_2882,N_2809);
or U3250 (N_3250,N_2624,N_2834);
nor U3251 (N_3251,N_2868,N_2809);
and U3252 (N_3252,N_2708,N_2694);
xor U3253 (N_3253,N_2660,N_2896);
nand U3254 (N_3254,N_2979,N_2512);
or U3255 (N_3255,N_2512,N_2528);
and U3256 (N_3256,N_2716,N_2967);
nand U3257 (N_3257,N_2802,N_2966);
and U3258 (N_3258,N_2868,N_2817);
nor U3259 (N_3259,N_2809,N_2952);
nor U3260 (N_3260,N_2636,N_2778);
nor U3261 (N_3261,N_2644,N_2657);
nand U3262 (N_3262,N_2930,N_2681);
xor U3263 (N_3263,N_2738,N_2658);
and U3264 (N_3264,N_2748,N_2739);
or U3265 (N_3265,N_2685,N_2619);
or U3266 (N_3266,N_2882,N_2780);
xnor U3267 (N_3267,N_2706,N_2722);
or U3268 (N_3268,N_2534,N_2903);
and U3269 (N_3269,N_2643,N_2585);
nand U3270 (N_3270,N_2949,N_2905);
or U3271 (N_3271,N_2535,N_2703);
or U3272 (N_3272,N_2793,N_2833);
or U3273 (N_3273,N_2773,N_2826);
nand U3274 (N_3274,N_2856,N_2966);
or U3275 (N_3275,N_2932,N_2527);
nand U3276 (N_3276,N_2533,N_2863);
nor U3277 (N_3277,N_2822,N_2806);
or U3278 (N_3278,N_2739,N_2905);
nand U3279 (N_3279,N_2803,N_2830);
and U3280 (N_3280,N_2994,N_2640);
xnor U3281 (N_3281,N_2511,N_2979);
and U3282 (N_3282,N_2790,N_2612);
and U3283 (N_3283,N_2887,N_2609);
xnor U3284 (N_3284,N_2993,N_2700);
and U3285 (N_3285,N_2902,N_2716);
nor U3286 (N_3286,N_2886,N_2680);
nand U3287 (N_3287,N_2700,N_2546);
or U3288 (N_3288,N_2844,N_2872);
xor U3289 (N_3289,N_2853,N_2980);
nor U3290 (N_3290,N_2973,N_2783);
nand U3291 (N_3291,N_2992,N_2576);
xor U3292 (N_3292,N_2902,N_2923);
or U3293 (N_3293,N_2917,N_2762);
nor U3294 (N_3294,N_2962,N_2898);
nor U3295 (N_3295,N_2964,N_2991);
xnor U3296 (N_3296,N_2575,N_2756);
or U3297 (N_3297,N_2770,N_2680);
or U3298 (N_3298,N_2833,N_2874);
nor U3299 (N_3299,N_2883,N_2561);
or U3300 (N_3300,N_2635,N_2890);
nand U3301 (N_3301,N_2569,N_2594);
nor U3302 (N_3302,N_2732,N_2754);
nor U3303 (N_3303,N_2637,N_2612);
nor U3304 (N_3304,N_2524,N_2771);
nor U3305 (N_3305,N_2755,N_2700);
and U3306 (N_3306,N_2903,N_2716);
or U3307 (N_3307,N_2978,N_2931);
and U3308 (N_3308,N_2514,N_2826);
xor U3309 (N_3309,N_2528,N_2670);
nor U3310 (N_3310,N_2801,N_2535);
nor U3311 (N_3311,N_2709,N_2875);
nand U3312 (N_3312,N_2858,N_2747);
or U3313 (N_3313,N_2933,N_2684);
or U3314 (N_3314,N_2932,N_2640);
nand U3315 (N_3315,N_2601,N_2959);
nand U3316 (N_3316,N_2971,N_2973);
xnor U3317 (N_3317,N_2828,N_2844);
and U3318 (N_3318,N_2842,N_2882);
or U3319 (N_3319,N_2817,N_2666);
and U3320 (N_3320,N_2900,N_2873);
xor U3321 (N_3321,N_2887,N_2668);
and U3322 (N_3322,N_2893,N_2600);
and U3323 (N_3323,N_2673,N_2969);
or U3324 (N_3324,N_2705,N_2677);
nand U3325 (N_3325,N_2602,N_2900);
or U3326 (N_3326,N_2952,N_2689);
xnor U3327 (N_3327,N_2875,N_2823);
or U3328 (N_3328,N_2935,N_2620);
nor U3329 (N_3329,N_2834,N_2554);
and U3330 (N_3330,N_2978,N_2805);
xor U3331 (N_3331,N_2734,N_2865);
or U3332 (N_3332,N_2851,N_2930);
nor U3333 (N_3333,N_2948,N_2782);
and U3334 (N_3334,N_2558,N_2869);
nand U3335 (N_3335,N_2540,N_2871);
and U3336 (N_3336,N_2860,N_2699);
nor U3337 (N_3337,N_2807,N_2572);
nand U3338 (N_3338,N_2537,N_2720);
nor U3339 (N_3339,N_2795,N_2748);
nor U3340 (N_3340,N_2745,N_2843);
and U3341 (N_3341,N_2654,N_2972);
nand U3342 (N_3342,N_2616,N_2560);
nor U3343 (N_3343,N_2734,N_2500);
or U3344 (N_3344,N_2962,N_2567);
xnor U3345 (N_3345,N_2611,N_2522);
nor U3346 (N_3346,N_2642,N_2682);
nor U3347 (N_3347,N_2503,N_2715);
nor U3348 (N_3348,N_2849,N_2872);
nor U3349 (N_3349,N_2741,N_2597);
and U3350 (N_3350,N_2964,N_2819);
nand U3351 (N_3351,N_2822,N_2989);
or U3352 (N_3352,N_2994,N_2938);
and U3353 (N_3353,N_2966,N_2884);
nor U3354 (N_3354,N_2984,N_2718);
and U3355 (N_3355,N_2731,N_2853);
nor U3356 (N_3356,N_2744,N_2723);
nand U3357 (N_3357,N_2818,N_2638);
nand U3358 (N_3358,N_2726,N_2809);
xor U3359 (N_3359,N_2893,N_2884);
xnor U3360 (N_3360,N_2676,N_2910);
or U3361 (N_3361,N_2628,N_2930);
and U3362 (N_3362,N_2907,N_2733);
xnor U3363 (N_3363,N_2990,N_2554);
xor U3364 (N_3364,N_2719,N_2789);
or U3365 (N_3365,N_2522,N_2748);
nor U3366 (N_3366,N_2794,N_2831);
and U3367 (N_3367,N_2636,N_2845);
xor U3368 (N_3368,N_2573,N_2688);
nand U3369 (N_3369,N_2735,N_2731);
nor U3370 (N_3370,N_2916,N_2580);
nor U3371 (N_3371,N_2664,N_2508);
xnor U3372 (N_3372,N_2975,N_2771);
nor U3373 (N_3373,N_2759,N_2552);
nand U3374 (N_3374,N_2748,N_2980);
nand U3375 (N_3375,N_2772,N_2573);
nor U3376 (N_3376,N_2939,N_2916);
or U3377 (N_3377,N_2594,N_2562);
and U3378 (N_3378,N_2681,N_2856);
and U3379 (N_3379,N_2905,N_2868);
nand U3380 (N_3380,N_2902,N_2524);
nor U3381 (N_3381,N_2890,N_2965);
or U3382 (N_3382,N_2734,N_2511);
nor U3383 (N_3383,N_2587,N_2855);
and U3384 (N_3384,N_2581,N_2548);
and U3385 (N_3385,N_2542,N_2963);
xnor U3386 (N_3386,N_2572,N_2554);
nand U3387 (N_3387,N_2875,N_2753);
nand U3388 (N_3388,N_2620,N_2858);
xnor U3389 (N_3389,N_2902,N_2993);
and U3390 (N_3390,N_2721,N_2966);
and U3391 (N_3391,N_2551,N_2958);
nand U3392 (N_3392,N_2551,N_2968);
or U3393 (N_3393,N_2729,N_2989);
nor U3394 (N_3394,N_2910,N_2573);
nand U3395 (N_3395,N_2946,N_2758);
and U3396 (N_3396,N_2642,N_2554);
nand U3397 (N_3397,N_2619,N_2887);
nand U3398 (N_3398,N_2958,N_2980);
nand U3399 (N_3399,N_2623,N_2704);
and U3400 (N_3400,N_2561,N_2694);
nand U3401 (N_3401,N_2601,N_2677);
nand U3402 (N_3402,N_2617,N_2976);
nand U3403 (N_3403,N_2734,N_2716);
nor U3404 (N_3404,N_2915,N_2914);
xnor U3405 (N_3405,N_2666,N_2789);
nand U3406 (N_3406,N_2754,N_2824);
xnor U3407 (N_3407,N_2955,N_2602);
nand U3408 (N_3408,N_2567,N_2648);
nand U3409 (N_3409,N_2715,N_2565);
nor U3410 (N_3410,N_2980,N_2650);
nor U3411 (N_3411,N_2826,N_2884);
or U3412 (N_3412,N_2804,N_2862);
nor U3413 (N_3413,N_2928,N_2526);
nor U3414 (N_3414,N_2784,N_2872);
nor U3415 (N_3415,N_2697,N_2816);
xor U3416 (N_3416,N_2780,N_2805);
nand U3417 (N_3417,N_2801,N_2967);
xor U3418 (N_3418,N_2648,N_2849);
and U3419 (N_3419,N_2755,N_2702);
nor U3420 (N_3420,N_2837,N_2770);
nand U3421 (N_3421,N_2625,N_2848);
xor U3422 (N_3422,N_2511,N_2663);
nand U3423 (N_3423,N_2797,N_2910);
nor U3424 (N_3424,N_2517,N_2731);
and U3425 (N_3425,N_2679,N_2589);
nor U3426 (N_3426,N_2772,N_2709);
xor U3427 (N_3427,N_2955,N_2997);
or U3428 (N_3428,N_2808,N_2561);
nand U3429 (N_3429,N_2915,N_2630);
nor U3430 (N_3430,N_2820,N_2881);
nor U3431 (N_3431,N_2712,N_2914);
or U3432 (N_3432,N_2900,N_2902);
nor U3433 (N_3433,N_2695,N_2524);
nand U3434 (N_3434,N_2789,N_2883);
or U3435 (N_3435,N_2691,N_2584);
nor U3436 (N_3436,N_2876,N_2901);
xor U3437 (N_3437,N_2566,N_2648);
nor U3438 (N_3438,N_2542,N_2616);
and U3439 (N_3439,N_2630,N_2891);
xnor U3440 (N_3440,N_2804,N_2708);
xor U3441 (N_3441,N_2975,N_2871);
xor U3442 (N_3442,N_2906,N_2931);
nand U3443 (N_3443,N_2544,N_2893);
and U3444 (N_3444,N_2645,N_2847);
and U3445 (N_3445,N_2824,N_2715);
and U3446 (N_3446,N_2907,N_2595);
nor U3447 (N_3447,N_2742,N_2656);
nor U3448 (N_3448,N_2905,N_2971);
nor U3449 (N_3449,N_2675,N_2881);
nor U3450 (N_3450,N_2971,N_2995);
nand U3451 (N_3451,N_2703,N_2908);
xor U3452 (N_3452,N_2837,N_2833);
nor U3453 (N_3453,N_2812,N_2726);
and U3454 (N_3454,N_2687,N_2544);
nand U3455 (N_3455,N_2619,N_2575);
and U3456 (N_3456,N_2622,N_2827);
nand U3457 (N_3457,N_2625,N_2514);
or U3458 (N_3458,N_2510,N_2512);
and U3459 (N_3459,N_2729,N_2695);
and U3460 (N_3460,N_2882,N_2511);
and U3461 (N_3461,N_2869,N_2919);
or U3462 (N_3462,N_2719,N_2795);
and U3463 (N_3463,N_2602,N_2899);
xor U3464 (N_3464,N_2624,N_2515);
or U3465 (N_3465,N_2545,N_2629);
or U3466 (N_3466,N_2662,N_2962);
nor U3467 (N_3467,N_2573,N_2782);
nand U3468 (N_3468,N_2949,N_2924);
xnor U3469 (N_3469,N_2614,N_2960);
xor U3470 (N_3470,N_2707,N_2642);
nand U3471 (N_3471,N_2895,N_2692);
nand U3472 (N_3472,N_2815,N_2739);
nand U3473 (N_3473,N_2733,N_2701);
nor U3474 (N_3474,N_2732,N_2916);
and U3475 (N_3475,N_2538,N_2525);
nor U3476 (N_3476,N_2969,N_2920);
nor U3477 (N_3477,N_2774,N_2517);
and U3478 (N_3478,N_2952,N_2787);
nor U3479 (N_3479,N_2893,N_2929);
and U3480 (N_3480,N_2854,N_2818);
nand U3481 (N_3481,N_2913,N_2544);
nand U3482 (N_3482,N_2882,N_2796);
xor U3483 (N_3483,N_2812,N_2819);
xnor U3484 (N_3484,N_2892,N_2885);
nand U3485 (N_3485,N_2510,N_2671);
nor U3486 (N_3486,N_2688,N_2779);
nor U3487 (N_3487,N_2940,N_2857);
nand U3488 (N_3488,N_2897,N_2753);
and U3489 (N_3489,N_2998,N_2868);
or U3490 (N_3490,N_2621,N_2501);
xor U3491 (N_3491,N_2678,N_2672);
nand U3492 (N_3492,N_2859,N_2793);
nor U3493 (N_3493,N_2804,N_2624);
nor U3494 (N_3494,N_2706,N_2730);
and U3495 (N_3495,N_2783,N_2707);
and U3496 (N_3496,N_2514,N_2702);
or U3497 (N_3497,N_2511,N_2646);
and U3498 (N_3498,N_2562,N_2882);
nand U3499 (N_3499,N_2946,N_2887);
and U3500 (N_3500,N_3229,N_3006);
and U3501 (N_3501,N_3443,N_3078);
xor U3502 (N_3502,N_3479,N_3266);
xnor U3503 (N_3503,N_3273,N_3373);
nor U3504 (N_3504,N_3206,N_3114);
xnor U3505 (N_3505,N_3001,N_3246);
or U3506 (N_3506,N_3093,N_3157);
or U3507 (N_3507,N_3057,N_3103);
or U3508 (N_3508,N_3307,N_3065);
and U3509 (N_3509,N_3327,N_3277);
nor U3510 (N_3510,N_3461,N_3320);
or U3511 (N_3511,N_3488,N_3066);
and U3512 (N_3512,N_3007,N_3261);
nand U3513 (N_3513,N_3087,N_3298);
xor U3514 (N_3514,N_3036,N_3013);
xor U3515 (N_3515,N_3258,N_3015);
nand U3516 (N_3516,N_3043,N_3251);
xnor U3517 (N_3517,N_3364,N_3353);
xnor U3518 (N_3518,N_3077,N_3407);
nand U3519 (N_3519,N_3440,N_3199);
nor U3520 (N_3520,N_3357,N_3146);
xnor U3521 (N_3521,N_3347,N_3183);
nand U3522 (N_3522,N_3321,N_3310);
xor U3523 (N_3523,N_3299,N_3195);
nand U3524 (N_3524,N_3457,N_3463);
xor U3525 (N_3525,N_3159,N_3196);
nand U3526 (N_3526,N_3282,N_3305);
or U3527 (N_3527,N_3296,N_3014);
nand U3528 (N_3528,N_3331,N_3155);
xnor U3529 (N_3529,N_3056,N_3302);
xnor U3530 (N_3530,N_3371,N_3102);
or U3531 (N_3531,N_3030,N_3079);
xor U3532 (N_3532,N_3100,N_3227);
nor U3533 (N_3533,N_3374,N_3438);
xnor U3534 (N_3534,N_3050,N_3085);
or U3535 (N_3535,N_3274,N_3349);
and U3536 (N_3536,N_3329,N_3315);
and U3537 (N_3537,N_3492,N_3234);
xor U3538 (N_3538,N_3242,N_3301);
nand U3539 (N_3539,N_3460,N_3401);
or U3540 (N_3540,N_3108,N_3205);
nand U3541 (N_3541,N_3002,N_3420);
or U3542 (N_3542,N_3498,N_3414);
nor U3543 (N_3543,N_3263,N_3481);
xor U3544 (N_3544,N_3366,N_3252);
xor U3545 (N_3545,N_3083,N_3484);
nand U3546 (N_3546,N_3293,N_3496);
and U3547 (N_3547,N_3117,N_3419);
or U3548 (N_3548,N_3437,N_3126);
and U3549 (N_3549,N_3360,N_3179);
nand U3550 (N_3550,N_3431,N_3332);
xnor U3551 (N_3551,N_3335,N_3330);
or U3552 (N_3552,N_3323,N_3406);
and U3553 (N_3553,N_3225,N_3433);
xor U3554 (N_3554,N_3200,N_3230);
or U3555 (N_3555,N_3344,N_3156);
xnor U3556 (N_3556,N_3141,N_3280);
nand U3557 (N_3557,N_3037,N_3023);
or U3558 (N_3558,N_3226,N_3415);
nor U3559 (N_3559,N_3361,N_3129);
xor U3560 (N_3560,N_3368,N_3047);
xor U3561 (N_3561,N_3352,N_3005);
and U3562 (N_3562,N_3188,N_3107);
xor U3563 (N_3563,N_3018,N_3308);
or U3564 (N_3564,N_3418,N_3191);
and U3565 (N_3565,N_3203,N_3193);
nand U3566 (N_3566,N_3499,N_3459);
nor U3567 (N_3567,N_3041,N_3209);
nor U3568 (N_3568,N_3053,N_3283);
and U3569 (N_3569,N_3491,N_3091);
or U3570 (N_3570,N_3482,N_3094);
xor U3571 (N_3571,N_3120,N_3171);
and U3572 (N_3572,N_3092,N_3081);
and U3573 (N_3573,N_3121,N_3137);
xnor U3574 (N_3574,N_3376,N_3086);
and U3575 (N_3575,N_3370,N_3393);
or U3576 (N_3576,N_3149,N_3465);
and U3577 (N_3577,N_3113,N_3148);
xor U3578 (N_3578,N_3178,N_3428);
and U3579 (N_3579,N_3316,N_3430);
nand U3580 (N_3580,N_3343,N_3469);
and U3581 (N_3581,N_3319,N_3346);
nand U3582 (N_3582,N_3182,N_3445);
or U3583 (N_3583,N_3067,N_3217);
xor U3584 (N_3584,N_3221,N_3142);
nand U3585 (N_3585,N_3294,N_3236);
xnor U3586 (N_3586,N_3076,N_3351);
xor U3587 (N_3587,N_3424,N_3454);
xnor U3588 (N_3588,N_3204,N_3449);
nor U3589 (N_3589,N_3385,N_3048);
and U3590 (N_3590,N_3208,N_3304);
or U3591 (N_3591,N_3487,N_3413);
and U3592 (N_3592,N_3213,N_3281);
or U3593 (N_3593,N_3279,N_3003);
xnor U3594 (N_3594,N_3216,N_3004);
or U3595 (N_3595,N_3358,N_3309);
nor U3596 (N_3596,N_3444,N_3462);
nor U3597 (N_3597,N_3244,N_3400);
nor U3598 (N_3598,N_3333,N_3340);
nand U3599 (N_3599,N_3185,N_3426);
nor U3600 (N_3600,N_3019,N_3194);
or U3601 (N_3601,N_3485,N_3169);
nor U3602 (N_3602,N_3009,N_3378);
or U3603 (N_3603,N_3254,N_3220);
nand U3604 (N_3604,N_3134,N_3474);
and U3605 (N_3605,N_3324,N_3446);
or U3606 (N_3606,N_3029,N_3174);
and U3607 (N_3607,N_3231,N_3202);
nor U3608 (N_3608,N_3211,N_3034);
xnor U3609 (N_3609,N_3111,N_3365);
nand U3610 (N_3610,N_3466,N_3166);
nor U3611 (N_3611,N_3115,N_3161);
nand U3612 (N_3612,N_3441,N_3022);
nand U3613 (N_3613,N_3223,N_3212);
or U3614 (N_3614,N_3239,N_3033);
or U3615 (N_3615,N_3452,N_3080);
nand U3616 (N_3616,N_3247,N_3381);
or U3617 (N_3617,N_3038,N_3404);
nand U3618 (N_3618,N_3442,N_3396);
nor U3619 (N_3619,N_3044,N_3024);
xnor U3620 (N_3620,N_3417,N_3104);
and U3621 (N_3621,N_3132,N_3054);
nand U3622 (N_3622,N_3477,N_3032);
or U3623 (N_3623,N_3392,N_3164);
nand U3624 (N_3624,N_3110,N_3140);
xor U3625 (N_3625,N_3314,N_3421);
nor U3626 (N_3626,N_3153,N_3010);
nor U3627 (N_3627,N_3180,N_3342);
or U3628 (N_3628,N_3233,N_3160);
or U3629 (N_3629,N_3000,N_3362);
and U3630 (N_3630,N_3486,N_3040);
and U3631 (N_3631,N_3128,N_3409);
and U3632 (N_3632,N_3095,N_3173);
nor U3633 (N_3633,N_3399,N_3248);
xor U3634 (N_3634,N_3427,N_3215);
nand U3635 (N_3635,N_3028,N_3106);
nand U3636 (N_3636,N_3243,N_3434);
or U3637 (N_3637,N_3402,N_3397);
nor U3638 (N_3638,N_3354,N_3475);
or U3639 (N_3639,N_3101,N_3497);
or U3640 (N_3640,N_3058,N_3090);
and U3641 (N_3641,N_3326,N_3439);
nand U3642 (N_3642,N_3184,N_3493);
xor U3643 (N_3643,N_3175,N_3130);
and U3644 (N_3644,N_3168,N_3109);
xor U3645 (N_3645,N_3232,N_3272);
and U3646 (N_3646,N_3464,N_3025);
and U3647 (N_3647,N_3350,N_3412);
or U3648 (N_3648,N_3334,N_3060);
xnor U3649 (N_3649,N_3167,N_3453);
xor U3650 (N_3650,N_3312,N_3456);
or U3651 (N_3651,N_3388,N_3012);
and U3652 (N_3652,N_3467,N_3186);
xnor U3653 (N_3653,N_3097,N_3250);
nor U3654 (N_3654,N_3268,N_3386);
nor U3655 (N_3655,N_3139,N_3267);
xor U3656 (N_3656,N_3325,N_3295);
or U3657 (N_3657,N_3384,N_3145);
or U3658 (N_3658,N_3071,N_3235);
xor U3659 (N_3659,N_3472,N_3192);
nand U3660 (N_3660,N_3391,N_3069);
nand U3661 (N_3661,N_3099,N_3122);
xor U3662 (N_3662,N_3123,N_3483);
nor U3663 (N_3663,N_3152,N_3198);
xor U3664 (N_3664,N_3317,N_3422);
and U3665 (N_3665,N_3468,N_3052);
and U3666 (N_3666,N_3436,N_3218);
and U3667 (N_3667,N_3435,N_3318);
xor U3668 (N_3668,N_3133,N_3131);
nand U3669 (N_3669,N_3476,N_3098);
nand U3670 (N_3670,N_3119,N_3471);
nand U3671 (N_3671,N_3403,N_3031);
and U3672 (N_3672,N_3219,N_3458);
and U3673 (N_3673,N_3240,N_3292);
and U3674 (N_3674,N_3207,N_3395);
nor U3675 (N_3675,N_3494,N_3172);
nand U3676 (N_3676,N_3241,N_3062);
xor U3677 (N_3677,N_3398,N_3313);
and U3678 (N_3678,N_3075,N_3051);
or U3679 (N_3679,N_3027,N_3450);
nand U3680 (N_3680,N_3249,N_3214);
and U3681 (N_3681,N_3480,N_3070);
nand U3682 (N_3682,N_3288,N_3088);
and U3683 (N_3683,N_3377,N_3257);
xnor U3684 (N_3684,N_3064,N_3068);
nor U3685 (N_3685,N_3020,N_3336);
nor U3686 (N_3686,N_3016,N_3059);
nor U3687 (N_3687,N_3049,N_3238);
nand U3688 (N_3688,N_3394,N_3256);
nand U3689 (N_3689,N_3063,N_3181);
nand U3690 (N_3690,N_3228,N_3074);
nor U3691 (N_3691,N_3187,N_3408);
nor U3692 (N_3692,N_3447,N_3300);
nand U3693 (N_3693,N_3124,N_3303);
or U3694 (N_3694,N_3045,N_3008);
or U3695 (N_3695,N_3135,N_3410);
or U3696 (N_3696,N_3151,N_3286);
nor U3697 (N_3697,N_3432,N_3405);
xnor U3698 (N_3698,N_3262,N_3495);
or U3699 (N_3699,N_3337,N_3035);
and U3700 (N_3700,N_3253,N_3154);
or U3701 (N_3701,N_3042,N_3489);
nand U3702 (N_3702,N_3356,N_3285);
and U3703 (N_3703,N_3348,N_3383);
xnor U3704 (N_3704,N_3201,N_3072);
xor U3705 (N_3705,N_3189,N_3190);
nor U3706 (N_3706,N_3116,N_3306);
nand U3707 (N_3707,N_3278,N_3210);
xnor U3708 (N_3708,N_3150,N_3297);
and U3709 (N_3709,N_3237,N_3369);
xor U3710 (N_3710,N_3158,N_3411);
nand U3711 (N_3711,N_3136,N_3118);
nand U3712 (N_3712,N_3448,N_3287);
nor U3713 (N_3713,N_3138,N_3359);
and U3714 (N_3714,N_3473,N_3289);
nor U3715 (N_3715,N_3105,N_3291);
xor U3716 (N_3716,N_3423,N_3112);
and U3717 (N_3717,N_3176,N_3026);
nand U3718 (N_3718,N_3082,N_3355);
nor U3719 (N_3719,N_3162,N_3269);
xnor U3720 (N_3720,N_3276,N_3290);
and U3721 (N_3721,N_3084,N_3380);
and U3722 (N_3722,N_3017,N_3341);
and U3723 (N_3723,N_3478,N_3255);
xor U3724 (N_3724,N_3372,N_3021);
and U3725 (N_3725,N_3322,N_3073);
and U3726 (N_3726,N_3125,N_3451);
nor U3727 (N_3727,N_3165,N_3197);
and U3728 (N_3728,N_3061,N_3039);
nor U3729 (N_3729,N_3455,N_3470);
nand U3730 (N_3730,N_3367,N_3264);
or U3731 (N_3731,N_3375,N_3379);
nor U3732 (N_3732,N_3339,N_3143);
or U3733 (N_3733,N_3245,N_3259);
and U3734 (N_3734,N_3345,N_3265);
and U3735 (N_3735,N_3271,N_3338);
nand U3736 (N_3736,N_3390,N_3147);
nor U3737 (N_3737,N_3096,N_3144);
xnor U3738 (N_3738,N_3177,N_3382);
and U3739 (N_3739,N_3127,N_3387);
or U3740 (N_3740,N_3224,N_3163);
nor U3741 (N_3741,N_3429,N_3222);
nand U3742 (N_3742,N_3328,N_3311);
nand U3743 (N_3743,N_3425,N_3389);
nor U3744 (N_3744,N_3416,N_3490);
or U3745 (N_3745,N_3284,N_3089);
xor U3746 (N_3746,N_3363,N_3055);
and U3747 (N_3747,N_3275,N_3011);
nor U3748 (N_3748,N_3270,N_3170);
xnor U3749 (N_3749,N_3260,N_3046);
nand U3750 (N_3750,N_3020,N_3402);
nand U3751 (N_3751,N_3114,N_3413);
xnor U3752 (N_3752,N_3001,N_3030);
xor U3753 (N_3753,N_3156,N_3006);
or U3754 (N_3754,N_3240,N_3112);
and U3755 (N_3755,N_3263,N_3132);
xnor U3756 (N_3756,N_3233,N_3446);
and U3757 (N_3757,N_3446,N_3194);
nand U3758 (N_3758,N_3222,N_3294);
nor U3759 (N_3759,N_3374,N_3089);
and U3760 (N_3760,N_3101,N_3278);
nor U3761 (N_3761,N_3357,N_3124);
and U3762 (N_3762,N_3006,N_3277);
xnor U3763 (N_3763,N_3008,N_3088);
or U3764 (N_3764,N_3067,N_3470);
nand U3765 (N_3765,N_3129,N_3108);
xor U3766 (N_3766,N_3151,N_3280);
nor U3767 (N_3767,N_3191,N_3156);
nand U3768 (N_3768,N_3417,N_3115);
nand U3769 (N_3769,N_3478,N_3458);
or U3770 (N_3770,N_3145,N_3198);
nand U3771 (N_3771,N_3319,N_3260);
nand U3772 (N_3772,N_3018,N_3215);
nor U3773 (N_3773,N_3193,N_3306);
and U3774 (N_3774,N_3072,N_3420);
nand U3775 (N_3775,N_3442,N_3318);
and U3776 (N_3776,N_3010,N_3470);
nand U3777 (N_3777,N_3081,N_3173);
nor U3778 (N_3778,N_3229,N_3211);
xnor U3779 (N_3779,N_3227,N_3430);
xor U3780 (N_3780,N_3276,N_3419);
nand U3781 (N_3781,N_3206,N_3063);
nand U3782 (N_3782,N_3468,N_3258);
and U3783 (N_3783,N_3130,N_3391);
nor U3784 (N_3784,N_3380,N_3406);
nand U3785 (N_3785,N_3312,N_3265);
nor U3786 (N_3786,N_3376,N_3024);
and U3787 (N_3787,N_3426,N_3182);
or U3788 (N_3788,N_3438,N_3384);
xor U3789 (N_3789,N_3049,N_3145);
and U3790 (N_3790,N_3272,N_3337);
and U3791 (N_3791,N_3221,N_3235);
nand U3792 (N_3792,N_3360,N_3397);
nand U3793 (N_3793,N_3388,N_3445);
xnor U3794 (N_3794,N_3391,N_3185);
nand U3795 (N_3795,N_3096,N_3243);
nand U3796 (N_3796,N_3278,N_3297);
xnor U3797 (N_3797,N_3078,N_3419);
nor U3798 (N_3798,N_3213,N_3138);
xnor U3799 (N_3799,N_3312,N_3056);
or U3800 (N_3800,N_3349,N_3473);
nand U3801 (N_3801,N_3133,N_3417);
or U3802 (N_3802,N_3208,N_3095);
xnor U3803 (N_3803,N_3251,N_3417);
nand U3804 (N_3804,N_3411,N_3106);
or U3805 (N_3805,N_3073,N_3250);
nand U3806 (N_3806,N_3316,N_3393);
or U3807 (N_3807,N_3351,N_3408);
nor U3808 (N_3808,N_3396,N_3213);
or U3809 (N_3809,N_3110,N_3150);
nor U3810 (N_3810,N_3202,N_3137);
and U3811 (N_3811,N_3280,N_3490);
xor U3812 (N_3812,N_3319,N_3000);
nand U3813 (N_3813,N_3250,N_3396);
nor U3814 (N_3814,N_3154,N_3270);
or U3815 (N_3815,N_3474,N_3266);
or U3816 (N_3816,N_3076,N_3285);
nor U3817 (N_3817,N_3223,N_3411);
or U3818 (N_3818,N_3003,N_3394);
and U3819 (N_3819,N_3422,N_3250);
and U3820 (N_3820,N_3159,N_3422);
nor U3821 (N_3821,N_3010,N_3316);
or U3822 (N_3822,N_3383,N_3085);
xor U3823 (N_3823,N_3466,N_3246);
nor U3824 (N_3824,N_3259,N_3302);
and U3825 (N_3825,N_3267,N_3178);
and U3826 (N_3826,N_3414,N_3033);
xnor U3827 (N_3827,N_3383,N_3180);
and U3828 (N_3828,N_3319,N_3347);
nor U3829 (N_3829,N_3414,N_3003);
and U3830 (N_3830,N_3285,N_3440);
and U3831 (N_3831,N_3182,N_3338);
or U3832 (N_3832,N_3082,N_3158);
xnor U3833 (N_3833,N_3214,N_3493);
or U3834 (N_3834,N_3366,N_3182);
and U3835 (N_3835,N_3054,N_3114);
or U3836 (N_3836,N_3391,N_3290);
xor U3837 (N_3837,N_3182,N_3490);
xor U3838 (N_3838,N_3158,N_3042);
nand U3839 (N_3839,N_3119,N_3429);
and U3840 (N_3840,N_3084,N_3054);
xnor U3841 (N_3841,N_3235,N_3358);
nand U3842 (N_3842,N_3460,N_3237);
and U3843 (N_3843,N_3005,N_3476);
nor U3844 (N_3844,N_3214,N_3262);
nor U3845 (N_3845,N_3323,N_3100);
xor U3846 (N_3846,N_3077,N_3349);
or U3847 (N_3847,N_3177,N_3496);
nor U3848 (N_3848,N_3408,N_3171);
and U3849 (N_3849,N_3165,N_3168);
nor U3850 (N_3850,N_3224,N_3120);
nand U3851 (N_3851,N_3078,N_3369);
and U3852 (N_3852,N_3113,N_3319);
or U3853 (N_3853,N_3097,N_3126);
or U3854 (N_3854,N_3261,N_3242);
xnor U3855 (N_3855,N_3457,N_3210);
or U3856 (N_3856,N_3231,N_3183);
or U3857 (N_3857,N_3414,N_3157);
or U3858 (N_3858,N_3362,N_3168);
or U3859 (N_3859,N_3179,N_3265);
nor U3860 (N_3860,N_3421,N_3285);
nor U3861 (N_3861,N_3496,N_3152);
nor U3862 (N_3862,N_3269,N_3437);
or U3863 (N_3863,N_3230,N_3400);
nand U3864 (N_3864,N_3368,N_3153);
and U3865 (N_3865,N_3491,N_3131);
or U3866 (N_3866,N_3490,N_3045);
nand U3867 (N_3867,N_3431,N_3083);
and U3868 (N_3868,N_3186,N_3175);
and U3869 (N_3869,N_3334,N_3117);
or U3870 (N_3870,N_3025,N_3060);
xnor U3871 (N_3871,N_3190,N_3090);
and U3872 (N_3872,N_3353,N_3073);
xnor U3873 (N_3873,N_3373,N_3093);
or U3874 (N_3874,N_3383,N_3408);
and U3875 (N_3875,N_3305,N_3361);
or U3876 (N_3876,N_3113,N_3437);
nor U3877 (N_3877,N_3394,N_3494);
and U3878 (N_3878,N_3259,N_3314);
nand U3879 (N_3879,N_3059,N_3174);
nand U3880 (N_3880,N_3232,N_3243);
nand U3881 (N_3881,N_3353,N_3159);
or U3882 (N_3882,N_3002,N_3059);
nand U3883 (N_3883,N_3164,N_3497);
xnor U3884 (N_3884,N_3264,N_3153);
nor U3885 (N_3885,N_3205,N_3282);
and U3886 (N_3886,N_3114,N_3021);
or U3887 (N_3887,N_3347,N_3421);
nor U3888 (N_3888,N_3023,N_3214);
nand U3889 (N_3889,N_3297,N_3423);
or U3890 (N_3890,N_3464,N_3062);
nor U3891 (N_3891,N_3130,N_3318);
xnor U3892 (N_3892,N_3331,N_3242);
xnor U3893 (N_3893,N_3398,N_3087);
and U3894 (N_3894,N_3201,N_3285);
nand U3895 (N_3895,N_3275,N_3220);
or U3896 (N_3896,N_3102,N_3282);
or U3897 (N_3897,N_3331,N_3190);
or U3898 (N_3898,N_3492,N_3472);
or U3899 (N_3899,N_3366,N_3462);
or U3900 (N_3900,N_3362,N_3387);
nand U3901 (N_3901,N_3111,N_3153);
and U3902 (N_3902,N_3451,N_3004);
nor U3903 (N_3903,N_3485,N_3224);
and U3904 (N_3904,N_3146,N_3213);
nand U3905 (N_3905,N_3362,N_3241);
or U3906 (N_3906,N_3421,N_3342);
nand U3907 (N_3907,N_3365,N_3119);
nand U3908 (N_3908,N_3123,N_3051);
nor U3909 (N_3909,N_3311,N_3333);
xor U3910 (N_3910,N_3178,N_3208);
and U3911 (N_3911,N_3427,N_3126);
or U3912 (N_3912,N_3098,N_3113);
and U3913 (N_3913,N_3431,N_3214);
or U3914 (N_3914,N_3145,N_3354);
or U3915 (N_3915,N_3405,N_3444);
nand U3916 (N_3916,N_3287,N_3267);
nor U3917 (N_3917,N_3386,N_3053);
nand U3918 (N_3918,N_3484,N_3408);
and U3919 (N_3919,N_3453,N_3320);
xnor U3920 (N_3920,N_3096,N_3447);
nand U3921 (N_3921,N_3320,N_3004);
xnor U3922 (N_3922,N_3226,N_3015);
nor U3923 (N_3923,N_3208,N_3221);
nand U3924 (N_3924,N_3293,N_3413);
nor U3925 (N_3925,N_3046,N_3078);
nand U3926 (N_3926,N_3263,N_3006);
and U3927 (N_3927,N_3255,N_3482);
nor U3928 (N_3928,N_3152,N_3337);
nand U3929 (N_3929,N_3066,N_3182);
xnor U3930 (N_3930,N_3325,N_3279);
xnor U3931 (N_3931,N_3093,N_3246);
nor U3932 (N_3932,N_3255,N_3398);
nand U3933 (N_3933,N_3266,N_3194);
nand U3934 (N_3934,N_3197,N_3473);
xor U3935 (N_3935,N_3008,N_3070);
or U3936 (N_3936,N_3257,N_3341);
xor U3937 (N_3937,N_3059,N_3063);
and U3938 (N_3938,N_3450,N_3150);
xnor U3939 (N_3939,N_3012,N_3058);
nand U3940 (N_3940,N_3396,N_3486);
or U3941 (N_3941,N_3392,N_3379);
and U3942 (N_3942,N_3128,N_3212);
or U3943 (N_3943,N_3200,N_3296);
nor U3944 (N_3944,N_3311,N_3296);
and U3945 (N_3945,N_3144,N_3343);
nor U3946 (N_3946,N_3116,N_3073);
and U3947 (N_3947,N_3498,N_3066);
or U3948 (N_3948,N_3423,N_3315);
or U3949 (N_3949,N_3167,N_3243);
or U3950 (N_3950,N_3332,N_3397);
nand U3951 (N_3951,N_3432,N_3469);
and U3952 (N_3952,N_3231,N_3159);
or U3953 (N_3953,N_3014,N_3464);
nand U3954 (N_3954,N_3466,N_3105);
xnor U3955 (N_3955,N_3266,N_3471);
and U3956 (N_3956,N_3169,N_3079);
nand U3957 (N_3957,N_3200,N_3026);
or U3958 (N_3958,N_3325,N_3029);
xnor U3959 (N_3959,N_3485,N_3016);
or U3960 (N_3960,N_3055,N_3494);
and U3961 (N_3961,N_3469,N_3260);
xor U3962 (N_3962,N_3174,N_3495);
nand U3963 (N_3963,N_3330,N_3471);
xor U3964 (N_3964,N_3159,N_3359);
and U3965 (N_3965,N_3268,N_3029);
xor U3966 (N_3966,N_3492,N_3022);
xor U3967 (N_3967,N_3367,N_3488);
xor U3968 (N_3968,N_3246,N_3475);
xnor U3969 (N_3969,N_3483,N_3011);
nand U3970 (N_3970,N_3289,N_3265);
and U3971 (N_3971,N_3130,N_3127);
nor U3972 (N_3972,N_3390,N_3252);
nor U3973 (N_3973,N_3162,N_3430);
or U3974 (N_3974,N_3209,N_3348);
xor U3975 (N_3975,N_3261,N_3488);
xnor U3976 (N_3976,N_3060,N_3419);
nor U3977 (N_3977,N_3295,N_3123);
nor U3978 (N_3978,N_3117,N_3137);
and U3979 (N_3979,N_3327,N_3351);
nand U3980 (N_3980,N_3031,N_3266);
and U3981 (N_3981,N_3348,N_3342);
nand U3982 (N_3982,N_3393,N_3296);
nand U3983 (N_3983,N_3078,N_3195);
or U3984 (N_3984,N_3210,N_3084);
and U3985 (N_3985,N_3485,N_3243);
and U3986 (N_3986,N_3283,N_3259);
nor U3987 (N_3987,N_3271,N_3394);
and U3988 (N_3988,N_3395,N_3311);
or U3989 (N_3989,N_3092,N_3028);
and U3990 (N_3990,N_3137,N_3040);
or U3991 (N_3991,N_3209,N_3142);
nor U3992 (N_3992,N_3166,N_3138);
or U3993 (N_3993,N_3118,N_3479);
nand U3994 (N_3994,N_3410,N_3161);
nor U3995 (N_3995,N_3045,N_3420);
xnor U3996 (N_3996,N_3218,N_3337);
nor U3997 (N_3997,N_3421,N_3307);
or U3998 (N_3998,N_3264,N_3468);
xnor U3999 (N_3999,N_3432,N_3435);
xor U4000 (N_4000,N_3766,N_3929);
and U4001 (N_4001,N_3526,N_3851);
and U4002 (N_4002,N_3638,N_3806);
nand U4003 (N_4003,N_3558,N_3949);
xnor U4004 (N_4004,N_3898,N_3601);
or U4005 (N_4005,N_3504,N_3871);
xnor U4006 (N_4006,N_3826,N_3714);
or U4007 (N_4007,N_3562,N_3881);
nor U4008 (N_4008,N_3603,N_3663);
or U4009 (N_4009,N_3981,N_3625);
or U4010 (N_4010,N_3828,N_3692);
xnor U4011 (N_4011,N_3551,N_3676);
and U4012 (N_4012,N_3643,N_3689);
and U4013 (N_4013,N_3770,N_3564);
xor U4014 (N_4014,N_3545,N_3892);
and U4015 (N_4015,N_3712,N_3698);
nor U4016 (N_4016,N_3955,N_3668);
nand U4017 (N_4017,N_3715,N_3957);
xor U4018 (N_4018,N_3595,N_3758);
and U4019 (N_4019,N_3827,N_3612);
nand U4020 (N_4020,N_3855,N_3660);
nand U4021 (N_4021,N_3719,N_3598);
nor U4022 (N_4022,N_3838,N_3571);
xnor U4023 (N_4023,N_3756,N_3720);
or U4024 (N_4024,N_3535,N_3584);
nand U4025 (N_4025,N_3688,N_3619);
xor U4026 (N_4026,N_3975,N_3775);
xor U4027 (N_4027,N_3536,N_3730);
and U4028 (N_4028,N_3632,N_3729);
nand U4029 (N_4029,N_3800,N_3561);
or U4030 (N_4030,N_3780,N_3644);
or U4031 (N_4031,N_3565,N_3661);
nand U4032 (N_4032,N_3710,N_3938);
and U4033 (N_4033,N_3525,N_3646);
xnor U4034 (N_4034,N_3507,N_3925);
and U4035 (N_4035,N_3905,N_3534);
xor U4036 (N_4036,N_3736,N_3823);
nand U4037 (N_4037,N_3750,N_3718);
nor U4038 (N_4038,N_3642,N_3841);
xnor U4039 (N_4039,N_3967,N_3633);
nor U4040 (N_4040,N_3825,N_3793);
and U4041 (N_4041,N_3782,N_3917);
or U4042 (N_4042,N_3966,N_3749);
xor U4043 (N_4043,N_3690,N_3786);
and U4044 (N_4044,N_3854,N_3931);
and U4045 (N_4045,N_3735,N_3792);
xnor U4046 (N_4046,N_3997,N_3964);
xor U4047 (N_4047,N_3591,N_3909);
nand U4048 (N_4048,N_3654,N_3550);
nand U4049 (N_4049,N_3867,N_3670);
and U4050 (N_4050,N_3741,N_3830);
nor U4051 (N_4051,N_3728,N_3958);
nand U4052 (N_4052,N_3631,N_3563);
and U4053 (N_4053,N_3635,N_3748);
xor U4054 (N_4054,N_3559,N_3636);
xor U4055 (N_4055,N_3802,N_3916);
and U4056 (N_4056,N_3815,N_3685);
nand U4057 (N_4057,N_3989,N_3990);
nand U4058 (N_4058,N_3731,N_3543);
and U4059 (N_4059,N_3761,N_3896);
nor U4060 (N_4060,N_3502,N_3506);
xor U4061 (N_4061,N_3732,N_3940);
and U4062 (N_4062,N_3936,N_3512);
xnor U4063 (N_4063,N_3615,N_3983);
nand U4064 (N_4064,N_3653,N_3645);
nand U4065 (N_4065,N_3829,N_3546);
and U4066 (N_4066,N_3683,N_3878);
or U4067 (N_4067,N_3724,N_3630);
and U4068 (N_4068,N_3877,N_3888);
nand U4069 (N_4069,N_3999,N_3764);
or U4070 (N_4070,N_3751,N_3928);
or U4071 (N_4071,N_3529,N_3570);
nor U4072 (N_4072,N_3614,N_3588);
xor U4073 (N_4073,N_3589,N_3622);
nor U4074 (N_4074,N_3651,N_3921);
or U4075 (N_4075,N_3869,N_3807);
or U4076 (N_4076,N_3942,N_3795);
and U4077 (N_4077,N_3599,N_3585);
xnor U4078 (N_4078,N_3541,N_3693);
or U4079 (N_4079,N_3530,N_3824);
or U4080 (N_4080,N_3652,N_3608);
nand U4081 (N_4081,N_3560,N_3915);
or U4082 (N_4082,N_3518,N_3757);
or U4083 (N_4083,N_3734,N_3965);
nand U4084 (N_4084,N_3739,N_3717);
nand U4085 (N_4085,N_3620,N_3813);
or U4086 (N_4086,N_3796,N_3572);
or U4087 (N_4087,N_3821,N_3787);
or U4088 (N_4088,N_3863,N_3773);
nand U4089 (N_4089,N_3969,N_3771);
xor U4090 (N_4090,N_3658,N_3845);
nand U4091 (N_4091,N_3846,N_3567);
nand U4092 (N_4092,N_3575,N_3934);
nand U4093 (N_4093,N_3705,N_3686);
xnor U4094 (N_4094,N_3699,N_3850);
nand U4095 (N_4095,N_3669,N_3743);
and U4096 (N_4096,N_3860,N_3818);
nor U4097 (N_4097,N_3596,N_3948);
xnor U4098 (N_4098,N_3794,N_3656);
or U4099 (N_4099,N_3662,N_3856);
nand U4100 (N_4100,N_3779,N_3616);
nor U4101 (N_4101,N_3857,N_3996);
nor U4102 (N_4102,N_3994,N_3801);
or U4103 (N_4103,N_3872,N_3918);
nor U4104 (N_4104,N_3664,N_3944);
nand U4105 (N_4105,N_3959,N_3574);
nor U4106 (N_4106,N_3882,N_3726);
nand U4107 (N_4107,N_3820,N_3586);
and U4108 (N_4108,N_3709,N_3727);
nor U4109 (N_4109,N_3691,N_3680);
xor U4110 (N_4110,N_3523,N_3939);
or U4111 (N_4111,N_3703,N_3781);
nand U4112 (N_4112,N_3941,N_3597);
and U4113 (N_4113,N_3988,N_3557);
nor U4114 (N_4114,N_3763,N_3516);
xnor U4115 (N_4115,N_3890,N_3899);
or U4116 (N_4116,N_3903,N_3953);
nand U4117 (N_4117,N_3737,N_3665);
or U4118 (N_4118,N_3513,N_3627);
and U4119 (N_4119,N_3978,N_3870);
xor U4120 (N_4120,N_3935,N_3579);
or U4121 (N_4121,N_3687,N_3883);
nor U4122 (N_4122,N_3920,N_3681);
and U4123 (N_4123,N_3947,N_3992);
or U4124 (N_4124,N_3859,N_3666);
or U4125 (N_4125,N_3533,N_3522);
nor U4126 (N_4126,N_3640,N_3812);
nand U4127 (N_4127,N_3875,N_3865);
xor U4128 (N_4128,N_3626,N_3544);
nor U4129 (N_4129,N_3581,N_3832);
or U4130 (N_4130,N_3976,N_3623);
and U4131 (N_4131,N_3702,N_3887);
xnor U4132 (N_4132,N_3803,N_3776);
or U4133 (N_4133,N_3542,N_3836);
nor U4134 (N_4134,N_3503,N_3744);
xnor U4135 (N_4135,N_3943,N_3956);
nand U4136 (N_4136,N_3852,N_3907);
nand U4137 (N_4137,N_3667,N_3605);
nor U4138 (N_4138,N_3762,N_3884);
nand U4139 (N_4139,N_3962,N_3835);
and U4140 (N_4140,N_3606,N_3822);
and U4141 (N_4141,N_3540,N_3639);
nand U4142 (N_4142,N_3974,N_3704);
nor U4143 (N_4143,N_3675,N_3873);
xor U4144 (N_4144,N_3894,N_3924);
or U4145 (N_4145,N_3919,N_3985);
and U4146 (N_4146,N_3723,N_3747);
nor U4147 (N_4147,N_3991,N_3861);
nand U4148 (N_4148,N_3752,N_3611);
and U4149 (N_4149,N_3906,N_3696);
nor U4150 (N_4150,N_3628,N_3971);
xnor U4151 (N_4151,N_3922,N_3713);
nor U4152 (N_4152,N_3501,N_3509);
or U4153 (N_4153,N_3740,N_3582);
or U4154 (N_4154,N_3914,N_3798);
nand U4155 (N_4155,N_3811,N_3769);
xor U4156 (N_4156,N_3566,N_3848);
and U4157 (N_4157,N_3933,N_3609);
and U4158 (N_4158,N_3755,N_3908);
and U4159 (N_4159,N_3834,N_3746);
and U4160 (N_4160,N_3515,N_3897);
nand U4161 (N_4161,N_3604,N_3968);
and U4162 (N_4162,N_3514,N_3960);
xnor U4163 (N_4163,N_3538,N_3913);
nand U4164 (N_4164,N_3701,N_3594);
nor U4165 (N_4165,N_3785,N_3624);
or U4166 (N_4166,N_3765,N_3554);
or U4167 (N_4167,N_3952,N_3866);
xnor U4168 (N_4168,N_3926,N_3777);
and U4169 (N_4169,N_3977,N_3767);
nand U4170 (N_4170,N_3858,N_3521);
or U4171 (N_4171,N_3721,N_3874);
nor U4172 (N_4172,N_3553,N_3843);
xnor U4173 (N_4173,N_3982,N_3677);
nor U4174 (N_4174,N_3520,N_3549);
xor U4175 (N_4175,N_3912,N_3864);
nor U4176 (N_4176,N_3602,N_3984);
or U4177 (N_4177,N_3816,N_3814);
or U4178 (N_4178,N_3774,N_3634);
nand U4179 (N_4179,N_3946,N_3970);
xnor U4180 (N_4180,N_3568,N_3697);
xnor U4181 (N_4181,N_3986,N_3837);
nor U4182 (N_4182,N_3847,N_3706);
or U4183 (N_4183,N_3500,N_3784);
nand U4184 (N_4184,N_3862,N_3655);
and U4185 (N_4185,N_3517,N_3889);
or U4186 (N_4186,N_3694,N_3853);
and U4187 (N_4187,N_3556,N_3657);
nand U4188 (N_4188,N_3979,N_3754);
and U4189 (N_4189,N_3895,N_3760);
nor U4190 (N_4190,N_3911,N_3849);
and U4191 (N_4191,N_3539,N_3809);
or U4192 (N_4192,N_3617,N_3972);
xor U4193 (N_4193,N_3930,N_3537);
or U4194 (N_4194,N_3527,N_3711);
or U4195 (N_4195,N_3790,N_3548);
nand U4196 (N_4196,N_3842,N_3508);
or U4197 (N_4197,N_3954,N_3524);
xor U4198 (N_4198,N_3951,N_3844);
and U4199 (N_4199,N_3700,N_3901);
and U4200 (N_4200,N_3637,N_3886);
nand U4201 (N_4201,N_3650,N_3885);
xor U4202 (N_4202,N_3722,N_3641);
nor U4203 (N_4203,N_3839,N_3573);
or U4204 (N_4204,N_3945,N_3674);
nand U4205 (N_4205,N_3576,N_3745);
and U4206 (N_4206,N_3891,N_3902);
nand U4207 (N_4207,N_3980,N_3684);
and U4208 (N_4208,N_3613,N_3659);
or U4209 (N_4209,N_3950,N_3927);
nand U4210 (N_4210,N_3961,N_3932);
nor U4211 (N_4211,N_3995,N_3577);
nor U4212 (N_4212,N_3973,N_3511);
or U4213 (N_4213,N_3580,N_3552);
and U4214 (N_4214,N_3578,N_3868);
and U4215 (N_4215,N_3649,N_3587);
nor U4216 (N_4216,N_3679,N_3904);
or U4217 (N_4217,N_3778,N_3808);
or U4218 (N_4218,N_3592,N_3600);
nand U4219 (N_4219,N_3876,N_3629);
and U4220 (N_4220,N_3569,N_3768);
nand U4221 (N_4221,N_3607,N_3742);
or U4222 (N_4222,N_3831,N_3772);
nor U4223 (N_4223,N_3993,N_3618);
or U4224 (N_4224,N_3879,N_3532);
and U4225 (N_4225,N_3672,N_3840);
and U4226 (N_4226,N_3725,N_3733);
xnor U4227 (N_4227,N_3910,N_3519);
xor U4228 (N_4228,N_3810,N_3528);
nand U4229 (N_4229,N_3791,N_3673);
nor U4230 (N_4230,N_3788,N_3987);
nand U4231 (N_4231,N_3900,N_3783);
xor U4232 (N_4232,N_3759,N_3805);
xor U4233 (N_4233,N_3648,N_3695);
and U4234 (N_4234,N_3708,N_3671);
xor U4235 (N_4235,N_3799,N_3716);
nand U4236 (N_4236,N_3707,N_3583);
nor U4237 (N_4237,N_3531,N_3817);
and U4238 (N_4238,N_3833,N_3937);
nor U4239 (N_4239,N_3678,N_3621);
nor U4240 (N_4240,N_3998,N_3753);
and U4241 (N_4241,N_3547,N_3555);
or U4242 (N_4242,N_3510,N_3819);
and U4243 (N_4243,N_3893,N_3647);
and U4244 (N_4244,N_3923,N_3789);
nor U4245 (N_4245,N_3963,N_3682);
nand U4246 (N_4246,N_3804,N_3610);
and U4247 (N_4247,N_3505,N_3593);
xnor U4248 (N_4248,N_3797,N_3590);
xor U4249 (N_4249,N_3738,N_3880);
or U4250 (N_4250,N_3733,N_3795);
and U4251 (N_4251,N_3967,N_3642);
or U4252 (N_4252,N_3974,N_3821);
nand U4253 (N_4253,N_3546,N_3580);
or U4254 (N_4254,N_3514,N_3953);
nor U4255 (N_4255,N_3866,N_3735);
nand U4256 (N_4256,N_3814,N_3724);
nand U4257 (N_4257,N_3650,N_3848);
nand U4258 (N_4258,N_3905,N_3987);
or U4259 (N_4259,N_3597,N_3517);
or U4260 (N_4260,N_3802,N_3658);
nand U4261 (N_4261,N_3942,N_3519);
and U4262 (N_4262,N_3767,N_3533);
nor U4263 (N_4263,N_3662,N_3630);
or U4264 (N_4264,N_3591,N_3774);
xor U4265 (N_4265,N_3583,N_3714);
nand U4266 (N_4266,N_3576,N_3554);
nor U4267 (N_4267,N_3873,N_3646);
xor U4268 (N_4268,N_3736,N_3830);
or U4269 (N_4269,N_3874,N_3792);
nand U4270 (N_4270,N_3764,N_3591);
nor U4271 (N_4271,N_3500,N_3888);
xnor U4272 (N_4272,N_3686,N_3690);
nor U4273 (N_4273,N_3969,N_3735);
nor U4274 (N_4274,N_3928,N_3845);
and U4275 (N_4275,N_3754,N_3817);
xnor U4276 (N_4276,N_3949,N_3926);
nor U4277 (N_4277,N_3510,N_3704);
xnor U4278 (N_4278,N_3947,N_3741);
and U4279 (N_4279,N_3687,N_3722);
nor U4280 (N_4280,N_3796,N_3818);
nand U4281 (N_4281,N_3565,N_3820);
or U4282 (N_4282,N_3829,N_3662);
and U4283 (N_4283,N_3533,N_3669);
nor U4284 (N_4284,N_3928,N_3909);
nand U4285 (N_4285,N_3742,N_3653);
or U4286 (N_4286,N_3931,N_3671);
nor U4287 (N_4287,N_3564,N_3990);
nor U4288 (N_4288,N_3861,N_3539);
or U4289 (N_4289,N_3966,N_3771);
or U4290 (N_4290,N_3700,N_3588);
or U4291 (N_4291,N_3507,N_3784);
nor U4292 (N_4292,N_3635,N_3661);
nor U4293 (N_4293,N_3912,N_3517);
or U4294 (N_4294,N_3822,N_3780);
and U4295 (N_4295,N_3501,N_3631);
or U4296 (N_4296,N_3625,N_3529);
or U4297 (N_4297,N_3865,N_3623);
nor U4298 (N_4298,N_3698,N_3655);
or U4299 (N_4299,N_3768,N_3814);
or U4300 (N_4300,N_3582,N_3970);
xor U4301 (N_4301,N_3742,N_3790);
nor U4302 (N_4302,N_3897,N_3660);
xor U4303 (N_4303,N_3746,N_3845);
xnor U4304 (N_4304,N_3556,N_3536);
nand U4305 (N_4305,N_3952,N_3631);
xor U4306 (N_4306,N_3624,N_3610);
nor U4307 (N_4307,N_3761,N_3826);
or U4308 (N_4308,N_3717,N_3911);
nor U4309 (N_4309,N_3816,N_3766);
nor U4310 (N_4310,N_3521,N_3589);
nand U4311 (N_4311,N_3624,N_3872);
nor U4312 (N_4312,N_3669,N_3673);
or U4313 (N_4313,N_3679,N_3620);
nor U4314 (N_4314,N_3812,N_3843);
nor U4315 (N_4315,N_3713,N_3932);
nor U4316 (N_4316,N_3895,N_3835);
or U4317 (N_4317,N_3677,N_3901);
nand U4318 (N_4318,N_3683,N_3669);
xnor U4319 (N_4319,N_3826,N_3917);
or U4320 (N_4320,N_3837,N_3801);
or U4321 (N_4321,N_3962,N_3935);
nor U4322 (N_4322,N_3573,N_3922);
or U4323 (N_4323,N_3717,N_3843);
and U4324 (N_4324,N_3627,N_3950);
xnor U4325 (N_4325,N_3825,N_3706);
and U4326 (N_4326,N_3766,N_3991);
nand U4327 (N_4327,N_3672,N_3877);
and U4328 (N_4328,N_3781,N_3894);
and U4329 (N_4329,N_3621,N_3600);
nor U4330 (N_4330,N_3967,N_3703);
nand U4331 (N_4331,N_3722,N_3503);
nand U4332 (N_4332,N_3730,N_3874);
nand U4333 (N_4333,N_3836,N_3562);
and U4334 (N_4334,N_3549,N_3861);
nor U4335 (N_4335,N_3594,N_3804);
xor U4336 (N_4336,N_3660,N_3734);
xnor U4337 (N_4337,N_3966,N_3901);
nand U4338 (N_4338,N_3685,N_3769);
xnor U4339 (N_4339,N_3517,N_3893);
or U4340 (N_4340,N_3835,N_3552);
xnor U4341 (N_4341,N_3548,N_3904);
nand U4342 (N_4342,N_3696,N_3954);
nor U4343 (N_4343,N_3590,N_3997);
or U4344 (N_4344,N_3809,N_3665);
nand U4345 (N_4345,N_3514,N_3899);
nand U4346 (N_4346,N_3739,N_3942);
or U4347 (N_4347,N_3935,N_3505);
nand U4348 (N_4348,N_3615,N_3524);
or U4349 (N_4349,N_3872,N_3502);
nand U4350 (N_4350,N_3729,N_3615);
and U4351 (N_4351,N_3669,N_3827);
nor U4352 (N_4352,N_3914,N_3763);
and U4353 (N_4353,N_3776,N_3726);
and U4354 (N_4354,N_3793,N_3849);
nor U4355 (N_4355,N_3839,N_3590);
and U4356 (N_4356,N_3939,N_3559);
xnor U4357 (N_4357,N_3720,N_3655);
and U4358 (N_4358,N_3537,N_3877);
xor U4359 (N_4359,N_3684,N_3768);
xnor U4360 (N_4360,N_3632,N_3994);
nand U4361 (N_4361,N_3785,N_3925);
xor U4362 (N_4362,N_3929,N_3670);
nand U4363 (N_4363,N_3989,N_3886);
xnor U4364 (N_4364,N_3890,N_3597);
or U4365 (N_4365,N_3930,N_3560);
or U4366 (N_4366,N_3601,N_3522);
and U4367 (N_4367,N_3768,N_3501);
xnor U4368 (N_4368,N_3614,N_3996);
xnor U4369 (N_4369,N_3865,N_3985);
and U4370 (N_4370,N_3530,N_3539);
and U4371 (N_4371,N_3770,N_3864);
and U4372 (N_4372,N_3784,N_3748);
and U4373 (N_4373,N_3797,N_3617);
nor U4374 (N_4374,N_3824,N_3790);
nor U4375 (N_4375,N_3745,N_3775);
nor U4376 (N_4376,N_3801,N_3810);
nand U4377 (N_4377,N_3551,N_3627);
xor U4378 (N_4378,N_3847,N_3830);
and U4379 (N_4379,N_3885,N_3522);
or U4380 (N_4380,N_3744,N_3850);
and U4381 (N_4381,N_3599,N_3978);
nand U4382 (N_4382,N_3533,N_3879);
and U4383 (N_4383,N_3796,N_3917);
and U4384 (N_4384,N_3771,N_3981);
and U4385 (N_4385,N_3737,N_3686);
nand U4386 (N_4386,N_3926,N_3614);
and U4387 (N_4387,N_3788,N_3640);
xnor U4388 (N_4388,N_3885,N_3804);
nand U4389 (N_4389,N_3918,N_3954);
xnor U4390 (N_4390,N_3557,N_3603);
nor U4391 (N_4391,N_3957,N_3951);
nor U4392 (N_4392,N_3642,N_3884);
or U4393 (N_4393,N_3547,N_3741);
or U4394 (N_4394,N_3628,N_3972);
nand U4395 (N_4395,N_3903,N_3632);
nor U4396 (N_4396,N_3781,N_3765);
nand U4397 (N_4397,N_3855,N_3618);
or U4398 (N_4398,N_3991,N_3820);
and U4399 (N_4399,N_3573,N_3830);
or U4400 (N_4400,N_3901,N_3635);
nor U4401 (N_4401,N_3952,N_3678);
nand U4402 (N_4402,N_3500,N_3876);
nand U4403 (N_4403,N_3590,N_3623);
nand U4404 (N_4404,N_3877,N_3731);
and U4405 (N_4405,N_3642,N_3783);
nand U4406 (N_4406,N_3702,N_3695);
and U4407 (N_4407,N_3677,N_3539);
or U4408 (N_4408,N_3571,N_3661);
or U4409 (N_4409,N_3576,N_3681);
nand U4410 (N_4410,N_3848,N_3846);
or U4411 (N_4411,N_3765,N_3875);
or U4412 (N_4412,N_3656,N_3845);
xnor U4413 (N_4413,N_3643,N_3666);
xnor U4414 (N_4414,N_3774,N_3678);
and U4415 (N_4415,N_3889,N_3836);
nor U4416 (N_4416,N_3926,N_3730);
xor U4417 (N_4417,N_3586,N_3726);
xor U4418 (N_4418,N_3909,N_3559);
nand U4419 (N_4419,N_3611,N_3552);
nand U4420 (N_4420,N_3703,N_3790);
and U4421 (N_4421,N_3626,N_3943);
nor U4422 (N_4422,N_3733,N_3865);
or U4423 (N_4423,N_3931,N_3677);
nor U4424 (N_4424,N_3856,N_3840);
and U4425 (N_4425,N_3879,N_3526);
nand U4426 (N_4426,N_3822,N_3708);
and U4427 (N_4427,N_3532,N_3729);
nand U4428 (N_4428,N_3618,N_3533);
nand U4429 (N_4429,N_3999,N_3939);
xor U4430 (N_4430,N_3997,N_3557);
nor U4431 (N_4431,N_3928,N_3850);
nand U4432 (N_4432,N_3660,N_3786);
or U4433 (N_4433,N_3991,N_3858);
nand U4434 (N_4434,N_3919,N_3965);
nor U4435 (N_4435,N_3565,N_3531);
nor U4436 (N_4436,N_3634,N_3937);
xnor U4437 (N_4437,N_3669,N_3752);
nand U4438 (N_4438,N_3652,N_3570);
xor U4439 (N_4439,N_3506,N_3817);
nand U4440 (N_4440,N_3725,N_3662);
nand U4441 (N_4441,N_3635,N_3964);
xor U4442 (N_4442,N_3950,N_3519);
xnor U4443 (N_4443,N_3833,N_3981);
xnor U4444 (N_4444,N_3935,N_3898);
nand U4445 (N_4445,N_3704,N_3840);
and U4446 (N_4446,N_3999,N_3964);
and U4447 (N_4447,N_3855,N_3726);
and U4448 (N_4448,N_3675,N_3701);
xnor U4449 (N_4449,N_3662,N_3520);
xor U4450 (N_4450,N_3609,N_3602);
and U4451 (N_4451,N_3602,N_3737);
xnor U4452 (N_4452,N_3517,N_3790);
xnor U4453 (N_4453,N_3562,N_3620);
or U4454 (N_4454,N_3830,N_3934);
or U4455 (N_4455,N_3906,N_3624);
xnor U4456 (N_4456,N_3660,N_3917);
or U4457 (N_4457,N_3937,N_3562);
or U4458 (N_4458,N_3549,N_3602);
xnor U4459 (N_4459,N_3769,N_3957);
nor U4460 (N_4460,N_3688,N_3676);
nand U4461 (N_4461,N_3855,N_3806);
and U4462 (N_4462,N_3609,N_3914);
xor U4463 (N_4463,N_3694,N_3799);
or U4464 (N_4464,N_3505,N_3766);
or U4465 (N_4465,N_3882,N_3824);
and U4466 (N_4466,N_3885,N_3879);
xnor U4467 (N_4467,N_3619,N_3669);
and U4468 (N_4468,N_3805,N_3809);
or U4469 (N_4469,N_3956,N_3621);
xor U4470 (N_4470,N_3661,N_3888);
nor U4471 (N_4471,N_3953,N_3859);
xor U4472 (N_4472,N_3984,N_3506);
nor U4473 (N_4473,N_3703,N_3712);
or U4474 (N_4474,N_3595,N_3589);
xor U4475 (N_4475,N_3863,N_3848);
or U4476 (N_4476,N_3559,N_3711);
and U4477 (N_4477,N_3807,N_3826);
and U4478 (N_4478,N_3566,N_3986);
nand U4479 (N_4479,N_3980,N_3548);
and U4480 (N_4480,N_3775,N_3814);
or U4481 (N_4481,N_3873,N_3860);
nand U4482 (N_4482,N_3889,N_3817);
xor U4483 (N_4483,N_3673,N_3792);
nand U4484 (N_4484,N_3855,N_3710);
or U4485 (N_4485,N_3932,N_3885);
nor U4486 (N_4486,N_3569,N_3668);
or U4487 (N_4487,N_3781,N_3856);
and U4488 (N_4488,N_3658,N_3953);
nand U4489 (N_4489,N_3675,N_3673);
nand U4490 (N_4490,N_3999,N_3721);
nand U4491 (N_4491,N_3780,N_3748);
xor U4492 (N_4492,N_3513,N_3843);
or U4493 (N_4493,N_3584,N_3853);
or U4494 (N_4494,N_3814,N_3709);
xor U4495 (N_4495,N_3725,N_3819);
xor U4496 (N_4496,N_3537,N_3547);
and U4497 (N_4497,N_3846,N_3716);
and U4498 (N_4498,N_3653,N_3656);
xnor U4499 (N_4499,N_3643,N_3881);
and U4500 (N_4500,N_4377,N_4374);
xor U4501 (N_4501,N_4137,N_4498);
or U4502 (N_4502,N_4446,N_4259);
or U4503 (N_4503,N_4495,N_4460);
nand U4504 (N_4504,N_4131,N_4129);
xnor U4505 (N_4505,N_4272,N_4210);
nor U4506 (N_4506,N_4311,N_4300);
nand U4507 (N_4507,N_4345,N_4385);
and U4508 (N_4508,N_4242,N_4099);
nor U4509 (N_4509,N_4319,N_4497);
nor U4510 (N_4510,N_4478,N_4491);
or U4511 (N_4511,N_4083,N_4364);
nor U4512 (N_4512,N_4287,N_4053);
nor U4513 (N_4513,N_4321,N_4040);
or U4514 (N_4514,N_4017,N_4176);
and U4515 (N_4515,N_4089,N_4472);
nor U4516 (N_4516,N_4250,N_4270);
xor U4517 (N_4517,N_4235,N_4239);
nor U4518 (N_4518,N_4241,N_4370);
and U4519 (N_4519,N_4494,N_4014);
xnor U4520 (N_4520,N_4119,N_4147);
xor U4521 (N_4521,N_4171,N_4245);
nor U4522 (N_4522,N_4430,N_4406);
nor U4523 (N_4523,N_4379,N_4409);
nor U4524 (N_4524,N_4094,N_4304);
or U4525 (N_4525,N_4429,N_4323);
or U4526 (N_4526,N_4227,N_4400);
and U4527 (N_4527,N_4452,N_4246);
nand U4528 (N_4528,N_4381,N_4023);
nand U4529 (N_4529,N_4067,N_4393);
and U4530 (N_4530,N_4059,N_4139);
nand U4531 (N_4531,N_4154,N_4013);
nand U4532 (N_4532,N_4228,N_4063);
or U4533 (N_4533,N_4499,N_4149);
and U4534 (N_4534,N_4222,N_4218);
or U4535 (N_4535,N_4148,N_4316);
nor U4536 (N_4536,N_4141,N_4009);
or U4537 (N_4537,N_4484,N_4026);
xnor U4538 (N_4538,N_4344,N_4203);
or U4539 (N_4539,N_4248,N_4126);
nor U4540 (N_4540,N_4461,N_4180);
or U4541 (N_4541,N_4096,N_4035);
xnor U4542 (N_4542,N_4268,N_4281);
nor U4543 (N_4543,N_4032,N_4288);
nand U4544 (N_4544,N_4056,N_4209);
or U4545 (N_4545,N_4380,N_4293);
nor U4546 (N_4546,N_4136,N_4240);
and U4547 (N_4547,N_4016,N_4237);
and U4548 (N_4548,N_4284,N_4052);
nor U4549 (N_4549,N_4045,N_4388);
and U4550 (N_4550,N_4006,N_4042);
and U4551 (N_4551,N_4334,N_4039);
nand U4552 (N_4552,N_4010,N_4041);
nor U4553 (N_4553,N_4152,N_4140);
nor U4554 (N_4554,N_4118,N_4394);
and U4555 (N_4555,N_4111,N_4443);
or U4556 (N_4556,N_4213,N_4313);
xnor U4557 (N_4557,N_4405,N_4146);
and U4558 (N_4558,N_4093,N_4315);
or U4559 (N_4559,N_4266,N_4301);
or U4560 (N_4560,N_4269,N_4358);
nand U4561 (N_4561,N_4327,N_4464);
or U4562 (N_4562,N_4437,N_4167);
and U4563 (N_4563,N_4490,N_4106);
xor U4564 (N_4564,N_4387,N_4392);
and U4565 (N_4565,N_4476,N_4422);
xor U4566 (N_4566,N_4352,N_4351);
and U4567 (N_4567,N_4256,N_4424);
and U4568 (N_4568,N_4350,N_4465);
nor U4569 (N_4569,N_4254,N_4261);
nor U4570 (N_4570,N_4123,N_4453);
and U4571 (N_4571,N_4114,N_4399);
and U4572 (N_4572,N_4427,N_4031);
xnor U4573 (N_4573,N_4027,N_4365);
and U4574 (N_4574,N_4419,N_4279);
or U4575 (N_4575,N_4221,N_4277);
and U4576 (N_4576,N_4286,N_4356);
and U4577 (N_4577,N_4322,N_4265);
or U4578 (N_4578,N_4189,N_4431);
and U4579 (N_4579,N_4410,N_4463);
nand U4580 (N_4580,N_4208,N_4175);
and U4581 (N_4581,N_4054,N_4320);
or U4582 (N_4582,N_4366,N_4130);
nand U4583 (N_4583,N_4474,N_4193);
nor U4584 (N_4584,N_4011,N_4197);
or U4585 (N_4585,N_4361,N_4001);
xnor U4586 (N_4586,N_4191,N_4283);
xnor U4587 (N_4587,N_4244,N_4211);
nand U4588 (N_4588,N_4173,N_4289);
nor U4589 (N_4589,N_4090,N_4325);
and U4590 (N_4590,N_4165,N_4195);
nor U4591 (N_4591,N_4048,N_4481);
xnor U4592 (N_4592,N_4135,N_4003);
nand U4593 (N_4593,N_4447,N_4134);
nor U4594 (N_4594,N_4473,N_4426);
or U4595 (N_4595,N_4216,N_4187);
and U4596 (N_4596,N_4348,N_4445);
nor U4597 (N_4597,N_4024,N_4095);
nand U4598 (N_4598,N_4204,N_4368);
and U4599 (N_4599,N_4012,N_4098);
and U4600 (N_4600,N_4488,N_4205);
or U4601 (N_4601,N_4360,N_4333);
and U4602 (N_4602,N_4212,N_4477);
or U4603 (N_4603,N_4456,N_4029);
and U4604 (N_4604,N_4404,N_4375);
nor U4605 (N_4605,N_4415,N_4150);
nor U4606 (N_4606,N_4231,N_4076);
nand U4607 (N_4607,N_4182,N_4030);
xnor U4608 (N_4608,N_4233,N_4071);
and U4609 (N_4609,N_4072,N_4019);
nor U4610 (N_4610,N_4372,N_4143);
xor U4611 (N_4611,N_4338,N_4417);
nor U4612 (N_4612,N_4483,N_4201);
or U4613 (N_4613,N_4021,N_4274);
and U4614 (N_4614,N_4341,N_4047);
nor U4615 (N_4615,N_4342,N_4036);
nor U4616 (N_4616,N_4324,N_4060);
nor U4617 (N_4617,N_4064,N_4022);
or U4618 (N_4618,N_4421,N_4234);
xnor U4619 (N_4619,N_4184,N_4294);
and U4620 (N_4620,N_4340,N_4117);
nor U4621 (N_4621,N_4020,N_4258);
or U4622 (N_4622,N_4183,N_4363);
nor U4623 (N_4623,N_4467,N_4088);
xor U4624 (N_4624,N_4077,N_4262);
nand U4625 (N_4625,N_4051,N_4159);
and U4626 (N_4626,N_4223,N_4252);
nand U4627 (N_4627,N_4196,N_4219);
and U4628 (N_4628,N_4391,N_4110);
or U4629 (N_4629,N_4296,N_4309);
nand U4630 (N_4630,N_4257,N_4260);
and U4631 (N_4631,N_4492,N_4378);
xnor U4632 (N_4632,N_4493,N_4178);
nand U4633 (N_4633,N_4448,N_4438);
nand U4634 (N_4634,N_4367,N_4037);
nor U4635 (N_4635,N_4226,N_4275);
and U4636 (N_4636,N_4194,N_4157);
nand U4637 (N_4637,N_4395,N_4335);
or U4638 (N_4638,N_4075,N_4362);
xor U4639 (N_4639,N_4263,N_4229);
nand U4640 (N_4640,N_4232,N_4058);
nor U4641 (N_4641,N_4128,N_4408);
xor U4642 (N_4642,N_4120,N_4105);
nand U4643 (N_4643,N_4074,N_4202);
xnor U4644 (N_4644,N_4068,N_4065);
and U4645 (N_4645,N_4225,N_4423);
nand U4646 (N_4646,N_4444,N_4236);
nor U4647 (N_4647,N_4049,N_4170);
and U4648 (N_4648,N_4133,N_4081);
xor U4649 (N_4649,N_4185,N_4138);
nand U4650 (N_4650,N_4336,N_4145);
nand U4651 (N_4651,N_4092,N_4331);
and U4652 (N_4652,N_4057,N_4162);
nor U4653 (N_4653,N_4109,N_4295);
nor U4654 (N_4654,N_4034,N_4355);
nand U4655 (N_4655,N_4050,N_4144);
and U4656 (N_4656,N_4207,N_4471);
nand U4657 (N_4657,N_4346,N_4326);
xnor U4658 (N_4658,N_4329,N_4200);
nand U4659 (N_4659,N_4086,N_4121);
xnor U4660 (N_4660,N_4046,N_4310);
or U4661 (N_4661,N_4418,N_4238);
nand U4662 (N_4662,N_4115,N_4425);
nor U4663 (N_4663,N_4407,N_4215);
or U4664 (N_4664,N_4290,N_4302);
xor U4665 (N_4665,N_4280,N_4397);
nor U4666 (N_4666,N_4084,N_4091);
and U4667 (N_4667,N_4468,N_4420);
nand U4668 (N_4668,N_4396,N_4044);
or U4669 (N_4669,N_4299,N_4008);
xnor U4670 (N_4670,N_4217,N_4199);
xor U4671 (N_4671,N_4179,N_4282);
nand U4672 (N_4672,N_4442,N_4125);
or U4673 (N_4673,N_4354,N_4061);
nand U4674 (N_4674,N_4318,N_4455);
and U4675 (N_4675,N_4043,N_4033);
nand U4676 (N_4676,N_4398,N_4369);
or U4677 (N_4677,N_4155,N_4038);
nand U4678 (N_4678,N_4163,N_4332);
xor U4679 (N_4679,N_4271,N_4402);
or U4680 (N_4680,N_4214,N_4192);
nand U4681 (N_4681,N_4186,N_4161);
and U4682 (N_4682,N_4434,N_4103);
xor U4683 (N_4683,N_4018,N_4314);
nor U4684 (N_4684,N_4097,N_4328);
nand U4685 (N_4685,N_4383,N_4062);
nand U4686 (N_4686,N_4004,N_4306);
and U4687 (N_4687,N_4172,N_4116);
nand U4688 (N_4688,N_4458,N_4411);
nor U4689 (N_4689,N_4087,N_4108);
nor U4690 (N_4690,N_4292,N_4247);
xnor U4691 (N_4691,N_4353,N_4104);
nor U4692 (N_4692,N_4401,N_4132);
nor U4693 (N_4693,N_4337,N_4188);
nand U4694 (N_4694,N_4230,N_4428);
xnor U4695 (N_4695,N_4220,N_4475);
xnor U4696 (N_4696,N_4439,N_4079);
nand U4697 (N_4697,N_4459,N_4078);
xor U4698 (N_4698,N_4169,N_4181);
nand U4699 (N_4699,N_4317,N_4376);
nand U4700 (N_4700,N_4486,N_4454);
nand U4701 (N_4701,N_4413,N_4112);
nor U4702 (N_4702,N_4082,N_4305);
nand U4703 (N_4703,N_4470,N_4384);
nor U4704 (N_4704,N_4278,N_4449);
nor U4705 (N_4705,N_4005,N_4206);
xnor U4706 (N_4706,N_4291,N_4451);
nand U4707 (N_4707,N_4479,N_4276);
xnor U4708 (N_4708,N_4466,N_4142);
xnor U4709 (N_4709,N_4382,N_4253);
or U4710 (N_4710,N_4267,N_4158);
nand U4711 (N_4711,N_4264,N_4168);
and U4712 (N_4712,N_4462,N_4085);
nand U4713 (N_4713,N_4330,N_4174);
xnor U4714 (N_4714,N_4339,N_4070);
and U4715 (N_4715,N_4440,N_4273);
nor U4716 (N_4716,N_4343,N_4435);
xnor U4717 (N_4717,N_4100,N_4285);
or U4718 (N_4718,N_4482,N_4243);
nor U4719 (N_4719,N_4403,N_4113);
xnor U4720 (N_4720,N_4166,N_4312);
nand U4721 (N_4721,N_4457,N_4000);
and U4722 (N_4722,N_4297,N_4389);
xor U4723 (N_4723,N_4055,N_4007);
nor U4724 (N_4724,N_4066,N_4101);
and U4725 (N_4725,N_4496,N_4102);
xor U4726 (N_4726,N_4432,N_4414);
or U4727 (N_4727,N_4124,N_4107);
xor U4728 (N_4728,N_4489,N_4177);
and U4729 (N_4729,N_4357,N_4251);
nor U4730 (N_4730,N_4015,N_4436);
or U4731 (N_4731,N_4480,N_4469);
and U4732 (N_4732,N_4127,N_4156);
nor U4733 (N_4733,N_4069,N_4347);
nor U4734 (N_4734,N_4160,N_4028);
xor U4735 (N_4735,N_4122,N_4249);
or U4736 (N_4736,N_4359,N_4298);
nor U4737 (N_4737,N_4487,N_4416);
and U4738 (N_4738,N_4080,N_4224);
xor U4739 (N_4739,N_4025,N_4190);
nor U4740 (N_4740,N_4255,N_4198);
xnor U4741 (N_4741,N_4450,N_4349);
and U4742 (N_4742,N_4308,N_4164);
nor U4743 (N_4743,N_4151,N_4441);
or U4744 (N_4744,N_4412,N_4153);
nor U4745 (N_4745,N_4307,N_4485);
and U4746 (N_4746,N_4002,N_4371);
nand U4747 (N_4747,N_4373,N_4390);
nor U4748 (N_4748,N_4386,N_4433);
nor U4749 (N_4749,N_4303,N_4073);
and U4750 (N_4750,N_4380,N_4078);
nor U4751 (N_4751,N_4238,N_4345);
nand U4752 (N_4752,N_4295,N_4306);
and U4753 (N_4753,N_4041,N_4478);
xnor U4754 (N_4754,N_4200,N_4012);
nand U4755 (N_4755,N_4357,N_4417);
or U4756 (N_4756,N_4240,N_4043);
and U4757 (N_4757,N_4017,N_4138);
nor U4758 (N_4758,N_4281,N_4438);
nor U4759 (N_4759,N_4032,N_4237);
and U4760 (N_4760,N_4262,N_4302);
nand U4761 (N_4761,N_4152,N_4096);
nor U4762 (N_4762,N_4067,N_4498);
or U4763 (N_4763,N_4158,N_4208);
or U4764 (N_4764,N_4264,N_4267);
nand U4765 (N_4765,N_4380,N_4393);
and U4766 (N_4766,N_4459,N_4109);
and U4767 (N_4767,N_4486,N_4097);
nand U4768 (N_4768,N_4314,N_4115);
and U4769 (N_4769,N_4127,N_4270);
nand U4770 (N_4770,N_4242,N_4104);
nand U4771 (N_4771,N_4458,N_4442);
nor U4772 (N_4772,N_4117,N_4461);
and U4773 (N_4773,N_4085,N_4286);
or U4774 (N_4774,N_4325,N_4080);
xnor U4775 (N_4775,N_4344,N_4264);
and U4776 (N_4776,N_4110,N_4155);
and U4777 (N_4777,N_4221,N_4132);
and U4778 (N_4778,N_4447,N_4196);
and U4779 (N_4779,N_4092,N_4390);
or U4780 (N_4780,N_4291,N_4415);
nand U4781 (N_4781,N_4402,N_4105);
nand U4782 (N_4782,N_4366,N_4458);
and U4783 (N_4783,N_4172,N_4067);
or U4784 (N_4784,N_4349,N_4294);
nor U4785 (N_4785,N_4209,N_4484);
nand U4786 (N_4786,N_4349,N_4391);
xor U4787 (N_4787,N_4490,N_4113);
xor U4788 (N_4788,N_4209,N_4224);
nand U4789 (N_4789,N_4071,N_4052);
or U4790 (N_4790,N_4344,N_4265);
or U4791 (N_4791,N_4265,N_4496);
nand U4792 (N_4792,N_4422,N_4413);
xnor U4793 (N_4793,N_4406,N_4426);
nand U4794 (N_4794,N_4072,N_4125);
or U4795 (N_4795,N_4461,N_4416);
and U4796 (N_4796,N_4066,N_4495);
or U4797 (N_4797,N_4081,N_4057);
xor U4798 (N_4798,N_4463,N_4297);
xnor U4799 (N_4799,N_4022,N_4455);
or U4800 (N_4800,N_4190,N_4493);
nand U4801 (N_4801,N_4355,N_4052);
nor U4802 (N_4802,N_4029,N_4260);
and U4803 (N_4803,N_4324,N_4355);
or U4804 (N_4804,N_4489,N_4208);
nor U4805 (N_4805,N_4314,N_4034);
xnor U4806 (N_4806,N_4370,N_4108);
nand U4807 (N_4807,N_4053,N_4058);
nand U4808 (N_4808,N_4499,N_4266);
nand U4809 (N_4809,N_4479,N_4231);
nor U4810 (N_4810,N_4111,N_4278);
nand U4811 (N_4811,N_4051,N_4372);
nor U4812 (N_4812,N_4302,N_4195);
or U4813 (N_4813,N_4031,N_4448);
and U4814 (N_4814,N_4278,N_4465);
nand U4815 (N_4815,N_4342,N_4287);
nand U4816 (N_4816,N_4188,N_4393);
or U4817 (N_4817,N_4308,N_4493);
or U4818 (N_4818,N_4469,N_4247);
nand U4819 (N_4819,N_4356,N_4215);
nor U4820 (N_4820,N_4422,N_4167);
xor U4821 (N_4821,N_4301,N_4300);
nand U4822 (N_4822,N_4228,N_4020);
and U4823 (N_4823,N_4342,N_4253);
nor U4824 (N_4824,N_4061,N_4054);
xor U4825 (N_4825,N_4275,N_4245);
or U4826 (N_4826,N_4445,N_4005);
nand U4827 (N_4827,N_4472,N_4378);
xor U4828 (N_4828,N_4090,N_4119);
and U4829 (N_4829,N_4298,N_4284);
and U4830 (N_4830,N_4350,N_4364);
nor U4831 (N_4831,N_4001,N_4305);
xor U4832 (N_4832,N_4331,N_4193);
and U4833 (N_4833,N_4453,N_4265);
xnor U4834 (N_4834,N_4294,N_4350);
nand U4835 (N_4835,N_4112,N_4025);
xor U4836 (N_4836,N_4281,N_4300);
nand U4837 (N_4837,N_4113,N_4112);
or U4838 (N_4838,N_4413,N_4433);
nor U4839 (N_4839,N_4365,N_4008);
nor U4840 (N_4840,N_4403,N_4006);
xor U4841 (N_4841,N_4307,N_4327);
nand U4842 (N_4842,N_4219,N_4222);
and U4843 (N_4843,N_4033,N_4180);
xnor U4844 (N_4844,N_4454,N_4253);
or U4845 (N_4845,N_4164,N_4050);
or U4846 (N_4846,N_4283,N_4480);
and U4847 (N_4847,N_4173,N_4444);
and U4848 (N_4848,N_4106,N_4398);
or U4849 (N_4849,N_4256,N_4248);
or U4850 (N_4850,N_4321,N_4188);
and U4851 (N_4851,N_4267,N_4142);
and U4852 (N_4852,N_4428,N_4345);
or U4853 (N_4853,N_4090,N_4045);
and U4854 (N_4854,N_4389,N_4458);
nor U4855 (N_4855,N_4111,N_4264);
nor U4856 (N_4856,N_4038,N_4229);
and U4857 (N_4857,N_4407,N_4398);
nor U4858 (N_4858,N_4141,N_4330);
nor U4859 (N_4859,N_4037,N_4145);
and U4860 (N_4860,N_4403,N_4031);
and U4861 (N_4861,N_4477,N_4329);
or U4862 (N_4862,N_4418,N_4321);
or U4863 (N_4863,N_4291,N_4412);
xnor U4864 (N_4864,N_4330,N_4222);
xor U4865 (N_4865,N_4168,N_4092);
or U4866 (N_4866,N_4321,N_4035);
nor U4867 (N_4867,N_4474,N_4419);
or U4868 (N_4868,N_4354,N_4248);
nand U4869 (N_4869,N_4253,N_4034);
nand U4870 (N_4870,N_4497,N_4013);
and U4871 (N_4871,N_4138,N_4426);
nand U4872 (N_4872,N_4367,N_4035);
nor U4873 (N_4873,N_4329,N_4451);
and U4874 (N_4874,N_4137,N_4080);
xor U4875 (N_4875,N_4406,N_4303);
nand U4876 (N_4876,N_4253,N_4053);
xor U4877 (N_4877,N_4154,N_4094);
xor U4878 (N_4878,N_4476,N_4481);
nor U4879 (N_4879,N_4124,N_4434);
or U4880 (N_4880,N_4096,N_4192);
nand U4881 (N_4881,N_4483,N_4004);
nand U4882 (N_4882,N_4393,N_4223);
or U4883 (N_4883,N_4245,N_4268);
nand U4884 (N_4884,N_4437,N_4448);
nor U4885 (N_4885,N_4460,N_4285);
xnor U4886 (N_4886,N_4491,N_4240);
and U4887 (N_4887,N_4439,N_4482);
or U4888 (N_4888,N_4130,N_4224);
nor U4889 (N_4889,N_4254,N_4330);
xnor U4890 (N_4890,N_4192,N_4465);
or U4891 (N_4891,N_4194,N_4185);
xor U4892 (N_4892,N_4189,N_4342);
xor U4893 (N_4893,N_4469,N_4437);
nor U4894 (N_4894,N_4456,N_4000);
xnor U4895 (N_4895,N_4151,N_4478);
and U4896 (N_4896,N_4157,N_4050);
or U4897 (N_4897,N_4140,N_4489);
nor U4898 (N_4898,N_4093,N_4139);
and U4899 (N_4899,N_4258,N_4022);
nand U4900 (N_4900,N_4214,N_4082);
xor U4901 (N_4901,N_4016,N_4360);
nor U4902 (N_4902,N_4212,N_4127);
xnor U4903 (N_4903,N_4415,N_4155);
nor U4904 (N_4904,N_4493,N_4298);
nor U4905 (N_4905,N_4061,N_4318);
nand U4906 (N_4906,N_4260,N_4418);
nand U4907 (N_4907,N_4404,N_4365);
and U4908 (N_4908,N_4142,N_4094);
and U4909 (N_4909,N_4128,N_4456);
nand U4910 (N_4910,N_4281,N_4291);
xor U4911 (N_4911,N_4468,N_4368);
nor U4912 (N_4912,N_4062,N_4002);
or U4913 (N_4913,N_4133,N_4354);
or U4914 (N_4914,N_4271,N_4253);
nand U4915 (N_4915,N_4169,N_4078);
xnor U4916 (N_4916,N_4469,N_4200);
xnor U4917 (N_4917,N_4019,N_4347);
nand U4918 (N_4918,N_4474,N_4381);
nor U4919 (N_4919,N_4357,N_4149);
xnor U4920 (N_4920,N_4175,N_4200);
and U4921 (N_4921,N_4093,N_4044);
or U4922 (N_4922,N_4494,N_4186);
or U4923 (N_4923,N_4067,N_4218);
nor U4924 (N_4924,N_4196,N_4434);
xor U4925 (N_4925,N_4102,N_4456);
xnor U4926 (N_4926,N_4208,N_4497);
and U4927 (N_4927,N_4268,N_4095);
nor U4928 (N_4928,N_4193,N_4228);
or U4929 (N_4929,N_4073,N_4173);
nor U4930 (N_4930,N_4168,N_4336);
nand U4931 (N_4931,N_4171,N_4004);
nor U4932 (N_4932,N_4445,N_4282);
nor U4933 (N_4933,N_4301,N_4149);
nor U4934 (N_4934,N_4130,N_4333);
xnor U4935 (N_4935,N_4000,N_4460);
nor U4936 (N_4936,N_4331,N_4018);
or U4937 (N_4937,N_4490,N_4135);
nand U4938 (N_4938,N_4215,N_4231);
or U4939 (N_4939,N_4081,N_4358);
nor U4940 (N_4940,N_4286,N_4023);
or U4941 (N_4941,N_4304,N_4453);
nor U4942 (N_4942,N_4350,N_4485);
or U4943 (N_4943,N_4338,N_4091);
nor U4944 (N_4944,N_4292,N_4015);
or U4945 (N_4945,N_4408,N_4243);
or U4946 (N_4946,N_4013,N_4113);
nor U4947 (N_4947,N_4168,N_4247);
nor U4948 (N_4948,N_4363,N_4098);
and U4949 (N_4949,N_4289,N_4372);
or U4950 (N_4950,N_4115,N_4427);
and U4951 (N_4951,N_4317,N_4304);
xor U4952 (N_4952,N_4133,N_4003);
xnor U4953 (N_4953,N_4299,N_4104);
or U4954 (N_4954,N_4068,N_4441);
and U4955 (N_4955,N_4454,N_4132);
and U4956 (N_4956,N_4015,N_4117);
xnor U4957 (N_4957,N_4483,N_4097);
xor U4958 (N_4958,N_4104,N_4340);
xor U4959 (N_4959,N_4442,N_4118);
xnor U4960 (N_4960,N_4370,N_4185);
nor U4961 (N_4961,N_4007,N_4307);
nor U4962 (N_4962,N_4283,N_4393);
or U4963 (N_4963,N_4354,N_4081);
or U4964 (N_4964,N_4396,N_4354);
xnor U4965 (N_4965,N_4035,N_4146);
nand U4966 (N_4966,N_4376,N_4128);
or U4967 (N_4967,N_4427,N_4047);
nor U4968 (N_4968,N_4206,N_4125);
or U4969 (N_4969,N_4092,N_4335);
nor U4970 (N_4970,N_4316,N_4162);
xor U4971 (N_4971,N_4497,N_4086);
nor U4972 (N_4972,N_4151,N_4300);
or U4973 (N_4973,N_4240,N_4202);
nor U4974 (N_4974,N_4101,N_4002);
or U4975 (N_4975,N_4271,N_4032);
nand U4976 (N_4976,N_4166,N_4474);
or U4977 (N_4977,N_4198,N_4205);
nand U4978 (N_4978,N_4342,N_4350);
or U4979 (N_4979,N_4069,N_4222);
nand U4980 (N_4980,N_4339,N_4075);
and U4981 (N_4981,N_4027,N_4354);
xnor U4982 (N_4982,N_4402,N_4414);
or U4983 (N_4983,N_4146,N_4178);
nor U4984 (N_4984,N_4272,N_4143);
nor U4985 (N_4985,N_4139,N_4057);
and U4986 (N_4986,N_4146,N_4261);
or U4987 (N_4987,N_4371,N_4239);
nor U4988 (N_4988,N_4074,N_4046);
nand U4989 (N_4989,N_4426,N_4144);
or U4990 (N_4990,N_4032,N_4030);
or U4991 (N_4991,N_4396,N_4372);
nand U4992 (N_4992,N_4496,N_4061);
xnor U4993 (N_4993,N_4066,N_4412);
nand U4994 (N_4994,N_4065,N_4028);
nand U4995 (N_4995,N_4459,N_4096);
xor U4996 (N_4996,N_4461,N_4347);
and U4997 (N_4997,N_4047,N_4123);
nor U4998 (N_4998,N_4284,N_4185);
xnor U4999 (N_4999,N_4387,N_4027);
xor U5000 (N_5000,N_4500,N_4659);
nand U5001 (N_5001,N_4505,N_4936);
nand U5002 (N_5002,N_4653,N_4600);
nand U5003 (N_5003,N_4999,N_4805);
or U5004 (N_5004,N_4515,N_4526);
nor U5005 (N_5005,N_4713,N_4888);
nor U5006 (N_5006,N_4767,N_4572);
or U5007 (N_5007,N_4915,N_4528);
xor U5008 (N_5008,N_4913,N_4903);
and U5009 (N_5009,N_4670,N_4972);
nor U5010 (N_5010,N_4556,N_4871);
nand U5011 (N_5011,N_4583,N_4587);
nor U5012 (N_5012,N_4926,N_4584);
and U5013 (N_5013,N_4588,N_4763);
nor U5014 (N_5014,N_4567,N_4890);
and U5015 (N_5015,N_4754,N_4944);
or U5016 (N_5016,N_4712,N_4739);
nor U5017 (N_5017,N_4859,N_4563);
and U5018 (N_5018,N_4828,N_4909);
and U5019 (N_5019,N_4733,N_4994);
xor U5020 (N_5020,N_4882,N_4823);
nand U5021 (N_5021,N_4970,N_4801);
nor U5022 (N_5022,N_4605,N_4854);
xor U5023 (N_5023,N_4656,N_4917);
xor U5024 (N_5024,N_4965,N_4824);
nor U5025 (N_5025,N_4503,N_4596);
or U5026 (N_5026,N_4595,N_4960);
nor U5027 (N_5027,N_4535,N_4937);
nor U5028 (N_5028,N_4662,N_4778);
or U5029 (N_5029,N_4895,N_4790);
xor U5030 (N_5030,N_4615,N_4947);
nor U5031 (N_5031,N_4579,N_4610);
and U5032 (N_5032,N_4984,N_4938);
nor U5033 (N_5033,N_4773,N_4996);
and U5034 (N_5034,N_4811,N_4644);
nor U5035 (N_5035,N_4699,N_4869);
or U5036 (N_5036,N_4682,N_4919);
nor U5037 (N_5037,N_4930,N_4951);
xor U5038 (N_5038,N_4918,N_4940);
and U5039 (N_5039,N_4848,N_4537);
nand U5040 (N_5040,N_4525,N_4867);
nor U5041 (N_5041,N_4732,N_4643);
xnor U5042 (N_5042,N_4751,N_4845);
or U5043 (N_5043,N_4927,N_4928);
and U5044 (N_5044,N_4561,N_4623);
or U5045 (N_5045,N_4898,N_4568);
and U5046 (N_5046,N_4673,N_4973);
nor U5047 (N_5047,N_4706,N_4806);
or U5048 (N_5048,N_4862,N_4619);
xor U5049 (N_5049,N_4983,N_4648);
or U5050 (N_5050,N_4813,N_4880);
and U5051 (N_5051,N_4669,N_4672);
nor U5052 (N_5052,N_4746,N_4730);
and U5053 (N_5053,N_4594,N_4769);
nor U5054 (N_5054,N_4607,N_4993);
or U5055 (N_5055,N_4681,N_4818);
xor U5056 (N_5056,N_4814,N_4786);
nand U5057 (N_5057,N_4873,N_4618);
nand U5058 (N_5058,N_4765,N_4860);
nand U5059 (N_5059,N_4711,N_4633);
and U5060 (N_5060,N_4566,N_4534);
xnor U5061 (N_5061,N_4943,N_4830);
and U5062 (N_5062,N_4516,N_4784);
and U5063 (N_5063,N_4838,N_4597);
xnor U5064 (N_5064,N_4837,N_4952);
and U5065 (N_5065,N_4635,N_4771);
nand U5066 (N_5066,N_4536,N_4731);
nor U5067 (N_5067,N_4622,N_4742);
nor U5068 (N_5068,N_4961,N_4586);
or U5069 (N_5069,N_4887,N_4866);
xnor U5070 (N_5070,N_4690,N_4589);
or U5071 (N_5071,N_4708,N_4719);
xnor U5072 (N_5072,N_4743,N_4604);
or U5073 (N_5073,N_4570,N_4571);
xnor U5074 (N_5074,N_4950,N_4908);
nor U5075 (N_5075,N_4655,N_4901);
nand U5076 (N_5076,N_4522,N_4668);
xor U5077 (N_5077,N_4501,N_4540);
xnor U5078 (N_5078,N_4693,N_4544);
nand U5079 (N_5079,N_4781,N_4512);
nand U5080 (N_5080,N_4759,N_4585);
or U5081 (N_5081,N_4761,N_4510);
nand U5082 (N_5082,N_4612,N_4720);
xor U5083 (N_5083,N_4795,N_4640);
or U5084 (N_5084,N_4803,N_4636);
nand U5085 (N_5085,N_4911,N_4638);
xnor U5086 (N_5086,N_4735,N_4822);
nor U5087 (N_5087,N_4554,N_4722);
or U5088 (N_5088,N_4630,N_4709);
and U5089 (N_5089,N_4639,N_4542);
xor U5090 (N_5090,N_4920,N_4645);
or U5091 (N_5091,N_4617,N_4889);
nand U5092 (N_5092,N_4582,N_4881);
and U5093 (N_5093,N_4573,N_4502);
xor U5094 (N_5094,N_4817,N_4667);
nand U5095 (N_5095,N_4923,N_4691);
nand U5096 (N_5096,N_4853,N_4529);
and U5097 (N_5097,N_4997,N_4578);
nor U5098 (N_5098,N_4509,N_4872);
xor U5099 (N_5099,N_4728,N_4674);
nand U5100 (N_5100,N_4524,N_4948);
nand U5101 (N_5101,N_4995,N_4629);
xnor U5102 (N_5102,N_4552,N_4543);
xor U5103 (N_5103,N_4902,N_4760);
nand U5104 (N_5104,N_4885,N_4555);
xnor U5105 (N_5105,N_4967,N_4701);
and U5106 (N_5106,N_4721,N_4675);
and U5107 (N_5107,N_4812,N_4646);
xor U5108 (N_5108,N_4998,N_4593);
and U5109 (N_5109,N_4804,N_4521);
or U5110 (N_5110,N_4870,N_4530);
nor U5111 (N_5111,N_4832,N_4959);
xor U5112 (N_5112,N_4560,N_4748);
xnor U5113 (N_5113,N_4513,N_4694);
xnor U5114 (N_5114,N_4991,N_4851);
xnor U5115 (N_5115,N_4608,N_4780);
and U5116 (N_5116,N_4986,N_4798);
nor U5117 (N_5117,N_4546,N_4858);
nand U5118 (N_5118,N_4929,N_4657);
and U5119 (N_5119,N_4789,N_4723);
or U5120 (N_5120,N_4800,N_4856);
or U5121 (N_5121,N_4797,N_4963);
nor U5122 (N_5122,N_4831,N_4852);
and U5123 (N_5123,N_4686,N_4627);
or U5124 (N_5124,N_4621,N_4508);
nand U5125 (N_5125,N_4632,N_4504);
xor U5126 (N_5126,N_4857,N_4794);
nand U5127 (N_5127,N_4968,N_4978);
nand U5128 (N_5128,N_4520,N_4793);
nand U5129 (N_5129,N_4785,N_4792);
nand U5130 (N_5130,N_4865,N_4985);
xnor U5131 (N_5131,N_4874,N_4647);
nor U5132 (N_5132,N_4905,N_4533);
and U5133 (N_5133,N_4863,N_4727);
nand U5134 (N_5134,N_4819,N_4698);
xnor U5135 (N_5135,N_4922,N_4976);
nor U5136 (N_5136,N_4982,N_4841);
and U5137 (N_5137,N_4899,N_4807);
nor U5138 (N_5138,N_4749,N_4791);
nor U5139 (N_5139,N_4879,N_4966);
or U5140 (N_5140,N_4652,N_4599);
nor U5141 (N_5141,N_4736,N_4710);
xnor U5142 (N_5142,N_4833,N_4527);
nand U5143 (N_5143,N_4631,N_4897);
and U5144 (N_5144,N_4900,N_4684);
nor U5145 (N_5145,N_4810,N_4697);
and U5146 (N_5146,N_4741,N_4772);
and U5147 (N_5147,N_4839,N_4574);
and U5148 (N_5148,N_4715,N_4755);
nand U5149 (N_5149,N_4601,N_4849);
or U5150 (N_5150,N_4962,N_4843);
nand U5151 (N_5151,N_4891,N_4921);
xnor U5152 (N_5152,N_4569,N_4842);
xnor U5153 (N_5153,N_4990,N_4725);
xnor U5154 (N_5154,N_4689,N_4868);
or U5155 (N_5155,N_4992,N_4893);
or U5156 (N_5156,N_4906,N_4924);
and U5157 (N_5157,N_4934,N_4768);
nor U5158 (N_5158,N_4641,N_4775);
and U5159 (N_5159,N_4611,N_4762);
or U5160 (N_5160,N_4980,N_4606);
or U5161 (N_5161,N_4642,N_4941);
and U5162 (N_5162,N_4981,N_4703);
xor U5163 (N_5163,N_4931,N_4955);
and U5164 (N_5164,N_4676,N_4511);
xnor U5165 (N_5165,N_4756,N_4679);
nand U5166 (N_5166,N_4977,N_4942);
nor U5167 (N_5167,N_4827,N_4557);
or U5168 (N_5168,N_4989,N_4916);
nand U5169 (N_5169,N_4577,N_4750);
xor U5170 (N_5170,N_4753,N_4687);
nor U5171 (N_5171,N_4799,N_4660);
or U5172 (N_5172,N_4576,N_4957);
nor U5173 (N_5173,N_4883,N_4592);
nand U5174 (N_5174,N_4783,N_4816);
and U5175 (N_5175,N_4726,N_4558);
or U5176 (N_5176,N_4663,N_4809);
nor U5177 (N_5177,N_4729,N_4704);
nor U5178 (N_5178,N_4892,N_4815);
or U5179 (N_5179,N_4825,N_4779);
nor U5180 (N_5180,N_4696,N_4766);
and U5181 (N_5181,N_4737,N_4764);
nor U5182 (N_5182,N_4724,N_4747);
and U5183 (N_5183,N_4734,N_4796);
and U5184 (N_5184,N_4683,N_4626);
nand U5185 (N_5185,N_4770,N_4802);
nand U5186 (N_5186,N_4575,N_4717);
and U5187 (N_5187,N_4884,N_4894);
xor U5188 (N_5188,N_4776,N_4846);
nand U5189 (N_5189,N_4666,N_4532);
xnor U5190 (N_5190,N_4878,N_4861);
or U5191 (N_5191,N_4548,N_4598);
or U5192 (N_5192,N_4547,N_4840);
xor U5193 (N_5193,N_4954,N_4688);
nand U5194 (N_5194,N_4620,N_4877);
nand U5195 (N_5195,N_4519,N_4692);
and U5196 (N_5196,N_4820,N_4650);
xnor U5197 (N_5197,N_4559,N_4616);
and U5198 (N_5198,N_4700,N_4506);
nand U5199 (N_5199,N_4651,N_4671);
or U5200 (N_5200,N_4949,N_4553);
and U5201 (N_5201,N_4680,N_4539);
nor U5202 (N_5202,N_4896,N_4603);
nor U5203 (N_5203,N_4538,N_4945);
or U5204 (N_5204,N_4514,N_4581);
nand U5205 (N_5205,N_4987,N_4609);
nor U5206 (N_5206,N_4912,N_4550);
and U5207 (N_5207,N_4562,N_4757);
or U5208 (N_5208,N_4958,N_4718);
xnor U5209 (N_5209,N_4971,N_4834);
nor U5210 (N_5210,N_4507,N_4740);
nand U5211 (N_5211,N_4695,N_4886);
or U5212 (N_5212,N_4614,N_4602);
nand U5213 (N_5213,N_4932,N_4752);
and U5214 (N_5214,N_4774,N_4613);
and U5215 (N_5215,N_4975,N_4551);
nor U5216 (N_5216,N_4744,N_4517);
nand U5217 (N_5217,N_4714,N_4829);
nor U5218 (N_5218,N_4565,N_4836);
nor U5219 (N_5219,N_4545,N_4591);
nor U5220 (N_5220,N_4624,N_4678);
or U5221 (N_5221,N_4531,N_4661);
and U5222 (N_5222,N_4988,N_4523);
nand U5223 (N_5223,N_4541,N_4518);
nand U5224 (N_5224,N_4956,N_4549);
or U5225 (N_5225,N_4758,N_4787);
or U5226 (N_5226,N_4964,N_4974);
and U5227 (N_5227,N_4777,N_4625);
nand U5228 (N_5228,N_4782,N_4634);
and U5229 (N_5229,N_4637,N_4910);
or U5230 (N_5230,N_4658,N_4907);
nand U5231 (N_5231,N_4580,N_4664);
or U5232 (N_5232,N_4979,N_4933);
xor U5233 (N_5233,N_4705,N_4969);
xor U5234 (N_5234,N_4953,N_4935);
nor U5235 (N_5235,N_4864,N_4939);
xnor U5236 (N_5236,N_4685,N_4835);
nand U5237 (N_5237,N_4946,N_4925);
xor U5238 (N_5238,N_4707,N_4564);
or U5239 (N_5239,N_4821,N_4738);
nand U5240 (N_5240,N_4654,N_4788);
nor U5241 (N_5241,N_4677,N_4808);
and U5242 (N_5242,N_4590,N_4904);
or U5243 (N_5243,N_4826,N_4847);
nor U5244 (N_5244,N_4875,N_4649);
or U5245 (N_5245,N_4850,N_4628);
nor U5246 (N_5246,N_4914,N_4876);
xor U5247 (N_5247,N_4665,N_4745);
and U5248 (N_5248,N_4702,N_4844);
or U5249 (N_5249,N_4716,N_4855);
and U5250 (N_5250,N_4643,N_4549);
xor U5251 (N_5251,N_4809,N_4747);
xor U5252 (N_5252,N_4631,N_4628);
xor U5253 (N_5253,N_4988,N_4593);
and U5254 (N_5254,N_4984,N_4749);
nor U5255 (N_5255,N_4721,N_4934);
and U5256 (N_5256,N_4802,N_4531);
nand U5257 (N_5257,N_4593,N_4921);
and U5258 (N_5258,N_4629,N_4703);
nand U5259 (N_5259,N_4921,N_4854);
nor U5260 (N_5260,N_4576,N_4704);
nor U5261 (N_5261,N_4719,N_4950);
nand U5262 (N_5262,N_4690,N_4670);
xor U5263 (N_5263,N_4921,N_4610);
nor U5264 (N_5264,N_4592,N_4961);
nand U5265 (N_5265,N_4901,N_4586);
xnor U5266 (N_5266,N_4916,N_4708);
or U5267 (N_5267,N_4943,N_4669);
or U5268 (N_5268,N_4882,N_4886);
or U5269 (N_5269,N_4587,N_4896);
or U5270 (N_5270,N_4941,N_4547);
and U5271 (N_5271,N_4651,N_4594);
nor U5272 (N_5272,N_4980,N_4670);
xor U5273 (N_5273,N_4846,N_4542);
or U5274 (N_5274,N_4701,N_4969);
nand U5275 (N_5275,N_4629,N_4967);
or U5276 (N_5276,N_4691,N_4762);
nor U5277 (N_5277,N_4971,N_4939);
xnor U5278 (N_5278,N_4830,N_4647);
xor U5279 (N_5279,N_4781,N_4923);
nand U5280 (N_5280,N_4854,N_4968);
nor U5281 (N_5281,N_4989,N_4505);
and U5282 (N_5282,N_4558,N_4595);
nand U5283 (N_5283,N_4977,N_4623);
nor U5284 (N_5284,N_4784,N_4815);
nor U5285 (N_5285,N_4965,N_4818);
nor U5286 (N_5286,N_4520,N_4557);
nand U5287 (N_5287,N_4503,N_4603);
and U5288 (N_5288,N_4980,N_4876);
xor U5289 (N_5289,N_4671,N_4880);
and U5290 (N_5290,N_4545,N_4669);
and U5291 (N_5291,N_4819,N_4673);
xnor U5292 (N_5292,N_4799,N_4558);
nand U5293 (N_5293,N_4635,N_4624);
or U5294 (N_5294,N_4510,N_4716);
nor U5295 (N_5295,N_4522,N_4970);
xor U5296 (N_5296,N_4634,N_4643);
nand U5297 (N_5297,N_4783,N_4859);
nand U5298 (N_5298,N_4653,N_4985);
nand U5299 (N_5299,N_4758,N_4591);
xor U5300 (N_5300,N_4794,N_4740);
xor U5301 (N_5301,N_4652,N_4503);
nand U5302 (N_5302,N_4514,N_4977);
and U5303 (N_5303,N_4944,N_4865);
nor U5304 (N_5304,N_4534,N_4543);
nor U5305 (N_5305,N_4740,N_4904);
and U5306 (N_5306,N_4703,N_4667);
nor U5307 (N_5307,N_4967,N_4891);
nor U5308 (N_5308,N_4893,N_4954);
xnor U5309 (N_5309,N_4726,N_4970);
or U5310 (N_5310,N_4754,N_4849);
nand U5311 (N_5311,N_4895,N_4750);
nand U5312 (N_5312,N_4817,N_4803);
nor U5313 (N_5313,N_4761,N_4805);
or U5314 (N_5314,N_4783,N_4537);
or U5315 (N_5315,N_4504,N_4619);
or U5316 (N_5316,N_4810,N_4962);
nor U5317 (N_5317,N_4805,N_4637);
nand U5318 (N_5318,N_4572,N_4695);
nor U5319 (N_5319,N_4589,N_4976);
nor U5320 (N_5320,N_4788,N_4540);
and U5321 (N_5321,N_4975,N_4804);
and U5322 (N_5322,N_4537,N_4536);
xnor U5323 (N_5323,N_4561,N_4775);
xnor U5324 (N_5324,N_4501,N_4663);
xnor U5325 (N_5325,N_4777,N_4952);
nor U5326 (N_5326,N_4914,N_4521);
and U5327 (N_5327,N_4675,N_4780);
xor U5328 (N_5328,N_4796,N_4608);
and U5329 (N_5329,N_4934,N_4539);
nand U5330 (N_5330,N_4727,N_4587);
or U5331 (N_5331,N_4729,N_4763);
xnor U5332 (N_5332,N_4961,N_4763);
nand U5333 (N_5333,N_4582,N_4902);
or U5334 (N_5334,N_4905,N_4918);
nand U5335 (N_5335,N_4865,N_4770);
nor U5336 (N_5336,N_4534,N_4500);
xnor U5337 (N_5337,N_4649,N_4524);
nor U5338 (N_5338,N_4897,N_4715);
xor U5339 (N_5339,N_4598,N_4724);
nand U5340 (N_5340,N_4570,N_4601);
nor U5341 (N_5341,N_4542,N_4888);
nand U5342 (N_5342,N_4984,N_4920);
nor U5343 (N_5343,N_4881,N_4818);
and U5344 (N_5344,N_4997,N_4568);
nand U5345 (N_5345,N_4716,N_4944);
xor U5346 (N_5346,N_4802,N_4966);
and U5347 (N_5347,N_4892,N_4900);
or U5348 (N_5348,N_4551,N_4860);
xnor U5349 (N_5349,N_4574,N_4528);
and U5350 (N_5350,N_4926,N_4991);
or U5351 (N_5351,N_4851,N_4957);
nor U5352 (N_5352,N_4768,N_4634);
or U5353 (N_5353,N_4762,N_4773);
or U5354 (N_5354,N_4987,N_4887);
or U5355 (N_5355,N_4599,N_4720);
and U5356 (N_5356,N_4847,N_4940);
or U5357 (N_5357,N_4698,N_4596);
and U5358 (N_5358,N_4636,N_4643);
and U5359 (N_5359,N_4741,N_4656);
nor U5360 (N_5360,N_4789,N_4768);
or U5361 (N_5361,N_4837,N_4871);
xnor U5362 (N_5362,N_4807,N_4528);
and U5363 (N_5363,N_4832,N_4762);
nand U5364 (N_5364,N_4816,N_4946);
nand U5365 (N_5365,N_4798,N_4603);
xor U5366 (N_5366,N_4769,N_4952);
nor U5367 (N_5367,N_4738,N_4758);
or U5368 (N_5368,N_4753,N_4780);
xor U5369 (N_5369,N_4784,N_4584);
nor U5370 (N_5370,N_4619,N_4960);
and U5371 (N_5371,N_4848,N_4590);
xor U5372 (N_5372,N_4532,N_4647);
xnor U5373 (N_5373,N_4736,N_4884);
xor U5374 (N_5374,N_4712,N_4638);
and U5375 (N_5375,N_4812,N_4840);
nor U5376 (N_5376,N_4941,N_4765);
or U5377 (N_5377,N_4793,N_4698);
and U5378 (N_5378,N_4566,N_4894);
and U5379 (N_5379,N_4986,N_4559);
nand U5380 (N_5380,N_4715,N_4574);
or U5381 (N_5381,N_4721,N_4872);
xor U5382 (N_5382,N_4960,N_4730);
nor U5383 (N_5383,N_4610,N_4744);
nand U5384 (N_5384,N_4975,N_4689);
nor U5385 (N_5385,N_4527,N_4992);
nor U5386 (N_5386,N_4970,N_4866);
or U5387 (N_5387,N_4781,N_4921);
nand U5388 (N_5388,N_4667,N_4807);
or U5389 (N_5389,N_4778,N_4754);
xor U5390 (N_5390,N_4567,N_4970);
nand U5391 (N_5391,N_4590,N_4714);
and U5392 (N_5392,N_4829,N_4673);
xnor U5393 (N_5393,N_4842,N_4501);
and U5394 (N_5394,N_4626,N_4822);
and U5395 (N_5395,N_4766,N_4946);
or U5396 (N_5396,N_4782,N_4823);
xnor U5397 (N_5397,N_4986,N_4695);
or U5398 (N_5398,N_4796,N_4570);
xor U5399 (N_5399,N_4685,N_4528);
nor U5400 (N_5400,N_4560,N_4804);
and U5401 (N_5401,N_4649,N_4685);
or U5402 (N_5402,N_4870,N_4711);
and U5403 (N_5403,N_4564,N_4858);
xor U5404 (N_5404,N_4992,N_4863);
xnor U5405 (N_5405,N_4651,N_4528);
nor U5406 (N_5406,N_4965,N_4975);
xor U5407 (N_5407,N_4578,N_4600);
nand U5408 (N_5408,N_4994,N_4903);
and U5409 (N_5409,N_4689,N_4989);
and U5410 (N_5410,N_4741,N_4753);
or U5411 (N_5411,N_4795,N_4703);
nor U5412 (N_5412,N_4794,N_4755);
nor U5413 (N_5413,N_4976,N_4781);
nor U5414 (N_5414,N_4663,N_4856);
xor U5415 (N_5415,N_4920,N_4595);
nand U5416 (N_5416,N_4642,N_4983);
or U5417 (N_5417,N_4697,N_4922);
and U5418 (N_5418,N_4645,N_4936);
or U5419 (N_5419,N_4863,N_4781);
nor U5420 (N_5420,N_4782,N_4764);
nor U5421 (N_5421,N_4567,N_4520);
nand U5422 (N_5422,N_4502,N_4818);
xnor U5423 (N_5423,N_4617,N_4708);
and U5424 (N_5424,N_4638,N_4583);
nand U5425 (N_5425,N_4667,N_4606);
or U5426 (N_5426,N_4944,N_4780);
nand U5427 (N_5427,N_4914,N_4734);
xnor U5428 (N_5428,N_4711,N_4688);
nor U5429 (N_5429,N_4629,N_4887);
nand U5430 (N_5430,N_4649,N_4568);
or U5431 (N_5431,N_4700,N_4620);
and U5432 (N_5432,N_4640,N_4989);
nor U5433 (N_5433,N_4589,N_4626);
or U5434 (N_5434,N_4598,N_4581);
and U5435 (N_5435,N_4526,N_4568);
or U5436 (N_5436,N_4903,N_4695);
nor U5437 (N_5437,N_4528,N_4704);
xor U5438 (N_5438,N_4821,N_4675);
nand U5439 (N_5439,N_4860,N_4761);
xor U5440 (N_5440,N_4997,N_4502);
nor U5441 (N_5441,N_4903,N_4848);
xor U5442 (N_5442,N_4831,N_4536);
xnor U5443 (N_5443,N_4900,N_4611);
nand U5444 (N_5444,N_4833,N_4834);
nand U5445 (N_5445,N_4781,N_4930);
nor U5446 (N_5446,N_4879,N_4882);
xnor U5447 (N_5447,N_4976,N_4646);
and U5448 (N_5448,N_4517,N_4817);
or U5449 (N_5449,N_4998,N_4909);
nor U5450 (N_5450,N_4948,N_4959);
xnor U5451 (N_5451,N_4875,N_4897);
nand U5452 (N_5452,N_4982,N_4978);
nor U5453 (N_5453,N_4774,N_4979);
xnor U5454 (N_5454,N_4817,N_4890);
or U5455 (N_5455,N_4617,N_4984);
nand U5456 (N_5456,N_4668,N_4564);
nor U5457 (N_5457,N_4785,N_4514);
nor U5458 (N_5458,N_4870,N_4856);
nor U5459 (N_5459,N_4637,N_4554);
or U5460 (N_5460,N_4817,N_4867);
nor U5461 (N_5461,N_4914,N_4866);
nor U5462 (N_5462,N_4691,N_4908);
and U5463 (N_5463,N_4862,N_4906);
nand U5464 (N_5464,N_4614,N_4584);
or U5465 (N_5465,N_4890,N_4580);
or U5466 (N_5466,N_4650,N_4769);
nor U5467 (N_5467,N_4912,N_4661);
and U5468 (N_5468,N_4831,N_4505);
and U5469 (N_5469,N_4986,N_4668);
nand U5470 (N_5470,N_4830,N_4836);
and U5471 (N_5471,N_4822,N_4906);
and U5472 (N_5472,N_4759,N_4543);
xnor U5473 (N_5473,N_4570,N_4873);
nor U5474 (N_5474,N_4606,N_4504);
xnor U5475 (N_5475,N_4557,N_4550);
nand U5476 (N_5476,N_4766,N_4718);
or U5477 (N_5477,N_4552,N_4845);
nor U5478 (N_5478,N_4593,N_4575);
xor U5479 (N_5479,N_4699,N_4647);
or U5480 (N_5480,N_4813,N_4971);
and U5481 (N_5481,N_4864,N_4823);
nand U5482 (N_5482,N_4634,N_4620);
nand U5483 (N_5483,N_4776,N_4534);
or U5484 (N_5484,N_4934,N_4841);
nor U5485 (N_5485,N_4677,N_4858);
xor U5486 (N_5486,N_4973,N_4527);
xnor U5487 (N_5487,N_4630,N_4568);
and U5488 (N_5488,N_4651,N_4968);
nor U5489 (N_5489,N_4591,N_4815);
nand U5490 (N_5490,N_4850,N_4847);
nor U5491 (N_5491,N_4606,N_4858);
and U5492 (N_5492,N_4645,N_4715);
and U5493 (N_5493,N_4948,N_4541);
xnor U5494 (N_5494,N_4994,N_4954);
nor U5495 (N_5495,N_4556,N_4718);
nand U5496 (N_5496,N_4984,N_4879);
or U5497 (N_5497,N_4952,N_4671);
xor U5498 (N_5498,N_4806,N_4753);
and U5499 (N_5499,N_4876,N_4649);
nand U5500 (N_5500,N_5364,N_5217);
nor U5501 (N_5501,N_5324,N_5281);
or U5502 (N_5502,N_5186,N_5034);
xnor U5503 (N_5503,N_5295,N_5124);
nand U5504 (N_5504,N_5042,N_5294);
or U5505 (N_5505,N_5086,N_5134);
nand U5506 (N_5506,N_5396,N_5398);
or U5507 (N_5507,N_5017,N_5403);
xor U5508 (N_5508,N_5141,N_5147);
or U5509 (N_5509,N_5193,N_5122);
or U5510 (N_5510,N_5103,N_5130);
or U5511 (N_5511,N_5444,N_5374);
nor U5512 (N_5512,N_5464,N_5190);
xor U5513 (N_5513,N_5388,N_5430);
and U5514 (N_5514,N_5454,N_5062);
and U5515 (N_5515,N_5325,N_5437);
and U5516 (N_5516,N_5219,N_5225);
nand U5517 (N_5517,N_5336,N_5126);
nor U5518 (N_5518,N_5076,N_5263);
xor U5519 (N_5519,N_5303,N_5249);
or U5520 (N_5520,N_5256,N_5288);
nor U5521 (N_5521,N_5253,N_5316);
nand U5522 (N_5522,N_5381,N_5467);
nand U5523 (N_5523,N_5347,N_5280);
or U5524 (N_5524,N_5428,N_5269);
xor U5525 (N_5525,N_5414,N_5239);
xor U5526 (N_5526,N_5333,N_5262);
xor U5527 (N_5527,N_5450,N_5004);
nor U5528 (N_5528,N_5125,N_5290);
or U5529 (N_5529,N_5453,N_5440);
xnor U5530 (N_5530,N_5421,N_5093);
xnor U5531 (N_5531,N_5348,N_5349);
xor U5532 (N_5532,N_5418,N_5174);
or U5533 (N_5533,N_5088,N_5242);
or U5534 (N_5534,N_5244,N_5455);
or U5535 (N_5535,N_5267,N_5476);
nor U5536 (N_5536,N_5328,N_5479);
nand U5537 (N_5537,N_5304,N_5429);
nor U5538 (N_5538,N_5461,N_5060);
nand U5539 (N_5539,N_5458,N_5350);
xnor U5540 (N_5540,N_5240,N_5298);
nand U5541 (N_5541,N_5439,N_5268);
nor U5542 (N_5542,N_5023,N_5118);
xnor U5543 (N_5543,N_5010,N_5462);
nor U5544 (N_5544,N_5145,N_5206);
nand U5545 (N_5545,N_5137,N_5059);
nor U5546 (N_5546,N_5386,N_5053);
xor U5547 (N_5547,N_5344,N_5278);
nor U5548 (N_5548,N_5040,N_5265);
nand U5549 (N_5549,N_5291,N_5205);
xor U5550 (N_5550,N_5255,N_5358);
xor U5551 (N_5551,N_5431,N_5433);
and U5552 (N_5552,N_5412,N_5419);
xnor U5553 (N_5553,N_5299,N_5260);
nor U5554 (N_5554,N_5317,N_5334);
nand U5555 (N_5555,N_5071,N_5471);
nor U5556 (N_5556,N_5046,N_5183);
xor U5557 (N_5557,N_5377,N_5097);
and U5558 (N_5558,N_5150,N_5413);
xnor U5559 (N_5559,N_5153,N_5441);
or U5560 (N_5560,N_5084,N_5068);
or U5561 (N_5561,N_5109,N_5089);
xor U5562 (N_5562,N_5391,N_5101);
xor U5563 (N_5563,N_5104,N_5443);
and U5564 (N_5564,N_5392,N_5156);
and U5565 (N_5565,N_5445,N_5085);
nand U5566 (N_5566,N_5251,N_5436);
or U5567 (N_5567,N_5223,N_5468);
nand U5568 (N_5568,N_5070,N_5013);
and U5569 (N_5569,N_5169,N_5371);
nor U5570 (N_5570,N_5259,N_5207);
nor U5571 (N_5571,N_5230,N_5056);
and U5572 (N_5572,N_5360,N_5382);
and U5573 (N_5573,N_5138,N_5228);
and U5574 (N_5574,N_5055,N_5438);
nor U5575 (N_5575,N_5006,N_5490);
nor U5576 (N_5576,N_5261,N_5050);
nor U5577 (N_5577,N_5315,N_5110);
or U5578 (N_5578,N_5401,N_5483);
or U5579 (N_5579,N_5029,N_5338);
xor U5580 (N_5580,N_5319,N_5459);
xor U5581 (N_5581,N_5424,N_5170);
xnor U5582 (N_5582,N_5387,N_5111);
and U5583 (N_5583,N_5250,N_5065);
and U5584 (N_5584,N_5181,N_5289);
or U5585 (N_5585,N_5243,N_5200);
and U5586 (N_5586,N_5275,N_5102);
and U5587 (N_5587,N_5485,N_5066);
or U5588 (N_5588,N_5128,N_5486);
nand U5589 (N_5589,N_5305,N_5131);
and U5590 (N_5590,N_5033,N_5481);
nor U5591 (N_5591,N_5422,N_5273);
nand U5592 (N_5592,N_5359,N_5173);
nand U5593 (N_5593,N_5460,N_5079);
xor U5594 (N_5594,N_5044,N_5301);
xor U5595 (N_5595,N_5139,N_5376);
and U5596 (N_5596,N_5456,N_5083);
nor U5597 (N_5597,N_5494,N_5064);
xor U5598 (N_5598,N_5411,N_5195);
nor U5599 (N_5599,N_5340,N_5312);
xnor U5600 (N_5600,N_5287,N_5005);
nand U5601 (N_5601,N_5077,N_5149);
and U5602 (N_5602,N_5172,N_5451);
xor U5603 (N_5603,N_5368,N_5107);
nand U5604 (N_5604,N_5274,N_5321);
or U5605 (N_5605,N_5354,N_5492);
nor U5606 (N_5606,N_5096,N_5212);
xnor U5607 (N_5607,N_5361,N_5480);
xor U5608 (N_5608,N_5416,N_5166);
nand U5609 (N_5609,N_5277,N_5235);
nand U5610 (N_5610,N_5072,N_5318);
nor U5611 (N_5611,N_5427,N_5188);
xnor U5612 (N_5612,N_5018,N_5353);
and U5613 (N_5613,N_5308,N_5367);
xnor U5614 (N_5614,N_5435,N_5165);
or U5615 (N_5615,N_5108,N_5189);
nor U5616 (N_5616,N_5246,N_5270);
xor U5617 (N_5617,N_5393,N_5365);
nor U5618 (N_5618,N_5496,N_5432);
nor U5619 (N_5619,N_5081,N_5322);
nor U5620 (N_5620,N_5120,N_5495);
and U5621 (N_5621,N_5341,N_5178);
or U5622 (N_5622,N_5356,N_5221);
nand U5623 (N_5623,N_5168,N_5397);
and U5624 (N_5624,N_5019,N_5400);
nand U5625 (N_5625,N_5203,N_5241);
and U5626 (N_5626,N_5216,N_5497);
xor U5627 (N_5627,N_5293,N_5075);
nand U5628 (N_5628,N_5369,N_5067);
xnor U5629 (N_5629,N_5123,N_5475);
or U5630 (N_5630,N_5409,N_5048);
nor U5631 (N_5631,N_5208,N_5335);
xnor U5632 (N_5632,N_5320,N_5119);
and U5633 (N_5633,N_5478,N_5231);
and U5634 (N_5634,N_5129,N_5425);
and U5635 (N_5635,N_5488,N_5213);
nand U5636 (N_5636,N_5282,N_5405);
nand U5637 (N_5637,N_5373,N_5314);
nand U5638 (N_5638,N_5449,N_5284);
or U5639 (N_5639,N_5027,N_5021);
and U5640 (N_5640,N_5082,N_5390);
or U5641 (N_5641,N_5470,N_5226);
xnor U5642 (N_5642,N_5326,N_5002);
or U5643 (N_5643,N_5346,N_5052);
xor U5644 (N_5644,N_5136,N_5229);
nand U5645 (N_5645,N_5025,N_5035);
and U5646 (N_5646,N_5191,N_5041);
xnor U5647 (N_5647,N_5306,N_5198);
or U5648 (N_5648,N_5155,N_5000);
xor U5649 (N_5649,N_5484,N_5296);
and U5650 (N_5650,N_5215,N_5463);
nor U5651 (N_5651,N_5003,N_5473);
or U5652 (N_5652,N_5327,N_5420);
nand U5653 (N_5653,N_5252,N_5204);
nand U5654 (N_5654,N_5307,N_5133);
or U5655 (N_5655,N_5051,N_5469);
or U5656 (N_5656,N_5112,N_5161);
xnor U5657 (N_5657,N_5031,N_5127);
xnor U5658 (N_5658,N_5163,N_5266);
or U5659 (N_5659,N_5465,N_5415);
and U5660 (N_5660,N_5254,N_5448);
nand U5661 (N_5661,N_5264,N_5487);
and U5662 (N_5662,N_5043,N_5389);
nand U5663 (N_5663,N_5121,N_5383);
or U5664 (N_5664,N_5257,N_5047);
nand U5665 (N_5665,N_5489,N_5016);
nor U5666 (N_5666,N_5032,N_5297);
xor U5667 (N_5667,N_5045,N_5037);
nor U5668 (N_5668,N_5362,N_5012);
nand U5669 (N_5669,N_5247,N_5148);
nor U5670 (N_5670,N_5140,N_5406);
nor U5671 (N_5671,N_5074,N_5143);
nand U5672 (N_5672,N_5452,N_5009);
nand U5673 (N_5673,N_5114,N_5054);
or U5674 (N_5674,N_5309,N_5442);
and U5675 (N_5675,N_5423,N_5310);
nor U5676 (N_5676,N_5194,N_5345);
xnor U5677 (N_5677,N_5493,N_5026);
or U5678 (N_5678,N_5238,N_5106);
xnor U5679 (N_5679,N_5222,N_5185);
nand U5680 (N_5680,N_5337,N_5022);
xnor U5681 (N_5681,N_5008,N_5209);
xnor U5682 (N_5682,N_5285,N_5434);
or U5683 (N_5683,N_5248,N_5159);
nand U5684 (N_5684,N_5038,N_5020);
nor U5685 (N_5685,N_5329,N_5342);
and U5686 (N_5686,N_5176,N_5446);
and U5687 (N_5687,N_5302,N_5098);
and U5688 (N_5688,N_5196,N_5457);
xnor U5689 (N_5689,N_5152,N_5171);
nand U5690 (N_5690,N_5095,N_5224);
and U5691 (N_5691,N_5498,N_5036);
and U5692 (N_5692,N_5091,N_5132);
nor U5693 (N_5693,N_5323,N_5292);
nand U5694 (N_5694,N_5039,N_5482);
xor U5695 (N_5695,N_5007,N_5339);
xor U5696 (N_5696,N_5408,N_5179);
xor U5697 (N_5697,N_5258,N_5162);
nor U5698 (N_5698,N_5113,N_5061);
nor U5699 (N_5699,N_5151,N_5232);
nand U5700 (N_5700,N_5370,N_5366);
nand U5701 (N_5701,N_5447,N_5384);
nand U5702 (N_5702,N_5466,N_5426);
or U5703 (N_5703,N_5199,N_5491);
and U5704 (N_5704,N_5211,N_5363);
or U5705 (N_5705,N_5375,N_5201);
nor U5706 (N_5706,N_5144,N_5407);
or U5707 (N_5707,N_5214,N_5351);
nor U5708 (N_5708,N_5395,N_5117);
nor U5709 (N_5709,N_5014,N_5276);
xor U5710 (N_5710,N_5164,N_5202);
and U5711 (N_5711,N_5057,N_5245);
and U5712 (N_5712,N_5094,N_5099);
nor U5713 (N_5713,N_5028,N_5080);
nand U5714 (N_5714,N_5154,N_5343);
nand U5715 (N_5715,N_5157,N_5220);
or U5716 (N_5716,N_5499,N_5311);
or U5717 (N_5717,N_5146,N_5378);
xnor U5718 (N_5718,N_5286,N_5078);
nor U5719 (N_5719,N_5184,N_5063);
nand U5720 (N_5720,N_5001,N_5069);
nor U5721 (N_5721,N_5087,N_5355);
or U5722 (N_5722,N_5180,N_5399);
nand U5723 (N_5723,N_5227,N_5158);
nand U5724 (N_5724,N_5234,N_5218);
xnor U5725 (N_5725,N_5192,N_5187);
or U5726 (N_5726,N_5160,N_5474);
or U5727 (N_5727,N_5385,N_5300);
nand U5728 (N_5728,N_5116,N_5352);
nand U5729 (N_5729,N_5210,N_5233);
nor U5730 (N_5730,N_5417,N_5331);
nor U5731 (N_5731,N_5357,N_5379);
nand U5732 (N_5732,N_5404,N_5135);
nor U5733 (N_5733,N_5279,N_5090);
xor U5734 (N_5734,N_5410,N_5024);
nand U5735 (N_5735,N_5332,N_5271);
nor U5736 (N_5736,N_5175,N_5283);
xor U5737 (N_5737,N_5197,N_5030);
xor U5738 (N_5738,N_5115,N_5477);
or U5739 (N_5739,N_5011,N_5058);
or U5740 (N_5740,N_5177,N_5100);
xor U5741 (N_5741,N_5313,N_5073);
nor U5742 (N_5742,N_5380,N_5182);
or U5743 (N_5743,N_5015,N_5394);
nand U5744 (N_5744,N_5092,N_5372);
xnor U5745 (N_5745,N_5237,N_5236);
nand U5746 (N_5746,N_5049,N_5330);
nor U5747 (N_5747,N_5472,N_5402);
and U5748 (N_5748,N_5167,N_5142);
nor U5749 (N_5749,N_5105,N_5272);
nor U5750 (N_5750,N_5397,N_5439);
or U5751 (N_5751,N_5199,N_5069);
xor U5752 (N_5752,N_5426,N_5232);
nand U5753 (N_5753,N_5152,N_5145);
xnor U5754 (N_5754,N_5307,N_5326);
or U5755 (N_5755,N_5036,N_5280);
and U5756 (N_5756,N_5105,N_5143);
nor U5757 (N_5757,N_5105,N_5277);
and U5758 (N_5758,N_5121,N_5096);
nand U5759 (N_5759,N_5453,N_5221);
and U5760 (N_5760,N_5154,N_5025);
xor U5761 (N_5761,N_5182,N_5008);
nand U5762 (N_5762,N_5177,N_5339);
or U5763 (N_5763,N_5151,N_5361);
nor U5764 (N_5764,N_5358,N_5417);
nor U5765 (N_5765,N_5289,N_5276);
nor U5766 (N_5766,N_5195,N_5191);
nor U5767 (N_5767,N_5358,N_5335);
xor U5768 (N_5768,N_5171,N_5051);
nand U5769 (N_5769,N_5146,N_5244);
and U5770 (N_5770,N_5132,N_5310);
xnor U5771 (N_5771,N_5085,N_5309);
nor U5772 (N_5772,N_5158,N_5461);
xor U5773 (N_5773,N_5292,N_5469);
nor U5774 (N_5774,N_5217,N_5356);
nand U5775 (N_5775,N_5006,N_5137);
xor U5776 (N_5776,N_5124,N_5115);
nor U5777 (N_5777,N_5436,N_5403);
nand U5778 (N_5778,N_5325,N_5009);
nor U5779 (N_5779,N_5054,N_5276);
nand U5780 (N_5780,N_5332,N_5203);
nand U5781 (N_5781,N_5283,N_5119);
and U5782 (N_5782,N_5101,N_5068);
and U5783 (N_5783,N_5143,N_5354);
xnor U5784 (N_5784,N_5064,N_5389);
xor U5785 (N_5785,N_5291,N_5419);
nand U5786 (N_5786,N_5321,N_5299);
or U5787 (N_5787,N_5416,N_5492);
and U5788 (N_5788,N_5314,N_5090);
and U5789 (N_5789,N_5474,N_5099);
nor U5790 (N_5790,N_5169,N_5395);
nand U5791 (N_5791,N_5131,N_5326);
xnor U5792 (N_5792,N_5152,N_5388);
nand U5793 (N_5793,N_5440,N_5016);
nor U5794 (N_5794,N_5357,N_5375);
nor U5795 (N_5795,N_5391,N_5412);
xor U5796 (N_5796,N_5271,N_5238);
nand U5797 (N_5797,N_5359,N_5467);
or U5798 (N_5798,N_5093,N_5158);
nand U5799 (N_5799,N_5100,N_5080);
or U5800 (N_5800,N_5058,N_5100);
and U5801 (N_5801,N_5042,N_5337);
nand U5802 (N_5802,N_5263,N_5140);
and U5803 (N_5803,N_5242,N_5395);
and U5804 (N_5804,N_5391,N_5289);
nor U5805 (N_5805,N_5012,N_5486);
nand U5806 (N_5806,N_5201,N_5471);
and U5807 (N_5807,N_5132,N_5302);
and U5808 (N_5808,N_5048,N_5232);
or U5809 (N_5809,N_5425,N_5211);
xor U5810 (N_5810,N_5374,N_5465);
or U5811 (N_5811,N_5499,N_5235);
or U5812 (N_5812,N_5023,N_5295);
nand U5813 (N_5813,N_5295,N_5300);
nor U5814 (N_5814,N_5057,N_5024);
or U5815 (N_5815,N_5153,N_5234);
and U5816 (N_5816,N_5478,N_5109);
nand U5817 (N_5817,N_5174,N_5430);
or U5818 (N_5818,N_5404,N_5260);
nand U5819 (N_5819,N_5307,N_5355);
or U5820 (N_5820,N_5390,N_5278);
nor U5821 (N_5821,N_5157,N_5390);
or U5822 (N_5822,N_5132,N_5419);
and U5823 (N_5823,N_5039,N_5254);
and U5824 (N_5824,N_5428,N_5267);
xnor U5825 (N_5825,N_5431,N_5115);
nand U5826 (N_5826,N_5158,N_5345);
and U5827 (N_5827,N_5478,N_5020);
nor U5828 (N_5828,N_5460,N_5165);
and U5829 (N_5829,N_5303,N_5011);
or U5830 (N_5830,N_5157,N_5163);
nor U5831 (N_5831,N_5492,N_5322);
xor U5832 (N_5832,N_5099,N_5265);
or U5833 (N_5833,N_5464,N_5491);
or U5834 (N_5834,N_5083,N_5211);
xor U5835 (N_5835,N_5110,N_5140);
xor U5836 (N_5836,N_5401,N_5063);
and U5837 (N_5837,N_5064,N_5487);
and U5838 (N_5838,N_5473,N_5025);
or U5839 (N_5839,N_5445,N_5238);
or U5840 (N_5840,N_5107,N_5378);
xor U5841 (N_5841,N_5110,N_5017);
and U5842 (N_5842,N_5401,N_5083);
and U5843 (N_5843,N_5222,N_5482);
and U5844 (N_5844,N_5174,N_5472);
or U5845 (N_5845,N_5294,N_5216);
nand U5846 (N_5846,N_5051,N_5162);
nand U5847 (N_5847,N_5073,N_5353);
or U5848 (N_5848,N_5083,N_5333);
or U5849 (N_5849,N_5064,N_5079);
xor U5850 (N_5850,N_5231,N_5134);
xor U5851 (N_5851,N_5319,N_5281);
nor U5852 (N_5852,N_5372,N_5452);
nor U5853 (N_5853,N_5026,N_5060);
or U5854 (N_5854,N_5192,N_5166);
xnor U5855 (N_5855,N_5209,N_5380);
nand U5856 (N_5856,N_5187,N_5267);
or U5857 (N_5857,N_5446,N_5281);
or U5858 (N_5858,N_5360,N_5071);
or U5859 (N_5859,N_5006,N_5173);
nand U5860 (N_5860,N_5105,N_5005);
and U5861 (N_5861,N_5176,N_5206);
and U5862 (N_5862,N_5341,N_5238);
nor U5863 (N_5863,N_5114,N_5495);
nor U5864 (N_5864,N_5336,N_5177);
and U5865 (N_5865,N_5117,N_5473);
and U5866 (N_5866,N_5481,N_5069);
nor U5867 (N_5867,N_5421,N_5405);
nor U5868 (N_5868,N_5411,N_5104);
or U5869 (N_5869,N_5279,N_5223);
or U5870 (N_5870,N_5271,N_5140);
xor U5871 (N_5871,N_5201,N_5450);
or U5872 (N_5872,N_5303,N_5028);
nand U5873 (N_5873,N_5085,N_5415);
nor U5874 (N_5874,N_5282,N_5286);
nor U5875 (N_5875,N_5229,N_5059);
and U5876 (N_5876,N_5370,N_5421);
nand U5877 (N_5877,N_5359,N_5396);
nor U5878 (N_5878,N_5244,N_5015);
and U5879 (N_5879,N_5108,N_5093);
or U5880 (N_5880,N_5332,N_5441);
xnor U5881 (N_5881,N_5314,N_5334);
and U5882 (N_5882,N_5085,N_5286);
xnor U5883 (N_5883,N_5190,N_5221);
nor U5884 (N_5884,N_5039,N_5181);
xor U5885 (N_5885,N_5006,N_5476);
and U5886 (N_5886,N_5047,N_5250);
nand U5887 (N_5887,N_5358,N_5254);
nand U5888 (N_5888,N_5350,N_5451);
and U5889 (N_5889,N_5397,N_5293);
nand U5890 (N_5890,N_5339,N_5487);
or U5891 (N_5891,N_5263,N_5482);
xor U5892 (N_5892,N_5110,N_5161);
nor U5893 (N_5893,N_5352,N_5248);
nor U5894 (N_5894,N_5068,N_5058);
nor U5895 (N_5895,N_5121,N_5247);
or U5896 (N_5896,N_5275,N_5064);
nor U5897 (N_5897,N_5155,N_5193);
nand U5898 (N_5898,N_5003,N_5083);
nor U5899 (N_5899,N_5212,N_5077);
or U5900 (N_5900,N_5311,N_5016);
nor U5901 (N_5901,N_5192,N_5302);
and U5902 (N_5902,N_5101,N_5494);
and U5903 (N_5903,N_5069,N_5131);
xnor U5904 (N_5904,N_5240,N_5277);
or U5905 (N_5905,N_5327,N_5414);
nor U5906 (N_5906,N_5275,N_5364);
and U5907 (N_5907,N_5354,N_5423);
and U5908 (N_5908,N_5395,N_5377);
and U5909 (N_5909,N_5230,N_5241);
or U5910 (N_5910,N_5467,N_5363);
nor U5911 (N_5911,N_5255,N_5264);
xor U5912 (N_5912,N_5407,N_5203);
nor U5913 (N_5913,N_5469,N_5259);
or U5914 (N_5914,N_5496,N_5164);
and U5915 (N_5915,N_5026,N_5158);
and U5916 (N_5916,N_5394,N_5406);
and U5917 (N_5917,N_5235,N_5249);
xnor U5918 (N_5918,N_5015,N_5488);
and U5919 (N_5919,N_5013,N_5367);
xnor U5920 (N_5920,N_5237,N_5165);
nand U5921 (N_5921,N_5451,N_5049);
nor U5922 (N_5922,N_5294,N_5122);
nand U5923 (N_5923,N_5164,N_5435);
nor U5924 (N_5924,N_5099,N_5042);
nand U5925 (N_5925,N_5229,N_5449);
nand U5926 (N_5926,N_5039,N_5236);
nor U5927 (N_5927,N_5273,N_5276);
nand U5928 (N_5928,N_5251,N_5238);
xnor U5929 (N_5929,N_5167,N_5359);
nor U5930 (N_5930,N_5332,N_5300);
xnor U5931 (N_5931,N_5106,N_5009);
xor U5932 (N_5932,N_5451,N_5144);
or U5933 (N_5933,N_5179,N_5474);
xor U5934 (N_5934,N_5353,N_5418);
and U5935 (N_5935,N_5130,N_5223);
nor U5936 (N_5936,N_5029,N_5019);
or U5937 (N_5937,N_5416,N_5190);
xnor U5938 (N_5938,N_5283,N_5265);
nand U5939 (N_5939,N_5337,N_5297);
or U5940 (N_5940,N_5122,N_5365);
and U5941 (N_5941,N_5108,N_5442);
and U5942 (N_5942,N_5471,N_5041);
nor U5943 (N_5943,N_5210,N_5418);
nor U5944 (N_5944,N_5005,N_5268);
or U5945 (N_5945,N_5049,N_5263);
nor U5946 (N_5946,N_5481,N_5256);
nor U5947 (N_5947,N_5283,N_5064);
xor U5948 (N_5948,N_5092,N_5445);
and U5949 (N_5949,N_5280,N_5247);
xor U5950 (N_5950,N_5011,N_5421);
or U5951 (N_5951,N_5242,N_5134);
and U5952 (N_5952,N_5209,N_5315);
nand U5953 (N_5953,N_5469,N_5314);
nand U5954 (N_5954,N_5459,N_5218);
nor U5955 (N_5955,N_5333,N_5435);
and U5956 (N_5956,N_5377,N_5494);
nor U5957 (N_5957,N_5141,N_5265);
and U5958 (N_5958,N_5240,N_5035);
xor U5959 (N_5959,N_5242,N_5342);
nor U5960 (N_5960,N_5258,N_5377);
nor U5961 (N_5961,N_5263,N_5340);
nand U5962 (N_5962,N_5026,N_5370);
and U5963 (N_5963,N_5308,N_5013);
nor U5964 (N_5964,N_5311,N_5055);
xor U5965 (N_5965,N_5015,N_5284);
nand U5966 (N_5966,N_5336,N_5082);
nand U5967 (N_5967,N_5207,N_5205);
and U5968 (N_5968,N_5303,N_5157);
and U5969 (N_5969,N_5369,N_5119);
or U5970 (N_5970,N_5282,N_5311);
or U5971 (N_5971,N_5324,N_5386);
nand U5972 (N_5972,N_5404,N_5382);
nor U5973 (N_5973,N_5409,N_5232);
or U5974 (N_5974,N_5140,N_5387);
and U5975 (N_5975,N_5159,N_5409);
nand U5976 (N_5976,N_5041,N_5473);
and U5977 (N_5977,N_5157,N_5282);
nor U5978 (N_5978,N_5423,N_5308);
or U5979 (N_5979,N_5335,N_5299);
or U5980 (N_5980,N_5228,N_5165);
or U5981 (N_5981,N_5433,N_5014);
or U5982 (N_5982,N_5278,N_5196);
nand U5983 (N_5983,N_5294,N_5428);
or U5984 (N_5984,N_5168,N_5098);
nor U5985 (N_5985,N_5419,N_5280);
xnor U5986 (N_5986,N_5388,N_5319);
and U5987 (N_5987,N_5002,N_5361);
xnor U5988 (N_5988,N_5086,N_5199);
and U5989 (N_5989,N_5483,N_5056);
and U5990 (N_5990,N_5414,N_5141);
and U5991 (N_5991,N_5393,N_5179);
nor U5992 (N_5992,N_5416,N_5443);
xor U5993 (N_5993,N_5385,N_5129);
nand U5994 (N_5994,N_5141,N_5103);
xnor U5995 (N_5995,N_5261,N_5303);
nand U5996 (N_5996,N_5286,N_5334);
nand U5997 (N_5997,N_5134,N_5214);
xor U5998 (N_5998,N_5444,N_5311);
or U5999 (N_5999,N_5394,N_5260);
or U6000 (N_6000,N_5902,N_5742);
xnor U6001 (N_6001,N_5601,N_5644);
and U6002 (N_6002,N_5781,N_5619);
xor U6003 (N_6003,N_5567,N_5663);
xor U6004 (N_6004,N_5819,N_5778);
nand U6005 (N_6005,N_5706,N_5946);
or U6006 (N_6006,N_5981,N_5519);
xor U6007 (N_6007,N_5650,N_5647);
nor U6008 (N_6008,N_5598,N_5814);
and U6009 (N_6009,N_5585,N_5876);
nor U6010 (N_6010,N_5746,N_5556);
xnor U6011 (N_6011,N_5715,N_5530);
xor U6012 (N_6012,N_5827,N_5641);
and U6013 (N_6013,N_5994,N_5798);
nand U6014 (N_6014,N_5614,N_5793);
or U6015 (N_6015,N_5908,N_5990);
or U6016 (N_6016,N_5676,N_5504);
or U6017 (N_6017,N_5745,N_5751);
and U6018 (N_6018,N_5588,N_5978);
nand U6019 (N_6019,N_5979,N_5847);
or U6020 (N_6020,N_5924,N_5809);
nand U6021 (N_6021,N_5718,N_5666);
or U6022 (N_6022,N_5791,N_5917);
and U6023 (N_6023,N_5671,N_5905);
or U6024 (N_6024,N_5708,N_5702);
or U6025 (N_6025,N_5664,N_5865);
xor U6026 (N_6026,N_5531,N_5863);
nand U6027 (N_6027,N_5796,N_5823);
xor U6028 (N_6028,N_5941,N_5750);
or U6029 (N_6029,N_5563,N_5761);
xor U6030 (N_6030,N_5731,N_5872);
and U6031 (N_6031,N_5704,N_5557);
nor U6032 (N_6032,N_5998,N_5802);
or U6033 (N_6033,N_5717,N_5550);
nand U6034 (N_6034,N_5756,N_5696);
nor U6035 (N_6035,N_5995,N_5586);
or U6036 (N_6036,N_5501,N_5681);
or U6037 (N_6037,N_5707,N_5767);
and U6038 (N_6038,N_5965,N_5898);
and U6039 (N_6039,N_5669,N_5596);
xnor U6040 (N_6040,N_5901,N_5511);
nand U6041 (N_6041,N_5577,N_5535);
nor U6042 (N_6042,N_5513,N_5803);
and U6043 (N_6043,N_5560,N_5993);
xor U6044 (N_6044,N_5748,N_5942);
xnor U6045 (N_6045,N_5966,N_5839);
or U6046 (N_6046,N_5816,N_5939);
xor U6047 (N_6047,N_5688,N_5806);
or U6048 (N_6048,N_5616,N_5996);
nand U6049 (N_6049,N_5621,N_5777);
xnor U6050 (N_6050,N_5899,N_5655);
or U6051 (N_6051,N_5907,N_5575);
or U6052 (N_6052,N_5589,N_5953);
or U6053 (N_6053,N_5690,N_5852);
xor U6054 (N_6054,N_5507,N_5843);
xnor U6055 (N_6055,N_5785,N_5698);
nor U6056 (N_6056,N_5835,N_5721);
and U6057 (N_6057,N_5955,N_5515);
xnor U6058 (N_6058,N_5881,N_5730);
or U6059 (N_6059,N_5665,N_5738);
nor U6060 (N_6060,N_5684,N_5747);
nor U6061 (N_6061,N_5808,N_5739);
or U6062 (N_6062,N_5630,N_5913);
nor U6063 (N_6063,N_5574,N_5529);
and U6064 (N_6064,N_5562,N_5576);
and U6065 (N_6065,N_5735,N_5503);
nand U6066 (N_6066,N_5597,N_5769);
nor U6067 (N_6067,N_5672,N_5653);
nand U6068 (N_6068,N_5776,N_5879);
nand U6069 (N_6069,N_5697,N_5551);
or U6070 (N_6070,N_5635,N_5811);
nor U6071 (N_6071,N_5542,N_5555);
nand U6072 (N_6072,N_5935,N_5910);
or U6073 (N_6073,N_5593,N_5875);
xor U6074 (N_6074,N_5569,N_5667);
nor U6075 (N_6075,N_5895,N_5548);
nor U6076 (N_6076,N_5970,N_5631);
nand U6077 (N_6077,N_5537,N_5749);
nor U6078 (N_6078,N_5736,N_5645);
nor U6079 (N_6079,N_5932,N_5893);
xnor U6080 (N_6080,N_5991,N_5866);
nor U6081 (N_6081,N_5532,N_5741);
nand U6082 (N_6082,N_5662,N_5874);
and U6083 (N_6083,N_5716,N_5900);
and U6084 (N_6084,N_5976,N_5892);
and U6085 (N_6085,N_5817,N_5782);
or U6086 (N_6086,N_5982,N_5836);
or U6087 (N_6087,N_5595,N_5822);
xnor U6088 (N_6088,N_5643,N_5578);
nand U6089 (N_6089,N_5625,N_5760);
nor U6090 (N_6090,N_5714,N_5964);
or U6091 (N_6091,N_5624,N_5564);
nor U6092 (N_6092,N_5989,N_5915);
or U6093 (N_6093,N_5727,N_5558);
nor U6094 (N_6094,N_5612,N_5701);
or U6095 (N_6095,N_5694,N_5592);
and U6096 (N_6096,N_5607,N_5871);
or U6097 (N_6097,N_5768,N_5752);
and U6098 (N_6098,N_5617,N_5832);
xnor U6099 (N_6099,N_5544,N_5523);
nor U6100 (N_6100,N_5522,N_5547);
xor U6101 (N_6101,N_5825,N_5804);
nor U6102 (N_6102,N_5799,N_5784);
or U6103 (N_6103,N_5975,N_5772);
and U6104 (N_6104,N_5693,N_5897);
and U6105 (N_6105,N_5774,N_5923);
and U6106 (N_6106,N_5944,N_5658);
nand U6107 (N_6107,N_5830,N_5967);
xnor U6108 (N_6108,N_5849,N_5605);
or U6109 (N_6109,N_5673,N_5820);
nor U6110 (N_6110,N_5968,N_5733);
and U6111 (N_6111,N_5606,N_5985);
xnor U6112 (N_6112,N_5587,N_5510);
nand U6113 (N_6113,N_5566,N_5813);
nor U6114 (N_6114,N_5559,N_5512);
nand U6115 (N_6115,N_5660,N_5890);
nor U6116 (N_6116,N_5591,N_5980);
nor U6117 (N_6117,N_5831,N_5757);
or U6118 (N_6118,N_5930,N_5646);
xnor U6119 (N_6119,N_5807,N_5763);
or U6120 (N_6120,N_5922,N_5933);
and U6121 (N_6121,N_5695,N_5958);
and U6122 (N_6122,N_5634,N_5792);
nor U6123 (N_6123,N_5983,N_5710);
nand U6124 (N_6124,N_5740,N_5821);
xor U6125 (N_6125,N_5602,N_5801);
nand U6126 (N_6126,N_5858,N_5926);
and U6127 (N_6127,N_5561,N_5824);
nand U6128 (N_6128,N_5618,N_5581);
or U6129 (N_6129,N_5517,N_5845);
or U6130 (N_6130,N_5988,N_5584);
nand U6131 (N_6131,N_5580,N_5528);
nand U6132 (N_6132,N_5867,N_5686);
or U6133 (N_6133,N_5857,N_5683);
nand U6134 (N_6134,N_5670,N_5790);
nand U6135 (N_6135,N_5654,N_5565);
nand U6136 (N_6136,N_5725,N_5553);
and U6137 (N_6137,N_5947,N_5914);
nor U6138 (N_6138,N_5626,N_5709);
and U6139 (N_6139,N_5570,N_5868);
and U6140 (N_6140,N_5627,N_5909);
nand U6141 (N_6141,N_5508,N_5770);
nor U6142 (N_6142,N_5705,N_5974);
and U6143 (N_6143,N_5539,N_5853);
xnor U6144 (N_6144,N_5920,N_5755);
nand U6145 (N_6145,N_5734,N_5977);
nand U6146 (N_6146,N_5540,N_5579);
nand U6147 (N_6147,N_5744,N_5610);
and U6148 (N_6148,N_5885,N_5951);
and U6149 (N_6149,N_5894,N_5629);
nand U6150 (N_6150,N_5812,N_5961);
nand U6151 (N_6151,N_5877,N_5855);
or U6152 (N_6152,N_5838,N_5883);
and U6153 (N_6153,N_5640,N_5916);
nand U6154 (N_6154,N_5675,N_5516);
xnor U6155 (N_6155,N_5679,N_5687);
nor U6156 (N_6156,N_5795,N_5722);
or U6157 (N_6157,N_5657,N_5878);
and U6158 (N_6158,N_5963,N_5850);
nor U6159 (N_6159,N_5604,N_5903);
or U6160 (N_6160,N_5514,N_5729);
xor U6161 (N_6161,N_5632,N_5765);
xnor U6162 (N_6162,N_5904,N_5759);
nor U6163 (N_6163,N_5841,N_5919);
nand U6164 (N_6164,N_5954,N_5509);
xor U6165 (N_6165,N_5862,N_5789);
nor U6166 (N_6166,N_5712,N_5997);
nor U6167 (N_6167,N_5937,N_5959);
nand U6168 (N_6168,N_5940,N_5833);
nand U6169 (N_6169,N_5882,N_5753);
or U6170 (N_6170,N_5590,N_5689);
nor U6171 (N_6171,N_5928,N_5549);
xnor U6172 (N_6172,N_5794,N_5637);
and U6173 (N_6173,N_5956,N_5851);
nand U6174 (N_6174,N_5931,N_5828);
and U6175 (N_6175,N_5775,N_5805);
and U6176 (N_6176,N_5572,N_5525);
xor U6177 (N_6177,N_5886,N_5609);
xnor U6178 (N_6178,N_5620,N_5834);
or U6179 (N_6179,N_5987,N_5737);
or U6180 (N_6180,N_5538,N_5628);
and U6181 (N_6181,N_5533,N_5948);
nor U6182 (N_6182,N_5780,N_5674);
or U6183 (N_6183,N_5502,N_5613);
or U6184 (N_6184,N_5526,N_5927);
nor U6185 (N_6185,N_5552,N_5766);
or U6186 (N_6186,N_5639,N_5518);
nor U6187 (N_6187,N_5583,N_5728);
nand U6188 (N_6188,N_5615,N_5918);
nor U6189 (N_6189,N_5840,N_5659);
or U6190 (N_6190,N_5545,N_5668);
xnor U6191 (N_6191,N_5699,N_5906);
nor U6192 (N_6192,N_5788,N_5891);
nor U6193 (N_6193,N_5887,N_5743);
nand U6194 (N_6194,N_5711,N_5949);
or U6195 (N_6195,N_5929,N_5873);
and U6196 (N_6196,N_5723,N_5960);
nor U6197 (N_6197,N_5842,N_5732);
and U6198 (N_6198,N_5611,N_5859);
nor U6199 (N_6199,N_5636,N_5600);
nand U6200 (N_6200,N_5787,N_5888);
and U6201 (N_6201,N_5678,N_5884);
xor U6202 (N_6202,N_5505,N_5520);
or U6203 (N_6203,N_5934,N_5797);
nand U6204 (N_6204,N_5724,N_5726);
xnor U6205 (N_6205,N_5957,N_5962);
and U6206 (N_6206,N_5986,N_5758);
nor U6207 (N_6207,N_5762,N_5870);
and U6208 (N_6208,N_5971,N_5952);
or U6209 (N_6209,N_5783,N_5800);
or U6210 (N_6210,N_5677,N_5936);
nand U6211 (N_6211,N_5925,N_5568);
nand U6212 (N_6212,N_5656,N_5984);
or U6213 (N_6213,N_5911,N_5642);
and U6214 (N_6214,N_5764,N_5880);
nand U6215 (N_6215,N_5536,N_5573);
and U6216 (N_6216,N_5713,N_5912);
and U6217 (N_6217,N_5945,N_5869);
and U6218 (N_6218,N_5633,N_5844);
nand U6219 (N_6219,N_5571,N_5622);
nor U6220 (N_6220,N_5864,N_5719);
and U6221 (N_6221,N_5779,N_5829);
and U6222 (N_6222,N_5896,N_5524);
xnor U6223 (N_6223,N_5661,N_5623);
nor U6224 (N_6224,N_5856,N_5649);
xnor U6225 (N_6225,N_5854,N_5608);
nand U6226 (N_6226,N_5700,N_5603);
or U6227 (N_6227,N_5506,N_5771);
and U6228 (N_6228,N_5546,N_5543);
xor U6229 (N_6229,N_5691,N_5818);
and U6230 (N_6230,N_5950,N_5972);
nor U6231 (N_6231,N_5534,N_5599);
xor U6232 (N_6232,N_5861,N_5754);
and U6233 (N_6233,N_5582,N_5527);
and U6234 (N_6234,N_5938,N_5969);
and U6235 (N_6235,N_5773,N_5837);
xor U6236 (N_6236,N_5943,N_5720);
xnor U6237 (N_6237,N_5648,N_5999);
nor U6238 (N_6238,N_5594,N_5521);
and U6239 (N_6239,N_5815,N_5638);
nor U6240 (N_6240,N_5652,N_5703);
xor U6241 (N_6241,N_5889,N_5860);
and U6242 (N_6242,N_5973,N_5651);
nor U6243 (N_6243,N_5541,N_5554);
nand U6244 (N_6244,N_5786,N_5848);
xnor U6245 (N_6245,N_5685,N_5846);
nand U6246 (N_6246,N_5810,N_5692);
nor U6247 (N_6247,N_5992,N_5826);
nor U6248 (N_6248,N_5500,N_5680);
nand U6249 (N_6249,N_5921,N_5682);
or U6250 (N_6250,N_5552,N_5972);
xnor U6251 (N_6251,N_5821,N_5716);
or U6252 (N_6252,N_5993,N_5938);
nor U6253 (N_6253,N_5598,N_5926);
and U6254 (N_6254,N_5966,N_5947);
and U6255 (N_6255,N_5684,N_5588);
or U6256 (N_6256,N_5616,N_5946);
or U6257 (N_6257,N_5871,N_5792);
or U6258 (N_6258,N_5806,N_5738);
nor U6259 (N_6259,N_5598,N_5893);
nor U6260 (N_6260,N_5611,N_5630);
nand U6261 (N_6261,N_5662,N_5872);
nand U6262 (N_6262,N_5833,N_5627);
and U6263 (N_6263,N_5912,N_5893);
nand U6264 (N_6264,N_5791,N_5775);
and U6265 (N_6265,N_5640,N_5590);
nor U6266 (N_6266,N_5746,N_5689);
or U6267 (N_6267,N_5646,N_5733);
nand U6268 (N_6268,N_5840,N_5578);
nor U6269 (N_6269,N_5947,N_5888);
nand U6270 (N_6270,N_5677,N_5527);
nor U6271 (N_6271,N_5514,N_5972);
xnor U6272 (N_6272,N_5680,N_5954);
or U6273 (N_6273,N_5650,N_5845);
nand U6274 (N_6274,N_5808,N_5888);
and U6275 (N_6275,N_5633,N_5724);
nor U6276 (N_6276,N_5962,N_5921);
nor U6277 (N_6277,N_5632,N_5987);
nor U6278 (N_6278,N_5795,N_5993);
nor U6279 (N_6279,N_5512,N_5722);
nor U6280 (N_6280,N_5641,N_5820);
and U6281 (N_6281,N_5869,N_5517);
nor U6282 (N_6282,N_5597,N_5972);
xnor U6283 (N_6283,N_5557,N_5650);
nand U6284 (N_6284,N_5665,N_5503);
xnor U6285 (N_6285,N_5518,N_5793);
and U6286 (N_6286,N_5925,N_5688);
nor U6287 (N_6287,N_5837,N_5642);
xnor U6288 (N_6288,N_5899,N_5584);
or U6289 (N_6289,N_5806,N_5645);
nor U6290 (N_6290,N_5620,N_5617);
nand U6291 (N_6291,N_5896,N_5651);
nor U6292 (N_6292,N_5812,N_5535);
nor U6293 (N_6293,N_5739,N_5660);
nor U6294 (N_6294,N_5791,N_5576);
xnor U6295 (N_6295,N_5907,N_5871);
or U6296 (N_6296,N_5989,N_5604);
xor U6297 (N_6297,N_5803,N_5839);
and U6298 (N_6298,N_5712,N_5730);
or U6299 (N_6299,N_5653,N_5830);
nor U6300 (N_6300,N_5636,N_5638);
nor U6301 (N_6301,N_5923,N_5610);
or U6302 (N_6302,N_5728,N_5812);
xnor U6303 (N_6303,N_5995,N_5998);
nor U6304 (N_6304,N_5544,N_5539);
or U6305 (N_6305,N_5539,N_5943);
or U6306 (N_6306,N_5998,N_5892);
nor U6307 (N_6307,N_5637,N_5822);
xor U6308 (N_6308,N_5961,N_5983);
and U6309 (N_6309,N_5755,N_5922);
nand U6310 (N_6310,N_5816,N_5965);
or U6311 (N_6311,N_5755,N_5618);
and U6312 (N_6312,N_5993,N_5767);
xor U6313 (N_6313,N_5596,N_5733);
and U6314 (N_6314,N_5639,N_5726);
nand U6315 (N_6315,N_5641,N_5729);
xor U6316 (N_6316,N_5517,N_5745);
or U6317 (N_6317,N_5903,N_5742);
and U6318 (N_6318,N_5804,N_5712);
or U6319 (N_6319,N_5728,N_5776);
nor U6320 (N_6320,N_5890,N_5982);
nor U6321 (N_6321,N_5880,N_5507);
xor U6322 (N_6322,N_5543,N_5908);
nor U6323 (N_6323,N_5894,N_5707);
nand U6324 (N_6324,N_5840,N_5746);
xnor U6325 (N_6325,N_5511,N_5833);
and U6326 (N_6326,N_5687,N_5551);
nor U6327 (N_6327,N_5676,N_5636);
nor U6328 (N_6328,N_5706,N_5586);
xnor U6329 (N_6329,N_5774,N_5816);
nand U6330 (N_6330,N_5853,N_5585);
nand U6331 (N_6331,N_5581,N_5526);
xor U6332 (N_6332,N_5546,N_5640);
xor U6333 (N_6333,N_5635,N_5646);
or U6334 (N_6334,N_5703,N_5805);
xnor U6335 (N_6335,N_5667,N_5985);
nor U6336 (N_6336,N_5924,N_5548);
nor U6337 (N_6337,N_5681,N_5989);
xnor U6338 (N_6338,N_5596,N_5753);
nor U6339 (N_6339,N_5532,N_5659);
nor U6340 (N_6340,N_5662,N_5821);
xnor U6341 (N_6341,N_5668,N_5801);
nand U6342 (N_6342,N_5861,N_5908);
nand U6343 (N_6343,N_5706,N_5638);
nand U6344 (N_6344,N_5529,N_5910);
nor U6345 (N_6345,N_5768,N_5869);
nand U6346 (N_6346,N_5553,N_5597);
or U6347 (N_6347,N_5966,N_5618);
nand U6348 (N_6348,N_5885,N_5847);
and U6349 (N_6349,N_5606,N_5555);
xnor U6350 (N_6350,N_5515,N_5702);
nand U6351 (N_6351,N_5642,N_5822);
and U6352 (N_6352,N_5854,N_5686);
nor U6353 (N_6353,N_5834,N_5719);
or U6354 (N_6354,N_5857,N_5694);
nand U6355 (N_6355,N_5732,N_5521);
xor U6356 (N_6356,N_5923,N_5689);
xor U6357 (N_6357,N_5994,N_5582);
nor U6358 (N_6358,N_5811,N_5839);
nor U6359 (N_6359,N_5555,N_5547);
or U6360 (N_6360,N_5989,N_5804);
nand U6361 (N_6361,N_5938,N_5888);
and U6362 (N_6362,N_5559,N_5749);
or U6363 (N_6363,N_5649,N_5952);
nor U6364 (N_6364,N_5895,N_5539);
nor U6365 (N_6365,N_5721,N_5666);
nand U6366 (N_6366,N_5603,N_5673);
xor U6367 (N_6367,N_5762,N_5734);
or U6368 (N_6368,N_5611,N_5641);
and U6369 (N_6369,N_5527,N_5983);
xnor U6370 (N_6370,N_5648,N_5581);
or U6371 (N_6371,N_5833,N_5925);
or U6372 (N_6372,N_5642,N_5525);
nor U6373 (N_6373,N_5847,N_5729);
xor U6374 (N_6374,N_5737,N_5609);
and U6375 (N_6375,N_5511,N_5618);
xor U6376 (N_6376,N_5554,N_5888);
and U6377 (N_6377,N_5611,N_5915);
and U6378 (N_6378,N_5638,N_5926);
and U6379 (N_6379,N_5838,N_5666);
nor U6380 (N_6380,N_5617,N_5754);
nor U6381 (N_6381,N_5744,N_5984);
nor U6382 (N_6382,N_5541,N_5629);
and U6383 (N_6383,N_5540,N_5673);
xor U6384 (N_6384,N_5663,N_5697);
or U6385 (N_6385,N_5558,N_5963);
nor U6386 (N_6386,N_5844,N_5810);
nor U6387 (N_6387,N_5919,N_5924);
nand U6388 (N_6388,N_5874,N_5714);
nand U6389 (N_6389,N_5713,N_5632);
nand U6390 (N_6390,N_5909,N_5609);
nand U6391 (N_6391,N_5702,N_5634);
xor U6392 (N_6392,N_5812,N_5510);
or U6393 (N_6393,N_5678,N_5608);
xnor U6394 (N_6394,N_5781,N_5603);
and U6395 (N_6395,N_5796,N_5881);
or U6396 (N_6396,N_5953,N_5598);
xor U6397 (N_6397,N_5888,N_5575);
and U6398 (N_6398,N_5559,N_5744);
xor U6399 (N_6399,N_5762,N_5667);
and U6400 (N_6400,N_5630,N_5987);
or U6401 (N_6401,N_5601,N_5694);
or U6402 (N_6402,N_5972,N_5789);
or U6403 (N_6403,N_5563,N_5824);
xor U6404 (N_6404,N_5665,N_5816);
nand U6405 (N_6405,N_5846,N_5970);
nor U6406 (N_6406,N_5836,N_5741);
nor U6407 (N_6407,N_5954,N_5994);
nor U6408 (N_6408,N_5977,N_5644);
nor U6409 (N_6409,N_5713,N_5726);
xor U6410 (N_6410,N_5698,N_5828);
or U6411 (N_6411,N_5608,N_5719);
or U6412 (N_6412,N_5935,N_5591);
or U6413 (N_6413,N_5728,N_5677);
nor U6414 (N_6414,N_5757,N_5952);
and U6415 (N_6415,N_5874,N_5655);
or U6416 (N_6416,N_5787,N_5617);
nor U6417 (N_6417,N_5833,N_5567);
and U6418 (N_6418,N_5748,N_5995);
xor U6419 (N_6419,N_5872,N_5824);
or U6420 (N_6420,N_5533,N_5747);
or U6421 (N_6421,N_5945,N_5515);
and U6422 (N_6422,N_5972,N_5630);
or U6423 (N_6423,N_5743,N_5978);
nor U6424 (N_6424,N_5634,N_5946);
xnor U6425 (N_6425,N_5908,N_5789);
and U6426 (N_6426,N_5670,N_5805);
or U6427 (N_6427,N_5609,N_5612);
xor U6428 (N_6428,N_5968,N_5609);
or U6429 (N_6429,N_5784,N_5720);
nor U6430 (N_6430,N_5782,N_5707);
or U6431 (N_6431,N_5862,N_5513);
xor U6432 (N_6432,N_5996,N_5842);
xnor U6433 (N_6433,N_5814,N_5543);
and U6434 (N_6434,N_5778,N_5941);
and U6435 (N_6435,N_5752,N_5553);
xor U6436 (N_6436,N_5942,N_5664);
xnor U6437 (N_6437,N_5856,N_5717);
and U6438 (N_6438,N_5899,N_5530);
nor U6439 (N_6439,N_5653,N_5708);
xnor U6440 (N_6440,N_5557,N_5698);
or U6441 (N_6441,N_5716,N_5803);
and U6442 (N_6442,N_5677,N_5615);
nand U6443 (N_6443,N_5646,N_5919);
nor U6444 (N_6444,N_5542,N_5826);
xor U6445 (N_6445,N_5536,N_5647);
xor U6446 (N_6446,N_5536,N_5564);
or U6447 (N_6447,N_5662,N_5537);
or U6448 (N_6448,N_5883,N_5654);
nand U6449 (N_6449,N_5846,N_5895);
xor U6450 (N_6450,N_5569,N_5992);
xor U6451 (N_6451,N_5908,N_5825);
nand U6452 (N_6452,N_5528,N_5623);
or U6453 (N_6453,N_5835,N_5937);
nand U6454 (N_6454,N_5761,N_5800);
xor U6455 (N_6455,N_5731,N_5854);
or U6456 (N_6456,N_5716,N_5599);
xor U6457 (N_6457,N_5756,N_5993);
and U6458 (N_6458,N_5905,N_5702);
xor U6459 (N_6459,N_5650,N_5778);
xor U6460 (N_6460,N_5728,N_5991);
xnor U6461 (N_6461,N_5804,N_5597);
or U6462 (N_6462,N_5803,N_5722);
and U6463 (N_6463,N_5968,N_5933);
nor U6464 (N_6464,N_5524,N_5996);
xnor U6465 (N_6465,N_5786,N_5695);
nor U6466 (N_6466,N_5613,N_5665);
and U6467 (N_6467,N_5842,N_5828);
nand U6468 (N_6468,N_5894,N_5607);
nor U6469 (N_6469,N_5660,N_5849);
or U6470 (N_6470,N_5781,N_5521);
xnor U6471 (N_6471,N_5910,N_5738);
xnor U6472 (N_6472,N_5864,N_5949);
nor U6473 (N_6473,N_5866,N_5785);
xor U6474 (N_6474,N_5569,N_5577);
and U6475 (N_6475,N_5858,N_5841);
nor U6476 (N_6476,N_5864,N_5542);
nor U6477 (N_6477,N_5917,N_5785);
xor U6478 (N_6478,N_5524,N_5642);
nor U6479 (N_6479,N_5677,N_5693);
and U6480 (N_6480,N_5979,N_5737);
xnor U6481 (N_6481,N_5601,N_5548);
nor U6482 (N_6482,N_5805,N_5711);
or U6483 (N_6483,N_5734,N_5957);
or U6484 (N_6484,N_5565,N_5687);
nor U6485 (N_6485,N_5559,N_5636);
xor U6486 (N_6486,N_5937,N_5607);
or U6487 (N_6487,N_5906,N_5511);
xnor U6488 (N_6488,N_5647,N_5546);
xor U6489 (N_6489,N_5846,N_5560);
nor U6490 (N_6490,N_5842,N_5888);
nand U6491 (N_6491,N_5543,N_5753);
and U6492 (N_6492,N_5986,N_5544);
xnor U6493 (N_6493,N_5995,N_5773);
xnor U6494 (N_6494,N_5631,N_5509);
and U6495 (N_6495,N_5808,N_5908);
and U6496 (N_6496,N_5871,N_5764);
or U6497 (N_6497,N_5669,N_5745);
or U6498 (N_6498,N_5867,N_5703);
and U6499 (N_6499,N_5962,N_5994);
nor U6500 (N_6500,N_6308,N_6361);
nor U6501 (N_6501,N_6267,N_6149);
nand U6502 (N_6502,N_6192,N_6303);
or U6503 (N_6503,N_6489,N_6274);
nand U6504 (N_6504,N_6398,N_6029);
and U6505 (N_6505,N_6105,N_6247);
nand U6506 (N_6506,N_6455,N_6169);
nor U6507 (N_6507,N_6285,N_6134);
nand U6508 (N_6508,N_6337,N_6334);
and U6509 (N_6509,N_6041,N_6325);
nor U6510 (N_6510,N_6477,N_6332);
nor U6511 (N_6511,N_6025,N_6208);
nand U6512 (N_6512,N_6184,N_6294);
nand U6513 (N_6513,N_6392,N_6403);
nor U6514 (N_6514,N_6474,N_6152);
nor U6515 (N_6515,N_6087,N_6142);
xnor U6516 (N_6516,N_6250,N_6141);
nor U6517 (N_6517,N_6352,N_6387);
or U6518 (N_6518,N_6461,N_6377);
and U6519 (N_6519,N_6256,N_6206);
nor U6520 (N_6520,N_6435,N_6408);
and U6521 (N_6521,N_6157,N_6222);
nor U6522 (N_6522,N_6335,N_6226);
or U6523 (N_6523,N_6227,N_6073);
nand U6524 (N_6524,N_6101,N_6490);
xnor U6525 (N_6525,N_6263,N_6357);
xnor U6526 (N_6526,N_6478,N_6014);
nand U6527 (N_6527,N_6124,N_6034);
and U6528 (N_6528,N_6322,N_6447);
and U6529 (N_6529,N_6200,N_6004);
or U6530 (N_6530,N_6238,N_6095);
xor U6531 (N_6531,N_6363,N_6453);
nor U6532 (N_6532,N_6156,N_6469);
and U6533 (N_6533,N_6016,N_6472);
or U6534 (N_6534,N_6211,N_6033);
nor U6535 (N_6535,N_6243,N_6348);
xnor U6536 (N_6536,N_6049,N_6317);
or U6537 (N_6537,N_6107,N_6329);
xor U6538 (N_6538,N_6046,N_6019);
or U6539 (N_6539,N_6465,N_6341);
xnor U6540 (N_6540,N_6000,N_6035);
or U6541 (N_6541,N_6289,N_6082);
nand U6542 (N_6542,N_6462,N_6264);
or U6543 (N_6543,N_6383,N_6281);
xnor U6544 (N_6544,N_6470,N_6072);
nor U6545 (N_6545,N_6475,N_6254);
xor U6546 (N_6546,N_6103,N_6224);
xnor U6547 (N_6547,N_6452,N_6305);
or U6548 (N_6548,N_6297,N_6321);
or U6549 (N_6549,N_6293,N_6020);
or U6550 (N_6550,N_6189,N_6396);
and U6551 (N_6551,N_6302,N_6018);
nor U6552 (N_6552,N_6468,N_6121);
or U6553 (N_6553,N_6246,N_6145);
xnor U6554 (N_6554,N_6088,N_6032);
or U6555 (N_6555,N_6052,N_6413);
or U6556 (N_6556,N_6058,N_6292);
nand U6557 (N_6557,N_6146,N_6439);
or U6558 (N_6558,N_6013,N_6440);
nor U6559 (N_6559,N_6295,N_6170);
xnor U6560 (N_6560,N_6151,N_6111);
or U6561 (N_6561,N_6318,N_6068);
and U6562 (N_6562,N_6282,N_6312);
xor U6563 (N_6563,N_6081,N_6315);
and U6564 (N_6564,N_6060,N_6296);
xor U6565 (N_6565,N_6327,N_6011);
or U6566 (N_6566,N_6093,N_6045);
nor U6567 (N_6567,N_6126,N_6055);
and U6568 (N_6568,N_6009,N_6075);
nor U6569 (N_6569,N_6323,N_6186);
xnor U6570 (N_6570,N_6023,N_6185);
nand U6571 (N_6571,N_6333,N_6017);
and U6572 (N_6572,N_6027,N_6313);
or U6573 (N_6573,N_6493,N_6098);
and U6574 (N_6574,N_6195,N_6420);
nand U6575 (N_6575,N_6070,N_6172);
nor U6576 (N_6576,N_6237,N_6100);
nand U6577 (N_6577,N_6171,N_6063);
or U6578 (N_6578,N_6405,N_6175);
xor U6579 (N_6579,N_6492,N_6221);
nand U6580 (N_6580,N_6343,N_6463);
nor U6581 (N_6581,N_6319,N_6411);
nor U6582 (N_6582,N_6402,N_6300);
nand U6583 (N_6583,N_6229,N_6448);
nor U6584 (N_6584,N_6030,N_6154);
nand U6585 (N_6585,N_6129,N_6194);
and U6586 (N_6586,N_6230,N_6301);
nand U6587 (N_6587,N_6057,N_6407);
xor U6588 (N_6588,N_6132,N_6487);
xnor U6589 (N_6589,N_6048,N_6373);
nand U6590 (N_6590,N_6260,N_6423);
and U6591 (N_6591,N_6241,N_6012);
and U6592 (N_6592,N_6372,N_6273);
nand U6593 (N_6593,N_6473,N_6164);
nand U6594 (N_6594,N_6181,N_6066);
nor U6595 (N_6595,N_6042,N_6061);
nor U6596 (N_6596,N_6064,N_6249);
nand U6597 (N_6597,N_6133,N_6174);
and U6598 (N_6598,N_6375,N_6366);
nand U6599 (N_6599,N_6140,N_6476);
nor U6600 (N_6600,N_6320,N_6210);
xnor U6601 (N_6601,N_6094,N_6307);
and U6602 (N_6602,N_6125,N_6257);
or U6603 (N_6603,N_6284,N_6338);
and U6604 (N_6604,N_6431,N_6457);
and U6605 (N_6605,N_6397,N_6147);
nand U6606 (N_6606,N_6450,N_6117);
nor U6607 (N_6607,N_6481,N_6427);
nand U6608 (N_6608,N_6443,N_6269);
or U6609 (N_6609,N_6122,N_6110);
and U6610 (N_6610,N_6436,N_6471);
xor U6611 (N_6611,N_6374,N_6432);
or U6612 (N_6612,N_6090,N_6074);
and U6613 (N_6613,N_6173,N_6351);
or U6614 (N_6614,N_6022,N_6127);
xor U6615 (N_6615,N_6054,N_6290);
nor U6616 (N_6616,N_6008,N_6415);
xnor U6617 (N_6617,N_6028,N_6182);
and U6618 (N_6618,N_6135,N_6245);
xor U6619 (N_6619,N_6342,N_6310);
xor U6620 (N_6620,N_6119,N_6116);
nor U6621 (N_6621,N_6118,N_6409);
or U6622 (N_6622,N_6092,N_6456);
and U6623 (N_6623,N_6442,N_6165);
nor U6624 (N_6624,N_6039,N_6161);
nor U6625 (N_6625,N_6421,N_6038);
nor U6626 (N_6626,N_6277,N_6316);
and U6627 (N_6627,N_6414,N_6369);
or U6628 (N_6628,N_6219,N_6143);
or U6629 (N_6629,N_6479,N_6429);
and U6630 (N_6630,N_6158,N_6445);
nor U6631 (N_6631,N_6364,N_6391);
nand U6632 (N_6632,N_6040,N_6202);
and U6633 (N_6633,N_6144,N_6314);
and U6634 (N_6634,N_6253,N_6123);
nand U6635 (N_6635,N_6497,N_6089);
xor U6636 (N_6636,N_6485,N_6252);
nor U6637 (N_6637,N_6278,N_6036);
nand U6638 (N_6638,N_6499,N_6336);
nor U6639 (N_6639,N_6166,N_6390);
or U6640 (N_6640,N_6113,N_6153);
nand U6641 (N_6641,N_6223,N_6083);
or U6642 (N_6642,N_6464,N_6261);
and U6643 (N_6643,N_6367,N_6215);
and U6644 (N_6644,N_6422,N_6370);
and U6645 (N_6645,N_6104,N_6137);
nand U6646 (N_6646,N_6276,N_6044);
nand U6647 (N_6647,N_6209,N_6214);
xor U6648 (N_6648,N_6388,N_6062);
and U6649 (N_6649,N_6109,N_6031);
xnor U6650 (N_6650,N_6395,N_6394);
nor U6651 (N_6651,N_6309,N_6015);
or U6652 (N_6652,N_6085,N_6371);
nor U6653 (N_6653,N_6380,N_6003);
or U6654 (N_6654,N_6483,N_6345);
nor U6655 (N_6655,N_6331,N_6356);
nand U6656 (N_6656,N_6242,N_6212);
and U6657 (N_6657,N_6024,N_6159);
nand U6658 (N_6658,N_6381,N_6437);
nor U6659 (N_6659,N_6433,N_6205);
nand U6660 (N_6660,N_6270,N_6287);
or U6661 (N_6661,N_6275,N_6418);
and U6662 (N_6662,N_6138,N_6393);
or U6663 (N_6663,N_6136,N_6271);
and U6664 (N_6664,N_6350,N_6163);
or U6665 (N_6665,N_6291,N_6071);
and U6666 (N_6666,N_6021,N_6339);
nor U6667 (N_6667,N_6444,N_6176);
xor U6668 (N_6668,N_6378,N_6076);
or U6669 (N_6669,N_6106,N_6262);
or U6670 (N_6670,N_6283,N_6449);
xnor U6671 (N_6671,N_6428,N_6235);
and U6672 (N_6672,N_6268,N_6196);
nor U6673 (N_6673,N_6178,N_6412);
and U6674 (N_6674,N_6162,N_6150);
nand U6675 (N_6675,N_6078,N_6426);
xor U6676 (N_6676,N_6239,N_6197);
xnor U6677 (N_6677,N_6346,N_6096);
and U6678 (N_6678,N_6179,N_6190);
xor U6679 (N_6679,N_6494,N_6099);
xnor U6680 (N_6680,N_6353,N_6191);
and U6681 (N_6681,N_6005,N_6037);
nand U6682 (N_6682,N_6486,N_6446);
and U6683 (N_6683,N_6458,N_6355);
and U6684 (N_6684,N_6059,N_6386);
nand U6685 (N_6685,N_6160,N_6244);
or U6686 (N_6686,N_6399,N_6410);
xor U6687 (N_6687,N_6139,N_6376);
or U6688 (N_6688,N_6177,N_6077);
nand U6689 (N_6689,N_6183,N_6401);
and U6690 (N_6690,N_6467,N_6091);
nand U6691 (N_6691,N_6199,N_6218);
and U6692 (N_6692,N_6203,N_6050);
or U6693 (N_6693,N_6299,N_6417);
nand U6694 (N_6694,N_6451,N_6220);
and U6695 (N_6695,N_6404,N_6259);
nand U6696 (N_6696,N_6347,N_6498);
xor U6697 (N_6697,N_6384,N_6382);
and U6698 (N_6698,N_6217,N_6187);
xor U6699 (N_6699,N_6349,N_6488);
nor U6700 (N_6700,N_6379,N_6438);
nand U6701 (N_6701,N_6288,N_6459);
xor U6702 (N_6702,N_6047,N_6360);
xor U6703 (N_6703,N_6010,N_6430);
and U6704 (N_6704,N_6280,N_6051);
nor U6705 (N_6705,N_6067,N_6255);
nand U6706 (N_6706,N_6080,N_6419);
and U6707 (N_6707,N_6201,N_6265);
xor U6708 (N_6708,N_6007,N_6006);
nor U6709 (N_6709,N_6495,N_6326);
nor U6710 (N_6710,N_6228,N_6168);
nand U6711 (N_6711,N_6359,N_6454);
and U6712 (N_6712,N_6155,N_6231);
nand U6713 (N_6713,N_6114,N_6354);
nor U6714 (N_6714,N_6416,N_6328);
nor U6715 (N_6715,N_6258,N_6365);
or U6716 (N_6716,N_6102,N_6198);
xor U6717 (N_6717,N_6460,N_6232);
nand U6718 (N_6718,N_6484,N_6188);
xor U6719 (N_6719,N_6233,N_6400);
and U6720 (N_6720,N_6112,N_6148);
and U6721 (N_6721,N_6385,N_6079);
xnor U6722 (N_6722,N_6491,N_6425);
and U6723 (N_6723,N_6266,N_6234);
or U6724 (N_6724,N_6434,N_6108);
nor U6725 (N_6725,N_6368,N_6207);
xnor U6726 (N_6726,N_6306,N_6389);
and U6727 (N_6727,N_6279,N_6424);
xor U6728 (N_6728,N_6358,N_6496);
nand U6729 (N_6729,N_6340,N_6406);
and U6730 (N_6730,N_6120,N_6286);
or U6731 (N_6731,N_6311,N_6130);
nand U6732 (N_6732,N_6272,N_6056);
xnor U6733 (N_6733,N_6236,N_6240);
or U6734 (N_6734,N_6131,N_6086);
or U6735 (N_6735,N_6330,N_6441);
and U6736 (N_6736,N_6298,N_6002);
xnor U6737 (N_6737,N_6482,N_6480);
nor U6738 (N_6738,N_6053,N_6084);
and U6739 (N_6739,N_6204,N_6216);
xor U6740 (N_6740,N_6069,N_6362);
nand U6741 (N_6741,N_6213,N_6180);
or U6742 (N_6742,N_6065,N_6043);
nand U6743 (N_6743,N_6466,N_6128);
nor U6744 (N_6744,N_6304,N_6225);
and U6745 (N_6745,N_6251,N_6344);
xor U6746 (N_6746,N_6026,N_6324);
xnor U6747 (N_6747,N_6167,N_6193);
xnor U6748 (N_6748,N_6001,N_6097);
and U6749 (N_6749,N_6115,N_6248);
nor U6750 (N_6750,N_6015,N_6358);
nor U6751 (N_6751,N_6172,N_6246);
nor U6752 (N_6752,N_6172,N_6237);
and U6753 (N_6753,N_6170,N_6015);
xnor U6754 (N_6754,N_6277,N_6162);
and U6755 (N_6755,N_6034,N_6126);
xor U6756 (N_6756,N_6079,N_6433);
xnor U6757 (N_6757,N_6429,N_6008);
nor U6758 (N_6758,N_6047,N_6474);
and U6759 (N_6759,N_6470,N_6407);
and U6760 (N_6760,N_6028,N_6461);
or U6761 (N_6761,N_6001,N_6161);
nand U6762 (N_6762,N_6211,N_6278);
nor U6763 (N_6763,N_6068,N_6239);
and U6764 (N_6764,N_6209,N_6205);
xnor U6765 (N_6765,N_6463,N_6065);
nor U6766 (N_6766,N_6070,N_6237);
or U6767 (N_6767,N_6404,N_6346);
nor U6768 (N_6768,N_6111,N_6428);
xor U6769 (N_6769,N_6373,N_6093);
nor U6770 (N_6770,N_6055,N_6148);
nand U6771 (N_6771,N_6384,N_6120);
xnor U6772 (N_6772,N_6268,N_6191);
nand U6773 (N_6773,N_6056,N_6430);
xor U6774 (N_6774,N_6110,N_6298);
xnor U6775 (N_6775,N_6233,N_6106);
or U6776 (N_6776,N_6383,N_6325);
xnor U6777 (N_6777,N_6045,N_6076);
nor U6778 (N_6778,N_6372,N_6247);
or U6779 (N_6779,N_6210,N_6319);
and U6780 (N_6780,N_6208,N_6262);
nor U6781 (N_6781,N_6031,N_6389);
nand U6782 (N_6782,N_6251,N_6254);
nand U6783 (N_6783,N_6097,N_6312);
nand U6784 (N_6784,N_6490,N_6311);
or U6785 (N_6785,N_6195,N_6243);
nor U6786 (N_6786,N_6483,N_6297);
nand U6787 (N_6787,N_6389,N_6012);
xnor U6788 (N_6788,N_6395,N_6482);
and U6789 (N_6789,N_6429,N_6394);
nand U6790 (N_6790,N_6178,N_6355);
or U6791 (N_6791,N_6006,N_6199);
nor U6792 (N_6792,N_6250,N_6268);
or U6793 (N_6793,N_6421,N_6015);
or U6794 (N_6794,N_6087,N_6422);
or U6795 (N_6795,N_6461,N_6093);
xnor U6796 (N_6796,N_6494,N_6488);
xor U6797 (N_6797,N_6248,N_6361);
nand U6798 (N_6798,N_6156,N_6405);
xor U6799 (N_6799,N_6171,N_6274);
and U6800 (N_6800,N_6462,N_6221);
nor U6801 (N_6801,N_6453,N_6446);
xnor U6802 (N_6802,N_6252,N_6021);
and U6803 (N_6803,N_6027,N_6236);
nand U6804 (N_6804,N_6347,N_6005);
nor U6805 (N_6805,N_6087,N_6178);
or U6806 (N_6806,N_6404,N_6186);
or U6807 (N_6807,N_6387,N_6105);
and U6808 (N_6808,N_6428,N_6263);
xnor U6809 (N_6809,N_6375,N_6081);
nor U6810 (N_6810,N_6343,N_6114);
and U6811 (N_6811,N_6056,N_6478);
nor U6812 (N_6812,N_6381,N_6044);
xnor U6813 (N_6813,N_6324,N_6288);
or U6814 (N_6814,N_6373,N_6024);
or U6815 (N_6815,N_6404,N_6263);
or U6816 (N_6816,N_6070,N_6121);
nor U6817 (N_6817,N_6293,N_6009);
or U6818 (N_6818,N_6070,N_6031);
nand U6819 (N_6819,N_6066,N_6106);
nand U6820 (N_6820,N_6105,N_6351);
or U6821 (N_6821,N_6254,N_6231);
and U6822 (N_6822,N_6195,N_6284);
xnor U6823 (N_6823,N_6274,N_6251);
or U6824 (N_6824,N_6134,N_6224);
nand U6825 (N_6825,N_6304,N_6449);
and U6826 (N_6826,N_6027,N_6471);
and U6827 (N_6827,N_6372,N_6286);
nand U6828 (N_6828,N_6180,N_6205);
nor U6829 (N_6829,N_6352,N_6409);
nor U6830 (N_6830,N_6188,N_6356);
or U6831 (N_6831,N_6253,N_6160);
or U6832 (N_6832,N_6298,N_6403);
or U6833 (N_6833,N_6385,N_6498);
and U6834 (N_6834,N_6429,N_6155);
nor U6835 (N_6835,N_6096,N_6281);
nand U6836 (N_6836,N_6383,N_6428);
nor U6837 (N_6837,N_6346,N_6196);
or U6838 (N_6838,N_6221,N_6365);
xnor U6839 (N_6839,N_6198,N_6187);
nor U6840 (N_6840,N_6131,N_6384);
xor U6841 (N_6841,N_6488,N_6465);
nand U6842 (N_6842,N_6025,N_6220);
and U6843 (N_6843,N_6339,N_6205);
nand U6844 (N_6844,N_6011,N_6435);
or U6845 (N_6845,N_6322,N_6110);
or U6846 (N_6846,N_6299,N_6480);
and U6847 (N_6847,N_6278,N_6496);
and U6848 (N_6848,N_6365,N_6350);
xnor U6849 (N_6849,N_6403,N_6093);
or U6850 (N_6850,N_6148,N_6175);
xnor U6851 (N_6851,N_6309,N_6174);
and U6852 (N_6852,N_6357,N_6092);
or U6853 (N_6853,N_6298,N_6135);
and U6854 (N_6854,N_6199,N_6167);
and U6855 (N_6855,N_6214,N_6345);
nor U6856 (N_6856,N_6264,N_6266);
xor U6857 (N_6857,N_6197,N_6115);
and U6858 (N_6858,N_6142,N_6462);
or U6859 (N_6859,N_6115,N_6070);
or U6860 (N_6860,N_6079,N_6088);
nand U6861 (N_6861,N_6475,N_6493);
and U6862 (N_6862,N_6020,N_6204);
xor U6863 (N_6863,N_6495,N_6491);
nor U6864 (N_6864,N_6326,N_6146);
or U6865 (N_6865,N_6188,N_6194);
and U6866 (N_6866,N_6286,N_6304);
and U6867 (N_6867,N_6165,N_6216);
and U6868 (N_6868,N_6042,N_6315);
and U6869 (N_6869,N_6018,N_6351);
xor U6870 (N_6870,N_6277,N_6307);
or U6871 (N_6871,N_6309,N_6327);
xnor U6872 (N_6872,N_6260,N_6232);
or U6873 (N_6873,N_6065,N_6351);
and U6874 (N_6874,N_6388,N_6102);
and U6875 (N_6875,N_6269,N_6301);
nor U6876 (N_6876,N_6322,N_6325);
nor U6877 (N_6877,N_6084,N_6050);
xnor U6878 (N_6878,N_6452,N_6443);
and U6879 (N_6879,N_6072,N_6262);
nand U6880 (N_6880,N_6333,N_6022);
or U6881 (N_6881,N_6323,N_6045);
nor U6882 (N_6882,N_6114,N_6439);
or U6883 (N_6883,N_6434,N_6158);
nor U6884 (N_6884,N_6052,N_6145);
and U6885 (N_6885,N_6338,N_6394);
xor U6886 (N_6886,N_6140,N_6087);
nor U6887 (N_6887,N_6158,N_6076);
or U6888 (N_6888,N_6310,N_6273);
xor U6889 (N_6889,N_6052,N_6397);
nor U6890 (N_6890,N_6296,N_6078);
nor U6891 (N_6891,N_6035,N_6251);
nor U6892 (N_6892,N_6023,N_6195);
xnor U6893 (N_6893,N_6450,N_6246);
and U6894 (N_6894,N_6270,N_6445);
and U6895 (N_6895,N_6496,N_6439);
xor U6896 (N_6896,N_6097,N_6339);
and U6897 (N_6897,N_6252,N_6217);
nor U6898 (N_6898,N_6229,N_6335);
or U6899 (N_6899,N_6036,N_6022);
xnor U6900 (N_6900,N_6427,N_6108);
nand U6901 (N_6901,N_6026,N_6199);
nor U6902 (N_6902,N_6135,N_6147);
xor U6903 (N_6903,N_6293,N_6076);
nor U6904 (N_6904,N_6158,N_6191);
and U6905 (N_6905,N_6412,N_6066);
and U6906 (N_6906,N_6179,N_6426);
and U6907 (N_6907,N_6205,N_6367);
xor U6908 (N_6908,N_6075,N_6498);
xor U6909 (N_6909,N_6112,N_6311);
and U6910 (N_6910,N_6093,N_6302);
nand U6911 (N_6911,N_6002,N_6085);
nand U6912 (N_6912,N_6396,N_6436);
nand U6913 (N_6913,N_6058,N_6043);
xnor U6914 (N_6914,N_6179,N_6099);
and U6915 (N_6915,N_6026,N_6394);
and U6916 (N_6916,N_6192,N_6051);
and U6917 (N_6917,N_6154,N_6281);
xor U6918 (N_6918,N_6214,N_6189);
and U6919 (N_6919,N_6321,N_6325);
and U6920 (N_6920,N_6460,N_6018);
and U6921 (N_6921,N_6328,N_6161);
xor U6922 (N_6922,N_6329,N_6452);
nor U6923 (N_6923,N_6093,N_6299);
or U6924 (N_6924,N_6459,N_6447);
and U6925 (N_6925,N_6050,N_6139);
nand U6926 (N_6926,N_6198,N_6464);
or U6927 (N_6927,N_6408,N_6124);
nand U6928 (N_6928,N_6135,N_6423);
nand U6929 (N_6929,N_6211,N_6478);
nor U6930 (N_6930,N_6182,N_6263);
and U6931 (N_6931,N_6418,N_6038);
and U6932 (N_6932,N_6067,N_6263);
xnor U6933 (N_6933,N_6161,N_6085);
and U6934 (N_6934,N_6195,N_6090);
nor U6935 (N_6935,N_6474,N_6497);
or U6936 (N_6936,N_6008,N_6204);
and U6937 (N_6937,N_6233,N_6351);
nor U6938 (N_6938,N_6197,N_6262);
or U6939 (N_6939,N_6138,N_6231);
or U6940 (N_6940,N_6432,N_6260);
nor U6941 (N_6941,N_6006,N_6292);
nand U6942 (N_6942,N_6245,N_6440);
xor U6943 (N_6943,N_6281,N_6493);
nand U6944 (N_6944,N_6169,N_6280);
nand U6945 (N_6945,N_6378,N_6271);
nand U6946 (N_6946,N_6304,N_6187);
and U6947 (N_6947,N_6124,N_6260);
xor U6948 (N_6948,N_6407,N_6413);
nor U6949 (N_6949,N_6155,N_6195);
nand U6950 (N_6950,N_6335,N_6078);
nand U6951 (N_6951,N_6254,N_6389);
xor U6952 (N_6952,N_6430,N_6218);
nor U6953 (N_6953,N_6319,N_6006);
nor U6954 (N_6954,N_6395,N_6071);
nand U6955 (N_6955,N_6484,N_6458);
nand U6956 (N_6956,N_6230,N_6140);
or U6957 (N_6957,N_6249,N_6247);
and U6958 (N_6958,N_6343,N_6472);
xnor U6959 (N_6959,N_6492,N_6011);
nor U6960 (N_6960,N_6166,N_6060);
nand U6961 (N_6961,N_6436,N_6490);
and U6962 (N_6962,N_6383,N_6050);
and U6963 (N_6963,N_6252,N_6090);
nand U6964 (N_6964,N_6107,N_6204);
xor U6965 (N_6965,N_6130,N_6380);
nor U6966 (N_6966,N_6468,N_6135);
and U6967 (N_6967,N_6335,N_6029);
or U6968 (N_6968,N_6288,N_6310);
nor U6969 (N_6969,N_6367,N_6206);
nand U6970 (N_6970,N_6423,N_6127);
or U6971 (N_6971,N_6161,N_6330);
and U6972 (N_6972,N_6422,N_6167);
nor U6973 (N_6973,N_6329,N_6340);
or U6974 (N_6974,N_6252,N_6191);
and U6975 (N_6975,N_6353,N_6384);
nor U6976 (N_6976,N_6337,N_6429);
and U6977 (N_6977,N_6028,N_6225);
xnor U6978 (N_6978,N_6083,N_6264);
nor U6979 (N_6979,N_6236,N_6239);
nor U6980 (N_6980,N_6409,N_6410);
xnor U6981 (N_6981,N_6031,N_6414);
xnor U6982 (N_6982,N_6064,N_6316);
nor U6983 (N_6983,N_6427,N_6339);
nand U6984 (N_6984,N_6212,N_6126);
nor U6985 (N_6985,N_6324,N_6187);
or U6986 (N_6986,N_6417,N_6493);
xor U6987 (N_6987,N_6120,N_6075);
nand U6988 (N_6988,N_6351,N_6000);
xnor U6989 (N_6989,N_6172,N_6339);
xor U6990 (N_6990,N_6433,N_6194);
nor U6991 (N_6991,N_6271,N_6072);
and U6992 (N_6992,N_6422,N_6304);
and U6993 (N_6993,N_6216,N_6345);
and U6994 (N_6994,N_6048,N_6370);
xor U6995 (N_6995,N_6010,N_6002);
nand U6996 (N_6996,N_6132,N_6373);
nor U6997 (N_6997,N_6421,N_6288);
or U6998 (N_6998,N_6417,N_6495);
or U6999 (N_6999,N_6233,N_6454);
nor U7000 (N_7000,N_6945,N_6590);
and U7001 (N_7001,N_6989,N_6511);
xnor U7002 (N_7002,N_6826,N_6707);
and U7003 (N_7003,N_6628,N_6812);
nor U7004 (N_7004,N_6746,N_6916);
nor U7005 (N_7005,N_6768,N_6575);
nor U7006 (N_7006,N_6674,N_6983);
xnor U7007 (N_7007,N_6977,N_6809);
nand U7008 (N_7008,N_6885,N_6718);
nor U7009 (N_7009,N_6778,N_6640);
nor U7010 (N_7010,N_6741,N_6864);
xor U7011 (N_7011,N_6815,N_6634);
nor U7012 (N_7012,N_6609,N_6642);
or U7013 (N_7013,N_6997,N_6570);
and U7014 (N_7014,N_6537,N_6793);
and U7015 (N_7015,N_6940,N_6528);
and U7016 (N_7016,N_6935,N_6743);
nand U7017 (N_7017,N_6973,N_6587);
nor U7018 (N_7018,N_6858,N_6664);
and U7019 (N_7019,N_6623,N_6870);
nor U7020 (N_7020,N_6810,N_6950);
nor U7021 (N_7021,N_6644,N_6569);
or U7022 (N_7022,N_6899,N_6593);
and U7023 (N_7023,N_6777,N_6712);
nor U7024 (N_7024,N_6912,N_6941);
or U7025 (N_7025,N_6592,N_6536);
nand U7026 (N_7026,N_6748,N_6747);
nor U7027 (N_7027,N_6626,N_6907);
nand U7028 (N_7028,N_6524,N_6556);
and U7029 (N_7029,N_6995,N_6959);
nor U7030 (N_7030,N_6595,N_6848);
nor U7031 (N_7031,N_6790,N_6866);
nor U7032 (N_7032,N_6629,N_6632);
nor U7033 (N_7033,N_6561,N_6521);
and U7034 (N_7034,N_6739,N_6759);
and U7035 (N_7035,N_6695,N_6606);
xnor U7036 (N_7036,N_6863,N_6913);
nor U7037 (N_7037,N_6688,N_6651);
nor U7038 (N_7038,N_6734,N_6641);
nor U7039 (N_7039,N_6976,N_6986);
or U7040 (N_7040,N_6534,N_6517);
nand U7041 (N_7041,N_6689,N_6670);
xor U7042 (N_7042,N_6615,N_6836);
xor U7043 (N_7043,N_6729,N_6657);
or U7044 (N_7044,N_6714,N_6849);
nor U7045 (N_7045,N_6591,N_6868);
and U7046 (N_7046,N_6779,N_6539);
nor U7047 (N_7047,N_6920,N_6926);
nand U7048 (N_7048,N_6614,N_6830);
or U7049 (N_7049,N_6783,N_6699);
and U7050 (N_7050,N_6785,N_6869);
xnor U7051 (N_7051,N_6875,N_6512);
and U7052 (N_7052,N_6789,N_6597);
and U7053 (N_7053,N_6563,N_6622);
or U7054 (N_7054,N_6607,N_6543);
nand U7055 (N_7055,N_6904,N_6661);
xor U7056 (N_7056,N_6513,N_6672);
and U7057 (N_7057,N_6716,N_6525);
nor U7058 (N_7058,N_6558,N_6909);
xor U7059 (N_7059,N_6658,N_6829);
or U7060 (N_7060,N_6711,N_6946);
nor U7061 (N_7061,N_6805,N_6683);
or U7062 (N_7062,N_6884,N_6857);
or U7063 (N_7063,N_6667,N_6506);
nand U7064 (N_7064,N_6553,N_6838);
xor U7065 (N_7065,N_6673,N_6599);
or U7066 (N_7066,N_6668,N_6965);
and U7067 (N_7067,N_6881,N_6598);
or U7068 (N_7068,N_6839,N_6618);
xor U7069 (N_7069,N_6931,N_6705);
nor U7070 (N_7070,N_6948,N_6763);
nand U7071 (N_7071,N_6687,N_6765);
and U7072 (N_7072,N_6538,N_6760);
nand U7073 (N_7073,N_6723,N_6691);
or U7074 (N_7074,N_6800,N_6696);
or U7075 (N_7075,N_6555,N_6704);
nor U7076 (N_7076,N_6742,N_6727);
nand U7077 (N_7077,N_6862,N_6596);
nor U7078 (N_7078,N_6604,N_6933);
nand U7079 (N_7079,N_6533,N_6542);
or U7080 (N_7080,N_6730,N_6713);
nand U7081 (N_7081,N_6996,N_6566);
nand U7082 (N_7082,N_6717,N_6514);
or U7083 (N_7083,N_6828,N_6822);
or U7084 (N_7084,N_6625,N_6823);
xor U7085 (N_7085,N_6987,N_6821);
nor U7086 (N_7086,N_6720,N_6504);
xnor U7087 (N_7087,N_6740,N_6797);
nor U7088 (N_7088,N_6934,N_6663);
and U7089 (N_7089,N_6993,N_6865);
nand U7090 (N_7090,N_6613,N_6770);
or U7091 (N_7091,N_6649,N_6859);
or U7092 (N_7092,N_6682,N_6662);
nand U7093 (N_7093,N_6677,N_6549);
or U7094 (N_7094,N_6584,N_6999);
xnor U7095 (N_7095,N_6835,N_6580);
or U7096 (N_7096,N_6833,N_6841);
nor U7097 (N_7097,N_6726,N_6895);
nand U7098 (N_7098,N_6820,N_6627);
or U7099 (N_7099,N_6654,N_6775);
xor U7100 (N_7100,N_6776,N_6501);
nand U7101 (N_7101,N_6792,N_6850);
nand U7102 (N_7102,N_6588,N_6560);
or U7103 (N_7103,N_6708,N_6974);
nor U7104 (N_7104,N_6751,N_6943);
nand U7105 (N_7105,N_6877,N_6917);
or U7106 (N_7106,N_6981,N_6801);
or U7107 (N_7107,N_6998,N_6867);
and U7108 (N_7108,N_6709,N_6550);
and U7109 (N_7109,N_6960,N_6900);
nand U7110 (N_7110,N_6559,N_6646);
nand U7111 (N_7111,N_6594,N_6722);
nand U7112 (N_7112,N_6978,N_6761);
nand U7113 (N_7113,N_6834,N_6854);
xnor U7114 (N_7114,N_6698,N_6970);
or U7115 (N_7115,N_6874,N_6611);
and U7116 (N_7116,N_6665,N_6637);
xor U7117 (N_7117,N_6749,N_6937);
and U7118 (N_7118,N_6897,N_6601);
and U7119 (N_7119,N_6788,N_6503);
nand U7120 (N_7120,N_6929,N_6660);
xnor U7121 (N_7121,N_6737,N_6888);
xnor U7122 (N_7122,N_6733,N_6652);
xor U7123 (N_7123,N_6845,N_6619);
and U7124 (N_7124,N_6639,N_6681);
or U7125 (N_7125,N_6939,N_6925);
or U7126 (N_7126,N_6612,N_6635);
xnor U7127 (N_7127,N_6980,N_6562);
nor U7128 (N_7128,N_6535,N_6958);
nand U7129 (N_7129,N_6798,N_6516);
and U7130 (N_7130,N_6557,N_6745);
and U7131 (N_7131,N_6919,N_6938);
nand U7132 (N_7132,N_6804,N_6924);
xnor U7133 (N_7133,N_6856,N_6735);
nor U7134 (N_7134,N_6582,N_6914);
and U7135 (N_7135,N_6586,N_6832);
xor U7136 (N_7136,N_6731,N_6564);
nand U7137 (N_7137,N_6971,N_6756);
nor U7138 (N_7138,N_6769,N_6780);
nand U7139 (N_7139,N_6507,N_6831);
xor U7140 (N_7140,N_6969,N_6650);
or U7141 (N_7141,N_6956,N_6990);
and U7142 (N_7142,N_6903,N_6605);
nor U7143 (N_7143,N_6936,N_6876);
xnor U7144 (N_7144,N_6719,N_6706);
or U7145 (N_7145,N_6906,N_6523);
nand U7146 (N_7146,N_6762,N_6819);
and U7147 (N_7147,N_6992,N_6522);
xor U7148 (N_7148,N_6690,N_6616);
or U7149 (N_7149,N_6715,N_6692);
nand U7150 (N_7150,N_6908,N_6898);
nand U7151 (N_7151,N_6872,N_6702);
or U7152 (N_7152,N_6851,N_6944);
nor U7153 (N_7153,N_6679,N_6530);
and U7154 (N_7154,N_6824,N_6781);
and U7155 (N_7155,N_6813,N_6942);
nand U7156 (N_7156,N_6979,N_6784);
nand U7157 (N_7157,N_6574,N_6724);
xnor U7158 (N_7158,N_6896,N_6518);
nor U7159 (N_7159,N_6581,N_6655);
xor U7160 (N_7160,N_6972,N_6589);
or U7161 (N_7161,N_6548,N_6546);
nand U7162 (N_7162,N_6802,N_6984);
nand U7163 (N_7163,N_6795,N_6985);
nor U7164 (N_7164,N_6957,N_6952);
or U7165 (N_7165,N_6578,N_6879);
nor U7166 (N_7166,N_6608,N_6827);
nor U7167 (N_7167,N_6922,N_6887);
xor U7168 (N_7168,N_6532,N_6721);
xnor U7169 (N_7169,N_6685,N_6928);
and U7170 (N_7170,N_6782,N_6527);
nor U7171 (N_7171,N_6728,N_6693);
nor U7172 (N_7172,N_6817,N_6764);
xor U7173 (N_7173,N_6852,N_6966);
xor U7174 (N_7174,N_6840,N_6918);
or U7175 (N_7175,N_6773,N_6855);
nand U7176 (N_7176,N_6624,N_6552);
nand U7177 (N_7177,N_6975,N_6738);
nor U7178 (N_7178,N_6791,N_6675);
xnor U7179 (N_7179,N_6901,N_6954);
and U7180 (N_7180,N_6882,N_6803);
nor U7181 (N_7181,N_6653,N_6767);
xnor U7182 (N_7182,N_6752,N_6921);
nand U7183 (N_7183,N_6703,N_6818);
and U7184 (N_7184,N_6825,N_6878);
nor U7185 (N_7185,N_6645,N_6930);
nor U7186 (N_7186,N_6853,N_6505);
or U7187 (N_7187,N_6531,N_6621);
xor U7188 (N_7188,N_6710,N_6529);
nand U7189 (N_7189,N_6947,N_6669);
nand U7190 (N_7190,N_6774,N_6571);
or U7191 (N_7191,N_6736,N_6794);
and U7192 (N_7192,N_6732,N_6932);
nand U7193 (N_7193,N_6554,N_6955);
or U7194 (N_7194,N_6541,N_6787);
xnor U7195 (N_7195,N_6540,N_6545);
or U7196 (N_7196,N_6579,N_6758);
nand U7197 (N_7197,N_6982,N_6771);
xor U7198 (N_7198,N_6636,N_6676);
or U7199 (N_7199,N_6610,N_6889);
or U7200 (N_7200,N_6515,N_6509);
xnor U7201 (N_7201,N_6766,N_6643);
and U7202 (N_7202,N_6894,N_6603);
or U7203 (N_7203,N_6951,N_6754);
nor U7204 (N_7204,N_6744,N_6567);
nor U7205 (N_7205,N_6583,N_6786);
xor U7206 (N_7206,N_6816,N_6755);
and U7207 (N_7207,N_6659,N_6510);
or U7208 (N_7208,N_6799,N_6600);
nand U7209 (N_7209,N_6750,N_6842);
and U7210 (N_7210,N_6671,N_6576);
xnor U7211 (N_7211,N_6886,N_6961);
or U7212 (N_7212,N_6620,N_6656);
nand U7213 (N_7213,N_6902,N_6638);
nor U7214 (N_7214,N_6502,N_6631);
or U7215 (N_7215,N_6573,N_6630);
nand U7216 (N_7216,N_6927,N_6551);
or U7217 (N_7217,N_6648,N_6963);
nor U7218 (N_7218,N_6991,N_6519);
or U7219 (N_7219,N_6680,N_6962);
or U7220 (N_7220,N_6814,N_6994);
and U7221 (N_7221,N_6544,N_6861);
nor U7222 (N_7222,N_6883,N_6967);
xor U7223 (N_7223,N_6880,N_6526);
and U7224 (N_7224,N_6892,N_6568);
or U7225 (N_7225,N_6949,N_6905);
xnor U7226 (N_7226,N_6968,N_6633);
or U7227 (N_7227,N_6988,N_6686);
xor U7228 (N_7228,N_6647,N_6860);
nor U7229 (N_7229,N_6772,N_6808);
nor U7230 (N_7230,N_6508,N_6520);
nand U7231 (N_7231,N_6565,N_6697);
or U7232 (N_7232,N_6500,N_6891);
and U7233 (N_7233,N_6964,N_6844);
and U7234 (N_7234,N_6837,N_6701);
xor U7235 (N_7235,N_6871,N_6811);
nand U7236 (N_7236,N_6893,N_6684);
and U7237 (N_7237,N_6953,N_6843);
xor U7238 (N_7238,N_6806,N_6577);
xor U7239 (N_7239,N_6890,N_6846);
or U7240 (N_7240,N_6873,N_6694);
and U7241 (N_7241,N_6807,N_6617);
xor U7242 (N_7242,N_6753,N_6700);
and U7243 (N_7243,N_6911,N_6547);
or U7244 (N_7244,N_6666,N_6915);
nor U7245 (N_7245,N_6910,N_6923);
or U7246 (N_7246,N_6678,N_6796);
nor U7247 (N_7247,N_6725,N_6585);
and U7248 (N_7248,N_6602,N_6572);
or U7249 (N_7249,N_6847,N_6757);
xor U7250 (N_7250,N_6734,N_6538);
or U7251 (N_7251,N_6695,N_6675);
nand U7252 (N_7252,N_6884,N_6598);
nand U7253 (N_7253,N_6532,N_6927);
xor U7254 (N_7254,N_6655,N_6617);
nand U7255 (N_7255,N_6805,N_6738);
nor U7256 (N_7256,N_6661,N_6997);
xor U7257 (N_7257,N_6991,N_6618);
or U7258 (N_7258,N_6915,N_6633);
xor U7259 (N_7259,N_6639,N_6696);
nor U7260 (N_7260,N_6533,N_6504);
or U7261 (N_7261,N_6799,N_6901);
nor U7262 (N_7262,N_6690,N_6799);
xnor U7263 (N_7263,N_6818,N_6695);
nand U7264 (N_7264,N_6964,N_6668);
or U7265 (N_7265,N_6833,N_6527);
nor U7266 (N_7266,N_6824,N_6862);
or U7267 (N_7267,N_6935,N_6825);
nor U7268 (N_7268,N_6833,N_6659);
nand U7269 (N_7269,N_6596,N_6928);
and U7270 (N_7270,N_6678,N_6794);
nor U7271 (N_7271,N_6905,N_6605);
and U7272 (N_7272,N_6548,N_6652);
nand U7273 (N_7273,N_6670,N_6986);
nor U7274 (N_7274,N_6564,N_6589);
and U7275 (N_7275,N_6962,N_6957);
and U7276 (N_7276,N_6711,N_6899);
xnor U7277 (N_7277,N_6831,N_6706);
and U7278 (N_7278,N_6532,N_6649);
nor U7279 (N_7279,N_6628,N_6866);
and U7280 (N_7280,N_6726,N_6756);
nor U7281 (N_7281,N_6664,N_6696);
and U7282 (N_7282,N_6606,N_6694);
nor U7283 (N_7283,N_6886,N_6903);
nor U7284 (N_7284,N_6804,N_6851);
nor U7285 (N_7285,N_6801,N_6842);
or U7286 (N_7286,N_6820,N_6766);
or U7287 (N_7287,N_6502,N_6567);
nand U7288 (N_7288,N_6959,N_6634);
xnor U7289 (N_7289,N_6654,N_6794);
nor U7290 (N_7290,N_6636,N_6986);
nand U7291 (N_7291,N_6642,N_6906);
xnor U7292 (N_7292,N_6694,N_6658);
xor U7293 (N_7293,N_6611,N_6718);
and U7294 (N_7294,N_6518,N_6610);
or U7295 (N_7295,N_6990,N_6570);
and U7296 (N_7296,N_6962,N_6545);
nand U7297 (N_7297,N_6932,N_6648);
nand U7298 (N_7298,N_6852,N_6705);
and U7299 (N_7299,N_6779,N_6706);
nor U7300 (N_7300,N_6591,N_6843);
nand U7301 (N_7301,N_6587,N_6563);
nor U7302 (N_7302,N_6714,N_6781);
xor U7303 (N_7303,N_6578,N_6599);
xor U7304 (N_7304,N_6768,N_6728);
or U7305 (N_7305,N_6638,N_6768);
nor U7306 (N_7306,N_6553,N_6998);
and U7307 (N_7307,N_6743,N_6938);
or U7308 (N_7308,N_6643,N_6962);
xnor U7309 (N_7309,N_6869,N_6965);
nand U7310 (N_7310,N_6622,N_6995);
nor U7311 (N_7311,N_6732,N_6664);
nand U7312 (N_7312,N_6726,N_6628);
nor U7313 (N_7313,N_6852,N_6925);
and U7314 (N_7314,N_6550,N_6662);
or U7315 (N_7315,N_6601,N_6672);
nor U7316 (N_7316,N_6934,N_6714);
and U7317 (N_7317,N_6641,N_6919);
nand U7318 (N_7318,N_6622,N_6513);
nand U7319 (N_7319,N_6987,N_6932);
nand U7320 (N_7320,N_6932,N_6682);
or U7321 (N_7321,N_6982,N_6843);
and U7322 (N_7322,N_6560,N_6851);
and U7323 (N_7323,N_6979,N_6931);
nor U7324 (N_7324,N_6583,N_6978);
or U7325 (N_7325,N_6733,N_6830);
or U7326 (N_7326,N_6597,N_6918);
nand U7327 (N_7327,N_6539,N_6560);
nand U7328 (N_7328,N_6578,N_6655);
nor U7329 (N_7329,N_6988,N_6914);
and U7330 (N_7330,N_6993,N_6676);
nand U7331 (N_7331,N_6897,N_6817);
nand U7332 (N_7332,N_6971,N_6543);
and U7333 (N_7333,N_6732,N_6956);
nor U7334 (N_7334,N_6863,N_6672);
and U7335 (N_7335,N_6825,N_6911);
nand U7336 (N_7336,N_6978,N_6869);
nor U7337 (N_7337,N_6775,N_6985);
nand U7338 (N_7338,N_6955,N_6741);
and U7339 (N_7339,N_6727,N_6954);
or U7340 (N_7340,N_6985,N_6504);
and U7341 (N_7341,N_6627,N_6590);
nand U7342 (N_7342,N_6839,N_6610);
xor U7343 (N_7343,N_6536,N_6809);
and U7344 (N_7344,N_6744,N_6943);
and U7345 (N_7345,N_6677,N_6643);
or U7346 (N_7346,N_6880,N_6593);
xor U7347 (N_7347,N_6687,N_6697);
or U7348 (N_7348,N_6752,N_6758);
nand U7349 (N_7349,N_6646,N_6568);
or U7350 (N_7350,N_6782,N_6719);
nor U7351 (N_7351,N_6897,N_6956);
or U7352 (N_7352,N_6709,N_6551);
nor U7353 (N_7353,N_6653,N_6750);
and U7354 (N_7354,N_6888,N_6810);
nor U7355 (N_7355,N_6727,N_6804);
nand U7356 (N_7356,N_6914,N_6999);
or U7357 (N_7357,N_6773,N_6595);
or U7358 (N_7358,N_6671,N_6763);
nand U7359 (N_7359,N_6544,N_6583);
nand U7360 (N_7360,N_6784,N_6788);
and U7361 (N_7361,N_6746,N_6506);
nor U7362 (N_7362,N_6647,N_6934);
xnor U7363 (N_7363,N_6601,N_6990);
xnor U7364 (N_7364,N_6777,N_6758);
nor U7365 (N_7365,N_6766,N_6736);
nor U7366 (N_7366,N_6554,N_6631);
or U7367 (N_7367,N_6717,N_6622);
xor U7368 (N_7368,N_6829,N_6660);
nor U7369 (N_7369,N_6818,N_6736);
and U7370 (N_7370,N_6875,N_6979);
or U7371 (N_7371,N_6811,N_6851);
nor U7372 (N_7372,N_6927,N_6700);
or U7373 (N_7373,N_6509,N_6982);
nor U7374 (N_7374,N_6907,N_6802);
and U7375 (N_7375,N_6921,N_6520);
or U7376 (N_7376,N_6963,N_6687);
and U7377 (N_7377,N_6933,N_6912);
nor U7378 (N_7378,N_6877,N_6813);
and U7379 (N_7379,N_6536,N_6733);
or U7380 (N_7380,N_6914,N_6742);
nor U7381 (N_7381,N_6792,N_6819);
or U7382 (N_7382,N_6524,N_6547);
or U7383 (N_7383,N_6759,N_6724);
or U7384 (N_7384,N_6892,N_6679);
and U7385 (N_7385,N_6855,N_6619);
nor U7386 (N_7386,N_6801,N_6550);
nor U7387 (N_7387,N_6569,N_6782);
nor U7388 (N_7388,N_6637,N_6976);
and U7389 (N_7389,N_6522,N_6532);
nor U7390 (N_7390,N_6515,N_6574);
or U7391 (N_7391,N_6850,N_6736);
nand U7392 (N_7392,N_6905,N_6754);
and U7393 (N_7393,N_6685,N_6738);
nand U7394 (N_7394,N_6976,N_6558);
and U7395 (N_7395,N_6581,N_6745);
xor U7396 (N_7396,N_6756,N_6591);
nand U7397 (N_7397,N_6643,N_6510);
and U7398 (N_7398,N_6842,N_6962);
xnor U7399 (N_7399,N_6688,N_6558);
nand U7400 (N_7400,N_6900,N_6929);
nand U7401 (N_7401,N_6901,N_6943);
nor U7402 (N_7402,N_6555,N_6848);
or U7403 (N_7403,N_6739,N_6733);
nor U7404 (N_7404,N_6734,N_6880);
nand U7405 (N_7405,N_6946,N_6524);
nor U7406 (N_7406,N_6946,N_6908);
xor U7407 (N_7407,N_6866,N_6849);
nand U7408 (N_7408,N_6733,N_6700);
nor U7409 (N_7409,N_6637,N_6662);
nand U7410 (N_7410,N_6890,N_6682);
and U7411 (N_7411,N_6715,N_6501);
and U7412 (N_7412,N_6987,N_6923);
nor U7413 (N_7413,N_6552,N_6727);
xor U7414 (N_7414,N_6780,N_6893);
and U7415 (N_7415,N_6904,N_6987);
or U7416 (N_7416,N_6954,N_6607);
xor U7417 (N_7417,N_6555,N_6962);
nand U7418 (N_7418,N_6614,N_6930);
xnor U7419 (N_7419,N_6592,N_6708);
nor U7420 (N_7420,N_6811,N_6939);
xnor U7421 (N_7421,N_6501,N_6707);
nor U7422 (N_7422,N_6535,N_6816);
or U7423 (N_7423,N_6759,N_6568);
and U7424 (N_7424,N_6585,N_6910);
and U7425 (N_7425,N_6862,N_6920);
nand U7426 (N_7426,N_6949,N_6901);
and U7427 (N_7427,N_6986,N_6756);
and U7428 (N_7428,N_6583,N_6923);
nand U7429 (N_7429,N_6593,N_6689);
xnor U7430 (N_7430,N_6600,N_6784);
and U7431 (N_7431,N_6677,N_6676);
nor U7432 (N_7432,N_6743,N_6595);
nand U7433 (N_7433,N_6755,N_6768);
nor U7434 (N_7434,N_6879,N_6735);
and U7435 (N_7435,N_6786,N_6862);
nor U7436 (N_7436,N_6539,N_6679);
nor U7437 (N_7437,N_6918,N_6634);
or U7438 (N_7438,N_6733,N_6955);
xor U7439 (N_7439,N_6831,N_6978);
nor U7440 (N_7440,N_6823,N_6518);
nor U7441 (N_7441,N_6568,N_6690);
and U7442 (N_7442,N_6507,N_6569);
or U7443 (N_7443,N_6879,N_6678);
nand U7444 (N_7444,N_6645,N_6933);
and U7445 (N_7445,N_6632,N_6542);
nand U7446 (N_7446,N_6915,N_6701);
nor U7447 (N_7447,N_6926,N_6803);
nand U7448 (N_7448,N_6661,N_6561);
and U7449 (N_7449,N_6523,N_6985);
nor U7450 (N_7450,N_6569,N_6814);
nor U7451 (N_7451,N_6529,N_6834);
and U7452 (N_7452,N_6802,N_6981);
xor U7453 (N_7453,N_6731,N_6581);
and U7454 (N_7454,N_6639,N_6756);
xnor U7455 (N_7455,N_6745,N_6564);
nor U7456 (N_7456,N_6602,N_6581);
and U7457 (N_7457,N_6680,N_6787);
nand U7458 (N_7458,N_6697,N_6752);
nand U7459 (N_7459,N_6850,N_6837);
nor U7460 (N_7460,N_6949,N_6733);
xnor U7461 (N_7461,N_6701,N_6672);
nor U7462 (N_7462,N_6954,N_6807);
or U7463 (N_7463,N_6742,N_6721);
xnor U7464 (N_7464,N_6858,N_6900);
nand U7465 (N_7465,N_6548,N_6648);
or U7466 (N_7466,N_6715,N_6733);
xnor U7467 (N_7467,N_6589,N_6821);
nor U7468 (N_7468,N_6845,N_6803);
or U7469 (N_7469,N_6868,N_6988);
nor U7470 (N_7470,N_6773,N_6677);
xnor U7471 (N_7471,N_6858,N_6928);
nor U7472 (N_7472,N_6903,N_6579);
or U7473 (N_7473,N_6735,N_6544);
nor U7474 (N_7474,N_6837,N_6654);
nor U7475 (N_7475,N_6566,N_6697);
or U7476 (N_7476,N_6764,N_6701);
nor U7477 (N_7477,N_6940,N_6608);
xor U7478 (N_7478,N_6725,N_6674);
xor U7479 (N_7479,N_6712,N_6655);
or U7480 (N_7480,N_6978,N_6526);
nand U7481 (N_7481,N_6620,N_6646);
or U7482 (N_7482,N_6782,N_6650);
nor U7483 (N_7483,N_6503,N_6822);
nand U7484 (N_7484,N_6651,N_6727);
nor U7485 (N_7485,N_6733,N_6664);
xnor U7486 (N_7486,N_6640,N_6853);
nor U7487 (N_7487,N_6832,N_6821);
nand U7488 (N_7488,N_6572,N_6610);
and U7489 (N_7489,N_6858,N_6731);
or U7490 (N_7490,N_6616,N_6793);
nand U7491 (N_7491,N_6538,N_6718);
nor U7492 (N_7492,N_6639,N_6613);
and U7493 (N_7493,N_6872,N_6636);
xor U7494 (N_7494,N_6576,N_6613);
or U7495 (N_7495,N_6802,N_6864);
nand U7496 (N_7496,N_6977,N_6996);
or U7497 (N_7497,N_6741,N_6879);
nor U7498 (N_7498,N_6835,N_6600);
nand U7499 (N_7499,N_6526,N_6903);
and U7500 (N_7500,N_7030,N_7264);
xor U7501 (N_7501,N_7241,N_7059);
nor U7502 (N_7502,N_7147,N_7289);
or U7503 (N_7503,N_7384,N_7334);
and U7504 (N_7504,N_7421,N_7278);
nand U7505 (N_7505,N_7313,N_7470);
and U7506 (N_7506,N_7416,N_7284);
or U7507 (N_7507,N_7315,N_7231);
and U7508 (N_7508,N_7180,N_7006);
and U7509 (N_7509,N_7084,N_7129);
nand U7510 (N_7510,N_7145,N_7217);
nand U7511 (N_7511,N_7466,N_7350);
nor U7512 (N_7512,N_7149,N_7433);
nor U7513 (N_7513,N_7163,N_7279);
xor U7514 (N_7514,N_7302,N_7361);
nand U7515 (N_7515,N_7012,N_7082);
or U7516 (N_7516,N_7298,N_7010);
nor U7517 (N_7517,N_7423,N_7488);
or U7518 (N_7518,N_7045,N_7427);
nor U7519 (N_7519,N_7261,N_7176);
or U7520 (N_7520,N_7143,N_7036);
nor U7521 (N_7521,N_7085,N_7093);
and U7522 (N_7522,N_7251,N_7364);
xor U7523 (N_7523,N_7130,N_7424);
nand U7524 (N_7524,N_7357,N_7496);
nand U7525 (N_7525,N_7185,N_7151);
nor U7526 (N_7526,N_7223,N_7401);
xor U7527 (N_7527,N_7015,N_7202);
nor U7528 (N_7528,N_7389,N_7436);
or U7529 (N_7529,N_7312,N_7139);
and U7530 (N_7530,N_7038,N_7493);
xor U7531 (N_7531,N_7055,N_7088);
or U7532 (N_7532,N_7294,N_7365);
nor U7533 (N_7533,N_7097,N_7075);
nor U7534 (N_7534,N_7249,N_7183);
nand U7535 (N_7535,N_7367,N_7308);
nand U7536 (N_7536,N_7451,N_7374);
xor U7537 (N_7537,N_7192,N_7058);
or U7538 (N_7538,N_7104,N_7268);
nor U7539 (N_7539,N_7325,N_7169);
nor U7540 (N_7540,N_7219,N_7062);
or U7541 (N_7541,N_7087,N_7109);
and U7542 (N_7542,N_7438,N_7195);
nand U7543 (N_7543,N_7118,N_7295);
nor U7544 (N_7544,N_7481,N_7177);
nor U7545 (N_7545,N_7162,N_7484);
nand U7546 (N_7546,N_7197,N_7076);
or U7547 (N_7547,N_7383,N_7378);
xor U7548 (N_7548,N_7098,N_7155);
xnor U7549 (N_7549,N_7121,N_7469);
nand U7550 (N_7550,N_7485,N_7429);
or U7551 (N_7551,N_7404,N_7462);
or U7552 (N_7552,N_7014,N_7126);
and U7553 (N_7553,N_7277,N_7276);
nand U7554 (N_7554,N_7051,N_7138);
nor U7555 (N_7555,N_7090,N_7105);
nor U7556 (N_7556,N_7200,N_7495);
nand U7557 (N_7557,N_7210,N_7100);
or U7558 (N_7558,N_7236,N_7280);
and U7559 (N_7559,N_7181,N_7405);
nor U7560 (N_7560,N_7052,N_7204);
or U7561 (N_7561,N_7040,N_7127);
nor U7562 (N_7562,N_7487,N_7330);
or U7563 (N_7563,N_7158,N_7246);
xor U7564 (N_7564,N_7336,N_7463);
xor U7565 (N_7565,N_7019,N_7234);
nand U7566 (N_7566,N_7193,N_7369);
nand U7567 (N_7567,N_7356,N_7304);
and U7568 (N_7568,N_7397,N_7140);
xnor U7569 (N_7569,N_7095,N_7086);
nor U7570 (N_7570,N_7159,N_7073);
and U7571 (N_7571,N_7199,N_7172);
nand U7572 (N_7572,N_7046,N_7492);
nor U7573 (N_7573,N_7170,N_7007);
and U7574 (N_7574,N_7081,N_7410);
nand U7575 (N_7575,N_7431,N_7293);
or U7576 (N_7576,N_7047,N_7273);
nand U7577 (N_7577,N_7443,N_7286);
or U7578 (N_7578,N_7125,N_7292);
xor U7579 (N_7579,N_7326,N_7164);
nor U7580 (N_7580,N_7187,N_7373);
or U7581 (N_7581,N_7362,N_7414);
nand U7582 (N_7582,N_7478,N_7178);
and U7583 (N_7583,N_7455,N_7189);
xnor U7584 (N_7584,N_7198,N_7135);
nand U7585 (N_7585,N_7395,N_7255);
or U7586 (N_7586,N_7324,N_7418);
nand U7587 (N_7587,N_7420,N_7123);
xor U7588 (N_7588,N_7445,N_7233);
nor U7589 (N_7589,N_7209,N_7238);
xor U7590 (N_7590,N_7283,N_7415);
and U7591 (N_7591,N_7477,N_7372);
xor U7592 (N_7592,N_7305,N_7347);
and U7593 (N_7593,N_7160,N_7224);
xor U7594 (N_7594,N_7068,N_7113);
nand U7595 (N_7595,N_7215,N_7027);
nand U7596 (N_7596,N_7323,N_7101);
nor U7597 (N_7597,N_7165,N_7343);
or U7598 (N_7598,N_7327,N_7386);
or U7599 (N_7599,N_7029,N_7461);
xnor U7600 (N_7600,N_7201,N_7182);
xor U7601 (N_7601,N_7077,N_7239);
xor U7602 (N_7602,N_7049,N_7321);
xnor U7603 (N_7603,N_7240,N_7375);
nand U7604 (N_7604,N_7366,N_7322);
or U7605 (N_7605,N_7426,N_7490);
nand U7606 (N_7606,N_7004,N_7031);
nand U7607 (N_7607,N_7154,N_7368);
nand U7608 (N_7608,N_7299,N_7498);
or U7609 (N_7609,N_7446,N_7002);
xor U7610 (N_7610,N_7385,N_7044);
nand U7611 (N_7611,N_7475,N_7403);
nand U7612 (N_7612,N_7069,N_7053);
nor U7613 (N_7613,N_7320,N_7107);
nor U7614 (N_7614,N_7467,N_7211);
nand U7615 (N_7615,N_7137,N_7434);
and U7616 (N_7616,N_7430,N_7017);
and U7617 (N_7617,N_7253,N_7071);
nand U7618 (N_7618,N_7023,N_7254);
nor U7619 (N_7619,N_7065,N_7442);
xnor U7620 (N_7620,N_7190,N_7341);
and U7621 (N_7621,N_7425,N_7479);
and U7622 (N_7622,N_7491,N_7063);
nor U7623 (N_7623,N_7370,N_7272);
and U7624 (N_7624,N_7344,N_7248);
nand U7625 (N_7625,N_7025,N_7440);
xor U7626 (N_7626,N_7232,N_7296);
and U7627 (N_7627,N_7022,N_7458);
and U7628 (N_7628,N_7106,N_7270);
nand U7629 (N_7629,N_7003,N_7342);
nor U7630 (N_7630,N_7252,N_7146);
and U7631 (N_7631,N_7194,N_7230);
nor U7632 (N_7632,N_7021,N_7290);
xor U7633 (N_7633,N_7400,N_7092);
nand U7634 (N_7634,N_7175,N_7256);
xnor U7635 (N_7635,N_7407,N_7242);
nand U7636 (N_7636,N_7437,N_7134);
and U7637 (N_7637,N_7124,N_7432);
or U7638 (N_7638,N_7285,N_7102);
xor U7639 (N_7639,N_7244,N_7474);
nor U7640 (N_7640,N_7141,N_7482);
nor U7641 (N_7641,N_7448,N_7131);
or U7642 (N_7642,N_7345,N_7480);
and U7643 (N_7643,N_7460,N_7243);
nor U7644 (N_7644,N_7225,N_7398);
and U7645 (N_7645,N_7060,N_7112);
nand U7646 (N_7646,N_7222,N_7396);
or U7647 (N_7647,N_7260,N_7303);
nand U7648 (N_7648,N_7377,N_7483);
xor U7649 (N_7649,N_7428,N_7360);
nand U7650 (N_7650,N_7444,N_7091);
nor U7651 (N_7651,N_7235,N_7351);
nor U7652 (N_7652,N_7381,N_7136);
nor U7653 (N_7653,N_7150,N_7096);
nor U7654 (N_7654,N_7390,N_7009);
and U7655 (N_7655,N_7489,N_7108);
nand U7656 (N_7656,N_7122,N_7417);
and U7657 (N_7657,N_7048,N_7346);
nand U7658 (N_7658,N_7392,N_7115);
or U7659 (N_7659,N_7000,N_7218);
xnor U7660 (N_7660,N_7089,N_7228);
or U7661 (N_7661,N_7206,N_7173);
xor U7662 (N_7662,N_7291,N_7447);
xor U7663 (N_7663,N_7066,N_7376);
nor U7664 (N_7664,N_7161,N_7456);
nand U7665 (N_7665,N_7337,N_7083);
xor U7666 (N_7666,N_7499,N_7335);
or U7667 (N_7667,N_7250,N_7454);
nand U7668 (N_7668,N_7465,N_7494);
or U7669 (N_7669,N_7018,N_7412);
and U7670 (N_7670,N_7110,N_7166);
nor U7671 (N_7671,N_7033,N_7382);
or U7672 (N_7672,N_7354,N_7363);
and U7673 (N_7673,N_7316,N_7117);
or U7674 (N_7674,N_7457,N_7056);
or U7675 (N_7675,N_7358,N_7039);
nor U7676 (N_7676,N_7153,N_7037);
nor U7677 (N_7677,N_7453,N_7486);
nor U7678 (N_7678,N_7171,N_7352);
xnor U7679 (N_7679,N_7307,N_7080);
xor U7680 (N_7680,N_7057,N_7120);
nor U7681 (N_7681,N_7156,N_7409);
nor U7682 (N_7682,N_7314,N_7205);
nor U7683 (N_7683,N_7196,N_7203);
and U7684 (N_7684,N_7099,N_7042);
or U7685 (N_7685,N_7394,N_7245);
and U7686 (N_7686,N_7114,N_7310);
nor U7687 (N_7687,N_7464,N_7001);
or U7688 (N_7688,N_7449,N_7300);
nand U7689 (N_7689,N_7439,N_7471);
and U7690 (N_7690,N_7128,N_7262);
nand U7691 (N_7691,N_7317,N_7032);
nor U7692 (N_7692,N_7226,N_7028);
and U7693 (N_7693,N_7229,N_7258);
nor U7694 (N_7694,N_7331,N_7132);
or U7695 (N_7695,N_7338,N_7227);
nand U7696 (N_7696,N_7103,N_7034);
nand U7697 (N_7697,N_7328,N_7247);
nand U7698 (N_7698,N_7306,N_7349);
nand U7699 (N_7699,N_7266,N_7476);
nand U7700 (N_7700,N_7301,N_7274);
nand U7701 (N_7701,N_7297,N_7311);
nor U7702 (N_7702,N_7020,N_7207);
and U7703 (N_7703,N_7271,N_7216);
and U7704 (N_7704,N_7074,N_7359);
xnor U7705 (N_7705,N_7265,N_7067);
xnor U7706 (N_7706,N_7035,N_7275);
nand U7707 (N_7707,N_7329,N_7168);
and U7708 (N_7708,N_7041,N_7353);
or U7709 (N_7709,N_7393,N_7497);
nand U7710 (N_7710,N_7435,N_7043);
nand U7711 (N_7711,N_7214,N_7333);
xnor U7712 (N_7712,N_7011,N_7072);
nor U7713 (N_7713,N_7111,N_7016);
nand U7714 (N_7714,N_7391,N_7287);
nor U7715 (N_7715,N_7078,N_7259);
nand U7716 (N_7716,N_7422,N_7282);
xor U7717 (N_7717,N_7379,N_7257);
or U7718 (N_7718,N_7473,N_7402);
or U7719 (N_7719,N_7413,N_7157);
or U7720 (N_7720,N_7450,N_7208);
and U7721 (N_7721,N_7340,N_7411);
nor U7722 (N_7722,N_7116,N_7064);
xnor U7723 (N_7723,N_7094,N_7148);
nand U7724 (N_7724,N_7388,N_7079);
nand U7725 (N_7725,N_7026,N_7380);
nand U7726 (N_7726,N_7061,N_7005);
xor U7727 (N_7727,N_7472,N_7179);
nand U7728 (N_7728,N_7070,N_7387);
nand U7729 (N_7729,N_7441,N_7468);
or U7730 (N_7730,N_7013,N_7406);
nor U7731 (N_7731,N_7191,N_7174);
nand U7732 (N_7732,N_7348,N_7188);
xnor U7733 (N_7733,N_7319,N_7399);
xor U7734 (N_7734,N_7186,N_7220);
xnor U7735 (N_7735,N_7355,N_7269);
nor U7736 (N_7736,N_7309,N_7212);
and U7737 (N_7737,N_7288,N_7371);
or U7738 (N_7738,N_7142,N_7213);
xnor U7739 (N_7739,N_7267,N_7184);
nor U7740 (N_7740,N_7054,N_7281);
nand U7741 (N_7741,N_7008,N_7452);
or U7742 (N_7742,N_7050,N_7221);
and U7743 (N_7743,N_7152,N_7144);
nand U7744 (N_7744,N_7339,N_7459);
and U7745 (N_7745,N_7237,N_7167);
nor U7746 (N_7746,N_7318,N_7133);
and U7747 (N_7747,N_7408,N_7119);
nand U7748 (N_7748,N_7263,N_7024);
and U7749 (N_7749,N_7332,N_7419);
nor U7750 (N_7750,N_7344,N_7330);
xor U7751 (N_7751,N_7363,N_7272);
nor U7752 (N_7752,N_7257,N_7011);
nand U7753 (N_7753,N_7347,N_7150);
or U7754 (N_7754,N_7246,N_7242);
or U7755 (N_7755,N_7052,N_7082);
nand U7756 (N_7756,N_7188,N_7091);
nor U7757 (N_7757,N_7169,N_7269);
or U7758 (N_7758,N_7448,N_7203);
nor U7759 (N_7759,N_7375,N_7422);
and U7760 (N_7760,N_7023,N_7499);
nor U7761 (N_7761,N_7035,N_7039);
nand U7762 (N_7762,N_7365,N_7279);
and U7763 (N_7763,N_7262,N_7096);
xnor U7764 (N_7764,N_7206,N_7236);
xnor U7765 (N_7765,N_7360,N_7470);
and U7766 (N_7766,N_7359,N_7477);
xnor U7767 (N_7767,N_7061,N_7372);
nand U7768 (N_7768,N_7019,N_7241);
xnor U7769 (N_7769,N_7350,N_7134);
or U7770 (N_7770,N_7454,N_7057);
nand U7771 (N_7771,N_7016,N_7067);
xnor U7772 (N_7772,N_7029,N_7325);
xor U7773 (N_7773,N_7492,N_7206);
nor U7774 (N_7774,N_7345,N_7164);
xor U7775 (N_7775,N_7335,N_7397);
or U7776 (N_7776,N_7088,N_7246);
nor U7777 (N_7777,N_7418,N_7164);
and U7778 (N_7778,N_7336,N_7402);
xor U7779 (N_7779,N_7291,N_7109);
and U7780 (N_7780,N_7320,N_7090);
and U7781 (N_7781,N_7143,N_7419);
and U7782 (N_7782,N_7446,N_7411);
nor U7783 (N_7783,N_7497,N_7046);
xor U7784 (N_7784,N_7226,N_7256);
nor U7785 (N_7785,N_7354,N_7042);
or U7786 (N_7786,N_7112,N_7243);
and U7787 (N_7787,N_7138,N_7208);
nand U7788 (N_7788,N_7358,N_7015);
nand U7789 (N_7789,N_7247,N_7479);
or U7790 (N_7790,N_7235,N_7400);
or U7791 (N_7791,N_7281,N_7366);
nor U7792 (N_7792,N_7283,N_7214);
and U7793 (N_7793,N_7369,N_7173);
and U7794 (N_7794,N_7088,N_7471);
and U7795 (N_7795,N_7024,N_7003);
or U7796 (N_7796,N_7446,N_7238);
nor U7797 (N_7797,N_7279,N_7472);
and U7798 (N_7798,N_7323,N_7446);
nor U7799 (N_7799,N_7256,N_7428);
and U7800 (N_7800,N_7005,N_7103);
and U7801 (N_7801,N_7070,N_7380);
nand U7802 (N_7802,N_7067,N_7056);
xor U7803 (N_7803,N_7267,N_7347);
nor U7804 (N_7804,N_7163,N_7180);
and U7805 (N_7805,N_7176,N_7293);
nand U7806 (N_7806,N_7136,N_7372);
or U7807 (N_7807,N_7184,N_7275);
xnor U7808 (N_7808,N_7218,N_7383);
xnor U7809 (N_7809,N_7370,N_7456);
nand U7810 (N_7810,N_7469,N_7429);
xor U7811 (N_7811,N_7484,N_7226);
xor U7812 (N_7812,N_7109,N_7478);
or U7813 (N_7813,N_7216,N_7401);
nor U7814 (N_7814,N_7002,N_7333);
or U7815 (N_7815,N_7148,N_7473);
nor U7816 (N_7816,N_7266,N_7128);
nor U7817 (N_7817,N_7443,N_7146);
nand U7818 (N_7818,N_7191,N_7029);
nand U7819 (N_7819,N_7490,N_7057);
or U7820 (N_7820,N_7046,N_7423);
or U7821 (N_7821,N_7062,N_7314);
and U7822 (N_7822,N_7430,N_7026);
nor U7823 (N_7823,N_7243,N_7444);
or U7824 (N_7824,N_7131,N_7045);
and U7825 (N_7825,N_7025,N_7485);
xor U7826 (N_7826,N_7206,N_7291);
xnor U7827 (N_7827,N_7479,N_7149);
nor U7828 (N_7828,N_7042,N_7319);
xnor U7829 (N_7829,N_7108,N_7478);
and U7830 (N_7830,N_7123,N_7233);
and U7831 (N_7831,N_7350,N_7175);
xor U7832 (N_7832,N_7471,N_7391);
or U7833 (N_7833,N_7318,N_7105);
nand U7834 (N_7834,N_7440,N_7109);
xnor U7835 (N_7835,N_7324,N_7102);
xor U7836 (N_7836,N_7008,N_7034);
and U7837 (N_7837,N_7343,N_7429);
and U7838 (N_7838,N_7065,N_7101);
nor U7839 (N_7839,N_7359,N_7239);
and U7840 (N_7840,N_7223,N_7490);
nor U7841 (N_7841,N_7131,N_7374);
or U7842 (N_7842,N_7137,N_7264);
xor U7843 (N_7843,N_7094,N_7462);
nor U7844 (N_7844,N_7006,N_7022);
nand U7845 (N_7845,N_7157,N_7455);
nor U7846 (N_7846,N_7267,N_7274);
nand U7847 (N_7847,N_7411,N_7495);
xnor U7848 (N_7848,N_7167,N_7104);
xor U7849 (N_7849,N_7194,N_7226);
and U7850 (N_7850,N_7354,N_7270);
or U7851 (N_7851,N_7326,N_7392);
and U7852 (N_7852,N_7386,N_7406);
or U7853 (N_7853,N_7236,N_7249);
and U7854 (N_7854,N_7008,N_7075);
and U7855 (N_7855,N_7437,N_7452);
and U7856 (N_7856,N_7180,N_7011);
nor U7857 (N_7857,N_7207,N_7130);
nand U7858 (N_7858,N_7229,N_7113);
nor U7859 (N_7859,N_7328,N_7072);
nor U7860 (N_7860,N_7254,N_7056);
nor U7861 (N_7861,N_7060,N_7263);
or U7862 (N_7862,N_7080,N_7279);
xnor U7863 (N_7863,N_7472,N_7329);
nand U7864 (N_7864,N_7434,N_7249);
xor U7865 (N_7865,N_7390,N_7162);
or U7866 (N_7866,N_7454,N_7011);
nor U7867 (N_7867,N_7484,N_7430);
or U7868 (N_7868,N_7494,N_7178);
and U7869 (N_7869,N_7403,N_7120);
or U7870 (N_7870,N_7143,N_7022);
xnor U7871 (N_7871,N_7039,N_7189);
and U7872 (N_7872,N_7127,N_7130);
xnor U7873 (N_7873,N_7122,N_7105);
nand U7874 (N_7874,N_7101,N_7111);
and U7875 (N_7875,N_7107,N_7106);
xnor U7876 (N_7876,N_7107,N_7031);
xor U7877 (N_7877,N_7423,N_7479);
xor U7878 (N_7878,N_7389,N_7042);
nand U7879 (N_7879,N_7337,N_7169);
nor U7880 (N_7880,N_7176,N_7483);
and U7881 (N_7881,N_7190,N_7467);
or U7882 (N_7882,N_7412,N_7284);
and U7883 (N_7883,N_7189,N_7100);
and U7884 (N_7884,N_7444,N_7108);
and U7885 (N_7885,N_7090,N_7233);
or U7886 (N_7886,N_7374,N_7407);
xor U7887 (N_7887,N_7318,N_7359);
nand U7888 (N_7888,N_7004,N_7293);
and U7889 (N_7889,N_7115,N_7166);
nand U7890 (N_7890,N_7271,N_7207);
or U7891 (N_7891,N_7292,N_7227);
and U7892 (N_7892,N_7291,N_7238);
or U7893 (N_7893,N_7365,N_7042);
nand U7894 (N_7894,N_7439,N_7369);
nor U7895 (N_7895,N_7297,N_7143);
and U7896 (N_7896,N_7276,N_7005);
nor U7897 (N_7897,N_7016,N_7024);
xor U7898 (N_7898,N_7052,N_7308);
xor U7899 (N_7899,N_7127,N_7003);
xnor U7900 (N_7900,N_7365,N_7071);
and U7901 (N_7901,N_7296,N_7463);
xor U7902 (N_7902,N_7372,N_7453);
nor U7903 (N_7903,N_7360,N_7393);
nor U7904 (N_7904,N_7161,N_7412);
xor U7905 (N_7905,N_7005,N_7377);
or U7906 (N_7906,N_7195,N_7208);
nand U7907 (N_7907,N_7339,N_7383);
nor U7908 (N_7908,N_7052,N_7201);
nand U7909 (N_7909,N_7299,N_7086);
xnor U7910 (N_7910,N_7331,N_7445);
xor U7911 (N_7911,N_7339,N_7172);
or U7912 (N_7912,N_7205,N_7096);
nand U7913 (N_7913,N_7422,N_7127);
nand U7914 (N_7914,N_7223,N_7422);
nand U7915 (N_7915,N_7134,N_7483);
and U7916 (N_7916,N_7160,N_7301);
nand U7917 (N_7917,N_7091,N_7327);
or U7918 (N_7918,N_7034,N_7260);
xor U7919 (N_7919,N_7212,N_7272);
nand U7920 (N_7920,N_7376,N_7410);
and U7921 (N_7921,N_7106,N_7145);
nand U7922 (N_7922,N_7375,N_7364);
nor U7923 (N_7923,N_7160,N_7380);
nor U7924 (N_7924,N_7442,N_7495);
nor U7925 (N_7925,N_7203,N_7285);
nor U7926 (N_7926,N_7040,N_7377);
or U7927 (N_7927,N_7218,N_7445);
and U7928 (N_7928,N_7242,N_7475);
nand U7929 (N_7929,N_7483,N_7111);
or U7930 (N_7930,N_7417,N_7487);
xnor U7931 (N_7931,N_7076,N_7476);
or U7932 (N_7932,N_7455,N_7089);
nand U7933 (N_7933,N_7445,N_7249);
nand U7934 (N_7934,N_7076,N_7213);
nand U7935 (N_7935,N_7231,N_7356);
and U7936 (N_7936,N_7283,N_7356);
nor U7937 (N_7937,N_7429,N_7251);
nand U7938 (N_7938,N_7210,N_7086);
and U7939 (N_7939,N_7335,N_7003);
nor U7940 (N_7940,N_7429,N_7345);
or U7941 (N_7941,N_7231,N_7393);
xor U7942 (N_7942,N_7056,N_7166);
xnor U7943 (N_7943,N_7221,N_7364);
nor U7944 (N_7944,N_7169,N_7321);
xor U7945 (N_7945,N_7142,N_7413);
nor U7946 (N_7946,N_7015,N_7181);
nand U7947 (N_7947,N_7330,N_7451);
nand U7948 (N_7948,N_7412,N_7048);
nor U7949 (N_7949,N_7214,N_7218);
xnor U7950 (N_7950,N_7479,N_7129);
or U7951 (N_7951,N_7409,N_7162);
or U7952 (N_7952,N_7083,N_7154);
xnor U7953 (N_7953,N_7429,N_7418);
xor U7954 (N_7954,N_7060,N_7056);
and U7955 (N_7955,N_7180,N_7269);
nor U7956 (N_7956,N_7300,N_7359);
nand U7957 (N_7957,N_7381,N_7310);
nor U7958 (N_7958,N_7426,N_7467);
nand U7959 (N_7959,N_7364,N_7332);
nor U7960 (N_7960,N_7234,N_7367);
or U7961 (N_7961,N_7461,N_7012);
nor U7962 (N_7962,N_7464,N_7196);
nand U7963 (N_7963,N_7486,N_7228);
nor U7964 (N_7964,N_7448,N_7190);
or U7965 (N_7965,N_7306,N_7482);
xnor U7966 (N_7966,N_7152,N_7076);
and U7967 (N_7967,N_7296,N_7338);
nand U7968 (N_7968,N_7230,N_7015);
or U7969 (N_7969,N_7327,N_7418);
nand U7970 (N_7970,N_7421,N_7190);
nor U7971 (N_7971,N_7144,N_7298);
nor U7972 (N_7972,N_7443,N_7197);
xor U7973 (N_7973,N_7307,N_7288);
or U7974 (N_7974,N_7442,N_7459);
nand U7975 (N_7975,N_7419,N_7491);
xnor U7976 (N_7976,N_7131,N_7139);
and U7977 (N_7977,N_7046,N_7104);
or U7978 (N_7978,N_7040,N_7287);
or U7979 (N_7979,N_7146,N_7077);
and U7980 (N_7980,N_7368,N_7497);
nor U7981 (N_7981,N_7086,N_7467);
nor U7982 (N_7982,N_7251,N_7384);
nor U7983 (N_7983,N_7225,N_7340);
xor U7984 (N_7984,N_7364,N_7115);
xnor U7985 (N_7985,N_7283,N_7367);
or U7986 (N_7986,N_7095,N_7282);
xnor U7987 (N_7987,N_7096,N_7475);
nor U7988 (N_7988,N_7134,N_7071);
and U7989 (N_7989,N_7430,N_7079);
nand U7990 (N_7990,N_7408,N_7247);
nor U7991 (N_7991,N_7262,N_7199);
xnor U7992 (N_7992,N_7332,N_7248);
nand U7993 (N_7993,N_7499,N_7141);
or U7994 (N_7994,N_7264,N_7450);
xnor U7995 (N_7995,N_7154,N_7110);
or U7996 (N_7996,N_7484,N_7184);
or U7997 (N_7997,N_7410,N_7293);
xor U7998 (N_7998,N_7195,N_7361);
nor U7999 (N_7999,N_7015,N_7217);
nor U8000 (N_8000,N_7896,N_7883);
and U8001 (N_8001,N_7942,N_7962);
xor U8002 (N_8002,N_7867,N_7843);
and U8003 (N_8003,N_7506,N_7807);
nand U8004 (N_8004,N_7860,N_7939);
nand U8005 (N_8005,N_7610,N_7816);
and U8006 (N_8006,N_7967,N_7877);
nand U8007 (N_8007,N_7830,N_7837);
xnor U8008 (N_8008,N_7707,N_7679);
xor U8009 (N_8009,N_7954,N_7663);
or U8010 (N_8010,N_7561,N_7509);
xor U8011 (N_8011,N_7848,N_7670);
nand U8012 (N_8012,N_7640,N_7990);
or U8013 (N_8013,N_7888,N_7559);
nand U8014 (N_8014,N_7935,N_7708);
nand U8015 (N_8015,N_7534,N_7572);
and U8016 (N_8016,N_7932,N_7842);
and U8017 (N_8017,N_7682,N_7982);
nand U8018 (N_8018,N_7975,N_7964);
xnor U8019 (N_8019,N_7740,N_7666);
or U8020 (N_8020,N_7931,N_7518);
or U8021 (N_8021,N_7858,N_7621);
or U8022 (N_8022,N_7828,N_7758);
nand U8023 (N_8023,N_7531,N_7700);
or U8024 (N_8024,N_7529,N_7885);
or U8025 (N_8025,N_7716,N_7871);
and U8026 (N_8026,N_7650,N_7766);
xnor U8027 (N_8027,N_7907,N_7944);
xor U8028 (N_8028,N_7732,N_7624);
nor U8029 (N_8029,N_7702,N_7738);
xnor U8030 (N_8030,N_7676,N_7511);
nor U8031 (N_8031,N_7917,N_7839);
or U8032 (N_8032,N_7956,N_7642);
and U8033 (N_8033,N_7609,N_7668);
nor U8034 (N_8034,N_7587,N_7535);
and U8035 (N_8035,N_7512,N_7585);
xnor U8036 (N_8036,N_7524,N_7983);
and U8037 (N_8037,N_7658,N_7909);
nand U8038 (N_8038,N_7664,N_7746);
nor U8039 (N_8039,N_7965,N_7603);
and U8040 (N_8040,N_7892,N_7915);
and U8041 (N_8041,N_7726,N_7544);
or U8042 (N_8042,N_7796,N_7783);
and U8043 (N_8043,N_7699,N_7602);
xnor U8044 (N_8044,N_7825,N_7671);
or U8045 (N_8045,N_7727,N_7513);
or U8046 (N_8046,N_7763,N_7813);
xnor U8047 (N_8047,N_7593,N_7951);
nor U8048 (N_8048,N_7734,N_7757);
nand U8049 (N_8049,N_7645,N_7594);
or U8050 (N_8050,N_7809,N_7576);
and U8051 (N_8051,N_7681,N_7779);
nor U8052 (N_8052,N_7634,N_7874);
and U8053 (N_8053,N_7919,N_7749);
nor U8054 (N_8054,N_7756,N_7514);
nand U8055 (N_8055,N_7993,N_7966);
nand U8056 (N_8056,N_7865,N_7656);
nor U8057 (N_8057,N_7523,N_7748);
xnor U8058 (N_8058,N_7810,N_7998);
and U8059 (N_8059,N_7520,N_7550);
xor U8060 (N_8060,N_7677,N_7627);
nand U8061 (N_8061,N_7596,N_7856);
nand U8062 (N_8062,N_7969,N_7878);
xnor U8063 (N_8063,N_7555,N_7882);
or U8064 (N_8064,N_7979,N_7799);
nor U8065 (N_8065,N_7695,N_7884);
xor U8066 (N_8066,N_7812,N_7925);
nand U8067 (N_8067,N_7918,N_7741);
or U8068 (N_8068,N_7521,N_7597);
nor U8069 (N_8069,N_7687,N_7669);
and U8070 (N_8070,N_7528,N_7934);
and U8071 (N_8071,N_7978,N_7920);
nor U8072 (N_8072,N_7971,N_7833);
and U8073 (N_8073,N_7836,N_7557);
and U8074 (N_8074,N_7532,N_7914);
or U8075 (N_8075,N_7853,N_7973);
or U8076 (N_8076,N_7548,N_7578);
nor U8077 (N_8077,N_7575,N_7729);
nand U8078 (N_8078,N_7601,N_7968);
and U8079 (N_8079,N_7751,N_7846);
xor U8080 (N_8080,N_7859,N_7814);
nor U8081 (N_8081,N_7824,N_7574);
and U8082 (N_8082,N_7673,N_7893);
xnor U8083 (N_8083,N_7835,N_7818);
nand U8084 (N_8084,N_7780,N_7616);
xor U8085 (N_8085,N_7921,N_7902);
nor U8086 (N_8086,N_7988,N_7733);
nor U8087 (N_8087,N_7831,N_7638);
and U8088 (N_8088,N_7622,N_7866);
nor U8089 (N_8089,N_7963,N_7996);
nand U8090 (N_8090,N_7887,N_7592);
or U8091 (N_8091,N_7554,N_7560);
nor U8092 (N_8092,N_7608,N_7643);
and U8093 (N_8093,N_7999,N_7569);
and U8094 (N_8094,N_7916,N_7797);
nand U8095 (N_8095,N_7898,N_7508);
nand U8096 (N_8096,N_7644,N_7754);
nor U8097 (N_8097,N_7675,N_7957);
and U8098 (N_8098,N_7713,N_7654);
nand U8099 (N_8099,N_7568,N_7693);
and U8100 (N_8100,N_7571,N_7581);
xnor U8101 (N_8101,N_7960,N_7501);
nand U8102 (N_8102,N_7720,N_7595);
nor U8103 (N_8103,N_7728,N_7753);
or U8104 (N_8104,N_7995,N_7649);
nand U8105 (N_8105,N_7948,N_7742);
nor U8106 (N_8106,N_7710,N_7690);
and U8107 (N_8107,N_7913,N_7847);
xnor U8108 (N_8108,N_7667,N_7771);
or U8109 (N_8109,N_7547,N_7564);
nand U8110 (N_8110,N_7538,N_7850);
nand U8111 (N_8111,N_7711,N_7591);
and U8112 (N_8112,N_7773,N_7541);
and U8113 (N_8113,N_7970,N_7905);
and U8114 (N_8114,N_7659,N_7972);
nand U8115 (N_8115,N_7864,N_7803);
and U8116 (N_8116,N_7718,N_7684);
and U8117 (N_8117,N_7890,N_7764);
or U8118 (N_8118,N_7619,N_7778);
nand U8119 (N_8119,N_7792,N_7774);
nor U8120 (N_8120,N_7721,N_7976);
nand U8121 (N_8121,N_7891,N_7840);
xnor U8122 (N_8122,N_7857,N_7683);
or U8123 (N_8123,N_7637,N_7961);
or U8124 (N_8124,N_7689,N_7904);
nor U8125 (N_8125,N_7895,N_7873);
nand U8126 (N_8126,N_7827,N_7685);
and U8127 (N_8127,N_7519,N_7747);
and U8128 (N_8128,N_7991,N_7879);
or U8129 (N_8129,N_7768,N_7940);
and U8130 (N_8130,N_7880,N_7632);
xnor U8131 (N_8131,N_7826,N_7566);
nand U8132 (N_8132,N_7545,N_7722);
nand U8133 (N_8133,N_7854,N_7906);
and U8134 (N_8134,N_7698,N_7928);
xnor U8135 (N_8135,N_7787,N_7605);
nor U8136 (N_8136,N_7823,N_7974);
nor U8137 (N_8137,N_7762,N_7717);
or U8138 (N_8138,N_7706,N_7598);
nand U8139 (N_8139,N_7793,N_7789);
or U8140 (N_8140,N_7869,N_7556);
nor U8141 (N_8141,N_7590,N_7929);
nand U8142 (N_8142,N_7530,N_7903);
and U8143 (N_8143,N_7811,N_7577);
and U8144 (N_8144,N_7505,N_7750);
and U8145 (N_8145,N_7626,N_7977);
xnor U8146 (N_8146,N_7943,N_7703);
nand U8147 (N_8147,N_7949,N_7984);
xor U8148 (N_8148,N_7985,N_7776);
xnor U8149 (N_8149,N_7772,N_7736);
xor U8150 (N_8150,N_7760,N_7573);
nand U8151 (N_8151,N_7510,N_7938);
and U8152 (N_8152,N_7705,N_7950);
xnor U8153 (N_8153,N_7933,N_7817);
or U8154 (N_8154,N_7770,N_7875);
xor U8155 (N_8155,N_7997,N_7565);
and U8156 (N_8156,N_7680,N_7986);
xor U8157 (N_8157,N_7697,N_7820);
and U8158 (N_8158,N_7923,N_7522);
nor U8159 (N_8159,N_7543,N_7688);
and U8160 (N_8160,N_7936,N_7661);
or U8161 (N_8161,N_7562,N_7804);
or U8162 (N_8162,N_7502,N_7730);
or U8163 (N_8163,N_7795,N_7994);
nor U8164 (N_8164,N_7694,N_7635);
nand U8165 (N_8165,N_7805,N_7852);
nand U8166 (N_8166,N_7737,N_7712);
or U8167 (N_8167,N_7980,N_7719);
and U8168 (N_8168,N_7724,N_7525);
nand U8169 (N_8169,N_7924,N_7855);
and U8170 (N_8170,N_7822,N_7582);
nand U8171 (N_8171,N_7589,N_7851);
nor U8172 (N_8172,N_7900,N_7775);
nand U8173 (N_8173,N_7686,N_7715);
nor U8174 (N_8174,N_7662,N_7629);
xnor U8175 (N_8175,N_7870,N_7819);
nand U8176 (N_8176,N_7672,N_7539);
xnor U8177 (N_8177,N_7692,N_7526);
nand U8178 (N_8178,N_7861,N_7798);
and U8179 (N_8179,N_7599,N_7517);
and U8180 (N_8180,N_7714,N_7500);
and U8181 (N_8181,N_7911,N_7755);
or U8182 (N_8182,N_7845,N_7604);
or U8183 (N_8183,N_7647,N_7941);
nor U8184 (N_8184,N_7612,N_7946);
and U8185 (N_8185,N_7745,N_7927);
xnor U8186 (N_8186,N_7551,N_7868);
nand U8187 (N_8187,N_7841,N_7785);
nor U8188 (N_8188,N_7641,N_7584);
nand U8189 (N_8189,N_7801,N_7701);
nor U8190 (N_8190,N_7665,N_7926);
xor U8191 (N_8191,N_7953,N_7503);
xor U8192 (N_8192,N_7583,N_7876);
or U8193 (N_8193,N_7782,N_7735);
nand U8194 (N_8194,N_7646,N_7691);
nand U8195 (N_8195,N_7981,N_7633);
xnor U8196 (N_8196,N_7628,N_7617);
and U8197 (N_8197,N_7533,N_7655);
nor U8198 (N_8198,N_7800,N_7897);
xnor U8199 (N_8199,N_7791,N_7908);
xnor U8200 (N_8200,N_7821,N_7636);
and U8201 (N_8201,N_7955,N_7777);
nor U8202 (N_8202,N_7704,N_7886);
nor U8203 (N_8203,N_7849,N_7579);
nand U8204 (N_8204,N_7515,N_7620);
or U8205 (N_8205,N_7838,N_7794);
nand U8206 (N_8206,N_7652,N_7537);
nor U8207 (N_8207,N_7606,N_7678);
xor U8208 (N_8208,N_7613,N_7930);
or U8209 (N_8209,N_7657,N_7651);
and U8210 (N_8210,N_7786,N_7992);
or U8211 (N_8211,N_7922,N_7989);
or U8212 (N_8212,N_7894,N_7546);
nor U8213 (N_8213,N_7784,N_7731);
nand U8214 (N_8214,N_7947,N_7630);
or U8215 (N_8215,N_7536,N_7781);
xnor U8216 (N_8216,N_7912,N_7586);
and U8217 (N_8217,N_7767,N_7567);
xnor U8218 (N_8218,N_7611,N_7834);
nand U8219 (N_8219,N_7563,N_7618);
and U8220 (N_8220,N_7802,N_7844);
nor U8221 (N_8221,N_7872,N_7552);
nor U8222 (N_8222,N_7769,N_7881);
and U8223 (N_8223,N_7507,N_7901);
nand U8224 (N_8224,N_7945,N_7765);
or U8225 (N_8225,N_7542,N_7527);
and U8226 (N_8226,N_7549,N_7959);
nand U8227 (N_8227,N_7653,N_7615);
and U8228 (N_8228,N_7504,N_7660);
nand U8229 (N_8229,N_7987,N_7600);
and U8230 (N_8230,N_7614,N_7806);
xnor U8231 (N_8231,N_7623,N_7832);
nand U8232 (N_8232,N_7744,N_7580);
and U8233 (N_8233,N_7739,N_7588);
xor U8234 (N_8234,N_7743,N_7607);
and U8235 (N_8235,N_7790,N_7752);
or U8236 (N_8236,N_7761,N_7815);
nand U8237 (N_8237,N_7829,N_7889);
and U8238 (N_8238,N_7696,N_7553);
nor U8239 (N_8239,N_7674,N_7625);
xor U8240 (N_8240,N_7899,N_7862);
nor U8241 (N_8241,N_7952,N_7570);
nor U8242 (N_8242,N_7910,N_7725);
and U8243 (N_8243,N_7723,N_7648);
or U8244 (N_8244,N_7516,N_7937);
and U8245 (N_8245,N_7540,N_7558);
nor U8246 (N_8246,N_7788,N_7639);
xnor U8247 (N_8247,N_7709,N_7631);
xor U8248 (N_8248,N_7958,N_7863);
nand U8249 (N_8249,N_7808,N_7759);
xnor U8250 (N_8250,N_7745,N_7990);
nand U8251 (N_8251,N_7877,N_7671);
or U8252 (N_8252,N_7518,N_7662);
xnor U8253 (N_8253,N_7556,N_7910);
and U8254 (N_8254,N_7541,N_7817);
nor U8255 (N_8255,N_7618,N_7699);
nor U8256 (N_8256,N_7574,N_7571);
and U8257 (N_8257,N_7928,N_7833);
nor U8258 (N_8258,N_7617,N_7662);
nand U8259 (N_8259,N_7677,N_7906);
and U8260 (N_8260,N_7922,N_7614);
nor U8261 (N_8261,N_7887,N_7832);
nor U8262 (N_8262,N_7849,N_7867);
nor U8263 (N_8263,N_7891,N_7733);
xor U8264 (N_8264,N_7779,N_7829);
and U8265 (N_8265,N_7984,N_7982);
nand U8266 (N_8266,N_7822,N_7510);
nor U8267 (N_8267,N_7591,N_7516);
and U8268 (N_8268,N_7505,N_7845);
xor U8269 (N_8269,N_7633,N_7818);
nor U8270 (N_8270,N_7658,N_7579);
nand U8271 (N_8271,N_7620,N_7650);
nor U8272 (N_8272,N_7541,N_7885);
or U8273 (N_8273,N_7933,N_7855);
or U8274 (N_8274,N_7942,N_7670);
nor U8275 (N_8275,N_7864,N_7627);
nand U8276 (N_8276,N_7748,N_7605);
xnor U8277 (N_8277,N_7845,N_7740);
xnor U8278 (N_8278,N_7737,N_7786);
nand U8279 (N_8279,N_7661,N_7690);
xor U8280 (N_8280,N_7618,N_7734);
nor U8281 (N_8281,N_7537,N_7831);
and U8282 (N_8282,N_7795,N_7894);
xor U8283 (N_8283,N_7510,N_7722);
nand U8284 (N_8284,N_7856,N_7699);
or U8285 (N_8285,N_7694,N_7733);
xor U8286 (N_8286,N_7941,N_7971);
or U8287 (N_8287,N_7752,N_7979);
or U8288 (N_8288,N_7521,N_7835);
xnor U8289 (N_8289,N_7854,N_7795);
and U8290 (N_8290,N_7591,N_7503);
nand U8291 (N_8291,N_7510,N_7799);
xor U8292 (N_8292,N_7903,N_7816);
or U8293 (N_8293,N_7619,N_7970);
xor U8294 (N_8294,N_7998,N_7884);
nand U8295 (N_8295,N_7962,N_7996);
nand U8296 (N_8296,N_7741,N_7946);
nor U8297 (N_8297,N_7512,N_7972);
nor U8298 (N_8298,N_7722,N_7859);
and U8299 (N_8299,N_7515,N_7578);
xnor U8300 (N_8300,N_7588,N_7590);
nor U8301 (N_8301,N_7613,N_7913);
xnor U8302 (N_8302,N_7738,N_7700);
xor U8303 (N_8303,N_7846,N_7875);
or U8304 (N_8304,N_7858,N_7963);
or U8305 (N_8305,N_7779,N_7600);
xnor U8306 (N_8306,N_7608,N_7808);
nand U8307 (N_8307,N_7880,N_7942);
xnor U8308 (N_8308,N_7640,N_7870);
nand U8309 (N_8309,N_7938,N_7841);
xnor U8310 (N_8310,N_7841,N_7668);
nor U8311 (N_8311,N_7625,N_7677);
xnor U8312 (N_8312,N_7877,N_7542);
and U8313 (N_8313,N_7951,N_7584);
nor U8314 (N_8314,N_7645,N_7679);
nand U8315 (N_8315,N_7910,N_7878);
and U8316 (N_8316,N_7758,N_7692);
xnor U8317 (N_8317,N_7735,N_7660);
nand U8318 (N_8318,N_7568,N_7852);
or U8319 (N_8319,N_7680,N_7647);
and U8320 (N_8320,N_7931,N_7949);
and U8321 (N_8321,N_7949,N_7544);
xnor U8322 (N_8322,N_7528,N_7653);
and U8323 (N_8323,N_7809,N_7782);
and U8324 (N_8324,N_7888,N_7986);
nand U8325 (N_8325,N_7598,N_7571);
xor U8326 (N_8326,N_7627,N_7517);
nand U8327 (N_8327,N_7856,N_7958);
nand U8328 (N_8328,N_7604,N_7828);
nand U8329 (N_8329,N_7925,N_7536);
and U8330 (N_8330,N_7711,N_7948);
xor U8331 (N_8331,N_7712,N_7870);
or U8332 (N_8332,N_7768,N_7634);
nor U8333 (N_8333,N_7942,N_7641);
xnor U8334 (N_8334,N_7626,N_7648);
nand U8335 (N_8335,N_7503,N_7993);
nand U8336 (N_8336,N_7778,N_7573);
xnor U8337 (N_8337,N_7534,N_7634);
and U8338 (N_8338,N_7621,N_7724);
xnor U8339 (N_8339,N_7961,N_7835);
nor U8340 (N_8340,N_7848,N_7573);
nor U8341 (N_8341,N_7767,N_7648);
or U8342 (N_8342,N_7503,N_7543);
or U8343 (N_8343,N_7704,N_7774);
or U8344 (N_8344,N_7716,N_7947);
xnor U8345 (N_8345,N_7648,N_7555);
or U8346 (N_8346,N_7995,N_7733);
nor U8347 (N_8347,N_7955,N_7758);
and U8348 (N_8348,N_7742,N_7708);
and U8349 (N_8349,N_7973,N_7627);
nand U8350 (N_8350,N_7768,N_7851);
or U8351 (N_8351,N_7630,N_7775);
and U8352 (N_8352,N_7787,N_7748);
or U8353 (N_8353,N_7745,N_7877);
nand U8354 (N_8354,N_7982,N_7995);
nor U8355 (N_8355,N_7574,N_7768);
xor U8356 (N_8356,N_7960,N_7889);
or U8357 (N_8357,N_7557,N_7957);
nand U8358 (N_8358,N_7615,N_7964);
and U8359 (N_8359,N_7701,N_7595);
or U8360 (N_8360,N_7766,N_7964);
or U8361 (N_8361,N_7587,N_7527);
xnor U8362 (N_8362,N_7854,N_7504);
and U8363 (N_8363,N_7902,N_7971);
and U8364 (N_8364,N_7850,N_7743);
nand U8365 (N_8365,N_7809,N_7983);
and U8366 (N_8366,N_7979,N_7609);
and U8367 (N_8367,N_7575,N_7564);
xor U8368 (N_8368,N_7562,N_7632);
xor U8369 (N_8369,N_7553,N_7518);
nor U8370 (N_8370,N_7894,N_7545);
xnor U8371 (N_8371,N_7517,N_7776);
xnor U8372 (N_8372,N_7864,N_7669);
or U8373 (N_8373,N_7603,N_7756);
and U8374 (N_8374,N_7855,N_7626);
or U8375 (N_8375,N_7876,N_7531);
or U8376 (N_8376,N_7567,N_7971);
nand U8377 (N_8377,N_7806,N_7913);
nor U8378 (N_8378,N_7909,N_7582);
nand U8379 (N_8379,N_7610,N_7674);
and U8380 (N_8380,N_7536,N_7686);
xnor U8381 (N_8381,N_7964,N_7721);
xor U8382 (N_8382,N_7645,N_7543);
nand U8383 (N_8383,N_7967,N_7998);
and U8384 (N_8384,N_7787,N_7552);
nand U8385 (N_8385,N_7625,N_7936);
xor U8386 (N_8386,N_7848,N_7936);
or U8387 (N_8387,N_7968,N_7552);
or U8388 (N_8388,N_7925,N_7606);
xor U8389 (N_8389,N_7776,N_7827);
xnor U8390 (N_8390,N_7824,N_7736);
nand U8391 (N_8391,N_7892,N_7761);
nor U8392 (N_8392,N_7503,N_7852);
nand U8393 (N_8393,N_7862,N_7988);
and U8394 (N_8394,N_7913,N_7840);
and U8395 (N_8395,N_7624,N_7940);
nor U8396 (N_8396,N_7642,N_7544);
xnor U8397 (N_8397,N_7981,N_7962);
nand U8398 (N_8398,N_7535,N_7944);
xor U8399 (N_8399,N_7694,N_7644);
nor U8400 (N_8400,N_7923,N_7581);
and U8401 (N_8401,N_7946,N_7743);
xnor U8402 (N_8402,N_7520,N_7870);
nor U8403 (N_8403,N_7730,N_7591);
xor U8404 (N_8404,N_7714,N_7692);
and U8405 (N_8405,N_7962,N_7818);
and U8406 (N_8406,N_7833,N_7987);
or U8407 (N_8407,N_7531,N_7897);
xor U8408 (N_8408,N_7563,N_7746);
or U8409 (N_8409,N_7616,N_7893);
and U8410 (N_8410,N_7927,N_7903);
xor U8411 (N_8411,N_7803,N_7684);
nor U8412 (N_8412,N_7547,N_7697);
nor U8413 (N_8413,N_7526,N_7620);
nor U8414 (N_8414,N_7530,N_7844);
xnor U8415 (N_8415,N_7825,N_7857);
or U8416 (N_8416,N_7744,N_7849);
and U8417 (N_8417,N_7947,N_7941);
and U8418 (N_8418,N_7865,N_7780);
and U8419 (N_8419,N_7968,N_7982);
or U8420 (N_8420,N_7665,N_7539);
or U8421 (N_8421,N_7602,N_7752);
nand U8422 (N_8422,N_7551,N_7785);
xor U8423 (N_8423,N_7622,N_7777);
nor U8424 (N_8424,N_7560,N_7892);
or U8425 (N_8425,N_7984,N_7733);
or U8426 (N_8426,N_7685,N_7933);
and U8427 (N_8427,N_7574,N_7546);
or U8428 (N_8428,N_7799,N_7939);
nand U8429 (N_8429,N_7651,N_7840);
or U8430 (N_8430,N_7779,N_7546);
nand U8431 (N_8431,N_7600,N_7847);
xor U8432 (N_8432,N_7703,N_7583);
and U8433 (N_8433,N_7923,N_7869);
nor U8434 (N_8434,N_7525,N_7651);
or U8435 (N_8435,N_7670,N_7944);
xnor U8436 (N_8436,N_7722,N_7962);
nor U8437 (N_8437,N_7593,N_7578);
or U8438 (N_8438,N_7935,N_7887);
or U8439 (N_8439,N_7723,N_7824);
nand U8440 (N_8440,N_7809,N_7568);
nand U8441 (N_8441,N_7612,N_7715);
xnor U8442 (N_8442,N_7962,N_7776);
and U8443 (N_8443,N_7878,N_7746);
or U8444 (N_8444,N_7811,N_7749);
xnor U8445 (N_8445,N_7544,N_7772);
and U8446 (N_8446,N_7533,N_7633);
or U8447 (N_8447,N_7662,N_7824);
or U8448 (N_8448,N_7804,N_7650);
nand U8449 (N_8449,N_7623,N_7704);
nand U8450 (N_8450,N_7709,N_7554);
nand U8451 (N_8451,N_7541,N_7851);
xor U8452 (N_8452,N_7720,N_7678);
or U8453 (N_8453,N_7689,N_7651);
or U8454 (N_8454,N_7511,N_7726);
nor U8455 (N_8455,N_7936,N_7650);
nor U8456 (N_8456,N_7678,N_7666);
nor U8457 (N_8457,N_7509,N_7936);
xnor U8458 (N_8458,N_7928,N_7911);
or U8459 (N_8459,N_7793,N_7620);
or U8460 (N_8460,N_7563,N_7541);
nand U8461 (N_8461,N_7823,N_7955);
xnor U8462 (N_8462,N_7981,N_7891);
nand U8463 (N_8463,N_7551,N_7906);
and U8464 (N_8464,N_7536,N_7948);
and U8465 (N_8465,N_7896,N_7903);
xor U8466 (N_8466,N_7635,N_7801);
and U8467 (N_8467,N_7718,N_7986);
or U8468 (N_8468,N_7949,N_7792);
nand U8469 (N_8469,N_7997,N_7810);
and U8470 (N_8470,N_7868,N_7961);
xor U8471 (N_8471,N_7767,N_7875);
nand U8472 (N_8472,N_7741,N_7771);
xor U8473 (N_8473,N_7650,N_7556);
or U8474 (N_8474,N_7817,N_7833);
nand U8475 (N_8475,N_7686,N_7875);
and U8476 (N_8476,N_7565,N_7836);
nor U8477 (N_8477,N_7503,N_7602);
and U8478 (N_8478,N_7738,N_7581);
nand U8479 (N_8479,N_7803,N_7664);
nor U8480 (N_8480,N_7983,N_7537);
and U8481 (N_8481,N_7859,N_7579);
nor U8482 (N_8482,N_7974,N_7950);
and U8483 (N_8483,N_7556,N_7925);
nand U8484 (N_8484,N_7811,N_7689);
xnor U8485 (N_8485,N_7503,N_7821);
nor U8486 (N_8486,N_7520,N_7807);
nor U8487 (N_8487,N_7630,N_7882);
xor U8488 (N_8488,N_7938,N_7677);
nor U8489 (N_8489,N_7623,N_7569);
xor U8490 (N_8490,N_7864,N_7736);
or U8491 (N_8491,N_7815,N_7780);
or U8492 (N_8492,N_7716,N_7918);
nand U8493 (N_8493,N_7657,N_7626);
xnor U8494 (N_8494,N_7707,N_7722);
nand U8495 (N_8495,N_7852,N_7587);
and U8496 (N_8496,N_7856,N_7967);
or U8497 (N_8497,N_7642,N_7849);
xnor U8498 (N_8498,N_7673,N_7696);
nor U8499 (N_8499,N_7854,N_7519);
nor U8500 (N_8500,N_8407,N_8041);
and U8501 (N_8501,N_8215,N_8387);
xnor U8502 (N_8502,N_8152,N_8265);
nand U8503 (N_8503,N_8168,N_8287);
or U8504 (N_8504,N_8412,N_8175);
xnor U8505 (N_8505,N_8178,N_8472);
nand U8506 (N_8506,N_8317,N_8151);
or U8507 (N_8507,N_8065,N_8027);
xor U8508 (N_8508,N_8115,N_8224);
or U8509 (N_8509,N_8363,N_8286);
nand U8510 (N_8510,N_8309,N_8190);
nand U8511 (N_8511,N_8171,N_8100);
nand U8512 (N_8512,N_8433,N_8005);
nor U8513 (N_8513,N_8268,N_8052);
nand U8514 (N_8514,N_8166,N_8444);
xnor U8515 (N_8515,N_8495,N_8291);
nand U8516 (N_8516,N_8183,N_8246);
nor U8517 (N_8517,N_8223,N_8231);
nor U8518 (N_8518,N_8322,N_8455);
and U8519 (N_8519,N_8049,N_8182);
or U8520 (N_8520,N_8256,N_8149);
and U8521 (N_8521,N_8055,N_8457);
nor U8522 (N_8522,N_8078,N_8283);
xor U8523 (N_8523,N_8408,N_8478);
nor U8524 (N_8524,N_8276,N_8432);
nor U8525 (N_8525,N_8060,N_8150);
nand U8526 (N_8526,N_8260,N_8333);
or U8527 (N_8527,N_8370,N_8192);
or U8528 (N_8528,N_8430,N_8435);
nor U8529 (N_8529,N_8302,N_8127);
nor U8530 (N_8530,N_8353,N_8044);
nor U8531 (N_8531,N_8319,N_8138);
xnor U8532 (N_8532,N_8038,N_8063);
and U8533 (N_8533,N_8320,N_8101);
nand U8534 (N_8534,N_8311,N_8380);
or U8535 (N_8535,N_8070,N_8263);
nand U8536 (N_8536,N_8314,N_8419);
or U8537 (N_8537,N_8179,N_8176);
nand U8538 (N_8538,N_8146,N_8340);
nand U8539 (N_8539,N_8393,N_8219);
xnor U8540 (N_8540,N_8154,N_8191);
nand U8541 (N_8541,N_8185,N_8004);
xor U8542 (N_8542,N_8173,N_8446);
and U8543 (N_8543,N_8082,N_8274);
or U8544 (N_8544,N_8253,N_8003);
nand U8545 (N_8545,N_8037,N_8372);
and U8546 (N_8546,N_8139,N_8277);
nand U8547 (N_8547,N_8076,N_8424);
nand U8548 (N_8548,N_8418,N_8374);
nor U8549 (N_8549,N_8386,N_8232);
or U8550 (N_8550,N_8062,N_8362);
nor U8551 (N_8551,N_8259,N_8328);
or U8552 (N_8552,N_8463,N_8329);
nor U8553 (N_8553,N_8244,N_8261);
or U8554 (N_8554,N_8264,N_8066);
nand U8555 (N_8555,N_8343,N_8214);
or U8556 (N_8556,N_8113,N_8352);
or U8557 (N_8557,N_8327,N_8383);
or U8558 (N_8558,N_8085,N_8011);
nor U8559 (N_8559,N_8077,N_8258);
xnor U8560 (N_8560,N_8415,N_8434);
nor U8561 (N_8561,N_8459,N_8071);
nor U8562 (N_8562,N_8184,N_8417);
and U8563 (N_8563,N_8290,N_8086);
nand U8564 (N_8564,N_8394,N_8339);
or U8565 (N_8565,N_8292,N_8121);
xor U8566 (N_8566,N_8431,N_8324);
nor U8567 (N_8567,N_8491,N_8125);
and U8568 (N_8568,N_8451,N_8300);
xor U8569 (N_8569,N_8129,N_8002);
xor U8570 (N_8570,N_8306,N_8072);
and U8571 (N_8571,N_8046,N_8091);
or U8572 (N_8572,N_8128,N_8081);
nor U8573 (N_8573,N_8487,N_8064);
nand U8574 (N_8574,N_8198,N_8376);
nand U8575 (N_8575,N_8470,N_8388);
xor U8576 (N_8576,N_8498,N_8469);
nand U8577 (N_8577,N_8123,N_8104);
and U8578 (N_8578,N_8087,N_8272);
and U8579 (N_8579,N_8028,N_8405);
and U8580 (N_8580,N_8270,N_8172);
xnor U8581 (N_8581,N_8043,N_8134);
nand U8582 (N_8582,N_8426,N_8398);
or U8583 (N_8583,N_8341,N_8209);
nor U8584 (N_8584,N_8366,N_8312);
nand U8585 (N_8585,N_8102,N_8051);
nor U8586 (N_8586,N_8026,N_8120);
xor U8587 (N_8587,N_8437,N_8228);
nand U8588 (N_8588,N_8008,N_8109);
xnor U8589 (N_8589,N_8403,N_8156);
and U8590 (N_8590,N_8053,N_8461);
and U8591 (N_8591,N_8220,N_8203);
xnor U8592 (N_8592,N_8230,N_8036);
nand U8593 (N_8593,N_8337,N_8497);
xnor U8594 (N_8594,N_8208,N_8164);
and U8595 (N_8595,N_8323,N_8448);
nor U8596 (N_8596,N_8254,N_8089);
or U8597 (N_8597,N_8382,N_8019);
or U8598 (N_8598,N_8371,N_8465);
nor U8599 (N_8599,N_8217,N_8344);
or U8600 (N_8600,N_8480,N_8159);
xnor U8601 (N_8601,N_8474,N_8485);
and U8602 (N_8602,N_8092,N_8103);
nand U8603 (N_8603,N_8428,N_8143);
nand U8604 (N_8604,N_8169,N_8251);
nor U8605 (N_8605,N_8452,N_8356);
or U8606 (N_8606,N_8367,N_8385);
or U8607 (N_8607,N_8075,N_8117);
nand U8608 (N_8608,N_8464,N_8416);
or U8609 (N_8609,N_8364,N_8476);
nand U8610 (N_8610,N_8212,N_8449);
and U8611 (N_8611,N_8018,N_8155);
and U8612 (N_8612,N_8301,N_8310);
nor U8613 (N_8613,N_8048,N_8020);
xnor U8614 (N_8614,N_8330,N_8315);
nand U8615 (N_8615,N_8017,N_8069);
or U8616 (N_8616,N_8397,N_8411);
nand U8617 (N_8617,N_8378,N_8332);
nand U8618 (N_8618,N_8186,N_8074);
nand U8619 (N_8619,N_8318,N_8379);
nand U8620 (N_8620,N_8174,N_8181);
xnor U8621 (N_8621,N_8409,N_8458);
nor U8622 (N_8622,N_8079,N_8438);
xnor U8623 (N_8623,N_8357,N_8029);
nand U8624 (N_8624,N_8493,N_8222);
nand U8625 (N_8625,N_8421,N_8381);
and U8626 (N_8626,N_8250,N_8471);
and U8627 (N_8627,N_8110,N_8187);
nor U8628 (N_8628,N_8000,N_8450);
nand U8629 (N_8629,N_8006,N_8369);
or U8630 (N_8630,N_8202,N_8188);
or U8631 (N_8631,N_8278,N_8242);
nand U8632 (N_8632,N_8460,N_8475);
nand U8633 (N_8633,N_8249,N_8453);
nor U8634 (N_8634,N_8401,N_8289);
and U8635 (N_8635,N_8033,N_8130);
nor U8636 (N_8636,N_8090,N_8200);
xor U8637 (N_8637,N_8359,N_8294);
and U8638 (N_8638,N_8484,N_8167);
xnor U8639 (N_8639,N_8454,N_8210);
and U8640 (N_8640,N_8161,N_8269);
nor U8641 (N_8641,N_8482,N_8486);
and U8642 (N_8642,N_8271,N_8354);
xnor U8643 (N_8643,N_8410,N_8207);
or U8644 (N_8644,N_8084,N_8425);
nand U8645 (N_8645,N_8313,N_8299);
nand U8646 (N_8646,N_8334,N_8441);
and U8647 (N_8647,N_8439,N_8384);
or U8648 (N_8648,N_8336,N_8204);
nand U8649 (N_8649,N_8016,N_8023);
nor U8650 (N_8650,N_8132,N_8298);
nand U8651 (N_8651,N_8413,N_8481);
xor U8652 (N_8652,N_8377,N_8247);
and U8653 (N_8653,N_8050,N_8303);
or U8654 (N_8654,N_8427,N_8349);
nor U8655 (N_8655,N_8035,N_8494);
xnor U8656 (N_8656,N_8096,N_8236);
and U8657 (N_8657,N_8177,N_8348);
xnor U8658 (N_8658,N_8395,N_8252);
xnor U8659 (N_8659,N_8429,N_8281);
nor U8660 (N_8660,N_8248,N_8285);
and U8661 (N_8661,N_8282,N_8293);
and U8662 (N_8662,N_8373,N_8467);
and U8663 (N_8663,N_8124,N_8400);
or U8664 (N_8664,N_8445,N_8014);
and U8665 (N_8665,N_8045,N_8304);
nor U8666 (N_8666,N_8468,N_8047);
nor U8667 (N_8667,N_8153,N_8094);
or U8668 (N_8668,N_8447,N_8233);
nand U8669 (N_8669,N_8194,N_8034);
and U8670 (N_8670,N_8402,N_8201);
and U8671 (N_8671,N_8483,N_8114);
xor U8672 (N_8672,N_8112,N_8107);
or U8673 (N_8673,N_8158,N_8221);
or U8674 (N_8674,N_8105,N_8391);
or U8675 (N_8675,N_8197,N_8010);
or U8676 (N_8676,N_8142,N_8144);
nand U8677 (N_8677,N_8346,N_8414);
xnor U8678 (N_8678,N_8145,N_8466);
or U8679 (N_8679,N_8056,N_8436);
or U8680 (N_8680,N_8496,N_8307);
xor U8681 (N_8681,N_8406,N_8157);
nor U8682 (N_8682,N_8147,N_8245);
and U8683 (N_8683,N_8227,N_8325);
nor U8684 (N_8684,N_8342,N_8326);
or U8685 (N_8685,N_8358,N_8443);
or U8686 (N_8686,N_8226,N_8106);
nand U8687 (N_8687,N_8375,N_8235);
nand U8688 (N_8688,N_8073,N_8012);
and U8689 (N_8689,N_8141,N_8296);
and U8690 (N_8690,N_8135,N_8345);
or U8691 (N_8691,N_8279,N_8389);
and U8692 (N_8692,N_8030,N_8059);
and U8693 (N_8693,N_8039,N_8396);
nor U8694 (N_8694,N_8499,N_8473);
nor U8695 (N_8695,N_8390,N_8361);
nor U8696 (N_8696,N_8116,N_8237);
and U8697 (N_8697,N_8098,N_8218);
xor U8698 (N_8698,N_8392,N_8024);
and U8699 (N_8699,N_8133,N_8488);
nand U8700 (N_8700,N_8280,N_8216);
nand U8701 (N_8701,N_8067,N_8255);
or U8702 (N_8702,N_8288,N_8213);
nand U8703 (N_8703,N_8021,N_8351);
and U8704 (N_8704,N_8492,N_8308);
nor U8705 (N_8705,N_8205,N_8243);
nand U8706 (N_8706,N_8225,N_8399);
or U8707 (N_8707,N_8032,N_8331);
xnor U8708 (N_8708,N_8080,N_8119);
and U8709 (N_8709,N_8347,N_8099);
or U8710 (N_8710,N_8054,N_8257);
nand U8711 (N_8711,N_8489,N_8211);
and U8712 (N_8712,N_8097,N_8022);
or U8713 (N_8713,N_8316,N_8365);
nor U8714 (N_8714,N_8241,N_8058);
xnor U8715 (N_8715,N_8111,N_8170);
or U8716 (N_8716,N_8360,N_8136);
xnor U8717 (N_8717,N_8490,N_8015);
and U8718 (N_8718,N_8238,N_8338);
and U8719 (N_8719,N_8275,N_8462);
or U8720 (N_8720,N_8163,N_8456);
and U8721 (N_8721,N_8442,N_8042);
nand U8722 (N_8722,N_8189,N_8009);
nor U8723 (N_8723,N_8262,N_8355);
xor U8724 (N_8724,N_8126,N_8404);
xnor U8725 (N_8725,N_8479,N_8239);
nand U8726 (N_8726,N_8140,N_8148);
xor U8727 (N_8727,N_8165,N_8284);
or U8728 (N_8728,N_8093,N_8195);
nor U8729 (N_8729,N_8122,N_8013);
or U8730 (N_8730,N_8180,N_8321);
nor U8731 (N_8731,N_8083,N_8040);
and U8732 (N_8732,N_8422,N_8440);
nor U8733 (N_8733,N_8206,N_8108);
or U8734 (N_8734,N_8088,N_8229);
nor U8735 (N_8735,N_8335,N_8031);
and U8736 (N_8736,N_8267,N_8160);
xnor U8737 (N_8737,N_8137,N_8295);
or U8738 (N_8738,N_8007,N_8057);
nor U8739 (N_8739,N_8273,N_8350);
xnor U8740 (N_8740,N_8118,N_8068);
nand U8741 (N_8741,N_8001,N_8196);
and U8742 (N_8742,N_8266,N_8193);
and U8743 (N_8743,N_8368,N_8234);
xnor U8744 (N_8744,N_8162,N_8131);
and U8745 (N_8745,N_8297,N_8240);
nor U8746 (N_8746,N_8199,N_8095);
nor U8747 (N_8747,N_8061,N_8420);
and U8748 (N_8748,N_8477,N_8305);
nand U8749 (N_8749,N_8025,N_8423);
xnor U8750 (N_8750,N_8180,N_8027);
and U8751 (N_8751,N_8471,N_8273);
nor U8752 (N_8752,N_8156,N_8294);
xnor U8753 (N_8753,N_8421,N_8043);
or U8754 (N_8754,N_8410,N_8435);
and U8755 (N_8755,N_8435,N_8149);
and U8756 (N_8756,N_8448,N_8341);
nor U8757 (N_8757,N_8434,N_8195);
and U8758 (N_8758,N_8356,N_8234);
nor U8759 (N_8759,N_8084,N_8139);
and U8760 (N_8760,N_8201,N_8139);
and U8761 (N_8761,N_8289,N_8035);
nor U8762 (N_8762,N_8467,N_8345);
nor U8763 (N_8763,N_8209,N_8068);
and U8764 (N_8764,N_8491,N_8243);
and U8765 (N_8765,N_8364,N_8347);
nor U8766 (N_8766,N_8025,N_8037);
and U8767 (N_8767,N_8243,N_8272);
nor U8768 (N_8768,N_8352,N_8097);
nor U8769 (N_8769,N_8214,N_8062);
nor U8770 (N_8770,N_8363,N_8463);
nor U8771 (N_8771,N_8003,N_8098);
and U8772 (N_8772,N_8298,N_8059);
xor U8773 (N_8773,N_8304,N_8345);
nand U8774 (N_8774,N_8410,N_8192);
nor U8775 (N_8775,N_8452,N_8129);
nor U8776 (N_8776,N_8468,N_8358);
or U8777 (N_8777,N_8213,N_8241);
and U8778 (N_8778,N_8240,N_8002);
xor U8779 (N_8779,N_8137,N_8423);
nor U8780 (N_8780,N_8296,N_8143);
xnor U8781 (N_8781,N_8187,N_8244);
and U8782 (N_8782,N_8094,N_8308);
or U8783 (N_8783,N_8033,N_8153);
nor U8784 (N_8784,N_8300,N_8100);
nor U8785 (N_8785,N_8428,N_8134);
nor U8786 (N_8786,N_8425,N_8239);
nand U8787 (N_8787,N_8253,N_8389);
nand U8788 (N_8788,N_8228,N_8260);
and U8789 (N_8789,N_8164,N_8355);
nor U8790 (N_8790,N_8090,N_8035);
nand U8791 (N_8791,N_8358,N_8485);
nor U8792 (N_8792,N_8206,N_8165);
or U8793 (N_8793,N_8485,N_8147);
nor U8794 (N_8794,N_8356,N_8105);
xnor U8795 (N_8795,N_8380,N_8096);
and U8796 (N_8796,N_8390,N_8232);
or U8797 (N_8797,N_8309,N_8206);
or U8798 (N_8798,N_8143,N_8466);
xor U8799 (N_8799,N_8163,N_8353);
xor U8800 (N_8800,N_8169,N_8184);
nand U8801 (N_8801,N_8185,N_8403);
nand U8802 (N_8802,N_8104,N_8024);
nor U8803 (N_8803,N_8470,N_8011);
or U8804 (N_8804,N_8052,N_8408);
xnor U8805 (N_8805,N_8401,N_8415);
nor U8806 (N_8806,N_8338,N_8402);
and U8807 (N_8807,N_8449,N_8427);
or U8808 (N_8808,N_8103,N_8385);
nand U8809 (N_8809,N_8130,N_8073);
nand U8810 (N_8810,N_8154,N_8274);
xnor U8811 (N_8811,N_8188,N_8261);
xor U8812 (N_8812,N_8422,N_8441);
nor U8813 (N_8813,N_8398,N_8346);
and U8814 (N_8814,N_8013,N_8445);
or U8815 (N_8815,N_8451,N_8080);
and U8816 (N_8816,N_8083,N_8200);
and U8817 (N_8817,N_8034,N_8291);
nand U8818 (N_8818,N_8333,N_8446);
xnor U8819 (N_8819,N_8394,N_8487);
and U8820 (N_8820,N_8270,N_8108);
nand U8821 (N_8821,N_8335,N_8123);
and U8822 (N_8822,N_8254,N_8053);
or U8823 (N_8823,N_8372,N_8394);
or U8824 (N_8824,N_8198,N_8142);
or U8825 (N_8825,N_8132,N_8126);
xnor U8826 (N_8826,N_8349,N_8336);
nor U8827 (N_8827,N_8058,N_8228);
xnor U8828 (N_8828,N_8234,N_8376);
xnor U8829 (N_8829,N_8146,N_8174);
nor U8830 (N_8830,N_8312,N_8381);
or U8831 (N_8831,N_8246,N_8391);
nor U8832 (N_8832,N_8459,N_8358);
nor U8833 (N_8833,N_8099,N_8292);
and U8834 (N_8834,N_8395,N_8341);
nor U8835 (N_8835,N_8058,N_8213);
and U8836 (N_8836,N_8257,N_8358);
nor U8837 (N_8837,N_8355,N_8148);
and U8838 (N_8838,N_8309,N_8037);
xnor U8839 (N_8839,N_8088,N_8187);
or U8840 (N_8840,N_8288,N_8334);
nor U8841 (N_8841,N_8199,N_8083);
and U8842 (N_8842,N_8484,N_8122);
and U8843 (N_8843,N_8267,N_8132);
and U8844 (N_8844,N_8461,N_8475);
xnor U8845 (N_8845,N_8200,N_8019);
and U8846 (N_8846,N_8499,N_8317);
xnor U8847 (N_8847,N_8409,N_8434);
and U8848 (N_8848,N_8387,N_8062);
or U8849 (N_8849,N_8326,N_8124);
and U8850 (N_8850,N_8390,N_8278);
or U8851 (N_8851,N_8257,N_8425);
and U8852 (N_8852,N_8073,N_8499);
xnor U8853 (N_8853,N_8314,N_8214);
and U8854 (N_8854,N_8021,N_8203);
nor U8855 (N_8855,N_8326,N_8235);
nand U8856 (N_8856,N_8163,N_8157);
nand U8857 (N_8857,N_8397,N_8052);
or U8858 (N_8858,N_8179,N_8486);
xnor U8859 (N_8859,N_8242,N_8002);
nand U8860 (N_8860,N_8142,N_8197);
nor U8861 (N_8861,N_8046,N_8347);
nor U8862 (N_8862,N_8465,N_8102);
and U8863 (N_8863,N_8071,N_8159);
xnor U8864 (N_8864,N_8068,N_8165);
and U8865 (N_8865,N_8197,N_8333);
and U8866 (N_8866,N_8493,N_8263);
xnor U8867 (N_8867,N_8189,N_8253);
nor U8868 (N_8868,N_8309,N_8379);
nand U8869 (N_8869,N_8332,N_8132);
nor U8870 (N_8870,N_8308,N_8080);
nand U8871 (N_8871,N_8097,N_8310);
and U8872 (N_8872,N_8113,N_8205);
or U8873 (N_8873,N_8012,N_8136);
and U8874 (N_8874,N_8050,N_8079);
nand U8875 (N_8875,N_8139,N_8426);
or U8876 (N_8876,N_8004,N_8067);
or U8877 (N_8877,N_8466,N_8058);
nand U8878 (N_8878,N_8112,N_8029);
or U8879 (N_8879,N_8379,N_8337);
xnor U8880 (N_8880,N_8346,N_8131);
nor U8881 (N_8881,N_8457,N_8343);
or U8882 (N_8882,N_8282,N_8400);
and U8883 (N_8883,N_8420,N_8142);
nand U8884 (N_8884,N_8008,N_8389);
or U8885 (N_8885,N_8383,N_8106);
or U8886 (N_8886,N_8071,N_8016);
nor U8887 (N_8887,N_8498,N_8447);
or U8888 (N_8888,N_8035,N_8357);
nand U8889 (N_8889,N_8429,N_8046);
and U8890 (N_8890,N_8057,N_8375);
or U8891 (N_8891,N_8134,N_8009);
nor U8892 (N_8892,N_8388,N_8034);
nand U8893 (N_8893,N_8300,N_8488);
xor U8894 (N_8894,N_8040,N_8345);
and U8895 (N_8895,N_8150,N_8004);
or U8896 (N_8896,N_8015,N_8006);
xnor U8897 (N_8897,N_8368,N_8160);
xor U8898 (N_8898,N_8154,N_8088);
xnor U8899 (N_8899,N_8008,N_8334);
and U8900 (N_8900,N_8115,N_8158);
or U8901 (N_8901,N_8224,N_8450);
and U8902 (N_8902,N_8436,N_8307);
and U8903 (N_8903,N_8025,N_8135);
xor U8904 (N_8904,N_8015,N_8150);
xor U8905 (N_8905,N_8189,N_8345);
nor U8906 (N_8906,N_8455,N_8382);
nor U8907 (N_8907,N_8492,N_8272);
nor U8908 (N_8908,N_8135,N_8346);
nor U8909 (N_8909,N_8138,N_8352);
and U8910 (N_8910,N_8267,N_8381);
nor U8911 (N_8911,N_8430,N_8306);
nor U8912 (N_8912,N_8286,N_8235);
and U8913 (N_8913,N_8090,N_8102);
and U8914 (N_8914,N_8050,N_8296);
xor U8915 (N_8915,N_8281,N_8447);
nand U8916 (N_8916,N_8412,N_8398);
nor U8917 (N_8917,N_8432,N_8343);
and U8918 (N_8918,N_8483,N_8372);
nand U8919 (N_8919,N_8094,N_8231);
or U8920 (N_8920,N_8093,N_8146);
or U8921 (N_8921,N_8071,N_8039);
or U8922 (N_8922,N_8330,N_8309);
nand U8923 (N_8923,N_8363,N_8312);
or U8924 (N_8924,N_8168,N_8465);
and U8925 (N_8925,N_8081,N_8411);
or U8926 (N_8926,N_8170,N_8419);
xor U8927 (N_8927,N_8269,N_8456);
or U8928 (N_8928,N_8272,N_8213);
or U8929 (N_8929,N_8190,N_8011);
or U8930 (N_8930,N_8215,N_8058);
nand U8931 (N_8931,N_8157,N_8385);
or U8932 (N_8932,N_8369,N_8321);
nor U8933 (N_8933,N_8488,N_8350);
nor U8934 (N_8934,N_8112,N_8494);
and U8935 (N_8935,N_8073,N_8332);
or U8936 (N_8936,N_8375,N_8089);
nand U8937 (N_8937,N_8174,N_8015);
nor U8938 (N_8938,N_8191,N_8010);
and U8939 (N_8939,N_8469,N_8128);
or U8940 (N_8940,N_8390,N_8309);
nand U8941 (N_8941,N_8478,N_8058);
xor U8942 (N_8942,N_8142,N_8153);
nor U8943 (N_8943,N_8351,N_8319);
xor U8944 (N_8944,N_8326,N_8194);
xor U8945 (N_8945,N_8248,N_8237);
nand U8946 (N_8946,N_8418,N_8278);
xor U8947 (N_8947,N_8144,N_8386);
or U8948 (N_8948,N_8308,N_8070);
nand U8949 (N_8949,N_8179,N_8436);
or U8950 (N_8950,N_8208,N_8289);
or U8951 (N_8951,N_8202,N_8012);
or U8952 (N_8952,N_8390,N_8360);
xor U8953 (N_8953,N_8194,N_8209);
xnor U8954 (N_8954,N_8432,N_8239);
and U8955 (N_8955,N_8328,N_8390);
nand U8956 (N_8956,N_8231,N_8035);
or U8957 (N_8957,N_8034,N_8051);
nand U8958 (N_8958,N_8377,N_8029);
and U8959 (N_8959,N_8173,N_8334);
and U8960 (N_8960,N_8185,N_8156);
and U8961 (N_8961,N_8386,N_8139);
and U8962 (N_8962,N_8417,N_8143);
nand U8963 (N_8963,N_8482,N_8096);
nor U8964 (N_8964,N_8357,N_8143);
or U8965 (N_8965,N_8046,N_8026);
and U8966 (N_8966,N_8244,N_8387);
nand U8967 (N_8967,N_8215,N_8027);
or U8968 (N_8968,N_8432,N_8458);
and U8969 (N_8969,N_8481,N_8483);
or U8970 (N_8970,N_8454,N_8219);
and U8971 (N_8971,N_8066,N_8051);
xnor U8972 (N_8972,N_8130,N_8306);
nor U8973 (N_8973,N_8062,N_8154);
or U8974 (N_8974,N_8253,N_8147);
and U8975 (N_8975,N_8063,N_8065);
nor U8976 (N_8976,N_8454,N_8003);
nor U8977 (N_8977,N_8291,N_8011);
and U8978 (N_8978,N_8062,N_8147);
nand U8979 (N_8979,N_8457,N_8485);
xor U8980 (N_8980,N_8075,N_8000);
or U8981 (N_8981,N_8038,N_8248);
or U8982 (N_8982,N_8120,N_8221);
and U8983 (N_8983,N_8406,N_8327);
nor U8984 (N_8984,N_8357,N_8285);
nor U8985 (N_8985,N_8462,N_8398);
nand U8986 (N_8986,N_8078,N_8387);
nor U8987 (N_8987,N_8298,N_8109);
or U8988 (N_8988,N_8288,N_8286);
xor U8989 (N_8989,N_8130,N_8243);
or U8990 (N_8990,N_8178,N_8374);
nand U8991 (N_8991,N_8164,N_8237);
xnor U8992 (N_8992,N_8065,N_8228);
xnor U8993 (N_8993,N_8032,N_8414);
and U8994 (N_8994,N_8304,N_8038);
nand U8995 (N_8995,N_8404,N_8040);
nand U8996 (N_8996,N_8098,N_8082);
nand U8997 (N_8997,N_8458,N_8496);
and U8998 (N_8998,N_8177,N_8077);
nand U8999 (N_8999,N_8167,N_8162);
nand U9000 (N_9000,N_8763,N_8503);
nand U9001 (N_9001,N_8741,N_8862);
nor U9002 (N_9002,N_8795,N_8976);
nand U9003 (N_9003,N_8875,N_8788);
xor U9004 (N_9004,N_8529,N_8905);
and U9005 (N_9005,N_8807,N_8874);
xnor U9006 (N_9006,N_8513,N_8797);
xor U9007 (N_9007,N_8951,N_8628);
nor U9008 (N_9008,N_8592,N_8991);
and U9009 (N_9009,N_8667,N_8773);
or U9010 (N_9010,N_8534,N_8754);
and U9011 (N_9011,N_8963,N_8656);
nor U9012 (N_9012,N_8954,N_8502);
xnor U9013 (N_9013,N_8708,N_8728);
and U9014 (N_9014,N_8915,N_8775);
nor U9015 (N_9015,N_8657,N_8641);
and U9016 (N_9016,N_8898,N_8742);
nor U9017 (N_9017,N_8556,N_8910);
and U9018 (N_9018,N_8601,N_8853);
or U9019 (N_9019,N_8899,N_8683);
xor U9020 (N_9020,N_8958,N_8509);
xor U9021 (N_9021,N_8888,N_8572);
or U9022 (N_9022,N_8518,N_8539);
nand U9023 (N_9023,N_8867,N_8917);
or U9024 (N_9024,N_8645,N_8765);
nand U9025 (N_9025,N_8597,N_8883);
nor U9026 (N_9026,N_8916,N_8887);
nand U9027 (N_9027,N_8663,N_8685);
nor U9028 (N_9028,N_8660,N_8880);
nor U9029 (N_9029,N_8543,N_8726);
or U9030 (N_9030,N_8909,N_8922);
and U9031 (N_9031,N_8893,N_8623);
or U9032 (N_9032,N_8671,N_8712);
nor U9033 (N_9033,N_8749,N_8508);
nand U9034 (N_9034,N_8659,N_8897);
nor U9035 (N_9035,N_8527,N_8674);
or U9036 (N_9036,N_8582,N_8658);
nand U9037 (N_9037,N_8619,N_8557);
or U9038 (N_9038,N_8966,N_8849);
and U9039 (N_9039,N_8739,N_8998);
xnor U9040 (N_9040,N_8974,N_8566);
or U9041 (N_9041,N_8877,N_8759);
xnor U9042 (N_9042,N_8673,N_8666);
nand U9043 (N_9043,N_8921,N_8819);
xnor U9044 (N_9044,N_8675,N_8850);
and U9045 (N_9045,N_8724,N_8770);
and U9046 (N_9046,N_8780,N_8719);
xor U9047 (N_9047,N_8734,N_8787);
or U9048 (N_9048,N_8711,N_8945);
or U9049 (N_9049,N_8885,N_8882);
xor U9050 (N_9050,N_8886,N_8701);
xor U9051 (N_9051,N_8953,N_8935);
nand U9052 (N_9052,N_8532,N_8722);
and U9053 (N_9053,N_8737,N_8638);
or U9054 (N_9054,N_8784,N_8962);
nor U9055 (N_9055,N_8696,N_8687);
and U9056 (N_9056,N_8812,N_8650);
nor U9057 (N_9057,N_8591,N_8738);
or U9058 (N_9058,N_8919,N_8594);
or U9059 (N_9059,N_8692,N_8871);
nor U9060 (N_9060,N_8567,N_8858);
or U9061 (N_9061,N_8570,N_8861);
xor U9062 (N_9062,N_8914,N_8528);
and U9063 (N_9063,N_8767,N_8830);
nand U9064 (N_9064,N_8635,N_8575);
nand U9065 (N_9065,N_8583,N_8776);
and U9066 (N_9066,N_8578,N_8747);
and U9067 (N_9067,N_8985,N_8670);
and U9068 (N_9068,N_8891,N_8744);
and U9069 (N_9069,N_8693,N_8806);
and U9070 (N_9070,N_8637,N_8978);
nor U9071 (N_9071,N_8878,N_8705);
nor U9072 (N_9072,N_8699,N_8992);
nor U9073 (N_9073,N_8824,N_8586);
nand U9074 (N_9074,N_8766,N_8855);
or U9075 (N_9075,N_8621,N_8960);
or U9076 (N_9076,N_8729,N_8961);
nand U9077 (N_9077,N_8537,N_8545);
xnor U9078 (N_9078,N_8554,N_8504);
or U9079 (N_9079,N_8973,N_8615);
or U9080 (N_9080,N_8808,N_8600);
nor U9081 (N_9081,N_8533,N_8948);
xnor U9082 (N_9082,N_8792,N_8733);
xor U9083 (N_9083,N_8515,N_8967);
or U9084 (N_9084,N_8550,N_8941);
or U9085 (N_9085,N_8752,N_8818);
or U9086 (N_9086,N_8936,N_8987);
and U9087 (N_9087,N_8950,N_8559);
xnor U9088 (N_9088,N_8651,N_8803);
nand U9089 (N_9089,N_8714,N_8549);
nor U9090 (N_9090,N_8565,N_8720);
and U9091 (N_9091,N_8715,N_8736);
and U9092 (N_9092,N_8571,N_8869);
and U9093 (N_9093,N_8872,N_8965);
xnor U9094 (N_9094,N_8901,N_8932);
nor U9095 (N_9095,N_8852,N_8541);
xor U9096 (N_9096,N_8655,N_8895);
nor U9097 (N_9097,N_8717,N_8639);
nor U9098 (N_9098,N_8847,N_8611);
or U9099 (N_9099,N_8581,N_8688);
and U9100 (N_9100,N_8923,N_8800);
nand U9101 (N_9101,N_8512,N_8546);
or U9102 (N_9102,N_8760,N_8881);
nand U9103 (N_9103,N_8672,N_8616);
nor U9104 (N_9104,N_8979,N_8906);
xor U9105 (N_9105,N_8758,N_8939);
or U9106 (N_9106,N_8801,N_8614);
nand U9107 (N_9107,N_8704,N_8894);
xor U9108 (N_9108,N_8682,N_8779);
nor U9109 (N_9109,N_8725,N_8603);
nand U9110 (N_9110,N_8842,N_8802);
xnor U9111 (N_9111,N_8525,N_8661);
nand U9112 (N_9112,N_8892,N_8913);
or U9113 (N_9113,N_8846,N_8964);
nand U9114 (N_9114,N_8769,N_8561);
xor U9115 (N_9115,N_8632,N_8563);
or U9116 (N_9116,N_8646,N_8956);
nand U9117 (N_9117,N_8507,N_8520);
nor U9118 (N_9118,N_8957,N_8553);
or U9119 (N_9119,N_8721,N_8938);
xor U9120 (N_9120,N_8709,N_8774);
or U9121 (N_9121,N_8903,N_8786);
nor U9122 (N_9122,N_8564,N_8918);
or U9123 (N_9123,N_8573,N_8716);
xnor U9124 (N_9124,N_8924,N_8618);
xnor U9125 (N_9125,N_8653,N_8771);
nand U9126 (N_9126,N_8805,N_8691);
nand U9127 (N_9127,N_8835,N_8876);
nand U9128 (N_9128,N_8735,N_8652);
xnor U9129 (N_9129,N_8607,N_8562);
nor U9130 (N_9130,N_8997,N_8799);
nand U9131 (N_9131,N_8633,N_8505);
nand U9132 (N_9132,N_8702,N_8538);
nand U9133 (N_9133,N_8530,N_8925);
nor U9134 (N_9134,N_8926,N_8829);
nand U9135 (N_9135,N_8866,N_8501);
or U9136 (N_9136,N_8968,N_8755);
xnor U9137 (N_9137,N_8552,N_8854);
and U9138 (N_9138,N_8548,N_8605);
and U9139 (N_9139,N_8856,N_8713);
xnor U9140 (N_9140,N_8523,N_8514);
and U9141 (N_9141,N_8510,N_8524);
xor U9142 (N_9142,N_8697,N_8971);
nor U9143 (N_9143,N_8535,N_8983);
and U9144 (N_9144,N_8608,N_8560);
nor U9145 (N_9145,N_8588,N_8506);
nand U9146 (N_9146,N_8790,N_8904);
and U9147 (N_9147,N_8831,N_8860);
xnor U9148 (N_9148,N_8540,N_8838);
nand U9149 (N_9149,N_8868,N_8815);
and U9150 (N_9150,N_8519,N_8547);
or U9151 (N_9151,N_8890,N_8680);
xnor U9152 (N_9152,N_8946,N_8631);
xnor U9153 (N_9153,N_8940,N_8927);
or U9154 (N_9154,N_8865,N_8828);
xor U9155 (N_9155,N_8522,N_8649);
or U9156 (N_9156,N_8994,N_8959);
nand U9157 (N_9157,N_8606,N_8643);
nand U9158 (N_9158,N_8988,N_8848);
nor U9159 (N_9159,N_8664,N_8751);
nand U9160 (N_9160,N_8700,N_8827);
or U9161 (N_9161,N_8937,N_8589);
nor U9162 (N_9162,N_8745,N_8912);
xnor U9163 (N_9163,N_8996,N_8746);
or U9164 (N_9164,N_8781,N_8764);
nand U9165 (N_9165,N_8679,N_8977);
nor U9166 (N_9166,N_8689,N_8636);
xnor U9167 (N_9167,N_8995,N_8845);
and U9168 (N_9168,N_8896,N_8975);
nor U9169 (N_9169,N_8678,N_8785);
nand U9170 (N_9170,N_8943,N_8617);
nor U9171 (N_9171,N_8814,N_8695);
nand U9172 (N_9172,N_8604,N_8822);
nor U9173 (N_9173,N_8694,N_8836);
nand U9174 (N_9174,N_8947,N_8841);
nor U9175 (N_9175,N_8902,N_8718);
nor U9176 (N_9176,N_8710,N_8609);
and U9177 (N_9177,N_8930,N_8782);
or U9178 (N_9178,N_8762,N_8928);
nand U9179 (N_9179,N_8640,N_8684);
nand U9180 (N_9180,N_8654,N_8511);
xnor U9181 (N_9181,N_8984,N_8598);
or U9182 (N_9182,N_8864,N_8612);
and U9183 (N_9183,N_8844,N_8516);
or U9184 (N_9184,N_8740,N_8642);
and U9185 (N_9185,N_8840,N_8627);
nor U9186 (N_9186,N_8839,N_8952);
or U9187 (N_9187,N_8676,N_8870);
and U9188 (N_9188,N_8630,N_8778);
nor U9189 (N_9189,N_8796,N_8825);
xor U9190 (N_9190,N_8837,N_8521);
nand U9191 (N_9191,N_8593,N_8703);
or U9192 (N_9192,N_8727,N_8863);
nand U9193 (N_9193,N_8873,N_8933);
and U9194 (N_9194,N_8982,N_8558);
nand U9195 (N_9195,N_8580,N_8669);
nor U9196 (N_9196,N_8889,N_8622);
xor U9197 (N_9197,N_8686,N_8804);
nand U9198 (N_9198,N_8732,N_8730);
and U9199 (N_9199,N_8857,N_8579);
nor U9200 (N_9200,N_8810,N_8798);
nand U9201 (N_9201,N_8596,N_8753);
nor U9202 (N_9202,N_8625,N_8821);
and U9203 (N_9203,N_8681,N_8662);
nor U9204 (N_9204,N_8544,N_8907);
xor U9205 (N_9205,N_8900,N_8620);
xor U9206 (N_9206,N_8942,N_8536);
xor U9207 (N_9207,N_8599,N_8574);
nand U9208 (N_9208,N_8879,N_8809);
and U9209 (N_9209,N_8613,N_8944);
nor U9210 (N_9210,N_8955,N_8706);
nor U9211 (N_9211,N_8595,N_8833);
nand U9212 (N_9212,N_8629,N_8668);
and U9213 (N_9213,N_8634,N_8690);
nor U9214 (N_9214,N_8777,N_8990);
and U9215 (N_9215,N_8851,N_8931);
nand U9216 (N_9216,N_8587,N_8970);
or U9217 (N_9217,N_8789,N_8731);
or U9218 (N_9218,N_8748,N_8626);
and U9219 (N_9219,N_8568,N_8794);
and U9220 (N_9220,N_8743,N_8884);
xnor U9221 (N_9221,N_8817,N_8911);
xnor U9222 (N_9222,N_8768,N_8981);
and U9223 (N_9223,N_8989,N_8793);
nor U9224 (N_9224,N_8757,N_8761);
or U9225 (N_9225,N_8908,N_8624);
and U9226 (N_9226,N_8677,N_8813);
and U9227 (N_9227,N_8972,N_8823);
nor U9228 (N_9228,N_8500,N_8920);
or U9229 (N_9229,N_8811,N_8555);
nor U9230 (N_9230,N_8569,N_8834);
nand U9231 (N_9231,N_8644,N_8816);
nor U9232 (N_9232,N_8517,N_8602);
or U9233 (N_9233,N_8610,N_8542);
xnor U9234 (N_9234,N_8999,N_8707);
nor U9235 (N_9235,N_8783,N_8929);
nor U9236 (N_9236,N_8577,N_8820);
or U9237 (N_9237,N_8750,N_8969);
and U9238 (N_9238,N_8647,N_8590);
or U9239 (N_9239,N_8791,N_8980);
nand U9240 (N_9240,N_8648,N_8859);
or U9241 (N_9241,N_8526,N_8934);
nor U9242 (N_9242,N_8665,N_8698);
nand U9243 (N_9243,N_8585,N_8843);
nor U9244 (N_9244,N_8531,N_8551);
nor U9245 (N_9245,N_8756,N_8993);
nand U9246 (N_9246,N_8949,N_8826);
nand U9247 (N_9247,N_8772,N_8584);
xnor U9248 (N_9248,N_8576,N_8986);
xnor U9249 (N_9249,N_8723,N_8832);
nor U9250 (N_9250,N_8808,N_8873);
and U9251 (N_9251,N_8908,N_8736);
xnor U9252 (N_9252,N_8938,N_8878);
and U9253 (N_9253,N_8741,N_8984);
nand U9254 (N_9254,N_8999,N_8895);
and U9255 (N_9255,N_8589,N_8676);
nand U9256 (N_9256,N_8859,N_8658);
nand U9257 (N_9257,N_8706,N_8841);
and U9258 (N_9258,N_8820,N_8903);
or U9259 (N_9259,N_8904,N_8940);
xor U9260 (N_9260,N_8988,N_8606);
or U9261 (N_9261,N_8636,N_8966);
or U9262 (N_9262,N_8742,N_8970);
xor U9263 (N_9263,N_8508,N_8563);
nor U9264 (N_9264,N_8509,N_8548);
nor U9265 (N_9265,N_8757,N_8970);
nand U9266 (N_9266,N_8569,N_8904);
and U9267 (N_9267,N_8623,N_8833);
and U9268 (N_9268,N_8609,N_8706);
or U9269 (N_9269,N_8628,N_8502);
or U9270 (N_9270,N_8599,N_8668);
xor U9271 (N_9271,N_8733,N_8619);
and U9272 (N_9272,N_8680,N_8630);
nand U9273 (N_9273,N_8538,N_8644);
nor U9274 (N_9274,N_8893,N_8573);
xor U9275 (N_9275,N_8708,N_8859);
nor U9276 (N_9276,N_8739,N_8696);
nand U9277 (N_9277,N_8993,N_8815);
or U9278 (N_9278,N_8508,N_8556);
nand U9279 (N_9279,N_8920,N_8696);
nor U9280 (N_9280,N_8654,N_8515);
or U9281 (N_9281,N_8679,N_8786);
and U9282 (N_9282,N_8809,N_8793);
xor U9283 (N_9283,N_8883,N_8914);
xor U9284 (N_9284,N_8762,N_8820);
nand U9285 (N_9285,N_8510,N_8867);
and U9286 (N_9286,N_8673,N_8914);
nor U9287 (N_9287,N_8605,N_8907);
or U9288 (N_9288,N_8852,N_8768);
or U9289 (N_9289,N_8765,N_8826);
nor U9290 (N_9290,N_8529,N_8609);
nor U9291 (N_9291,N_8936,N_8648);
nand U9292 (N_9292,N_8635,N_8972);
and U9293 (N_9293,N_8609,N_8912);
nor U9294 (N_9294,N_8913,N_8881);
xnor U9295 (N_9295,N_8683,N_8603);
and U9296 (N_9296,N_8974,N_8891);
or U9297 (N_9297,N_8967,N_8531);
xor U9298 (N_9298,N_8943,N_8801);
or U9299 (N_9299,N_8621,N_8788);
xor U9300 (N_9300,N_8945,N_8768);
nor U9301 (N_9301,N_8597,N_8894);
nand U9302 (N_9302,N_8659,N_8770);
nor U9303 (N_9303,N_8619,N_8504);
or U9304 (N_9304,N_8580,N_8874);
xor U9305 (N_9305,N_8918,N_8879);
or U9306 (N_9306,N_8760,N_8866);
or U9307 (N_9307,N_8598,N_8842);
nor U9308 (N_9308,N_8560,N_8701);
and U9309 (N_9309,N_8846,N_8628);
xnor U9310 (N_9310,N_8552,N_8616);
and U9311 (N_9311,N_8765,N_8737);
nand U9312 (N_9312,N_8767,N_8678);
xor U9313 (N_9313,N_8980,N_8671);
or U9314 (N_9314,N_8896,N_8787);
xnor U9315 (N_9315,N_8526,N_8779);
and U9316 (N_9316,N_8626,N_8983);
or U9317 (N_9317,N_8949,N_8918);
nor U9318 (N_9318,N_8779,N_8825);
xnor U9319 (N_9319,N_8581,N_8873);
xnor U9320 (N_9320,N_8967,N_8891);
xor U9321 (N_9321,N_8960,N_8643);
nor U9322 (N_9322,N_8999,N_8923);
nor U9323 (N_9323,N_8921,N_8824);
nor U9324 (N_9324,N_8604,N_8830);
nand U9325 (N_9325,N_8807,N_8804);
and U9326 (N_9326,N_8721,N_8814);
xor U9327 (N_9327,N_8764,N_8699);
nor U9328 (N_9328,N_8743,N_8534);
nand U9329 (N_9329,N_8622,N_8550);
or U9330 (N_9330,N_8679,N_8546);
xor U9331 (N_9331,N_8759,N_8937);
or U9332 (N_9332,N_8955,N_8843);
xor U9333 (N_9333,N_8605,N_8736);
nand U9334 (N_9334,N_8764,N_8675);
nor U9335 (N_9335,N_8817,N_8756);
and U9336 (N_9336,N_8657,N_8723);
and U9337 (N_9337,N_8832,N_8791);
or U9338 (N_9338,N_8717,N_8933);
xnor U9339 (N_9339,N_8584,N_8826);
nor U9340 (N_9340,N_8795,N_8737);
xnor U9341 (N_9341,N_8518,N_8981);
nor U9342 (N_9342,N_8693,N_8823);
and U9343 (N_9343,N_8836,N_8751);
xor U9344 (N_9344,N_8537,N_8811);
or U9345 (N_9345,N_8890,N_8925);
nand U9346 (N_9346,N_8929,N_8587);
or U9347 (N_9347,N_8722,N_8744);
nor U9348 (N_9348,N_8630,N_8770);
xnor U9349 (N_9349,N_8529,N_8878);
xnor U9350 (N_9350,N_8750,N_8949);
xnor U9351 (N_9351,N_8767,N_8865);
or U9352 (N_9352,N_8753,N_8513);
and U9353 (N_9353,N_8735,N_8657);
nor U9354 (N_9354,N_8740,N_8601);
and U9355 (N_9355,N_8756,N_8546);
xnor U9356 (N_9356,N_8894,N_8857);
and U9357 (N_9357,N_8969,N_8807);
nor U9358 (N_9358,N_8685,N_8720);
nand U9359 (N_9359,N_8601,N_8949);
xor U9360 (N_9360,N_8842,N_8593);
or U9361 (N_9361,N_8801,N_8510);
and U9362 (N_9362,N_8793,N_8762);
nand U9363 (N_9363,N_8881,N_8827);
and U9364 (N_9364,N_8995,N_8675);
nand U9365 (N_9365,N_8730,N_8809);
xnor U9366 (N_9366,N_8836,N_8899);
or U9367 (N_9367,N_8506,N_8743);
nor U9368 (N_9368,N_8732,N_8517);
nand U9369 (N_9369,N_8591,N_8600);
and U9370 (N_9370,N_8547,N_8502);
or U9371 (N_9371,N_8934,N_8720);
and U9372 (N_9372,N_8924,N_8730);
nor U9373 (N_9373,N_8937,N_8564);
and U9374 (N_9374,N_8900,N_8997);
nand U9375 (N_9375,N_8976,N_8652);
and U9376 (N_9376,N_8666,N_8753);
nand U9377 (N_9377,N_8858,N_8551);
nand U9378 (N_9378,N_8913,N_8808);
or U9379 (N_9379,N_8952,N_8744);
nand U9380 (N_9380,N_8582,N_8914);
nor U9381 (N_9381,N_8917,N_8724);
xnor U9382 (N_9382,N_8971,N_8635);
xnor U9383 (N_9383,N_8505,N_8817);
nor U9384 (N_9384,N_8581,N_8547);
and U9385 (N_9385,N_8638,N_8557);
or U9386 (N_9386,N_8506,N_8599);
nor U9387 (N_9387,N_8891,N_8982);
nand U9388 (N_9388,N_8949,N_8705);
nor U9389 (N_9389,N_8540,N_8590);
xor U9390 (N_9390,N_8554,N_8887);
xor U9391 (N_9391,N_8841,N_8951);
and U9392 (N_9392,N_8587,N_8891);
nand U9393 (N_9393,N_8521,N_8655);
xnor U9394 (N_9394,N_8570,N_8738);
xnor U9395 (N_9395,N_8530,N_8912);
nand U9396 (N_9396,N_8766,N_8682);
or U9397 (N_9397,N_8942,N_8512);
and U9398 (N_9398,N_8663,N_8581);
nor U9399 (N_9399,N_8535,N_8659);
xor U9400 (N_9400,N_8873,N_8591);
nor U9401 (N_9401,N_8806,N_8832);
xor U9402 (N_9402,N_8529,N_8781);
or U9403 (N_9403,N_8713,N_8616);
nand U9404 (N_9404,N_8740,N_8770);
nor U9405 (N_9405,N_8504,N_8649);
xnor U9406 (N_9406,N_8546,N_8744);
nor U9407 (N_9407,N_8520,N_8699);
nor U9408 (N_9408,N_8853,N_8703);
nor U9409 (N_9409,N_8908,N_8596);
nor U9410 (N_9410,N_8825,N_8950);
xor U9411 (N_9411,N_8629,N_8503);
or U9412 (N_9412,N_8515,N_8771);
nor U9413 (N_9413,N_8519,N_8528);
or U9414 (N_9414,N_8767,N_8554);
nand U9415 (N_9415,N_8628,N_8877);
or U9416 (N_9416,N_8784,N_8675);
and U9417 (N_9417,N_8677,N_8690);
nor U9418 (N_9418,N_8686,N_8710);
xor U9419 (N_9419,N_8621,N_8860);
nand U9420 (N_9420,N_8585,N_8538);
and U9421 (N_9421,N_8861,N_8781);
nand U9422 (N_9422,N_8976,N_8630);
xnor U9423 (N_9423,N_8981,N_8505);
xnor U9424 (N_9424,N_8566,N_8901);
nand U9425 (N_9425,N_8730,N_8706);
xnor U9426 (N_9426,N_8538,N_8727);
nand U9427 (N_9427,N_8773,N_8967);
nand U9428 (N_9428,N_8943,N_8513);
nor U9429 (N_9429,N_8645,N_8716);
nand U9430 (N_9430,N_8809,N_8980);
xnor U9431 (N_9431,N_8773,N_8606);
xnor U9432 (N_9432,N_8897,N_8611);
nand U9433 (N_9433,N_8923,N_8865);
nand U9434 (N_9434,N_8940,N_8864);
and U9435 (N_9435,N_8740,N_8952);
or U9436 (N_9436,N_8956,N_8850);
nor U9437 (N_9437,N_8935,N_8884);
xor U9438 (N_9438,N_8635,N_8874);
and U9439 (N_9439,N_8574,N_8597);
and U9440 (N_9440,N_8743,N_8725);
nand U9441 (N_9441,N_8960,N_8749);
and U9442 (N_9442,N_8865,N_8994);
nor U9443 (N_9443,N_8598,N_8828);
nand U9444 (N_9444,N_8540,N_8544);
or U9445 (N_9445,N_8874,N_8972);
xnor U9446 (N_9446,N_8859,N_8531);
xor U9447 (N_9447,N_8948,N_8946);
nand U9448 (N_9448,N_8542,N_8521);
xnor U9449 (N_9449,N_8720,N_8543);
or U9450 (N_9450,N_8560,N_8735);
nand U9451 (N_9451,N_8763,N_8790);
xor U9452 (N_9452,N_8737,N_8541);
or U9453 (N_9453,N_8668,N_8681);
nor U9454 (N_9454,N_8752,N_8811);
nand U9455 (N_9455,N_8679,N_8916);
nor U9456 (N_9456,N_8501,N_8721);
and U9457 (N_9457,N_8615,N_8884);
or U9458 (N_9458,N_8506,N_8672);
and U9459 (N_9459,N_8572,N_8609);
nor U9460 (N_9460,N_8778,N_8911);
xor U9461 (N_9461,N_8802,N_8518);
or U9462 (N_9462,N_8751,N_8950);
and U9463 (N_9463,N_8639,N_8550);
nand U9464 (N_9464,N_8764,N_8585);
or U9465 (N_9465,N_8905,N_8897);
nand U9466 (N_9466,N_8933,N_8997);
or U9467 (N_9467,N_8899,N_8594);
and U9468 (N_9468,N_8524,N_8595);
nand U9469 (N_9469,N_8994,N_8580);
nand U9470 (N_9470,N_8913,N_8945);
nor U9471 (N_9471,N_8522,N_8777);
nand U9472 (N_9472,N_8823,N_8759);
nand U9473 (N_9473,N_8671,N_8670);
or U9474 (N_9474,N_8859,N_8500);
nand U9475 (N_9475,N_8823,N_8979);
xnor U9476 (N_9476,N_8973,N_8561);
nand U9477 (N_9477,N_8702,N_8731);
nand U9478 (N_9478,N_8777,N_8789);
and U9479 (N_9479,N_8654,N_8505);
xor U9480 (N_9480,N_8614,N_8635);
nand U9481 (N_9481,N_8954,N_8911);
nor U9482 (N_9482,N_8704,N_8654);
nor U9483 (N_9483,N_8789,N_8995);
nor U9484 (N_9484,N_8908,N_8969);
xnor U9485 (N_9485,N_8626,N_8694);
nor U9486 (N_9486,N_8953,N_8857);
or U9487 (N_9487,N_8532,N_8892);
and U9488 (N_9488,N_8860,N_8791);
or U9489 (N_9489,N_8634,N_8909);
xnor U9490 (N_9490,N_8756,N_8535);
nor U9491 (N_9491,N_8593,N_8600);
nor U9492 (N_9492,N_8530,N_8502);
or U9493 (N_9493,N_8667,N_8559);
nand U9494 (N_9494,N_8503,N_8594);
or U9495 (N_9495,N_8533,N_8811);
nor U9496 (N_9496,N_8682,N_8931);
xor U9497 (N_9497,N_8961,N_8813);
or U9498 (N_9498,N_8686,N_8742);
or U9499 (N_9499,N_8590,N_8644);
nor U9500 (N_9500,N_9438,N_9339);
nand U9501 (N_9501,N_9368,N_9324);
or U9502 (N_9502,N_9065,N_9040);
or U9503 (N_9503,N_9044,N_9402);
nor U9504 (N_9504,N_9170,N_9135);
nand U9505 (N_9505,N_9495,N_9046);
nor U9506 (N_9506,N_9228,N_9022);
and U9507 (N_9507,N_9471,N_9246);
and U9508 (N_9508,N_9155,N_9034);
and U9509 (N_9509,N_9197,N_9395);
and U9510 (N_9510,N_9026,N_9355);
nand U9511 (N_9511,N_9442,N_9434);
nand U9512 (N_9512,N_9115,N_9164);
nand U9513 (N_9513,N_9312,N_9499);
nand U9514 (N_9514,N_9095,N_9107);
nor U9515 (N_9515,N_9353,N_9089);
nand U9516 (N_9516,N_9371,N_9012);
or U9517 (N_9517,N_9243,N_9459);
nor U9518 (N_9518,N_9343,N_9458);
or U9519 (N_9519,N_9340,N_9413);
nand U9520 (N_9520,N_9112,N_9225);
nor U9521 (N_9521,N_9150,N_9049);
or U9522 (N_9522,N_9494,N_9311);
nor U9523 (N_9523,N_9336,N_9364);
nand U9524 (N_9524,N_9420,N_9140);
and U9525 (N_9525,N_9131,N_9293);
xor U9526 (N_9526,N_9329,N_9249);
or U9527 (N_9527,N_9305,N_9271);
or U9528 (N_9528,N_9110,N_9377);
nor U9529 (N_9529,N_9393,N_9153);
nor U9530 (N_9530,N_9488,N_9453);
xor U9531 (N_9531,N_9027,N_9177);
nand U9532 (N_9532,N_9174,N_9361);
xnor U9533 (N_9533,N_9075,N_9380);
and U9534 (N_9534,N_9412,N_9354);
nor U9535 (N_9535,N_9190,N_9073);
and U9536 (N_9536,N_9423,N_9138);
nor U9537 (N_9537,N_9320,N_9024);
xor U9538 (N_9538,N_9121,N_9268);
and U9539 (N_9539,N_9242,N_9461);
nand U9540 (N_9540,N_9373,N_9141);
and U9541 (N_9541,N_9403,N_9345);
xnor U9542 (N_9542,N_9408,N_9326);
nor U9543 (N_9543,N_9222,N_9032);
xnor U9544 (N_9544,N_9008,N_9129);
nand U9545 (N_9545,N_9234,N_9261);
nand U9546 (N_9546,N_9106,N_9422);
nand U9547 (N_9547,N_9194,N_9430);
xor U9548 (N_9548,N_9376,N_9133);
nand U9549 (N_9549,N_9172,N_9160);
or U9550 (N_9550,N_9143,N_9233);
or U9551 (N_9551,N_9030,N_9196);
or U9552 (N_9552,N_9436,N_9229);
nor U9553 (N_9553,N_9010,N_9079);
nand U9554 (N_9554,N_9415,N_9045);
xor U9555 (N_9555,N_9314,N_9016);
and U9556 (N_9556,N_9317,N_9433);
nor U9557 (N_9557,N_9206,N_9451);
nor U9558 (N_9558,N_9241,N_9255);
nand U9559 (N_9559,N_9168,N_9295);
or U9560 (N_9560,N_9029,N_9148);
or U9561 (N_9561,N_9344,N_9021);
or U9562 (N_9562,N_9178,N_9257);
and U9563 (N_9563,N_9286,N_9464);
and U9564 (N_9564,N_9439,N_9493);
nor U9565 (N_9565,N_9267,N_9357);
nand U9566 (N_9566,N_9417,N_9158);
nor U9567 (N_9567,N_9485,N_9446);
or U9568 (N_9568,N_9122,N_9309);
or U9569 (N_9569,N_9479,N_9210);
or U9570 (N_9570,N_9327,N_9483);
or U9571 (N_9571,N_9189,N_9192);
xor U9572 (N_9572,N_9104,N_9059);
and U9573 (N_9573,N_9039,N_9342);
nand U9574 (N_9574,N_9328,N_9139);
and U9575 (N_9575,N_9318,N_9467);
and U9576 (N_9576,N_9202,N_9244);
or U9577 (N_9577,N_9369,N_9020);
or U9578 (N_9578,N_9088,N_9404);
xnor U9579 (N_9579,N_9047,N_9247);
or U9580 (N_9580,N_9449,N_9332);
nand U9581 (N_9581,N_9183,N_9350);
xnor U9582 (N_9582,N_9260,N_9279);
and U9583 (N_9583,N_9273,N_9308);
xnor U9584 (N_9584,N_9048,N_9252);
nand U9585 (N_9585,N_9217,N_9060);
nor U9586 (N_9586,N_9452,N_9013);
nand U9587 (N_9587,N_9203,N_9391);
nand U9588 (N_9588,N_9208,N_9390);
and U9589 (N_9589,N_9227,N_9297);
nor U9590 (N_9590,N_9066,N_9477);
or U9591 (N_9591,N_9341,N_9062);
xnor U9592 (N_9592,N_9410,N_9482);
nor U9593 (N_9593,N_9173,N_9416);
nand U9594 (N_9594,N_9157,N_9383);
and U9595 (N_9595,N_9057,N_9082);
or U9596 (N_9596,N_9292,N_9090);
or U9597 (N_9597,N_9447,N_9084);
and U9598 (N_9598,N_9374,N_9251);
nor U9599 (N_9599,N_9041,N_9035);
nand U9600 (N_9600,N_9205,N_9238);
nand U9601 (N_9601,N_9180,N_9386);
nand U9602 (N_9602,N_9108,N_9322);
xnor U9603 (N_9603,N_9262,N_9366);
nand U9604 (N_9604,N_9136,N_9080);
nor U9605 (N_9605,N_9018,N_9419);
xor U9606 (N_9606,N_9333,N_9359);
or U9607 (N_9607,N_9248,N_9487);
and U9608 (N_9608,N_9071,N_9437);
xor U9609 (N_9609,N_9389,N_9282);
nor U9610 (N_9610,N_9443,N_9492);
xor U9611 (N_9611,N_9280,N_9193);
nor U9612 (N_9612,N_9315,N_9111);
xnor U9613 (N_9613,N_9382,N_9239);
nand U9614 (N_9614,N_9074,N_9414);
nor U9615 (N_9615,N_9278,N_9171);
or U9616 (N_9616,N_9213,N_9220);
and U9617 (N_9617,N_9457,N_9067);
nand U9618 (N_9618,N_9161,N_9052);
nand U9619 (N_9619,N_9085,N_9011);
nor U9620 (N_9620,N_9211,N_9226);
and U9621 (N_9621,N_9159,N_9272);
and U9622 (N_9622,N_9000,N_9236);
nand U9623 (N_9623,N_9288,N_9137);
or U9624 (N_9624,N_9102,N_9269);
or U9625 (N_9625,N_9421,N_9091);
nor U9626 (N_9626,N_9166,N_9113);
nor U9627 (N_9627,N_9431,N_9496);
and U9628 (N_9628,N_9004,N_9142);
nand U9629 (N_9629,N_9147,N_9425);
and U9630 (N_9630,N_9463,N_9294);
and U9631 (N_9631,N_9209,N_9025);
or U9632 (N_9632,N_9491,N_9188);
xnor U9633 (N_9633,N_9235,N_9219);
nand U9634 (N_9634,N_9385,N_9175);
or U9635 (N_9635,N_9033,N_9154);
nor U9636 (N_9636,N_9145,N_9237);
and U9637 (N_9637,N_9378,N_9116);
xnor U9638 (N_9638,N_9440,N_9043);
nor U9639 (N_9639,N_9017,N_9214);
xnor U9640 (N_9640,N_9289,N_9117);
xor U9641 (N_9641,N_9475,N_9195);
and U9642 (N_9642,N_9253,N_9019);
nor U9643 (N_9643,N_9156,N_9298);
nand U9644 (N_9644,N_9381,N_9375);
nand U9645 (N_9645,N_9128,N_9151);
nor U9646 (N_9646,N_9384,N_9042);
nor U9647 (N_9647,N_9358,N_9306);
xor U9648 (N_9648,N_9006,N_9388);
nand U9649 (N_9649,N_9401,N_9335);
xor U9650 (N_9650,N_9127,N_9152);
and U9651 (N_9651,N_9363,N_9392);
xnor U9652 (N_9652,N_9037,N_9356);
nand U9653 (N_9653,N_9338,N_9299);
nor U9654 (N_9654,N_9283,N_9321);
and U9655 (N_9655,N_9015,N_9093);
xor U9656 (N_9656,N_9334,N_9448);
xnor U9657 (N_9657,N_9184,N_9124);
nand U9658 (N_9658,N_9303,N_9103);
nor U9659 (N_9659,N_9284,N_9435);
nand U9660 (N_9660,N_9456,N_9365);
or U9661 (N_9661,N_9346,N_9096);
xor U9662 (N_9662,N_9497,N_9256);
nor U9663 (N_9663,N_9411,N_9486);
nand U9664 (N_9664,N_9064,N_9187);
nor U9665 (N_9665,N_9360,N_9351);
nor U9666 (N_9666,N_9051,N_9460);
nand U9667 (N_9667,N_9455,N_9405);
and U9668 (N_9668,N_9218,N_9474);
xor U9669 (N_9669,N_9325,N_9407);
nor U9670 (N_9670,N_9428,N_9216);
nor U9671 (N_9671,N_9319,N_9231);
or U9672 (N_9672,N_9167,N_9396);
nor U9673 (N_9673,N_9304,N_9296);
or U9674 (N_9674,N_9441,N_9083);
and U9675 (N_9675,N_9480,N_9086);
or U9676 (N_9676,N_9061,N_9200);
nand U9677 (N_9677,N_9290,N_9254);
xnor U9678 (N_9678,N_9277,N_9427);
nand U9679 (N_9679,N_9069,N_9007);
or U9680 (N_9680,N_9201,N_9215);
nand U9681 (N_9681,N_9031,N_9038);
xnor U9682 (N_9682,N_9444,N_9212);
nand U9683 (N_9683,N_9399,N_9418);
nor U9684 (N_9684,N_9469,N_9109);
and U9685 (N_9685,N_9259,N_9182);
nand U9686 (N_9686,N_9274,N_9094);
nand U9687 (N_9687,N_9023,N_9300);
nand U9688 (N_9688,N_9331,N_9123);
or U9689 (N_9689,N_9165,N_9470);
and U9690 (N_9690,N_9005,N_9367);
xor U9691 (N_9691,N_9379,N_9070);
or U9692 (N_9692,N_9287,N_9149);
xor U9693 (N_9693,N_9001,N_9068);
nor U9694 (N_9694,N_9281,N_9207);
xor U9695 (N_9695,N_9489,N_9264);
xnor U9696 (N_9696,N_9054,N_9498);
and U9697 (N_9697,N_9307,N_9199);
or U9698 (N_9698,N_9092,N_9406);
nand U9699 (N_9699,N_9078,N_9323);
nor U9700 (N_9700,N_9204,N_9330);
or U9701 (N_9701,N_9348,N_9310);
nand U9702 (N_9702,N_9105,N_9424);
nand U9703 (N_9703,N_9191,N_9481);
xnor U9704 (N_9704,N_9473,N_9445);
and U9705 (N_9705,N_9362,N_9432);
xor U9706 (N_9706,N_9014,N_9198);
or U9707 (N_9707,N_9462,N_9466);
or U9708 (N_9708,N_9186,N_9270);
and U9709 (N_9709,N_9099,N_9125);
nand U9710 (N_9710,N_9397,N_9301);
nand U9711 (N_9711,N_9224,N_9370);
nand U9712 (N_9712,N_9050,N_9245);
xnor U9713 (N_9713,N_9176,N_9101);
xor U9714 (N_9714,N_9098,N_9400);
or U9715 (N_9715,N_9429,N_9185);
nor U9716 (N_9716,N_9120,N_9276);
and U9717 (N_9717,N_9053,N_9002);
xnor U9718 (N_9718,N_9003,N_9472);
nor U9719 (N_9719,N_9132,N_9398);
xnor U9720 (N_9720,N_9162,N_9394);
xor U9721 (N_9721,N_9036,N_9221);
xor U9722 (N_9722,N_9258,N_9028);
or U9723 (N_9723,N_9181,N_9114);
or U9724 (N_9724,N_9087,N_9076);
nand U9725 (N_9725,N_9240,N_9266);
nor U9726 (N_9726,N_9163,N_9056);
nor U9727 (N_9727,N_9250,N_9223);
xor U9728 (N_9728,N_9454,N_9372);
nand U9729 (N_9729,N_9265,N_9476);
or U9730 (N_9730,N_9468,N_9426);
xor U9731 (N_9731,N_9349,N_9179);
xnor U9732 (N_9732,N_9490,N_9081);
xnor U9733 (N_9733,N_9063,N_9337);
nor U9734 (N_9734,N_9144,N_9009);
xor U9735 (N_9735,N_9291,N_9232);
nand U9736 (N_9736,N_9275,N_9263);
nand U9737 (N_9737,N_9387,N_9100);
nor U9738 (N_9738,N_9465,N_9134);
and U9739 (N_9739,N_9058,N_9478);
or U9740 (N_9740,N_9072,N_9097);
xor U9741 (N_9741,N_9077,N_9130);
nor U9742 (N_9742,N_9316,N_9126);
xnor U9743 (N_9743,N_9285,N_9169);
nor U9744 (N_9744,N_9313,N_9055);
and U9745 (N_9745,N_9146,N_9230);
nor U9746 (N_9746,N_9118,N_9347);
nor U9747 (N_9747,N_9450,N_9484);
nor U9748 (N_9748,N_9409,N_9302);
xor U9749 (N_9749,N_9119,N_9352);
nand U9750 (N_9750,N_9147,N_9326);
nor U9751 (N_9751,N_9454,N_9386);
xnor U9752 (N_9752,N_9035,N_9257);
and U9753 (N_9753,N_9426,N_9420);
nor U9754 (N_9754,N_9261,N_9411);
and U9755 (N_9755,N_9060,N_9134);
nand U9756 (N_9756,N_9293,N_9063);
nor U9757 (N_9757,N_9488,N_9265);
or U9758 (N_9758,N_9403,N_9233);
and U9759 (N_9759,N_9327,N_9454);
nor U9760 (N_9760,N_9365,N_9016);
and U9761 (N_9761,N_9368,N_9319);
or U9762 (N_9762,N_9405,N_9325);
nand U9763 (N_9763,N_9016,N_9499);
xor U9764 (N_9764,N_9381,N_9287);
or U9765 (N_9765,N_9206,N_9367);
and U9766 (N_9766,N_9395,N_9034);
nand U9767 (N_9767,N_9129,N_9130);
nor U9768 (N_9768,N_9297,N_9353);
and U9769 (N_9769,N_9455,N_9102);
and U9770 (N_9770,N_9184,N_9222);
nand U9771 (N_9771,N_9120,N_9149);
or U9772 (N_9772,N_9340,N_9462);
or U9773 (N_9773,N_9391,N_9171);
or U9774 (N_9774,N_9359,N_9020);
nand U9775 (N_9775,N_9472,N_9301);
and U9776 (N_9776,N_9122,N_9130);
or U9777 (N_9777,N_9125,N_9084);
xor U9778 (N_9778,N_9435,N_9469);
and U9779 (N_9779,N_9452,N_9471);
xnor U9780 (N_9780,N_9031,N_9166);
nand U9781 (N_9781,N_9365,N_9092);
nand U9782 (N_9782,N_9131,N_9165);
or U9783 (N_9783,N_9389,N_9065);
or U9784 (N_9784,N_9110,N_9458);
and U9785 (N_9785,N_9061,N_9299);
or U9786 (N_9786,N_9296,N_9113);
xnor U9787 (N_9787,N_9309,N_9135);
and U9788 (N_9788,N_9243,N_9058);
nor U9789 (N_9789,N_9394,N_9241);
nor U9790 (N_9790,N_9442,N_9405);
and U9791 (N_9791,N_9237,N_9239);
nand U9792 (N_9792,N_9243,N_9423);
xnor U9793 (N_9793,N_9273,N_9401);
nand U9794 (N_9794,N_9350,N_9080);
and U9795 (N_9795,N_9156,N_9052);
xnor U9796 (N_9796,N_9064,N_9389);
nor U9797 (N_9797,N_9412,N_9190);
xnor U9798 (N_9798,N_9488,N_9284);
nor U9799 (N_9799,N_9352,N_9221);
or U9800 (N_9800,N_9117,N_9276);
and U9801 (N_9801,N_9393,N_9200);
xnor U9802 (N_9802,N_9282,N_9459);
and U9803 (N_9803,N_9250,N_9327);
nand U9804 (N_9804,N_9251,N_9350);
nor U9805 (N_9805,N_9470,N_9298);
xnor U9806 (N_9806,N_9442,N_9335);
or U9807 (N_9807,N_9406,N_9187);
nand U9808 (N_9808,N_9043,N_9143);
nand U9809 (N_9809,N_9369,N_9470);
or U9810 (N_9810,N_9359,N_9326);
nand U9811 (N_9811,N_9356,N_9253);
or U9812 (N_9812,N_9315,N_9238);
nor U9813 (N_9813,N_9219,N_9182);
or U9814 (N_9814,N_9059,N_9249);
or U9815 (N_9815,N_9486,N_9063);
nor U9816 (N_9816,N_9296,N_9074);
nand U9817 (N_9817,N_9437,N_9166);
xnor U9818 (N_9818,N_9028,N_9422);
nand U9819 (N_9819,N_9178,N_9478);
xor U9820 (N_9820,N_9299,N_9170);
nand U9821 (N_9821,N_9087,N_9095);
nand U9822 (N_9822,N_9224,N_9344);
or U9823 (N_9823,N_9354,N_9443);
or U9824 (N_9824,N_9485,N_9498);
nand U9825 (N_9825,N_9014,N_9395);
nand U9826 (N_9826,N_9492,N_9346);
or U9827 (N_9827,N_9397,N_9195);
and U9828 (N_9828,N_9098,N_9041);
or U9829 (N_9829,N_9129,N_9065);
or U9830 (N_9830,N_9359,N_9142);
nor U9831 (N_9831,N_9309,N_9216);
and U9832 (N_9832,N_9090,N_9143);
and U9833 (N_9833,N_9099,N_9451);
nor U9834 (N_9834,N_9310,N_9288);
and U9835 (N_9835,N_9136,N_9211);
nand U9836 (N_9836,N_9321,N_9049);
nand U9837 (N_9837,N_9033,N_9015);
and U9838 (N_9838,N_9222,N_9131);
xor U9839 (N_9839,N_9033,N_9262);
xnor U9840 (N_9840,N_9031,N_9451);
xor U9841 (N_9841,N_9428,N_9246);
or U9842 (N_9842,N_9195,N_9108);
nand U9843 (N_9843,N_9457,N_9432);
nand U9844 (N_9844,N_9260,N_9015);
nand U9845 (N_9845,N_9072,N_9215);
nor U9846 (N_9846,N_9129,N_9051);
or U9847 (N_9847,N_9312,N_9009);
nor U9848 (N_9848,N_9268,N_9464);
or U9849 (N_9849,N_9153,N_9180);
xor U9850 (N_9850,N_9411,N_9355);
nor U9851 (N_9851,N_9196,N_9104);
xor U9852 (N_9852,N_9074,N_9272);
xnor U9853 (N_9853,N_9054,N_9220);
nand U9854 (N_9854,N_9364,N_9211);
nor U9855 (N_9855,N_9318,N_9347);
nor U9856 (N_9856,N_9499,N_9143);
or U9857 (N_9857,N_9184,N_9329);
and U9858 (N_9858,N_9392,N_9426);
or U9859 (N_9859,N_9091,N_9209);
xor U9860 (N_9860,N_9053,N_9191);
xor U9861 (N_9861,N_9177,N_9072);
nor U9862 (N_9862,N_9174,N_9408);
xnor U9863 (N_9863,N_9191,N_9258);
and U9864 (N_9864,N_9101,N_9497);
nand U9865 (N_9865,N_9250,N_9020);
nor U9866 (N_9866,N_9027,N_9028);
or U9867 (N_9867,N_9060,N_9087);
nor U9868 (N_9868,N_9240,N_9188);
and U9869 (N_9869,N_9085,N_9082);
xor U9870 (N_9870,N_9140,N_9410);
xnor U9871 (N_9871,N_9224,N_9055);
nand U9872 (N_9872,N_9461,N_9287);
nand U9873 (N_9873,N_9127,N_9488);
xor U9874 (N_9874,N_9434,N_9146);
or U9875 (N_9875,N_9100,N_9242);
nand U9876 (N_9876,N_9241,N_9485);
and U9877 (N_9877,N_9398,N_9386);
xor U9878 (N_9878,N_9459,N_9359);
and U9879 (N_9879,N_9027,N_9130);
nand U9880 (N_9880,N_9003,N_9411);
xnor U9881 (N_9881,N_9321,N_9063);
xnor U9882 (N_9882,N_9275,N_9233);
and U9883 (N_9883,N_9482,N_9459);
and U9884 (N_9884,N_9040,N_9359);
or U9885 (N_9885,N_9034,N_9013);
xnor U9886 (N_9886,N_9412,N_9052);
xor U9887 (N_9887,N_9041,N_9205);
or U9888 (N_9888,N_9494,N_9254);
nand U9889 (N_9889,N_9073,N_9334);
nor U9890 (N_9890,N_9388,N_9311);
nor U9891 (N_9891,N_9094,N_9246);
or U9892 (N_9892,N_9485,N_9279);
and U9893 (N_9893,N_9169,N_9437);
nand U9894 (N_9894,N_9084,N_9296);
and U9895 (N_9895,N_9116,N_9381);
or U9896 (N_9896,N_9127,N_9068);
nor U9897 (N_9897,N_9490,N_9038);
and U9898 (N_9898,N_9453,N_9298);
or U9899 (N_9899,N_9139,N_9179);
and U9900 (N_9900,N_9368,N_9278);
nand U9901 (N_9901,N_9210,N_9430);
or U9902 (N_9902,N_9221,N_9313);
xor U9903 (N_9903,N_9296,N_9372);
and U9904 (N_9904,N_9247,N_9447);
xor U9905 (N_9905,N_9239,N_9492);
or U9906 (N_9906,N_9325,N_9174);
xnor U9907 (N_9907,N_9068,N_9165);
xnor U9908 (N_9908,N_9202,N_9133);
and U9909 (N_9909,N_9378,N_9357);
xor U9910 (N_9910,N_9093,N_9483);
nand U9911 (N_9911,N_9175,N_9389);
nor U9912 (N_9912,N_9459,N_9206);
nor U9913 (N_9913,N_9254,N_9273);
or U9914 (N_9914,N_9114,N_9284);
nand U9915 (N_9915,N_9196,N_9164);
xor U9916 (N_9916,N_9416,N_9482);
nand U9917 (N_9917,N_9174,N_9001);
xnor U9918 (N_9918,N_9263,N_9123);
and U9919 (N_9919,N_9068,N_9016);
or U9920 (N_9920,N_9496,N_9083);
nand U9921 (N_9921,N_9497,N_9428);
nor U9922 (N_9922,N_9336,N_9092);
xnor U9923 (N_9923,N_9035,N_9334);
nand U9924 (N_9924,N_9191,N_9285);
nor U9925 (N_9925,N_9142,N_9311);
or U9926 (N_9926,N_9436,N_9429);
or U9927 (N_9927,N_9109,N_9104);
or U9928 (N_9928,N_9207,N_9171);
nand U9929 (N_9929,N_9115,N_9035);
or U9930 (N_9930,N_9435,N_9402);
xnor U9931 (N_9931,N_9396,N_9039);
or U9932 (N_9932,N_9177,N_9453);
or U9933 (N_9933,N_9479,N_9097);
nor U9934 (N_9934,N_9181,N_9421);
nor U9935 (N_9935,N_9040,N_9300);
nand U9936 (N_9936,N_9446,N_9180);
xnor U9937 (N_9937,N_9423,N_9056);
or U9938 (N_9938,N_9106,N_9366);
nand U9939 (N_9939,N_9371,N_9017);
xor U9940 (N_9940,N_9010,N_9179);
xor U9941 (N_9941,N_9256,N_9356);
or U9942 (N_9942,N_9472,N_9032);
xor U9943 (N_9943,N_9061,N_9439);
and U9944 (N_9944,N_9444,N_9422);
xnor U9945 (N_9945,N_9132,N_9189);
nand U9946 (N_9946,N_9392,N_9272);
xnor U9947 (N_9947,N_9393,N_9495);
nor U9948 (N_9948,N_9179,N_9260);
xnor U9949 (N_9949,N_9460,N_9214);
or U9950 (N_9950,N_9384,N_9138);
nand U9951 (N_9951,N_9146,N_9109);
nor U9952 (N_9952,N_9411,N_9185);
and U9953 (N_9953,N_9336,N_9443);
nor U9954 (N_9954,N_9319,N_9069);
or U9955 (N_9955,N_9186,N_9487);
nor U9956 (N_9956,N_9167,N_9060);
or U9957 (N_9957,N_9363,N_9124);
nor U9958 (N_9958,N_9149,N_9044);
or U9959 (N_9959,N_9163,N_9052);
or U9960 (N_9960,N_9114,N_9118);
xnor U9961 (N_9961,N_9071,N_9356);
or U9962 (N_9962,N_9073,N_9012);
nor U9963 (N_9963,N_9316,N_9442);
or U9964 (N_9964,N_9145,N_9415);
nand U9965 (N_9965,N_9093,N_9116);
nor U9966 (N_9966,N_9007,N_9351);
xor U9967 (N_9967,N_9155,N_9158);
nor U9968 (N_9968,N_9069,N_9484);
nand U9969 (N_9969,N_9000,N_9470);
xor U9970 (N_9970,N_9425,N_9045);
nor U9971 (N_9971,N_9388,N_9351);
xnor U9972 (N_9972,N_9074,N_9395);
or U9973 (N_9973,N_9219,N_9205);
and U9974 (N_9974,N_9306,N_9498);
xnor U9975 (N_9975,N_9401,N_9043);
and U9976 (N_9976,N_9325,N_9417);
and U9977 (N_9977,N_9441,N_9494);
and U9978 (N_9978,N_9448,N_9028);
nor U9979 (N_9979,N_9210,N_9163);
nor U9980 (N_9980,N_9497,N_9081);
and U9981 (N_9981,N_9294,N_9214);
or U9982 (N_9982,N_9397,N_9256);
or U9983 (N_9983,N_9416,N_9243);
xnor U9984 (N_9984,N_9094,N_9383);
and U9985 (N_9985,N_9411,N_9375);
and U9986 (N_9986,N_9199,N_9061);
nand U9987 (N_9987,N_9305,N_9367);
or U9988 (N_9988,N_9023,N_9304);
nor U9989 (N_9989,N_9459,N_9354);
xnor U9990 (N_9990,N_9120,N_9331);
and U9991 (N_9991,N_9245,N_9418);
nor U9992 (N_9992,N_9291,N_9359);
xor U9993 (N_9993,N_9101,N_9420);
or U9994 (N_9994,N_9211,N_9080);
xor U9995 (N_9995,N_9393,N_9404);
and U9996 (N_9996,N_9180,N_9062);
and U9997 (N_9997,N_9230,N_9272);
nand U9998 (N_9998,N_9348,N_9289);
xor U9999 (N_9999,N_9492,N_9069);
and U10000 (N_10000,N_9904,N_9597);
or U10001 (N_10001,N_9771,N_9880);
or U10002 (N_10002,N_9945,N_9815);
nand U10003 (N_10003,N_9690,N_9654);
and U10004 (N_10004,N_9641,N_9881);
and U10005 (N_10005,N_9850,N_9606);
and U10006 (N_10006,N_9914,N_9998);
nand U10007 (N_10007,N_9609,N_9896);
nor U10008 (N_10008,N_9522,N_9991);
xnor U10009 (N_10009,N_9842,N_9649);
or U10010 (N_10010,N_9915,N_9903);
and U10011 (N_10011,N_9767,N_9770);
and U10012 (N_10012,N_9584,N_9685);
nand U10013 (N_10013,N_9849,N_9604);
nor U10014 (N_10014,N_9612,N_9683);
nor U10015 (N_10015,N_9553,N_9673);
nand U10016 (N_10016,N_9759,N_9986);
and U10017 (N_10017,N_9530,N_9971);
xor U10018 (N_10018,N_9718,N_9885);
or U10019 (N_10019,N_9941,N_9708);
or U10020 (N_10020,N_9848,N_9954);
or U10021 (N_10021,N_9669,N_9982);
xor U10022 (N_10022,N_9875,N_9811);
nand U10023 (N_10023,N_9660,N_9816);
xnor U10024 (N_10024,N_9961,N_9664);
nand U10025 (N_10025,N_9934,N_9587);
nor U10026 (N_10026,N_9514,N_9826);
or U10027 (N_10027,N_9720,N_9761);
or U10028 (N_10028,N_9920,N_9916);
xnor U10029 (N_10029,N_9800,N_9756);
nor U10030 (N_10030,N_9861,N_9699);
and U10031 (N_10031,N_9693,N_9882);
xor U10032 (N_10032,N_9924,N_9860);
or U10033 (N_10033,N_9837,N_9757);
or U10034 (N_10034,N_9653,N_9758);
or U10035 (N_10035,N_9959,N_9547);
xnor U10036 (N_10036,N_9824,N_9626);
xnor U10037 (N_10037,N_9561,N_9675);
nor U10038 (N_10038,N_9734,N_9859);
xnor U10039 (N_10039,N_9987,N_9972);
and U10040 (N_10040,N_9546,N_9878);
xnor U10041 (N_10041,N_9802,N_9732);
or U10042 (N_10042,N_9817,N_9872);
nand U10043 (N_10043,N_9554,N_9648);
nor U10044 (N_10044,N_9864,N_9845);
xnor U10045 (N_10045,N_9764,N_9911);
or U10046 (N_10046,N_9936,N_9957);
and U10047 (N_10047,N_9948,N_9536);
and U10048 (N_10048,N_9605,N_9560);
or U10049 (N_10049,N_9651,N_9777);
xor U10050 (N_10050,N_9836,N_9969);
or U10051 (N_10051,N_9960,N_9712);
or U10052 (N_10052,N_9978,N_9659);
nand U10053 (N_10053,N_9611,N_9939);
nor U10054 (N_10054,N_9766,N_9876);
and U10055 (N_10055,N_9567,N_9899);
nand U10056 (N_10056,N_9863,N_9513);
nand U10057 (N_10057,N_9932,N_9588);
nand U10058 (N_10058,N_9517,N_9744);
or U10059 (N_10059,N_9794,N_9602);
nor U10060 (N_10060,N_9773,N_9974);
xnor U10061 (N_10061,N_9727,N_9776);
xnor U10062 (N_10062,N_9716,N_9742);
or U10063 (N_10063,N_9753,N_9599);
or U10064 (N_10064,N_9698,N_9938);
and U10065 (N_10065,N_9964,N_9709);
and U10066 (N_10066,N_9990,N_9804);
or U10067 (N_10067,N_9821,N_9722);
or U10068 (N_10068,N_9857,N_9908);
or U10069 (N_10069,N_9928,N_9502);
xor U10070 (N_10070,N_9607,N_9565);
xnor U10071 (N_10071,N_9970,N_9680);
and U10072 (N_10072,N_9900,N_9687);
xor U10073 (N_10073,N_9563,N_9595);
nand U10074 (N_10074,N_9894,N_9645);
xor U10075 (N_10075,N_9762,N_9585);
nand U10076 (N_10076,N_9644,N_9573);
xor U10077 (N_10077,N_9737,N_9786);
and U10078 (N_10078,N_9576,N_9636);
nand U10079 (N_10079,N_9862,N_9510);
and U10080 (N_10080,N_9662,N_9808);
or U10081 (N_10081,N_9608,N_9877);
or U10082 (N_10082,N_9526,N_9858);
and U10083 (N_10083,N_9840,N_9906);
or U10084 (N_10084,N_9593,N_9754);
xor U10085 (N_10085,N_9844,N_9962);
or U10086 (N_10086,N_9634,N_9729);
or U10087 (N_10087,N_9516,N_9967);
xnor U10088 (N_10088,N_9582,N_9600);
and U10089 (N_10089,N_9658,N_9571);
xor U10090 (N_10090,N_9772,N_9704);
xnor U10091 (N_10091,N_9854,N_9806);
xnor U10092 (N_10092,N_9999,N_9968);
nand U10093 (N_10093,N_9851,N_9639);
nand U10094 (N_10094,N_9796,N_9705);
or U10095 (N_10095,N_9801,N_9839);
nand U10096 (N_10096,N_9763,N_9564);
and U10097 (N_10097,N_9784,N_9622);
and U10098 (N_10098,N_9689,N_9907);
and U10099 (N_10099,N_9694,N_9581);
or U10100 (N_10100,N_9993,N_9696);
or U10101 (N_10101,N_9892,N_9966);
xor U10102 (N_10102,N_9504,N_9943);
xor U10103 (N_10103,N_9765,N_9655);
xor U10104 (N_10104,N_9549,N_9615);
xor U10105 (N_10105,N_9511,N_9621);
nand U10106 (N_10106,N_9995,N_9681);
or U10107 (N_10107,N_9719,N_9871);
and U10108 (N_10108,N_9847,N_9527);
or U10109 (N_10109,N_9782,N_9726);
or U10110 (N_10110,N_9623,N_9569);
or U10111 (N_10111,N_9556,N_9975);
or U10112 (N_10112,N_9503,N_9515);
or U10113 (N_10113,N_9724,N_9946);
nand U10114 (N_10114,N_9947,N_9852);
or U10115 (N_10115,N_9632,N_9937);
xor U10116 (N_10116,N_9702,N_9940);
and U10117 (N_10117,N_9520,N_9787);
and U10118 (N_10118,N_9890,N_9665);
xnor U10119 (N_10119,N_9614,N_9559);
xor U10120 (N_10120,N_9731,N_9883);
and U10121 (N_10121,N_9671,N_9925);
and U10122 (N_10122,N_9829,N_9589);
nor U10123 (N_10123,N_9867,N_9590);
nor U10124 (N_10124,N_9919,N_9538);
and U10125 (N_10125,N_9841,N_9843);
and U10126 (N_10126,N_9524,N_9578);
and U10127 (N_10127,N_9596,N_9679);
nand U10128 (N_10128,N_9898,N_9748);
xnor U10129 (N_10129,N_9952,N_9781);
or U10130 (N_10130,N_9501,N_9789);
nor U10131 (N_10131,N_9778,N_9783);
xor U10132 (N_10132,N_9973,N_9977);
or U10133 (N_10133,N_9529,N_9713);
nand U10134 (N_10134,N_9544,N_9834);
or U10135 (N_10135,N_9523,N_9631);
and U10136 (N_10136,N_9535,N_9942);
and U10137 (N_10137,N_9979,N_9785);
nand U10138 (N_10138,N_9819,N_9537);
xnor U10139 (N_10139,N_9927,N_9682);
nor U10140 (N_10140,N_9506,N_9820);
xor U10141 (N_10141,N_9674,N_9981);
nor U10142 (N_10142,N_9901,N_9886);
nand U10143 (N_10143,N_9656,N_9566);
and U10144 (N_10144,N_9574,N_9628);
nand U10145 (N_10145,N_9629,N_9866);
or U10146 (N_10146,N_9846,N_9598);
or U10147 (N_10147,N_9638,N_9805);
nand U10148 (N_10148,N_9730,N_9921);
and U10149 (N_10149,N_9933,N_9521);
xor U10150 (N_10150,N_9795,N_9922);
nor U10151 (N_10151,N_9743,N_9775);
nand U10152 (N_10152,N_9518,N_9617);
xnor U10153 (N_10153,N_9684,N_9868);
or U10154 (N_10154,N_9910,N_9663);
xnor U10155 (N_10155,N_9799,N_9525);
nor U10156 (N_10156,N_9555,N_9642);
xor U10157 (N_10157,N_9780,N_9562);
nor U10158 (N_10158,N_9723,N_9703);
or U10159 (N_10159,N_9887,N_9838);
xor U10160 (N_10160,N_9616,N_9798);
nand U10161 (N_10161,N_9930,N_9706);
or U10162 (N_10162,N_9591,N_9953);
xor U10163 (N_10163,N_9958,N_9735);
xor U10164 (N_10164,N_9557,N_9640);
nor U10165 (N_10165,N_9989,N_9750);
nand U10166 (N_10166,N_9733,N_9893);
and U10167 (N_10167,N_9895,N_9779);
nor U10168 (N_10168,N_9650,N_9738);
xnor U10169 (N_10169,N_9740,N_9828);
nand U10170 (N_10170,N_9807,N_9913);
nand U10171 (N_10171,N_9539,N_9884);
nor U10172 (N_10172,N_9668,N_9984);
nand U10173 (N_10173,N_9902,N_9949);
and U10174 (N_10174,N_9630,N_9992);
nand U10175 (N_10175,N_9688,N_9749);
and U10176 (N_10176,N_9728,N_9792);
or U10177 (N_10177,N_9701,N_9646);
and U10178 (N_10178,N_9865,N_9586);
or U10179 (N_10179,N_9528,N_9714);
and U10180 (N_10180,N_9905,N_9545);
or U10181 (N_10181,N_9917,N_9980);
xnor U10182 (N_10182,N_9793,N_9620);
or U10183 (N_10183,N_9889,N_9739);
and U10184 (N_10184,N_9788,N_9583);
xnor U10185 (N_10185,N_9891,N_9822);
or U10186 (N_10186,N_9711,N_9963);
nor U10187 (N_10187,N_9831,N_9790);
nor U10188 (N_10188,N_9827,N_9552);
nor U10189 (N_10189,N_9580,N_9717);
nor U10190 (N_10190,N_9769,N_9951);
or U10191 (N_10191,N_9603,N_9570);
and U10192 (N_10192,N_9624,N_9736);
nor U10193 (N_10193,N_9768,N_9601);
xor U10194 (N_10194,N_9825,N_9677);
nand U10195 (N_10195,N_9550,N_9507);
and U10196 (N_10196,N_9809,N_9508);
or U10197 (N_10197,N_9558,N_9812);
nand U10198 (N_10198,N_9542,N_9613);
nand U10199 (N_10199,N_9814,N_9944);
and U10200 (N_10200,N_9707,N_9956);
or U10201 (N_10201,N_9912,N_9935);
nand U10202 (N_10202,N_9996,N_9965);
xor U10203 (N_10203,N_9803,N_9874);
nor U10204 (N_10204,N_9540,N_9647);
xnor U10205 (N_10205,N_9997,N_9592);
and U10206 (N_10206,N_9572,N_9519);
xnor U10207 (N_10207,N_9856,N_9746);
nor U10208 (N_10208,N_9879,N_9532);
nand U10209 (N_10209,N_9627,N_9985);
xnor U10210 (N_10210,N_9870,N_9994);
nand U10211 (N_10211,N_9512,N_9830);
or U10212 (N_10212,N_9618,N_9909);
or U10213 (N_10213,N_9551,N_9823);
or U10214 (N_10214,N_9509,N_9929);
nand U10215 (N_10215,N_9950,N_9751);
nand U10216 (N_10216,N_9594,N_9774);
nor U10217 (N_10217,N_9625,N_9752);
and U10218 (N_10218,N_9700,N_9923);
and U10219 (N_10219,N_9976,N_9855);
nand U10220 (N_10220,N_9721,N_9918);
nor U10221 (N_10221,N_9531,N_9575);
xor U10222 (N_10222,N_9619,N_9568);
and U10223 (N_10223,N_9813,N_9810);
and U10224 (N_10224,N_9633,N_9661);
nor U10225 (N_10225,N_9686,N_9797);
or U10226 (N_10226,N_9755,N_9931);
or U10227 (N_10227,N_9988,N_9505);
nand U10228 (N_10228,N_9741,N_9500);
and U10229 (N_10229,N_9637,N_9869);
and U10230 (N_10230,N_9543,N_9715);
xnor U10231 (N_10231,N_9791,N_9652);
nand U10232 (N_10232,N_9541,N_9853);
nor U10233 (N_10233,N_9533,N_9897);
nor U10234 (N_10234,N_9833,N_9818);
and U10235 (N_10235,N_9760,N_9725);
nor U10236 (N_10236,N_9534,N_9670);
nor U10237 (N_10237,N_9678,N_9548);
nor U10238 (N_10238,N_9747,N_9610);
nand U10239 (N_10239,N_9657,N_9697);
nor U10240 (N_10240,N_9832,N_9710);
and U10241 (N_10241,N_9745,N_9666);
nor U10242 (N_10242,N_9926,N_9643);
nor U10243 (N_10243,N_9579,N_9695);
nand U10244 (N_10244,N_9635,N_9672);
nor U10245 (N_10245,N_9873,N_9835);
or U10246 (N_10246,N_9692,N_9577);
and U10247 (N_10247,N_9676,N_9691);
nor U10248 (N_10248,N_9983,N_9888);
nor U10249 (N_10249,N_9955,N_9667);
and U10250 (N_10250,N_9958,N_9957);
nand U10251 (N_10251,N_9776,N_9831);
nor U10252 (N_10252,N_9891,N_9679);
xnor U10253 (N_10253,N_9672,N_9967);
or U10254 (N_10254,N_9646,N_9503);
or U10255 (N_10255,N_9583,N_9613);
nor U10256 (N_10256,N_9969,N_9800);
or U10257 (N_10257,N_9602,N_9907);
nand U10258 (N_10258,N_9993,N_9996);
xor U10259 (N_10259,N_9771,N_9608);
or U10260 (N_10260,N_9555,N_9672);
and U10261 (N_10261,N_9674,N_9588);
xor U10262 (N_10262,N_9939,N_9867);
and U10263 (N_10263,N_9685,N_9523);
nor U10264 (N_10264,N_9939,N_9995);
xor U10265 (N_10265,N_9694,N_9548);
or U10266 (N_10266,N_9666,N_9882);
xor U10267 (N_10267,N_9968,N_9949);
xor U10268 (N_10268,N_9647,N_9926);
nor U10269 (N_10269,N_9640,N_9948);
xor U10270 (N_10270,N_9728,N_9745);
or U10271 (N_10271,N_9552,N_9871);
nor U10272 (N_10272,N_9826,N_9707);
nand U10273 (N_10273,N_9504,N_9518);
nand U10274 (N_10274,N_9810,N_9614);
and U10275 (N_10275,N_9529,N_9574);
xnor U10276 (N_10276,N_9824,N_9616);
xnor U10277 (N_10277,N_9600,N_9768);
nand U10278 (N_10278,N_9958,N_9638);
and U10279 (N_10279,N_9878,N_9554);
nand U10280 (N_10280,N_9738,N_9775);
nor U10281 (N_10281,N_9828,N_9985);
xor U10282 (N_10282,N_9909,N_9900);
nor U10283 (N_10283,N_9773,N_9993);
or U10284 (N_10284,N_9966,N_9929);
and U10285 (N_10285,N_9880,N_9730);
or U10286 (N_10286,N_9764,N_9798);
nor U10287 (N_10287,N_9667,N_9856);
and U10288 (N_10288,N_9823,N_9905);
nor U10289 (N_10289,N_9813,N_9665);
or U10290 (N_10290,N_9657,N_9859);
nand U10291 (N_10291,N_9916,N_9898);
or U10292 (N_10292,N_9571,N_9964);
nor U10293 (N_10293,N_9527,N_9590);
and U10294 (N_10294,N_9992,N_9508);
or U10295 (N_10295,N_9692,N_9736);
or U10296 (N_10296,N_9516,N_9634);
nor U10297 (N_10297,N_9554,N_9502);
nor U10298 (N_10298,N_9988,N_9961);
and U10299 (N_10299,N_9996,N_9864);
and U10300 (N_10300,N_9749,N_9623);
nor U10301 (N_10301,N_9688,N_9647);
nand U10302 (N_10302,N_9755,N_9627);
or U10303 (N_10303,N_9785,N_9730);
nor U10304 (N_10304,N_9907,N_9546);
and U10305 (N_10305,N_9714,N_9720);
xor U10306 (N_10306,N_9634,N_9662);
nand U10307 (N_10307,N_9794,N_9643);
nor U10308 (N_10308,N_9656,N_9813);
nor U10309 (N_10309,N_9531,N_9630);
nand U10310 (N_10310,N_9745,N_9704);
and U10311 (N_10311,N_9747,N_9654);
nand U10312 (N_10312,N_9576,N_9560);
nor U10313 (N_10313,N_9593,N_9746);
xnor U10314 (N_10314,N_9640,N_9538);
or U10315 (N_10315,N_9794,N_9726);
and U10316 (N_10316,N_9843,N_9798);
xor U10317 (N_10317,N_9589,N_9714);
nor U10318 (N_10318,N_9948,N_9826);
or U10319 (N_10319,N_9763,N_9970);
nor U10320 (N_10320,N_9967,N_9841);
or U10321 (N_10321,N_9563,N_9507);
nand U10322 (N_10322,N_9793,N_9754);
or U10323 (N_10323,N_9864,N_9576);
xor U10324 (N_10324,N_9990,N_9770);
or U10325 (N_10325,N_9901,N_9683);
nor U10326 (N_10326,N_9917,N_9873);
xor U10327 (N_10327,N_9611,N_9509);
nand U10328 (N_10328,N_9547,N_9780);
xnor U10329 (N_10329,N_9971,N_9907);
xnor U10330 (N_10330,N_9782,N_9898);
nand U10331 (N_10331,N_9913,N_9562);
nand U10332 (N_10332,N_9545,N_9678);
and U10333 (N_10333,N_9748,N_9640);
and U10334 (N_10334,N_9967,N_9729);
or U10335 (N_10335,N_9950,N_9663);
nor U10336 (N_10336,N_9590,N_9832);
and U10337 (N_10337,N_9921,N_9851);
and U10338 (N_10338,N_9875,N_9742);
nor U10339 (N_10339,N_9759,N_9559);
nor U10340 (N_10340,N_9818,N_9961);
nand U10341 (N_10341,N_9977,N_9858);
nand U10342 (N_10342,N_9831,N_9876);
and U10343 (N_10343,N_9755,N_9543);
nand U10344 (N_10344,N_9917,N_9584);
nor U10345 (N_10345,N_9759,N_9817);
or U10346 (N_10346,N_9577,N_9612);
nand U10347 (N_10347,N_9834,N_9678);
xor U10348 (N_10348,N_9660,N_9511);
nand U10349 (N_10349,N_9570,N_9768);
xnor U10350 (N_10350,N_9585,N_9811);
nand U10351 (N_10351,N_9934,N_9828);
nor U10352 (N_10352,N_9901,N_9570);
and U10353 (N_10353,N_9676,N_9956);
nor U10354 (N_10354,N_9677,N_9914);
nor U10355 (N_10355,N_9792,N_9761);
nand U10356 (N_10356,N_9787,N_9626);
xnor U10357 (N_10357,N_9985,N_9782);
xor U10358 (N_10358,N_9896,N_9851);
nand U10359 (N_10359,N_9573,N_9795);
xor U10360 (N_10360,N_9693,N_9784);
nand U10361 (N_10361,N_9637,N_9729);
xor U10362 (N_10362,N_9765,N_9559);
xor U10363 (N_10363,N_9665,N_9905);
or U10364 (N_10364,N_9583,N_9618);
or U10365 (N_10365,N_9900,N_9734);
or U10366 (N_10366,N_9867,N_9519);
or U10367 (N_10367,N_9587,N_9592);
or U10368 (N_10368,N_9547,N_9607);
and U10369 (N_10369,N_9569,N_9627);
xor U10370 (N_10370,N_9624,N_9944);
nand U10371 (N_10371,N_9661,N_9585);
nand U10372 (N_10372,N_9628,N_9783);
nor U10373 (N_10373,N_9916,N_9562);
xnor U10374 (N_10374,N_9777,N_9760);
nand U10375 (N_10375,N_9613,N_9647);
and U10376 (N_10376,N_9674,N_9576);
nand U10377 (N_10377,N_9747,N_9745);
or U10378 (N_10378,N_9594,N_9694);
or U10379 (N_10379,N_9510,N_9725);
nor U10380 (N_10380,N_9757,N_9796);
nor U10381 (N_10381,N_9661,N_9723);
xnor U10382 (N_10382,N_9552,N_9733);
nor U10383 (N_10383,N_9743,N_9993);
nand U10384 (N_10384,N_9947,N_9654);
and U10385 (N_10385,N_9792,N_9845);
and U10386 (N_10386,N_9874,N_9956);
nand U10387 (N_10387,N_9946,N_9805);
and U10388 (N_10388,N_9798,N_9746);
and U10389 (N_10389,N_9857,N_9546);
nand U10390 (N_10390,N_9710,N_9609);
nor U10391 (N_10391,N_9517,N_9926);
nor U10392 (N_10392,N_9840,N_9757);
or U10393 (N_10393,N_9593,N_9898);
nand U10394 (N_10394,N_9524,N_9869);
nor U10395 (N_10395,N_9686,N_9862);
nand U10396 (N_10396,N_9791,N_9730);
or U10397 (N_10397,N_9778,N_9541);
or U10398 (N_10398,N_9897,N_9796);
and U10399 (N_10399,N_9519,N_9979);
nand U10400 (N_10400,N_9853,N_9658);
xnor U10401 (N_10401,N_9883,N_9689);
or U10402 (N_10402,N_9640,N_9910);
and U10403 (N_10403,N_9541,N_9532);
and U10404 (N_10404,N_9633,N_9960);
or U10405 (N_10405,N_9995,N_9770);
xnor U10406 (N_10406,N_9999,N_9734);
or U10407 (N_10407,N_9643,N_9683);
xor U10408 (N_10408,N_9656,N_9942);
nor U10409 (N_10409,N_9989,N_9953);
or U10410 (N_10410,N_9826,N_9537);
or U10411 (N_10411,N_9717,N_9879);
xnor U10412 (N_10412,N_9718,N_9545);
and U10413 (N_10413,N_9712,N_9747);
and U10414 (N_10414,N_9964,N_9986);
xor U10415 (N_10415,N_9681,N_9565);
and U10416 (N_10416,N_9881,N_9744);
nand U10417 (N_10417,N_9531,N_9860);
and U10418 (N_10418,N_9990,N_9994);
nand U10419 (N_10419,N_9522,N_9954);
and U10420 (N_10420,N_9854,N_9997);
nor U10421 (N_10421,N_9842,N_9639);
xnor U10422 (N_10422,N_9932,N_9990);
nor U10423 (N_10423,N_9735,N_9702);
xor U10424 (N_10424,N_9937,N_9755);
xor U10425 (N_10425,N_9979,N_9599);
nor U10426 (N_10426,N_9575,N_9987);
or U10427 (N_10427,N_9626,N_9865);
nand U10428 (N_10428,N_9995,N_9636);
nor U10429 (N_10429,N_9858,N_9922);
xnor U10430 (N_10430,N_9718,N_9605);
or U10431 (N_10431,N_9761,N_9717);
and U10432 (N_10432,N_9681,N_9974);
and U10433 (N_10433,N_9661,N_9644);
nand U10434 (N_10434,N_9649,N_9967);
and U10435 (N_10435,N_9688,N_9625);
or U10436 (N_10436,N_9936,N_9871);
nand U10437 (N_10437,N_9724,N_9559);
or U10438 (N_10438,N_9999,N_9858);
xnor U10439 (N_10439,N_9685,N_9822);
and U10440 (N_10440,N_9672,N_9984);
and U10441 (N_10441,N_9880,N_9940);
nand U10442 (N_10442,N_9777,N_9997);
xor U10443 (N_10443,N_9845,N_9821);
nor U10444 (N_10444,N_9981,N_9930);
and U10445 (N_10445,N_9645,N_9697);
or U10446 (N_10446,N_9751,N_9598);
xor U10447 (N_10447,N_9930,N_9788);
and U10448 (N_10448,N_9909,N_9641);
nor U10449 (N_10449,N_9637,N_9545);
nand U10450 (N_10450,N_9892,N_9534);
nor U10451 (N_10451,N_9661,N_9948);
xor U10452 (N_10452,N_9829,N_9655);
xor U10453 (N_10453,N_9867,N_9544);
nor U10454 (N_10454,N_9685,N_9962);
nand U10455 (N_10455,N_9944,N_9535);
xnor U10456 (N_10456,N_9837,N_9512);
and U10457 (N_10457,N_9782,N_9869);
nand U10458 (N_10458,N_9958,N_9605);
or U10459 (N_10459,N_9758,N_9636);
and U10460 (N_10460,N_9856,N_9878);
nand U10461 (N_10461,N_9974,N_9998);
and U10462 (N_10462,N_9586,N_9506);
xnor U10463 (N_10463,N_9945,N_9962);
nor U10464 (N_10464,N_9569,N_9923);
or U10465 (N_10465,N_9820,N_9635);
nor U10466 (N_10466,N_9524,N_9633);
xnor U10467 (N_10467,N_9632,N_9694);
nor U10468 (N_10468,N_9574,N_9800);
nor U10469 (N_10469,N_9695,N_9585);
nand U10470 (N_10470,N_9730,N_9969);
nand U10471 (N_10471,N_9821,N_9503);
and U10472 (N_10472,N_9871,N_9507);
and U10473 (N_10473,N_9792,N_9505);
or U10474 (N_10474,N_9717,N_9810);
and U10475 (N_10475,N_9938,N_9599);
nor U10476 (N_10476,N_9931,N_9725);
xor U10477 (N_10477,N_9508,N_9774);
xnor U10478 (N_10478,N_9646,N_9623);
and U10479 (N_10479,N_9559,N_9955);
and U10480 (N_10480,N_9946,N_9986);
xnor U10481 (N_10481,N_9751,N_9589);
nand U10482 (N_10482,N_9594,N_9610);
or U10483 (N_10483,N_9929,N_9794);
nor U10484 (N_10484,N_9898,N_9519);
xor U10485 (N_10485,N_9701,N_9692);
and U10486 (N_10486,N_9831,N_9596);
nand U10487 (N_10487,N_9856,N_9741);
xnor U10488 (N_10488,N_9637,N_9938);
and U10489 (N_10489,N_9501,N_9715);
nand U10490 (N_10490,N_9574,N_9920);
or U10491 (N_10491,N_9501,N_9547);
nand U10492 (N_10492,N_9724,N_9909);
nand U10493 (N_10493,N_9502,N_9567);
nand U10494 (N_10494,N_9838,N_9912);
nand U10495 (N_10495,N_9743,N_9924);
or U10496 (N_10496,N_9667,N_9839);
or U10497 (N_10497,N_9716,N_9567);
nor U10498 (N_10498,N_9657,N_9839);
nand U10499 (N_10499,N_9615,N_9777);
and U10500 (N_10500,N_10317,N_10249);
xnor U10501 (N_10501,N_10054,N_10238);
nor U10502 (N_10502,N_10177,N_10000);
and U10503 (N_10503,N_10481,N_10042);
or U10504 (N_10504,N_10183,N_10160);
nor U10505 (N_10505,N_10327,N_10422);
or U10506 (N_10506,N_10149,N_10028);
nand U10507 (N_10507,N_10113,N_10403);
or U10508 (N_10508,N_10460,N_10179);
and U10509 (N_10509,N_10125,N_10003);
and U10510 (N_10510,N_10118,N_10194);
xor U10511 (N_10511,N_10369,N_10310);
xnor U10512 (N_10512,N_10338,N_10137);
nor U10513 (N_10513,N_10409,N_10335);
xor U10514 (N_10514,N_10455,N_10474);
and U10515 (N_10515,N_10124,N_10260);
xor U10516 (N_10516,N_10464,N_10313);
and U10517 (N_10517,N_10389,N_10452);
or U10518 (N_10518,N_10448,N_10405);
and U10519 (N_10519,N_10371,N_10044);
and U10520 (N_10520,N_10312,N_10075);
or U10521 (N_10521,N_10127,N_10472);
or U10522 (N_10522,N_10341,N_10352);
or U10523 (N_10523,N_10357,N_10039);
and U10524 (N_10524,N_10411,N_10220);
or U10525 (N_10525,N_10202,N_10120);
xor U10526 (N_10526,N_10283,N_10100);
or U10527 (N_10527,N_10226,N_10138);
xnor U10528 (N_10528,N_10205,N_10081);
and U10529 (N_10529,N_10402,N_10478);
and U10530 (N_10530,N_10269,N_10439);
and U10531 (N_10531,N_10417,N_10350);
xnor U10532 (N_10532,N_10356,N_10180);
and U10533 (N_10533,N_10092,N_10461);
or U10534 (N_10534,N_10359,N_10107);
or U10535 (N_10535,N_10302,N_10366);
nor U10536 (N_10536,N_10032,N_10470);
and U10537 (N_10537,N_10383,N_10274);
nand U10538 (N_10538,N_10386,N_10395);
nand U10539 (N_10539,N_10372,N_10201);
and U10540 (N_10540,N_10326,N_10370);
or U10541 (N_10541,N_10355,N_10353);
nor U10542 (N_10542,N_10027,N_10459);
nand U10543 (N_10543,N_10303,N_10440);
xnor U10544 (N_10544,N_10024,N_10112);
and U10545 (N_10545,N_10189,N_10301);
xnor U10546 (N_10546,N_10408,N_10410);
nor U10547 (N_10547,N_10026,N_10047);
or U10548 (N_10548,N_10135,N_10190);
and U10549 (N_10549,N_10126,N_10087);
xor U10550 (N_10550,N_10074,N_10485);
xnor U10551 (N_10551,N_10421,N_10415);
nor U10552 (N_10552,N_10392,N_10334);
and U10553 (N_10553,N_10433,N_10157);
xnor U10554 (N_10554,N_10059,N_10367);
nand U10555 (N_10555,N_10017,N_10342);
or U10556 (N_10556,N_10099,N_10245);
nor U10557 (N_10557,N_10071,N_10469);
and U10558 (N_10558,N_10193,N_10022);
xnor U10559 (N_10559,N_10115,N_10178);
nand U10560 (N_10560,N_10451,N_10407);
nand U10561 (N_10561,N_10321,N_10045);
nor U10562 (N_10562,N_10465,N_10295);
xnor U10563 (N_10563,N_10457,N_10446);
xor U10564 (N_10564,N_10221,N_10218);
and U10565 (N_10565,N_10215,N_10288);
nor U10566 (N_10566,N_10234,N_10393);
and U10567 (N_10567,N_10311,N_10196);
or U10568 (N_10568,N_10363,N_10197);
xor U10569 (N_10569,N_10466,N_10148);
xnor U10570 (N_10570,N_10108,N_10060);
xnor U10571 (N_10571,N_10486,N_10299);
and U10572 (N_10572,N_10134,N_10235);
nand U10573 (N_10573,N_10094,N_10128);
xor U10574 (N_10574,N_10061,N_10257);
nand U10575 (N_10575,N_10471,N_10263);
nand U10576 (N_10576,N_10343,N_10225);
nand U10577 (N_10577,N_10067,N_10442);
nand U10578 (N_10578,N_10420,N_10033);
xor U10579 (N_10579,N_10462,N_10055);
nand U10580 (N_10580,N_10499,N_10058);
nand U10581 (N_10581,N_10449,N_10078);
nor U10582 (N_10582,N_10423,N_10318);
nor U10583 (N_10583,N_10289,N_10002);
xor U10584 (N_10584,N_10103,N_10139);
and U10585 (N_10585,N_10132,N_10144);
xor U10586 (N_10586,N_10337,N_10016);
or U10587 (N_10587,N_10390,N_10171);
or U10588 (N_10588,N_10043,N_10285);
xor U10589 (N_10589,N_10164,N_10019);
xor U10590 (N_10590,N_10004,N_10090);
nand U10591 (N_10591,N_10458,N_10111);
and U10592 (N_10592,N_10129,N_10314);
xnor U10593 (N_10593,N_10377,N_10438);
nor U10594 (N_10594,N_10426,N_10292);
and U10595 (N_10595,N_10276,N_10480);
or U10596 (N_10596,N_10354,N_10294);
and U10597 (N_10597,N_10162,N_10284);
nor U10598 (N_10598,N_10324,N_10007);
or U10599 (N_10599,N_10053,N_10333);
nor U10600 (N_10600,N_10089,N_10418);
and U10601 (N_10601,N_10040,N_10435);
nand U10602 (N_10602,N_10308,N_10203);
nand U10603 (N_10603,N_10241,N_10250);
or U10604 (N_10604,N_10325,N_10242);
nand U10605 (N_10605,N_10217,N_10315);
nand U10606 (N_10606,N_10101,N_10165);
nand U10607 (N_10607,N_10166,N_10271);
nor U10608 (N_10608,N_10298,N_10009);
nand U10609 (N_10609,N_10488,N_10006);
and U10610 (N_10610,N_10320,N_10484);
xnor U10611 (N_10611,N_10211,N_10419);
nand U10612 (N_10612,N_10198,N_10209);
xnor U10613 (N_10613,N_10114,N_10096);
nor U10614 (N_10614,N_10261,N_10041);
nand U10615 (N_10615,N_10265,N_10428);
nor U10616 (N_10616,N_10079,N_10098);
or U10617 (N_10617,N_10266,N_10191);
and U10618 (N_10618,N_10048,N_10012);
and U10619 (N_10619,N_10216,N_10210);
xnor U10620 (N_10620,N_10319,N_10119);
nand U10621 (N_10621,N_10330,N_10362);
nand U10622 (N_10622,N_10279,N_10391);
and U10623 (N_10623,N_10328,N_10412);
or U10624 (N_10624,N_10483,N_10181);
nor U10625 (N_10625,N_10093,N_10150);
xor U10626 (N_10626,N_10222,N_10429);
and U10627 (N_10627,N_10229,N_10404);
xnor U10628 (N_10628,N_10425,N_10256);
nor U10629 (N_10629,N_10175,N_10029);
or U10630 (N_10630,N_10495,N_10049);
xor U10631 (N_10631,N_10219,N_10456);
xor U10632 (N_10632,N_10168,N_10236);
xor U10633 (N_10633,N_10349,N_10035);
nor U10634 (N_10634,N_10116,N_10434);
nand U10635 (N_10635,N_10163,N_10212);
nand U10636 (N_10636,N_10489,N_10014);
nor U10637 (N_10637,N_10277,N_10368);
nor U10638 (N_10638,N_10316,N_10005);
xor U10639 (N_10639,N_10188,N_10104);
xnor U10640 (N_10640,N_10496,N_10036);
xor U10641 (N_10641,N_10056,N_10463);
xor U10642 (N_10642,N_10037,N_10167);
xor U10643 (N_10643,N_10381,N_10297);
and U10644 (N_10644,N_10063,N_10182);
xnor U10645 (N_10645,N_10070,N_10214);
nand U10646 (N_10646,N_10360,N_10291);
nand U10647 (N_10647,N_10254,N_10062);
or U10648 (N_10648,N_10145,N_10095);
or U10649 (N_10649,N_10482,N_10154);
nand U10650 (N_10650,N_10146,N_10185);
nor U10651 (N_10651,N_10388,N_10064);
nor U10652 (N_10652,N_10227,N_10228);
nand U10653 (N_10653,N_10244,N_10382);
nor U10654 (N_10654,N_10267,N_10153);
xor U10655 (N_10655,N_10176,N_10376);
nor U10656 (N_10656,N_10052,N_10130);
xor U10657 (N_10657,N_10020,N_10379);
nand U10658 (N_10658,N_10206,N_10172);
and U10659 (N_10659,N_10307,N_10348);
nand U10660 (N_10660,N_10290,N_10424);
nor U10661 (N_10661,N_10273,N_10258);
nand U10662 (N_10662,N_10230,N_10406);
nand U10663 (N_10663,N_10444,N_10268);
nand U10664 (N_10664,N_10492,N_10141);
or U10665 (N_10665,N_10140,N_10309);
xor U10666 (N_10666,N_10015,N_10246);
and U10667 (N_10667,N_10296,N_10476);
nand U10668 (N_10668,N_10468,N_10264);
nand U10669 (N_10669,N_10156,N_10477);
or U10670 (N_10670,N_10046,N_10432);
nor U10671 (N_10671,N_10394,N_10498);
and U10672 (N_10672,N_10018,N_10023);
nor U10673 (N_10673,N_10414,N_10339);
xnor U10674 (N_10674,N_10199,N_10497);
and U10675 (N_10675,N_10345,N_10322);
nor U10676 (N_10676,N_10122,N_10142);
nor U10677 (N_10677,N_10083,N_10192);
or U10678 (N_10678,N_10347,N_10011);
nor U10679 (N_10679,N_10281,N_10110);
or U10680 (N_10680,N_10231,N_10387);
xor U10681 (N_10681,N_10123,N_10025);
nor U10682 (N_10682,N_10385,N_10237);
and U10683 (N_10683,N_10332,N_10454);
or U10684 (N_10684,N_10323,N_10204);
and U10685 (N_10685,N_10151,N_10223);
nor U10686 (N_10686,N_10475,N_10427);
or U10687 (N_10687,N_10351,N_10155);
nand U10688 (N_10688,N_10365,N_10187);
or U10689 (N_10689,N_10300,N_10085);
or U10690 (N_10690,N_10051,N_10473);
nand U10691 (N_10691,N_10080,N_10255);
nor U10692 (N_10692,N_10293,N_10034);
and U10693 (N_10693,N_10340,N_10195);
or U10694 (N_10694,N_10270,N_10361);
or U10695 (N_10695,N_10329,N_10170);
nor U10696 (N_10696,N_10013,N_10494);
and U10697 (N_10697,N_10275,N_10068);
nand U10698 (N_10698,N_10010,N_10105);
or U10699 (N_10699,N_10375,N_10262);
nand U10700 (N_10700,N_10397,N_10431);
nand U10701 (N_10701,N_10253,N_10358);
nor U10702 (N_10702,N_10286,N_10186);
nor U10703 (N_10703,N_10437,N_10445);
and U10704 (N_10704,N_10280,N_10117);
or U10705 (N_10705,N_10443,N_10384);
nand U10706 (N_10706,N_10133,N_10084);
and U10707 (N_10707,N_10207,N_10493);
xor U10708 (N_10708,N_10436,N_10378);
nor U10709 (N_10709,N_10121,N_10441);
or U10710 (N_10710,N_10050,N_10008);
or U10711 (N_10711,N_10213,N_10380);
and U10712 (N_10712,N_10447,N_10416);
or U10713 (N_10713,N_10413,N_10467);
xor U10714 (N_10714,N_10072,N_10161);
nand U10715 (N_10715,N_10091,N_10224);
nand U10716 (N_10716,N_10159,N_10143);
nor U10717 (N_10717,N_10208,N_10396);
nand U10718 (N_10718,N_10305,N_10106);
nor U10719 (N_10719,N_10287,N_10248);
nand U10720 (N_10720,N_10374,N_10346);
nor U10721 (N_10721,N_10252,N_10247);
xnor U10722 (N_10722,N_10184,N_10239);
xnor U10723 (N_10723,N_10001,N_10152);
nand U10724 (N_10724,N_10282,N_10251);
nand U10725 (N_10725,N_10077,N_10073);
nor U10726 (N_10726,N_10200,N_10076);
nor U10727 (N_10727,N_10136,N_10259);
nor U10728 (N_10728,N_10147,N_10030);
or U10729 (N_10729,N_10174,N_10243);
xor U10730 (N_10730,N_10364,N_10088);
xor U10731 (N_10731,N_10400,N_10069);
and U10732 (N_10732,N_10373,N_10490);
nand U10733 (N_10733,N_10065,N_10344);
or U10734 (N_10734,N_10086,N_10278);
nor U10735 (N_10735,N_10399,N_10131);
xor U10736 (N_10736,N_10102,N_10097);
and U10737 (N_10737,N_10336,N_10082);
nor U10738 (N_10738,N_10487,N_10169);
xor U10739 (N_10739,N_10031,N_10272);
xor U10740 (N_10740,N_10158,N_10450);
nand U10741 (N_10741,N_10109,N_10240);
nand U10742 (N_10742,N_10331,N_10232);
xor U10743 (N_10743,N_10233,N_10479);
nor U10744 (N_10744,N_10398,N_10057);
and U10745 (N_10745,N_10491,N_10453);
or U10746 (N_10746,N_10430,N_10066);
and U10747 (N_10747,N_10304,N_10173);
or U10748 (N_10748,N_10021,N_10306);
xor U10749 (N_10749,N_10038,N_10401);
or U10750 (N_10750,N_10012,N_10296);
or U10751 (N_10751,N_10461,N_10454);
and U10752 (N_10752,N_10125,N_10032);
or U10753 (N_10753,N_10436,N_10189);
or U10754 (N_10754,N_10346,N_10277);
or U10755 (N_10755,N_10112,N_10032);
nand U10756 (N_10756,N_10259,N_10472);
nor U10757 (N_10757,N_10299,N_10465);
and U10758 (N_10758,N_10302,N_10050);
xor U10759 (N_10759,N_10062,N_10488);
and U10760 (N_10760,N_10477,N_10112);
nor U10761 (N_10761,N_10149,N_10270);
or U10762 (N_10762,N_10399,N_10172);
xnor U10763 (N_10763,N_10118,N_10214);
nor U10764 (N_10764,N_10460,N_10160);
or U10765 (N_10765,N_10460,N_10332);
nor U10766 (N_10766,N_10225,N_10020);
and U10767 (N_10767,N_10273,N_10224);
and U10768 (N_10768,N_10324,N_10497);
nor U10769 (N_10769,N_10076,N_10432);
nor U10770 (N_10770,N_10103,N_10485);
nand U10771 (N_10771,N_10428,N_10122);
nand U10772 (N_10772,N_10226,N_10326);
and U10773 (N_10773,N_10282,N_10453);
and U10774 (N_10774,N_10454,N_10180);
xor U10775 (N_10775,N_10298,N_10413);
and U10776 (N_10776,N_10364,N_10433);
and U10777 (N_10777,N_10147,N_10353);
nand U10778 (N_10778,N_10412,N_10243);
nand U10779 (N_10779,N_10117,N_10064);
or U10780 (N_10780,N_10339,N_10028);
nand U10781 (N_10781,N_10407,N_10174);
nor U10782 (N_10782,N_10164,N_10191);
xnor U10783 (N_10783,N_10441,N_10174);
nand U10784 (N_10784,N_10367,N_10437);
or U10785 (N_10785,N_10271,N_10424);
nor U10786 (N_10786,N_10165,N_10291);
nor U10787 (N_10787,N_10230,N_10494);
and U10788 (N_10788,N_10127,N_10356);
nand U10789 (N_10789,N_10486,N_10027);
nor U10790 (N_10790,N_10438,N_10085);
nor U10791 (N_10791,N_10415,N_10470);
or U10792 (N_10792,N_10044,N_10198);
xnor U10793 (N_10793,N_10296,N_10487);
or U10794 (N_10794,N_10008,N_10234);
and U10795 (N_10795,N_10140,N_10343);
xor U10796 (N_10796,N_10129,N_10201);
nand U10797 (N_10797,N_10328,N_10185);
or U10798 (N_10798,N_10085,N_10401);
xor U10799 (N_10799,N_10194,N_10440);
nand U10800 (N_10800,N_10297,N_10433);
xnor U10801 (N_10801,N_10037,N_10154);
and U10802 (N_10802,N_10493,N_10255);
or U10803 (N_10803,N_10143,N_10396);
or U10804 (N_10804,N_10380,N_10459);
nand U10805 (N_10805,N_10479,N_10368);
or U10806 (N_10806,N_10170,N_10392);
or U10807 (N_10807,N_10006,N_10419);
and U10808 (N_10808,N_10295,N_10069);
nand U10809 (N_10809,N_10199,N_10030);
xor U10810 (N_10810,N_10207,N_10106);
nor U10811 (N_10811,N_10363,N_10450);
nand U10812 (N_10812,N_10095,N_10342);
nand U10813 (N_10813,N_10406,N_10110);
nand U10814 (N_10814,N_10056,N_10413);
xnor U10815 (N_10815,N_10252,N_10345);
nor U10816 (N_10816,N_10127,N_10452);
nor U10817 (N_10817,N_10359,N_10221);
and U10818 (N_10818,N_10387,N_10276);
xor U10819 (N_10819,N_10499,N_10126);
xor U10820 (N_10820,N_10364,N_10146);
and U10821 (N_10821,N_10444,N_10046);
or U10822 (N_10822,N_10258,N_10262);
or U10823 (N_10823,N_10434,N_10158);
xnor U10824 (N_10824,N_10310,N_10476);
and U10825 (N_10825,N_10482,N_10323);
or U10826 (N_10826,N_10000,N_10006);
xor U10827 (N_10827,N_10440,N_10152);
or U10828 (N_10828,N_10152,N_10434);
or U10829 (N_10829,N_10363,N_10255);
or U10830 (N_10830,N_10015,N_10213);
nand U10831 (N_10831,N_10267,N_10371);
and U10832 (N_10832,N_10277,N_10492);
and U10833 (N_10833,N_10076,N_10376);
nand U10834 (N_10834,N_10142,N_10042);
nand U10835 (N_10835,N_10093,N_10159);
xnor U10836 (N_10836,N_10065,N_10135);
and U10837 (N_10837,N_10152,N_10294);
or U10838 (N_10838,N_10070,N_10186);
or U10839 (N_10839,N_10105,N_10358);
nor U10840 (N_10840,N_10340,N_10349);
nor U10841 (N_10841,N_10422,N_10008);
nand U10842 (N_10842,N_10339,N_10290);
and U10843 (N_10843,N_10261,N_10098);
or U10844 (N_10844,N_10245,N_10281);
xor U10845 (N_10845,N_10302,N_10016);
or U10846 (N_10846,N_10277,N_10332);
xor U10847 (N_10847,N_10200,N_10229);
nand U10848 (N_10848,N_10416,N_10426);
xnor U10849 (N_10849,N_10185,N_10222);
or U10850 (N_10850,N_10400,N_10357);
and U10851 (N_10851,N_10056,N_10241);
xnor U10852 (N_10852,N_10263,N_10158);
xor U10853 (N_10853,N_10030,N_10385);
and U10854 (N_10854,N_10017,N_10082);
nor U10855 (N_10855,N_10164,N_10470);
nand U10856 (N_10856,N_10365,N_10206);
xor U10857 (N_10857,N_10360,N_10337);
xnor U10858 (N_10858,N_10306,N_10407);
and U10859 (N_10859,N_10129,N_10222);
xor U10860 (N_10860,N_10285,N_10113);
and U10861 (N_10861,N_10458,N_10212);
nor U10862 (N_10862,N_10181,N_10149);
or U10863 (N_10863,N_10011,N_10323);
nor U10864 (N_10864,N_10333,N_10424);
xor U10865 (N_10865,N_10016,N_10463);
and U10866 (N_10866,N_10219,N_10161);
or U10867 (N_10867,N_10491,N_10173);
xor U10868 (N_10868,N_10268,N_10216);
or U10869 (N_10869,N_10111,N_10324);
and U10870 (N_10870,N_10397,N_10047);
or U10871 (N_10871,N_10036,N_10281);
xor U10872 (N_10872,N_10129,N_10217);
or U10873 (N_10873,N_10073,N_10214);
nor U10874 (N_10874,N_10442,N_10473);
xnor U10875 (N_10875,N_10232,N_10348);
or U10876 (N_10876,N_10332,N_10189);
xor U10877 (N_10877,N_10105,N_10437);
nand U10878 (N_10878,N_10140,N_10284);
nor U10879 (N_10879,N_10437,N_10381);
and U10880 (N_10880,N_10109,N_10221);
nand U10881 (N_10881,N_10101,N_10286);
nor U10882 (N_10882,N_10023,N_10091);
and U10883 (N_10883,N_10431,N_10065);
and U10884 (N_10884,N_10420,N_10085);
or U10885 (N_10885,N_10248,N_10490);
or U10886 (N_10886,N_10290,N_10484);
or U10887 (N_10887,N_10030,N_10064);
or U10888 (N_10888,N_10188,N_10055);
nor U10889 (N_10889,N_10297,N_10256);
nor U10890 (N_10890,N_10204,N_10337);
and U10891 (N_10891,N_10100,N_10451);
xor U10892 (N_10892,N_10026,N_10372);
nand U10893 (N_10893,N_10176,N_10181);
and U10894 (N_10894,N_10308,N_10122);
or U10895 (N_10895,N_10021,N_10026);
nor U10896 (N_10896,N_10356,N_10364);
or U10897 (N_10897,N_10283,N_10315);
nand U10898 (N_10898,N_10090,N_10429);
nand U10899 (N_10899,N_10317,N_10136);
and U10900 (N_10900,N_10339,N_10022);
or U10901 (N_10901,N_10457,N_10334);
and U10902 (N_10902,N_10023,N_10031);
nand U10903 (N_10903,N_10264,N_10358);
xor U10904 (N_10904,N_10076,N_10103);
xor U10905 (N_10905,N_10491,N_10269);
or U10906 (N_10906,N_10051,N_10245);
nor U10907 (N_10907,N_10334,N_10138);
or U10908 (N_10908,N_10139,N_10426);
nand U10909 (N_10909,N_10453,N_10098);
or U10910 (N_10910,N_10405,N_10495);
or U10911 (N_10911,N_10100,N_10083);
and U10912 (N_10912,N_10376,N_10400);
nand U10913 (N_10913,N_10027,N_10223);
nor U10914 (N_10914,N_10234,N_10119);
or U10915 (N_10915,N_10269,N_10148);
nor U10916 (N_10916,N_10383,N_10486);
xnor U10917 (N_10917,N_10238,N_10227);
or U10918 (N_10918,N_10357,N_10089);
nand U10919 (N_10919,N_10437,N_10460);
and U10920 (N_10920,N_10249,N_10182);
or U10921 (N_10921,N_10454,N_10375);
and U10922 (N_10922,N_10491,N_10287);
nor U10923 (N_10923,N_10019,N_10240);
nand U10924 (N_10924,N_10367,N_10206);
nand U10925 (N_10925,N_10448,N_10106);
xor U10926 (N_10926,N_10106,N_10258);
nor U10927 (N_10927,N_10450,N_10222);
and U10928 (N_10928,N_10363,N_10489);
or U10929 (N_10929,N_10151,N_10113);
nand U10930 (N_10930,N_10443,N_10396);
or U10931 (N_10931,N_10292,N_10093);
or U10932 (N_10932,N_10499,N_10332);
xor U10933 (N_10933,N_10038,N_10004);
xor U10934 (N_10934,N_10325,N_10204);
nand U10935 (N_10935,N_10445,N_10185);
xor U10936 (N_10936,N_10240,N_10009);
nand U10937 (N_10937,N_10208,N_10244);
xnor U10938 (N_10938,N_10041,N_10006);
nand U10939 (N_10939,N_10163,N_10437);
xnor U10940 (N_10940,N_10489,N_10047);
or U10941 (N_10941,N_10386,N_10428);
and U10942 (N_10942,N_10253,N_10256);
and U10943 (N_10943,N_10322,N_10191);
nand U10944 (N_10944,N_10404,N_10059);
and U10945 (N_10945,N_10186,N_10190);
or U10946 (N_10946,N_10405,N_10324);
and U10947 (N_10947,N_10429,N_10194);
nand U10948 (N_10948,N_10401,N_10419);
and U10949 (N_10949,N_10016,N_10068);
nand U10950 (N_10950,N_10259,N_10279);
nand U10951 (N_10951,N_10422,N_10146);
nor U10952 (N_10952,N_10265,N_10415);
and U10953 (N_10953,N_10184,N_10122);
or U10954 (N_10954,N_10372,N_10230);
or U10955 (N_10955,N_10178,N_10027);
or U10956 (N_10956,N_10231,N_10117);
or U10957 (N_10957,N_10344,N_10172);
or U10958 (N_10958,N_10470,N_10135);
xnor U10959 (N_10959,N_10031,N_10064);
nor U10960 (N_10960,N_10231,N_10366);
nor U10961 (N_10961,N_10378,N_10388);
nor U10962 (N_10962,N_10382,N_10452);
xor U10963 (N_10963,N_10310,N_10211);
xnor U10964 (N_10964,N_10177,N_10382);
or U10965 (N_10965,N_10376,N_10366);
nor U10966 (N_10966,N_10173,N_10440);
or U10967 (N_10967,N_10287,N_10425);
or U10968 (N_10968,N_10242,N_10385);
xor U10969 (N_10969,N_10280,N_10205);
nor U10970 (N_10970,N_10050,N_10282);
or U10971 (N_10971,N_10321,N_10429);
nor U10972 (N_10972,N_10116,N_10351);
nand U10973 (N_10973,N_10387,N_10122);
nand U10974 (N_10974,N_10349,N_10241);
nor U10975 (N_10975,N_10378,N_10396);
nor U10976 (N_10976,N_10231,N_10027);
nor U10977 (N_10977,N_10063,N_10347);
nor U10978 (N_10978,N_10329,N_10220);
and U10979 (N_10979,N_10281,N_10309);
and U10980 (N_10980,N_10243,N_10463);
nand U10981 (N_10981,N_10374,N_10165);
xor U10982 (N_10982,N_10384,N_10254);
nand U10983 (N_10983,N_10013,N_10258);
and U10984 (N_10984,N_10039,N_10478);
nand U10985 (N_10985,N_10115,N_10308);
and U10986 (N_10986,N_10193,N_10207);
xor U10987 (N_10987,N_10099,N_10179);
nand U10988 (N_10988,N_10436,N_10101);
and U10989 (N_10989,N_10006,N_10055);
nand U10990 (N_10990,N_10077,N_10028);
or U10991 (N_10991,N_10174,N_10114);
and U10992 (N_10992,N_10365,N_10077);
nand U10993 (N_10993,N_10476,N_10435);
xor U10994 (N_10994,N_10111,N_10314);
nor U10995 (N_10995,N_10184,N_10037);
or U10996 (N_10996,N_10410,N_10190);
nor U10997 (N_10997,N_10373,N_10252);
or U10998 (N_10998,N_10481,N_10026);
xor U10999 (N_10999,N_10155,N_10279);
xor U11000 (N_11000,N_10914,N_10567);
nor U11001 (N_11001,N_10563,N_10819);
or U11002 (N_11002,N_10513,N_10882);
and U11003 (N_11003,N_10821,N_10859);
and U11004 (N_11004,N_10793,N_10924);
nor U11005 (N_11005,N_10542,N_10686);
and U11006 (N_11006,N_10708,N_10776);
or U11007 (N_11007,N_10875,N_10811);
nand U11008 (N_11008,N_10705,N_10549);
and U11009 (N_11009,N_10537,N_10618);
nor U11010 (N_11010,N_10520,N_10511);
and U11011 (N_11011,N_10727,N_10990);
or U11012 (N_11012,N_10646,N_10901);
xor U11013 (N_11013,N_10608,N_10641);
nand U11014 (N_11014,N_10980,N_10896);
nand U11015 (N_11015,N_10621,N_10586);
nand U11016 (N_11016,N_10566,N_10868);
nand U11017 (N_11017,N_10570,N_10704);
nand U11018 (N_11018,N_10554,N_10594);
nor U11019 (N_11019,N_10956,N_10802);
and U11020 (N_11020,N_10611,N_10879);
and U11021 (N_11021,N_10625,N_10992);
and U11022 (N_11022,N_10562,N_10989);
xnor U11023 (N_11023,N_10753,N_10838);
xnor U11024 (N_11024,N_10984,N_10536);
and U11025 (N_11025,N_10770,N_10512);
nand U11026 (N_11026,N_10858,N_10905);
xnor U11027 (N_11027,N_10779,N_10650);
or U11028 (N_11028,N_10736,N_10794);
or U11029 (N_11029,N_10660,N_10789);
xor U11030 (N_11030,N_10517,N_10579);
or U11031 (N_11031,N_10503,N_10800);
and U11032 (N_11032,N_10857,N_10693);
or U11033 (N_11033,N_10718,N_10685);
nand U11034 (N_11034,N_10750,N_10778);
nand U11035 (N_11035,N_10599,N_10837);
xnor U11036 (N_11036,N_10583,N_10535);
xor U11037 (N_11037,N_10902,N_10762);
xor U11038 (N_11038,N_10795,N_10595);
and U11039 (N_11039,N_10523,N_10604);
or U11040 (N_11040,N_10585,N_10780);
or U11041 (N_11041,N_10756,N_10767);
nand U11042 (N_11042,N_10737,N_10950);
nor U11043 (N_11043,N_10827,N_10856);
xor U11044 (N_11044,N_10831,N_10713);
nand U11045 (N_11045,N_10777,N_10803);
and U11046 (N_11046,N_10926,N_10832);
nand U11047 (N_11047,N_10597,N_10741);
or U11048 (N_11048,N_10522,N_10689);
nor U11049 (N_11049,N_10936,N_10572);
xor U11050 (N_11050,N_10654,N_10612);
nor U11051 (N_11051,N_10904,N_10974);
or U11052 (N_11052,N_10889,N_10560);
nand U11053 (N_11053,N_10662,N_10561);
nand U11054 (N_11054,N_10573,N_10675);
nand U11055 (N_11055,N_10665,N_10640);
nor U11056 (N_11056,N_10518,N_10853);
and U11057 (N_11057,N_10922,N_10574);
xor U11058 (N_11058,N_10995,N_10748);
xnor U11059 (N_11059,N_10801,N_10623);
nand U11060 (N_11060,N_10528,N_10946);
nand U11061 (N_11061,N_10769,N_10526);
nor U11062 (N_11062,N_10601,N_10939);
nor U11063 (N_11063,N_10920,N_10697);
nor U11064 (N_11064,N_10724,N_10758);
nor U11065 (N_11065,N_10836,N_10867);
nand U11066 (N_11066,N_10533,N_10725);
nand U11067 (N_11067,N_10943,N_10696);
or U11068 (N_11068,N_10672,N_10988);
or U11069 (N_11069,N_10979,N_10861);
xor U11070 (N_11070,N_10516,N_10728);
nand U11071 (N_11071,N_10527,N_10541);
nand U11072 (N_11072,N_10847,N_10596);
xor U11073 (N_11073,N_10829,N_10531);
xor U11074 (N_11074,N_10695,N_10808);
nor U11075 (N_11075,N_10627,N_10547);
or U11076 (N_11076,N_10578,N_10783);
nand U11077 (N_11077,N_10830,N_10940);
xor U11078 (N_11078,N_10912,N_10701);
and U11079 (N_11079,N_10746,N_10894);
and U11080 (N_11080,N_10954,N_10655);
or U11081 (N_11081,N_10991,N_10900);
and U11082 (N_11082,N_10941,N_10949);
or U11083 (N_11083,N_10843,N_10993);
nand U11084 (N_11084,N_10898,N_10834);
or U11085 (N_11085,N_10809,N_10813);
nand U11086 (N_11086,N_10961,N_10607);
and U11087 (N_11087,N_10617,N_10507);
nand U11088 (N_11088,N_10973,N_10545);
nor U11089 (N_11089,N_10822,N_10917);
nand U11090 (N_11090,N_10791,N_10669);
and U11091 (N_11091,N_10616,N_10505);
nor U11092 (N_11092,N_10626,N_10878);
nor U11093 (N_11093,N_10987,N_10909);
nor U11094 (N_11094,N_10738,N_10722);
nand U11095 (N_11095,N_10732,N_10812);
or U11096 (N_11096,N_10622,N_10884);
and U11097 (N_11097,N_10862,N_10935);
or U11098 (N_11098,N_10807,N_10919);
nand U11099 (N_11099,N_10761,N_10958);
nor U11100 (N_11100,N_10624,N_10575);
or U11101 (N_11101,N_10872,N_10927);
nand U11102 (N_11102,N_10947,N_10698);
nand U11103 (N_11103,N_10735,N_10815);
xor U11104 (N_11104,N_10850,N_10907);
nand U11105 (N_11105,N_10757,N_10630);
nor U11106 (N_11106,N_10848,N_10967);
nor U11107 (N_11107,N_10886,N_10707);
or U11108 (N_11108,N_10982,N_10629);
and U11109 (N_11109,N_10681,N_10752);
xnor U11110 (N_11110,N_10983,N_10667);
xnor U11111 (N_11111,N_10582,N_10797);
and U11112 (N_11112,N_10703,N_10895);
and U11113 (N_11113,N_10508,N_10885);
nor U11114 (N_11114,N_10818,N_10814);
nand U11115 (N_11115,N_10500,N_10682);
nand U11116 (N_11116,N_10883,N_10931);
and U11117 (N_11117,N_10619,N_10871);
and U11118 (N_11118,N_10690,N_10564);
and U11119 (N_11119,N_10828,N_10955);
nor U11120 (N_11120,N_10798,N_10816);
nand U11121 (N_11121,N_10953,N_10580);
nor U11122 (N_11122,N_10606,N_10592);
xor U11123 (N_11123,N_10544,N_10986);
and U11124 (N_11124,N_10839,N_10951);
or U11125 (N_11125,N_10817,N_10581);
and U11126 (N_11126,N_10530,N_10659);
or U11127 (N_11127,N_10602,N_10893);
xnor U11128 (N_11128,N_10833,N_10658);
and U11129 (N_11129,N_10873,N_10589);
nor U11130 (N_11130,N_10740,N_10504);
nor U11131 (N_11131,N_10842,N_10768);
xnor U11132 (N_11132,N_10965,N_10845);
nand U11133 (N_11133,N_10666,N_10913);
nor U11134 (N_11134,N_10652,N_10598);
or U11135 (N_11135,N_10805,N_10790);
nor U11136 (N_11136,N_10590,N_10540);
or U11137 (N_11137,N_10944,N_10892);
nand U11138 (N_11138,N_10674,N_10806);
or U11139 (N_11139,N_10663,N_10639);
nor U11140 (N_11140,N_10706,N_10749);
xor U11141 (N_11141,N_10880,N_10632);
nor U11142 (N_11142,N_10835,N_10866);
xor U11143 (N_11143,N_10971,N_10964);
nor U11144 (N_11144,N_10937,N_10730);
xnor U11145 (N_11145,N_10911,N_10678);
and U11146 (N_11146,N_10636,N_10772);
xor U11147 (N_11147,N_10825,N_10899);
or U11148 (N_11148,N_10864,N_10710);
xnor U11149 (N_11149,N_10918,N_10890);
nor U11150 (N_11150,N_10925,N_10714);
and U11151 (N_11151,N_10700,N_10569);
or U11152 (N_11152,N_10521,N_10635);
or U11153 (N_11153,N_10824,N_10942);
nand U11154 (N_11154,N_10647,N_10774);
xor U11155 (N_11155,N_10796,N_10820);
xnor U11156 (N_11156,N_10933,N_10763);
nor U11157 (N_11157,N_10643,N_10903);
or U11158 (N_11158,N_10605,N_10711);
nor U11159 (N_11159,N_10677,N_10782);
and U11160 (N_11160,N_10760,N_10874);
xor U11161 (N_11161,N_10865,N_10870);
xnor U11162 (N_11162,N_10717,N_10787);
nor U11163 (N_11163,N_10534,N_10576);
xor U11164 (N_11164,N_10648,N_10957);
xnor U11165 (N_11165,N_10614,N_10519);
or U11166 (N_11166,N_10960,N_10719);
or U11167 (N_11167,N_10915,N_10591);
and U11168 (N_11168,N_10747,N_10551);
nor U11169 (N_11169,N_10600,N_10860);
and U11170 (N_11170,N_10754,N_10637);
or U11171 (N_11171,N_10593,N_10966);
nand U11172 (N_11172,N_10555,N_10588);
nor U11173 (N_11173,N_10683,N_10680);
xor U11174 (N_11174,N_10609,N_10876);
or U11175 (N_11175,N_10733,N_10745);
and U11176 (N_11176,N_10969,N_10620);
and U11177 (N_11177,N_10928,N_10502);
nand U11178 (N_11178,N_10851,N_10649);
and U11179 (N_11179,N_10906,N_10577);
nor U11180 (N_11180,N_10692,N_10981);
nand U11181 (N_11181,N_10657,N_10962);
xor U11182 (N_11182,N_10863,N_10932);
nor U11183 (N_11183,N_10877,N_10726);
nor U11184 (N_11184,N_10846,N_10997);
xnor U11185 (N_11185,N_10615,N_10720);
nor U11186 (N_11186,N_10687,N_10552);
and U11187 (N_11187,N_10653,N_10804);
and U11188 (N_11188,N_10688,N_10977);
nor U11189 (N_11189,N_10702,N_10952);
nor U11190 (N_11190,N_10849,N_10673);
or U11191 (N_11191,N_10510,N_10785);
xnor U11192 (N_11192,N_10742,N_10501);
nand U11193 (N_11193,N_10633,N_10645);
nor U11194 (N_11194,N_10841,N_10529);
xnor U11195 (N_11195,N_10691,N_10996);
nor U11196 (N_11196,N_10610,N_10603);
and U11197 (N_11197,N_10644,N_10679);
nor U11198 (N_11198,N_10810,N_10999);
xor U11199 (N_11199,N_10945,N_10743);
nor U11200 (N_11200,N_10712,N_10676);
or U11201 (N_11201,N_10799,N_10731);
nand U11202 (N_11202,N_10565,N_10921);
and U11203 (N_11203,N_10887,N_10908);
xnor U11204 (N_11204,N_10784,N_10998);
nand U11205 (N_11205,N_10923,N_10509);
xor U11206 (N_11206,N_10729,N_10525);
nor U11207 (N_11207,N_10938,N_10515);
nor U11208 (N_11208,N_10694,N_10584);
xnor U11209 (N_11209,N_10963,N_10897);
xnor U11210 (N_11210,N_10959,N_10930);
nand U11211 (N_11211,N_10631,N_10855);
nor U11212 (N_11212,N_10709,N_10514);
and U11213 (N_11213,N_10765,N_10755);
nand U11214 (N_11214,N_10587,N_10642);
nor U11215 (N_11215,N_10715,N_10670);
and U11216 (N_11216,N_10716,N_10881);
nor U11217 (N_11217,N_10869,N_10852);
nand U11218 (N_11218,N_10888,N_10985);
nor U11219 (N_11219,N_10557,N_10910);
nor U11220 (N_11220,N_10568,N_10543);
nand U11221 (N_11221,N_10550,N_10788);
nand U11222 (N_11222,N_10546,N_10751);
and U11223 (N_11223,N_10628,N_10775);
xor U11224 (N_11224,N_10723,N_10766);
nand U11225 (N_11225,N_10978,N_10972);
xnor U11226 (N_11226,N_10538,N_10968);
and U11227 (N_11227,N_10559,N_10840);
nor U11228 (N_11228,N_10651,N_10792);
nand U11229 (N_11229,N_10571,N_10759);
nor U11230 (N_11230,N_10823,N_10854);
nor U11231 (N_11231,N_10556,N_10773);
and U11232 (N_11232,N_10970,N_10668);
xnor U11233 (N_11233,N_10656,N_10634);
or U11234 (N_11234,N_10781,N_10661);
or U11235 (N_11235,N_10976,N_10539);
and U11236 (N_11236,N_10975,N_10934);
and U11237 (N_11237,N_10553,N_10524);
and U11238 (N_11238,N_10734,N_10844);
and U11239 (N_11239,N_10744,N_10506);
xnor U11240 (N_11240,N_10948,N_10721);
xnor U11241 (N_11241,N_10994,N_10664);
nand U11242 (N_11242,N_10699,N_10891);
nand U11243 (N_11243,N_10826,N_10684);
and U11244 (N_11244,N_10638,N_10771);
nand U11245 (N_11245,N_10929,N_10558);
or U11246 (N_11246,N_10764,N_10613);
xor U11247 (N_11247,N_10739,N_10671);
and U11248 (N_11248,N_10548,N_10786);
or U11249 (N_11249,N_10916,N_10532);
or U11250 (N_11250,N_10857,N_10974);
nor U11251 (N_11251,N_10831,N_10501);
nand U11252 (N_11252,N_10920,N_10713);
nor U11253 (N_11253,N_10756,N_10606);
and U11254 (N_11254,N_10735,N_10916);
xor U11255 (N_11255,N_10971,N_10926);
and U11256 (N_11256,N_10585,N_10733);
and U11257 (N_11257,N_10970,N_10692);
xor U11258 (N_11258,N_10863,N_10836);
nand U11259 (N_11259,N_10972,N_10500);
nand U11260 (N_11260,N_10582,N_10597);
and U11261 (N_11261,N_10821,N_10525);
nand U11262 (N_11262,N_10985,N_10959);
or U11263 (N_11263,N_10543,N_10610);
and U11264 (N_11264,N_10901,N_10876);
or U11265 (N_11265,N_10608,N_10519);
and U11266 (N_11266,N_10906,N_10760);
and U11267 (N_11267,N_10700,N_10501);
and U11268 (N_11268,N_10587,N_10807);
nand U11269 (N_11269,N_10932,N_10994);
xnor U11270 (N_11270,N_10841,N_10523);
xor U11271 (N_11271,N_10552,N_10786);
nand U11272 (N_11272,N_10667,N_10600);
xnor U11273 (N_11273,N_10772,N_10714);
or U11274 (N_11274,N_10911,N_10833);
nand U11275 (N_11275,N_10846,N_10683);
and U11276 (N_11276,N_10621,N_10598);
nor U11277 (N_11277,N_10899,N_10944);
or U11278 (N_11278,N_10732,N_10678);
and U11279 (N_11279,N_10676,N_10984);
xor U11280 (N_11280,N_10539,N_10575);
or U11281 (N_11281,N_10571,N_10613);
nor U11282 (N_11282,N_10731,N_10982);
or U11283 (N_11283,N_10910,N_10913);
nor U11284 (N_11284,N_10729,N_10514);
nor U11285 (N_11285,N_10745,N_10952);
or U11286 (N_11286,N_10891,N_10613);
nor U11287 (N_11287,N_10987,N_10570);
xnor U11288 (N_11288,N_10640,N_10692);
xnor U11289 (N_11289,N_10658,N_10805);
xnor U11290 (N_11290,N_10778,N_10741);
nand U11291 (N_11291,N_10622,N_10547);
nand U11292 (N_11292,N_10831,N_10615);
xnor U11293 (N_11293,N_10667,N_10510);
nand U11294 (N_11294,N_10832,N_10517);
nand U11295 (N_11295,N_10542,N_10584);
nand U11296 (N_11296,N_10968,N_10686);
or U11297 (N_11297,N_10621,N_10807);
nand U11298 (N_11298,N_10947,N_10646);
or U11299 (N_11299,N_10871,N_10837);
or U11300 (N_11300,N_10712,N_10962);
nor U11301 (N_11301,N_10808,N_10756);
and U11302 (N_11302,N_10936,N_10676);
nor U11303 (N_11303,N_10630,N_10900);
nor U11304 (N_11304,N_10830,N_10896);
xor U11305 (N_11305,N_10753,N_10936);
nor U11306 (N_11306,N_10922,N_10968);
or U11307 (N_11307,N_10947,N_10605);
nor U11308 (N_11308,N_10559,N_10541);
and U11309 (N_11309,N_10943,N_10563);
and U11310 (N_11310,N_10860,N_10605);
nor U11311 (N_11311,N_10908,N_10684);
nand U11312 (N_11312,N_10563,N_10685);
or U11313 (N_11313,N_10907,N_10723);
and U11314 (N_11314,N_10734,N_10681);
nor U11315 (N_11315,N_10678,N_10756);
nor U11316 (N_11316,N_10577,N_10946);
nor U11317 (N_11317,N_10618,N_10775);
nand U11318 (N_11318,N_10805,N_10539);
nand U11319 (N_11319,N_10513,N_10949);
nand U11320 (N_11320,N_10557,N_10958);
and U11321 (N_11321,N_10534,N_10809);
or U11322 (N_11322,N_10830,N_10867);
and U11323 (N_11323,N_10725,N_10658);
xnor U11324 (N_11324,N_10854,N_10638);
xor U11325 (N_11325,N_10729,N_10551);
nor U11326 (N_11326,N_10589,N_10904);
and U11327 (N_11327,N_10604,N_10521);
or U11328 (N_11328,N_10742,N_10843);
and U11329 (N_11329,N_10596,N_10544);
nand U11330 (N_11330,N_10618,N_10898);
or U11331 (N_11331,N_10970,N_10949);
and U11332 (N_11332,N_10558,N_10519);
and U11333 (N_11333,N_10698,N_10668);
nor U11334 (N_11334,N_10859,N_10593);
nor U11335 (N_11335,N_10679,N_10763);
and U11336 (N_11336,N_10949,N_10520);
nand U11337 (N_11337,N_10824,N_10807);
nor U11338 (N_11338,N_10500,N_10639);
xor U11339 (N_11339,N_10786,N_10893);
or U11340 (N_11340,N_10512,N_10767);
xnor U11341 (N_11341,N_10715,N_10806);
or U11342 (N_11342,N_10882,N_10945);
nand U11343 (N_11343,N_10985,N_10702);
nand U11344 (N_11344,N_10641,N_10675);
or U11345 (N_11345,N_10749,N_10978);
and U11346 (N_11346,N_10799,N_10592);
nand U11347 (N_11347,N_10555,N_10743);
and U11348 (N_11348,N_10945,N_10676);
or U11349 (N_11349,N_10528,N_10559);
nand U11350 (N_11350,N_10846,N_10970);
or U11351 (N_11351,N_10678,N_10709);
and U11352 (N_11352,N_10914,N_10850);
nand U11353 (N_11353,N_10678,N_10599);
nor U11354 (N_11354,N_10961,N_10710);
nand U11355 (N_11355,N_10720,N_10850);
xor U11356 (N_11356,N_10507,N_10675);
xor U11357 (N_11357,N_10569,N_10883);
and U11358 (N_11358,N_10964,N_10644);
nor U11359 (N_11359,N_10861,N_10980);
and U11360 (N_11360,N_10997,N_10646);
and U11361 (N_11361,N_10917,N_10812);
nor U11362 (N_11362,N_10728,N_10776);
nand U11363 (N_11363,N_10657,N_10697);
and U11364 (N_11364,N_10879,N_10638);
or U11365 (N_11365,N_10961,N_10855);
nor U11366 (N_11366,N_10582,N_10876);
nor U11367 (N_11367,N_10894,N_10880);
nand U11368 (N_11368,N_10833,N_10514);
and U11369 (N_11369,N_10823,N_10960);
or U11370 (N_11370,N_10524,N_10751);
nor U11371 (N_11371,N_10572,N_10679);
nor U11372 (N_11372,N_10705,N_10634);
or U11373 (N_11373,N_10936,N_10579);
nor U11374 (N_11374,N_10954,N_10713);
and U11375 (N_11375,N_10855,N_10680);
xnor U11376 (N_11376,N_10741,N_10726);
nand U11377 (N_11377,N_10942,N_10775);
nor U11378 (N_11378,N_10971,N_10540);
nor U11379 (N_11379,N_10623,N_10549);
or U11380 (N_11380,N_10542,N_10954);
nor U11381 (N_11381,N_10649,N_10827);
and U11382 (N_11382,N_10800,N_10808);
and U11383 (N_11383,N_10591,N_10660);
nor U11384 (N_11384,N_10504,N_10865);
and U11385 (N_11385,N_10597,N_10594);
nand U11386 (N_11386,N_10603,N_10598);
and U11387 (N_11387,N_10513,N_10716);
xnor U11388 (N_11388,N_10774,N_10607);
nand U11389 (N_11389,N_10594,N_10637);
nor U11390 (N_11390,N_10644,N_10618);
xnor U11391 (N_11391,N_10568,N_10793);
nor U11392 (N_11392,N_10679,N_10821);
nand U11393 (N_11393,N_10673,N_10953);
nor U11394 (N_11394,N_10940,N_10641);
xor U11395 (N_11395,N_10693,N_10870);
or U11396 (N_11396,N_10559,N_10866);
nand U11397 (N_11397,N_10863,N_10895);
nand U11398 (N_11398,N_10539,N_10641);
nand U11399 (N_11399,N_10759,N_10771);
nand U11400 (N_11400,N_10922,N_10957);
and U11401 (N_11401,N_10720,N_10739);
and U11402 (N_11402,N_10892,N_10700);
and U11403 (N_11403,N_10508,N_10571);
xnor U11404 (N_11404,N_10958,N_10984);
and U11405 (N_11405,N_10963,N_10752);
xor U11406 (N_11406,N_10519,N_10529);
nor U11407 (N_11407,N_10640,N_10951);
or U11408 (N_11408,N_10619,N_10706);
nor U11409 (N_11409,N_10909,N_10757);
xnor U11410 (N_11410,N_10890,N_10980);
or U11411 (N_11411,N_10749,N_10944);
or U11412 (N_11412,N_10791,N_10697);
and U11413 (N_11413,N_10799,N_10836);
nor U11414 (N_11414,N_10522,N_10573);
xnor U11415 (N_11415,N_10616,N_10664);
or U11416 (N_11416,N_10725,N_10578);
and U11417 (N_11417,N_10822,N_10991);
nor U11418 (N_11418,N_10913,N_10812);
nor U11419 (N_11419,N_10561,N_10987);
nor U11420 (N_11420,N_10785,N_10632);
xnor U11421 (N_11421,N_10761,N_10534);
nand U11422 (N_11422,N_10760,N_10911);
or U11423 (N_11423,N_10935,N_10834);
and U11424 (N_11424,N_10800,N_10683);
nor U11425 (N_11425,N_10907,N_10624);
or U11426 (N_11426,N_10972,N_10775);
and U11427 (N_11427,N_10852,N_10862);
and U11428 (N_11428,N_10961,N_10684);
nor U11429 (N_11429,N_10903,N_10987);
and U11430 (N_11430,N_10850,N_10902);
and U11431 (N_11431,N_10643,N_10763);
and U11432 (N_11432,N_10669,N_10865);
or U11433 (N_11433,N_10718,N_10763);
xnor U11434 (N_11434,N_10506,N_10562);
or U11435 (N_11435,N_10696,N_10972);
nor U11436 (N_11436,N_10921,N_10558);
and U11437 (N_11437,N_10970,N_10787);
and U11438 (N_11438,N_10932,N_10688);
nand U11439 (N_11439,N_10596,N_10705);
or U11440 (N_11440,N_10847,N_10595);
or U11441 (N_11441,N_10687,N_10996);
nor U11442 (N_11442,N_10906,N_10593);
and U11443 (N_11443,N_10731,N_10530);
and U11444 (N_11444,N_10680,N_10597);
and U11445 (N_11445,N_10614,N_10547);
nand U11446 (N_11446,N_10820,N_10937);
nand U11447 (N_11447,N_10830,N_10889);
nor U11448 (N_11448,N_10721,N_10937);
nand U11449 (N_11449,N_10608,N_10734);
xnor U11450 (N_11450,N_10566,N_10808);
and U11451 (N_11451,N_10665,N_10554);
and U11452 (N_11452,N_10978,N_10694);
and U11453 (N_11453,N_10905,N_10542);
nor U11454 (N_11454,N_10552,N_10767);
nand U11455 (N_11455,N_10628,N_10688);
nand U11456 (N_11456,N_10864,N_10610);
nor U11457 (N_11457,N_10779,N_10936);
or U11458 (N_11458,N_10837,N_10522);
nand U11459 (N_11459,N_10705,N_10663);
or U11460 (N_11460,N_10556,N_10885);
and U11461 (N_11461,N_10599,N_10727);
and U11462 (N_11462,N_10519,N_10692);
xor U11463 (N_11463,N_10799,N_10535);
xor U11464 (N_11464,N_10975,N_10726);
xor U11465 (N_11465,N_10870,N_10755);
nor U11466 (N_11466,N_10813,N_10829);
nor U11467 (N_11467,N_10557,N_10904);
nand U11468 (N_11468,N_10605,N_10616);
nor U11469 (N_11469,N_10816,N_10744);
and U11470 (N_11470,N_10709,N_10996);
and U11471 (N_11471,N_10629,N_10781);
nor U11472 (N_11472,N_10639,N_10521);
and U11473 (N_11473,N_10765,N_10697);
or U11474 (N_11474,N_10893,N_10772);
and U11475 (N_11475,N_10690,N_10647);
or U11476 (N_11476,N_10658,N_10943);
or U11477 (N_11477,N_10749,N_10958);
nor U11478 (N_11478,N_10522,N_10561);
nor U11479 (N_11479,N_10719,N_10851);
or U11480 (N_11480,N_10850,N_10554);
xor U11481 (N_11481,N_10549,N_10548);
nor U11482 (N_11482,N_10763,N_10886);
nor U11483 (N_11483,N_10803,N_10570);
nor U11484 (N_11484,N_10854,N_10994);
nand U11485 (N_11485,N_10600,N_10895);
nor U11486 (N_11486,N_10961,N_10871);
and U11487 (N_11487,N_10917,N_10891);
and U11488 (N_11488,N_10809,N_10559);
and U11489 (N_11489,N_10712,N_10711);
nand U11490 (N_11490,N_10502,N_10623);
or U11491 (N_11491,N_10740,N_10921);
nand U11492 (N_11492,N_10639,N_10984);
nor U11493 (N_11493,N_10950,N_10786);
nor U11494 (N_11494,N_10783,N_10797);
or U11495 (N_11495,N_10776,N_10525);
nor U11496 (N_11496,N_10915,N_10738);
xnor U11497 (N_11497,N_10781,N_10610);
and U11498 (N_11498,N_10780,N_10651);
xor U11499 (N_11499,N_10992,N_10556);
xnor U11500 (N_11500,N_11122,N_11447);
nand U11501 (N_11501,N_11465,N_11454);
xor U11502 (N_11502,N_11106,N_11479);
or U11503 (N_11503,N_11226,N_11087);
or U11504 (N_11504,N_11370,N_11260);
nor U11505 (N_11505,N_11333,N_11450);
or U11506 (N_11506,N_11012,N_11360);
or U11507 (N_11507,N_11064,N_11038);
xor U11508 (N_11508,N_11459,N_11267);
xor U11509 (N_11509,N_11388,N_11437);
nor U11510 (N_11510,N_11014,N_11468);
nand U11511 (N_11511,N_11434,N_11103);
nor U11512 (N_11512,N_11273,N_11149);
xor U11513 (N_11513,N_11111,N_11320);
and U11514 (N_11514,N_11299,N_11289);
nor U11515 (N_11515,N_11372,N_11290);
nand U11516 (N_11516,N_11195,N_11263);
nor U11517 (N_11517,N_11250,N_11209);
xnor U11518 (N_11518,N_11442,N_11377);
nand U11519 (N_11519,N_11379,N_11191);
and U11520 (N_11520,N_11008,N_11251);
and U11521 (N_11521,N_11252,N_11066);
xnor U11522 (N_11522,N_11295,N_11256);
xnor U11523 (N_11523,N_11239,N_11347);
or U11524 (N_11524,N_11194,N_11301);
or U11525 (N_11525,N_11444,N_11424);
xnor U11526 (N_11526,N_11351,N_11004);
nor U11527 (N_11527,N_11141,N_11349);
xor U11528 (N_11528,N_11027,N_11268);
or U11529 (N_11529,N_11018,N_11003);
nor U11530 (N_11530,N_11205,N_11086);
nor U11531 (N_11531,N_11146,N_11330);
or U11532 (N_11532,N_11096,N_11161);
or U11533 (N_11533,N_11002,N_11221);
nor U11534 (N_11534,N_11021,N_11053);
xor U11535 (N_11535,N_11387,N_11155);
nor U11536 (N_11536,N_11059,N_11190);
and U11537 (N_11537,N_11400,N_11361);
nand U11538 (N_11538,N_11325,N_11303);
and U11539 (N_11539,N_11030,N_11089);
nand U11540 (N_11540,N_11178,N_11117);
or U11541 (N_11541,N_11151,N_11298);
and U11542 (N_11542,N_11308,N_11331);
or U11543 (N_11543,N_11319,N_11133);
xor U11544 (N_11544,N_11156,N_11140);
and U11545 (N_11545,N_11382,N_11037);
nand U11546 (N_11546,N_11409,N_11475);
or U11547 (N_11547,N_11159,N_11040);
nor U11548 (N_11548,N_11310,N_11197);
xor U11549 (N_11549,N_11392,N_11481);
and U11550 (N_11550,N_11042,N_11296);
xnor U11551 (N_11551,N_11452,N_11085);
or U11552 (N_11552,N_11337,N_11408);
xor U11553 (N_11553,N_11274,N_11072);
nor U11554 (N_11554,N_11081,N_11000);
nand U11555 (N_11555,N_11160,N_11026);
nand U11556 (N_11556,N_11128,N_11054);
nor U11557 (N_11557,N_11150,N_11075);
xnor U11558 (N_11558,N_11234,N_11169);
nand U11559 (N_11559,N_11284,N_11316);
or U11560 (N_11560,N_11436,N_11184);
nand U11561 (N_11561,N_11098,N_11441);
nor U11562 (N_11562,N_11354,N_11300);
nand U11563 (N_11563,N_11204,N_11171);
nor U11564 (N_11564,N_11278,N_11246);
xor U11565 (N_11565,N_11068,N_11218);
nand U11566 (N_11566,N_11448,N_11243);
xor U11567 (N_11567,N_11463,N_11013);
nor U11568 (N_11568,N_11285,N_11126);
or U11569 (N_11569,N_11427,N_11244);
xor U11570 (N_11570,N_11217,N_11312);
xor U11571 (N_11571,N_11130,N_11374);
or U11572 (N_11572,N_11145,N_11074);
and U11573 (N_11573,N_11487,N_11367);
and U11574 (N_11574,N_11148,N_11462);
nand U11575 (N_11575,N_11152,N_11208);
or U11576 (N_11576,N_11467,N_11253);
and U11577 (N_11577,N_11005,N_11366);
xnor U11578 (N_11578,N_11426,N_11421);
and U11579 (N_11579,N_11491,N_11431);
or U11580 (N_11580,N_11332,N_11084);
xnor U11581 (N_11581,N_11136,N_11390);
or U11582 (N_11582,N_11201,N_11359);
nor U11583 (N_11583,N_11067,N_11286);
and U11584 (N_11584,N_11348,N_11439);
nor U11585 (N_11585,N_11193,N_11402);
and U11586 (N_11586,N_11214,N_11265);
nand U11587 (N_11587,N_11259,N_11153);
nand U11588 (N_11588,N_11093,N_11358);
xor U11589 (N_11589,N_11394,N_11187);
and U11590 (N_11590,N_11235,N_11416);
and U11591 (N_11591,N_11060,N_11464);
xnor U11592 (N_11592,N_11422,N_11488);
and U11593 (N_11593,N_11227,N_11174);
nand U11594 (N_11594,N_11228,N_11288);
nand U11595 (N_11595,N_11200,N_11199);
xnor U11596 (N_11596,N_11185,N_11485);
xor U11597 (N_11597,N_11183,N_11118);
and U11598 (N_11598,N_11025,N_11362);
xor U11599 (N_11599,N_11345,N_11119);
and U11600 (N_11600,N_11051,N_11034);
nand U11601 (N_11601,N_11486,N_11353);
and U11602 (N_11602,N_11469,N_11329);
or U11603 (N_11603,N_11473,N_11065);
nand U11604 (N_11604,N_11323,N_11180);
or U11605 (N_11605,N_11061,N_11283);
nor U11606 (N_11606,N_11062,N_11318);
and U11607 (N_11607,N_11079,N_11203);
or U11608 (N_11608,N_11466,N_11007);
and U11609 (N_11609,N_11045,N_11324);
nand U11610 (N_11610,N_11039,N_11429);
nor U11611 (N_11611,N_11175,N_11499);
nor U11612 (N_11612,N_11102,N_11438);
and U11613 (N_11613,N_11368,N_11369);
xor U11614 (N_11614,N_11346,N_11129);
or U11615 (N_11615,N_11032,N_11410);
and U11616 (N_11616,N_11154,N_11425);
and U11617 (N_11617,N_11317,N_11229);
xor U11618 (N_11618,N_11236,N_11188);
nor U11619 (N_11619,N_11046,N_11123);
nor U11620 (N_11620,N_11398,N_11456);
xor U11621 (N_11621,N_11498,N_11210);
and U11622 (N_11622,N_11406,N_11428);
or U11623 (N_11623,N_11326,N_11470);
xnor U11624 (N_11624,N_11177,N_11322);
or U11625 (N_11625,N_11321,N_11471);
xnor U11626 (N_11626,N_11272,N_11069);
and U11627 (N_11627,N_11137,N_11001);
nor U11628 (N_11628,N_11225,N_11385);
and U11629 (N_11629,N_11168,N_11440);
nand U11630 (N_11630,N_11076,N_11099);
nand U11631 (N_11631,N_11041,N_11355);
nor U11632 (N_11632,N_11092,N_11165);
nor U11633 (N_11633,N_11058,N_11248);
nor U11634 (N_11634,N_11457,N_11131);
xnor U11635 (N_11635,N_11478,N_11049);
xnor U11636 (N_11636,N_11472,N_11182);
or U11637 (N_11637,N_11413,N_11019);
xor U11638 (N_11638,N_11297,N_11024);
xnor U11639 (N_11639,N_11222,N_11373);
nor U11640 (N_11640,N_11423,N_11143);
and U11641 (N_11641,N_11121,N_11418);
or U11642 (N_11642,N_11474,N_11132);
nand U11643 (N_11643,N_11033,N_11455);
nand U11644 (N_11644,N_11264,N_11029);
nor U11645 (N_11645,N_11277,N_11052);
nor U11646 (N_11646,N_11271,N_11179);
nor U11647 (N_11647,N_11314,N_11022);
or U11648 (N_11648,N_11443,N_11449);
or U11649 (N_11649,N_11077,N_11309);
nand U11650 (N_11650,N_11224,N_11230);
nor U11651 (N_11651,N_11166,N_11335);
nor U11652 (N_11652,N_11281,N_11125);
or U11653 (N_11653,N_11202,N_11138);
xor U11654 (N_11654,N_11010,N_11057);
nand U11655 (N_11655,N_11453,N_11395);
nand U11656 (N_11656,N_11006,N_11334);
and U11657 (N_11657,N_11196,N_11080);
xnor U11658 (N_11658,N_11480,N_11241);
or U11659 (N_11659,N_11198,N_11167);
nor U11660 (N_11660,N_11280,N_11186);
xor U11661 (N_11661,N_11071,N_11258);
or U11662 (N_11662,N_11483,N_11381);
or U11663 (N_11663,N_11489,N_11164);
xor U11664 (N_11664,N_11477,N_11494);
or U11665 (N_11665,N_11420,N_11056);
nor U11666 (N_11666,N_11430,N_11015);
or U11667 (N_11667,N_11343,N_11375);
or U11668 (N_11668,N_11232,N_11115);
nand U11669 (N_11669,N_11233,N_11091);
or U11670 (N_11670,N_11484,N_11476);
nor U11671 (N_11671,N_11411,N_11100);
nor U11672 (N_11672,N_11294,N_11432);
nand U11673 (N_11673,N_11350,N_11142);
or U11674 (N_11674,N_11238,N_11393);
and U11675 (N_11675,N_11257,N_11082);
or U11676 (N_11676,N_11386,N_11269);
xnor U11677 (N_11677,N_11176,N_11108);
or U11678 (N_11678,N_11247,N_11352);
nor U11679 (N_11679,N_11254,N_11276);
and U11680 (N_11680,N_11011,N_11113);
xor U11681 (N_11681,N_11356,N_11212);
and U11682 (N_11682,N_11127,N_11105);
nand U11683 (N_11683,N_11088,N_11031);
and U11684 (N_11684,N_11163,N_11050);
and U11685 (N_11685,N_11495,N_11357);
nor U11686 (N_11686,N_11219,N_11028);
and U11687 (N_11687,N_11490,N_11315);
nand U11688 (N_11688,N_11407,N_11134);
xnor U11689 (N_11689,N_11223,N_11094);
or U11690 (N_11690,N_11399,N_11492);
nand U11691 (N_11691,N_11365,N_11497);
xor U11692 (N_11692,N_11192,N_11482);
xnor U11693 (N_11693,N_11270,N_11451);
nor U11694 (N_11694,N_11139,N_11173);
nand U11695 (N_11695,N_11339,N_11336);
xor U11696 (N_11696,N_11090,N_11097);
xnor U11697 (N_11697,N_11240,N_11048);
nand U11698 (N_11698,N_11404,N_11162);
nor U11699 (N_11699,N_11158,N_11433);
xor U11700 (N_11700,N_11157,N_11396);
nor U11701 (N_11701,N_11435,N_11047);
nand U11702 (N_11702,N_11083,N_11135);
and U11703 (N_11703,N_11262,N_11405);
nand U11704 (N_11704,N_11364,N_11237);
nor U11705 (N_11705,N_11242,N_11327);
nand U11706 (N_11706,N_11419,N_11101);
nand U11707 (N_11707,N_11383,N_11311);
nor U11708 (N_11708,N_11304,N_11144);
xnor U11709 (N_11709,N_11461,N_11170);
or U11710 (N_11710,N_11206,N_11109);
nor U11711 (N_11711,N_11384,N_11120);
or U11712 (N_11712,N_11095,N_11389);
and U11713 (N_11713,N_11016,N_11172);
and U11714 (N_11714,N_11044,N_11104);
or U11715 (N_11715,N_11255,N_11009);
nand U11716 (N_11716,N_11220,N_11376);
xor U11717 (N_11717,N_11073,N_11207);
nor U11718 (N_11718,N_11302,N_11292);
and U11719 (N_11719,N_11403,N_11445);
or U11720 (N_11720,N_11305,N_11231);
or U11721 (N_11721,N_11211,N_11078);
nand U11722 (N_11722,N_11110,N_11306);
nor U11723 (N_11723,N_11342,N_11415);
xor U11724 (N_11724,N_11460,N_11189);
nor U11725 (N_11725,N_11055,N_11293);
or U11726 (N_11726,N_11341,N_11291);
and U11727 (N_11727,N_11215,N_11401);
xor U11728 (N_11728,N_11391,N_11261);
or U11729 (N_11729,N_11279,N_11338);
nor U11730 (N_11730,N_11063,N_11344);
nand U11731 (N_11731,N_11070,N_11412);
xor U11732 (N_11732,N_11245,N_11147);
or U11733 (N_11733,N_11446,N_11124);
xor U11734 (N_11734,N_11036,N_11378);
and U11735 (N_11735,N_11043,N_11493);
xnor U11736 (N_11736,N_11371,N_11107);
or U11737 (N_11737,N_11213,N_11287);
or U11738 (N_11738,N_11112,N_11282);
or U11739 (N_11739,N_11020,N_11017);
xnor U11740 (N_11740,N_11340,N_11249);
nand U11741 (N_11741,N_11458,N_11380);
nor U11742 (N_11742,N_11266,N_11307);
and U11743 (N_11743,N_11114,N_11216);
and U11744 (N_11744,N_11023,N_11116);
xor U11745 (N_11745,N_11035,N_11328);
nor U11746 (N_11746,N_11397,N_11275);
and U11747 (N_11747,N_11181,N_11417);
nand U11748 (N_11748,N_11496,N_11414);
nand U11749 (N_11749,N_11363,N_11313);
and U11750 (N_11750,N_11441,N_11355);
nand U11751 (N_11751,N_11008,N_11252);
and U11752 (N_11752,N_11235,N_11392);
xnor U11753 (N_11753,N_11173,N_11436);
and U11754 (N_11754,N_11262,N_11162);
and U11755 (N_11755,N_11168,N_11219);
and U11756 (N_11756,N_11346,N_11021);
and U11757 (N_11757,N_11426,N_11270);
nor U11758 (N_11758,N_11165,N_11375);
and U11759 (N_11759,N_11080,N_11212);
nand U11760 (N_11760,N_11021,N_11078);
nand U11761 (N_11761,N_11007,N_11057);
xor U11762 (N_11762,N_11015,N_11422);
nor U11763 (N_11763,N_11218,N_11176);
or U11764 (N_11764,N_11162,N_11325);
and U11765 (N_11765,N_11094,N_11304);
nor U11766 (N_11766,N_11491,N_11306);
nor U11767 (N_11767,N_11241,N_11303);
xnor U11768 (N_11768,N_11154,N_11164);
or U11769 (N_11769,N_11491,N_11069);
nand U11770 (N_11770,N_11121,N_11228);
nand U11771 (N_11771,N_11159,N_11288);
xor U11772 (N_11772,N_11212,N_11475);
nor U11773 (N_11773,N_11178,N_11273);
or U11774 (N_11774,N_11288,N_11087);
and U11775 (N_11775,N_11429,N_11096);
or U11776 (N_11776,N_11307,N_11148);
xor U11777 (N_11777,N_11475,N_11336);
xor U11778 (N_11778,N_11402,N_11051);
xnor U11779 (N_11779,N_11202,N_11025);
xor U11780 (N_11780,N_11335,N_11226);
xnor U11781 (N_11781,N_11256,N_11292);
and U11782 (N_11782,N_11382,N_11090);
and U11783 (N_11783,N_11362,N_11115);
and U11784 (N_11784,N_11287,N_11170);
xor U11785 (N_11785,N_11376,N_11402);
and U11786 (N_11786,N_11023,N_11105);
and U11787 (N_11787,N_11257,N_11390);
and U11788 (N_11788,N_11331,N_11166);
xnor U11789 (N_11789,N_11024,N_11319);
nand U11790 (N_11790,N_11307,N_11144);
or U11791 (N_11791,N_11127,N_11352);
xnor U11792 (N_11792,N_11034,N_11430);
nand U11793 (N_11793,N_11402,N_11334);
nand U11794 (N_11794,N_11144,N_11080);
xnor U11795 (N_11795,N_11129,N_11091);
nand U11796 (N_11796,N_11152,N_11289);
and U11797 (N_11797,N_11444,N_11003);
nand U11798 (N_11798,N_11158,N_11301);
xnor U11799 (N_11799,N_11365,N_11386);
and U11800 (N_11800,N_11487,N_11325);
nor U11801 (N_11801,N_11489,N_11317);
and U11802 (N_11802,N_11371,N_11064);
nor U11803 (N_11803,N_11377,N_11099);
nand U11804 (N_11804,N_11094,N_11444);
and U11805 (N_11805,N_11185,N_11494);
and U11806 (N_11806,N_11333,N_11331);
xor U11807 (N_11807,N_11379,N_11371);
or U11808 (N_11808,N_11241,N_11052);
nor U11809 (N_11809,N_11435,N_11275);
nand U11810 (N_11810,N_11089,N_11464);
nand U11811 (N_11811,N_11306,N_11330);
nor U11812 (N_11812,N_11223,N_11113);
xor U11813 (N_11813,N_11213,N_11197);
and U11814 (N_11814,N_11011,N_11109);
or U11815 (N_11815,N_11028,N_11178);
nor U11816 (N_11816,N_11039,N_11466);
and U11817 (N_11817,N_11458,N_11247);
nor U11818 (N_11818,N_11326,N_11284);
xor U11819 (N_11819,N_11122,N_11024);
nand U11820 (N_11820,N_11185,N_11135);
nand U11821 (N_11821,N_11304,N_11275);
and U11822 (N_11822,N_11342,N_11300);
and U11823 (N_11823,N_11005,N_11375);
nor U11824 (N_11824,N_11071,N_11478);
nand U11825 (N_11825,N_11173,N_11468);
or U11826 (N_11826,N_11244,N_11003);
and U11827 (N_11827,N_11253,N_11453);
and U11828 (N_11828,N_11205,N_11264);
or U11829 (N_11829,N_11088,N_11015);
or U11830 (N_11830,N_11458,N_11306);
nand U11831 (N_11831,N_11253,N_11040);
xnor U11832 (N_11832,N_11461,N_11496);
and U11833 (N_11833,N_11015,N_11249);
and U11834 (N_11834,N_11334,N_11288);
and U11835 (N_11835,N_11292,N_11480);
nor U11836 (N_11836,N_11137,N_11318);
or U11837 (N_11837,N_11451,N_11398);
xor U11838 (N_11838,N_11281,N_11043);
xor U11839 (N_11839,N_11004,N_11173);
nor U11840 (N_11840,N_11177,N_11108);
nor U11841 (N_11841,N_11054,N_11326);
nor U11842 (N_11842,N_11330,N_11433);
or U11843 (N_11843,N_11435,N_11405);
xor U11844 (N_11844,N_11391,N_11029);
xor U11845 (N_11845,N_11416,N_11064);
nor U11846 (N_11846,N_11058,N_11362);
and U11847 (N_11847,N_11438,N_11012);
nor U11848 (N_11848,N_11097,N_11499);
nand U11849 (N_11849,N_11071,N_11170);
or U11850 (N_11850,N_11478,N_11457);
nand U11851 (N_11851,N_11480,N_11133);
or U11852 (N_11852,N_11147,N_11170);
nor U11853 (N_11853,N_11015,N_11315);
nor U11854 (N_11854,N_11454,N_11389);
nand U11855 (N_11855,N_11225,N_11056);
and U11856 (N_11856,N_11185,N_11448);
nor U11857 (N_11857,N_11066,N_11439);
and U11858 (N_11858,N_11304,N_11375);
and U11859 (N_11859,N_11358,N_11021);
xnor U11860 (N_11860,N_11273,N_11455);
and U11861 (N_11861,N_11458,N_11291);
and U11862 (N_11862,N_11405,N_11243);
xor U11863 (N_11863,N_11425,N_11118);
nor U11864 (N_11864,N_11037,N_11243);
nor U11865 (N_11865,N_11049,N_11494);
and U11866 (N_11866,N_11120,N_11009);
and U11867 (N_11867,N_11189,N_11371);
xor U11868 (N_11868,N_11093,N_11328);
and U11869 (N_11869,N_11490,N_11151);
nor U11870 (N_11870,N_11299,N_11122);
nand U11871 (N_11871,N_11344,N_11185);
nor U11872 (N_11872,N_11096,N_11125);
nand U11873 (N_11873,N_11324,N_11443);
xnor U11874 (N_11874,N_11140,N_11024);
xor U11875 (N_11875,N_11307,N_11097);
nand U11876 (N_11876,N_11339,N_11405);
and U11877 (N_11877,N_11317,N_11080);
nand U11878 (N_11878,N_11307,N_11242);
or U11879 (N_11879,N_11072,N_11175);
or U11880 (N_11880,N_11305,N_11112);
nand U11881 (N_11881,N_11483,N_11133);
xnor U11882 (N_11882,N_11164,N_11408);
nor U11883 (N_11883,N_11205,N_11122);
nor U11884 (N_11884,N_11469,N_11459);
xor U11885 (N_11885,N_11027,N_11093);
xnor U11886 (N_11886,N_11268,N_11393);
nor U11887 (N_11887,N_11048,N_11415);
nand U11888 (N_11888,N_11058,N_11016);
and U11889 (N_11889,N_11157,N_11236);
xor U11890 (N_11890,N_11353,N_11226);
and U11891 (N_11891,N_11336,N_11195);
nand U11892 (N_11892,N_11208,N_11270);
and U11893 (N_11893,N_11310,N_11041);
nor U11894 (N_11894,N_11123,N_11442);
xor U11895 (N_11895,N_11159,N_11129);
nor U11896 (N_11896,N_11096,N_11095);
nor U11897 (N_11897,N_11206,N_11128);
xnor U11898 (N_11898,N_11295,N_11026);
and U11899 (N_11899,N_11473,N_11189);
and U11900 (N_11900,N_11036,N_11469);
or U11901 (N_11901,N_11016,N_11365);
nand U11902 (N_11902,N_11348,N_11443);
and U11903 (N_11903,N_11024,N_11023);
nor U11904 (N_11904,N_11342,N_11361);
and U11905 (N_11905,N_11094,N_11100);
or U11906 (N_11906,N_11371,N_11491);
and U11907 (N_11907,N_11172,N_11092);
nand U11908 (N_11908,N_11316,N_11457);
nand U11909 (N_11909,N_11477,N_11248);
or U11910 (N_11910,N_11404,N_11220);
or U11911 (N_11911,N_11373,N_11043);
and U11912 (N_11912,N_11058,N_11487);
nand U11913 (N_11913,N_11241,N_11131);
xnor U11914 (N_11914,N_11337,N_11073);
nor U11915 (N_11915,N_11390,N_11197);
nor U11916 (N_11916,N_11331,N_11325);
nand U11917 (N_11917,N_11079,N_11245);
nor U11918 (N_11918,N_11133,N_11015);
or U11919 (N_11919,N_11463,N_11254);
and U11920 (N_11920,N_11442,N_11309);
nor U11921 (N_11921,N_11169,N_11353);
xor U11922 (N_11922,N_11150,N_11362);
nand U11923 (N_11923,N_11239,N_11455);
xor U11924 (N_11924,N_11287,N_11372);
or U11925 (N_11925,N_11269,N_11428);
and U11926 (N_11926,N_11206,N_11223);
or U11927 (N_11927,N_11362,N_11452);
and U11928 (N_11928,N_11187,N_11164);
and U11929 (N_11929,N_11323,N_11472);
nand U11930 (N_11930,N_11139,N_11061);
xnor U11931 (N_11931,N_11269,N_11328);
and U11932 (N_11932,N_11263,N_11249);
and U11933 (N_11933,N_11464,N_11127);
nand U11934 (N_11934,N_11197,N_11374);
and U11935 (N_11935,N_11396,N_11162);
xor U11936 (N_11936,N_11329,N_11298);
and U11937 (N_11937,N_11135,N_11428);
nor U11938 (N_11938,N_11284,N_11109);
nand U11939 (N_11939,N_11204,N_11143);
nor U11940 (N_11940,N_11042,N_11476);
nand U11941 (N_11941,N_11463,N_11332);
nor U11942 (N_11942,N_11116,N_11097);
nor U11943 (N_11943,N_11077,N_11224);
xor U11944 (N_11944,N_11266,N_11167);
xnor U11945 (N_11945,N_11021,N_11205);
nand U11946 (N_11946,N_11215,N_11167);
nand U11947 (N_11947,N_11203,N_11485);
nor U11948 (N_11948,N_11180,N_11486);
xor U11949 (N_11949,N_11302,N_11388);
nor U11950 (N_11950,N_11450,N_11459);
or U11951 (N_11951,N_11117,N_11317);
nor U11952 (N_11952,N_11136,N_11185);
nor U11953 (N_11953,N_11057,N_11061);
nand U11954 (N_11954,N_11033,N_11205);
xor U11955 (N_11955,N_11194,N_11479);
nand U11956 (N_11956,N_11230,N_11105);
xor U11957 (N_11957,N_11327,N_11473);
and U11958 (N_11958,N_11452,N_11392);
or U11959 (N_11959,N_11107,N_11086);
xor U11960 (N_11960,N_11015,N_11156);
nor U11961 (N_11961,N_11342,N_11440);
and U11962 (N_11962,N_11003,N_11273);
or U11963 (N_11963,N_11489,N_11106);
nor U11964 (N_11964,N_11012,N_11174);
xnor U11965 (N_11965,N_11054,N_11262);
xor U11966 (N_11966,N_11477,N_11099);
or U11967 (N_11967,N_11020,N_11431);
nor U11968 (N_11968,N_11235,N_11116);
nand U11969 (N_11969,N_11028,N_11478);
nor U11970 (N_11970,N_11289,N_11247);
or U11971 (N_11971,N_11006,N_11225);
nand U11972 (N_11972,N_11208,N_11433);
nand U11973 (N_11973,N_11424,N_11415);
nand U11974 (N_11974,N_11458,N_11353);
nor U11975 (N_11975,N_11172,N_11364);
and U11976 (N_11976,N_11259,N_11252);
xnor U11977 (N_11977,N_11459,N_11155);
nor U11978 (N_11978,N_11468,N_11390);
nand U11979 (N_11979,N_11244,N_11104);
and U11980 (N_11980,N_11352,N_11333);
xnor U11981 (N_11981,N_11232,N_11099);
and U11982 (N_11982,N_11397,N_11392);
nand U11983 (N_11983,N_11273,N_11385);
nand U11984 (N_11984,N_11348,N_11419);
nor U11985 (N_11985,N_11212,N_11453);
nand U11986 (N_11986,N_11379,N_11278);
xor U11987 (N_11987,N_11405,N_11005);
nor U11988 (N_11988,N_11164,N_11369);
and U11989 (N_11989,N_11061,N_11294);
or U11990 (N_11990,N_11162,N_11480);
or U11991 (N_11991,N_11150,N_11351);
xor U11992 (N_11992,N_11416,N_11439);
and U11993 (N_11993,N_11104,N_11096);
or U11994 (N_11994,N_11205,N_11126);
nor U11995 (N_11995,N_11079,N_11086);
nand U11996 (N_11996,N_11157,N_11202);
nand U11997 (N_11997,N_11303,N_11106);
nand U11998 (N_11998,N_11273,N_11040);
nand U11999 (N_11999,N_11224,N_11093);
and U12000 (N_12000,N_11855,N_11517);
nand U12001 (N_12001,N_11878,N_11745);
nor U12002 (N_12002,N_11894,N_11714);
xor U12003 (N_12003,N_11951,N_11567);
nand U12004 (N_12004,N_11725,N_11645);
nor U12005 (N_12005,N_11666,N_11932);
nor U12006 (N_12006,N_11710,N_11602);
xnor U12007 (N_12007,N_11763,N_11523);
or U12008 (N_12008,N_11586,N_11749);
nand U12009 (N_12009,N_11521,N_11513);
nor U12010 (N_12010,N_11698,N_11626);
or U12011 (N_12011,N_11885,N_11678);
nor U12012 (N_12012,N_11871,N_11802);
or U12013 (N_12013,N_11724,N_11667);
nor U12014 (N_12014,N_11590,N_11558);
and U12015 (N_12015,N_11840,N_11767);
nor U12016 (N_12016,N_11639,N_11524);
nand U12017 (N_12017,N_11575,N_11999);
or U12018 (N_12018,N_11832,N_11549);
and U12019 (N_12019,N_11861,N_11849);
nor U12020 (N_12020,N_11760,N_11801);
and U12021 (N_12021,N_11747,N_11653);
nand U12022 (N_12022,N_11778,N_11773);
or U12023 (N_12023,N_11550,N_11627);
nand U12024 (N_12024,N_11598,N_11620);
nand U12025 (N_12025,N_11704,N_11504);
or U12026 (N_12026,N_11930,N_11593);
or U12027 (N_12027,N_11670,N_11842);
or U12028 (N_12028,N_11957,N_11780);
or U12029 (N_12029,N_11883,N_11775);
or U12030 (N_12030,N_11764,N_11565);
nor U12031 (N_12031,N_11650,N_11969);
xor U12032 (N_12032,N_11755,N_11888);
nand U12033 (N_12033,N_11953,N_11881);
nand U12034 (N_12034,N_11975,N_11630);
and U12035 (N_12035,N_11908,N_11697);
xnor U12036 (N_12036,N_11891,N_11603);
or U12037 (N_12037,N_11604,N_11866);
nand U12038 (N_12038,N_11757,N_11948);
nand U12039 (N_12039,N_11737,N_11631);
or U12040 (N_12040,N_11945,N_11787);
nor U12041 (N_12041,N_11679,N_11587);
and U12042 (N_12042,N_11788,N_11560);
xnor U12043 (N_12043,N_11955,N_11858);
or U12044 (N_12044,N_11838,N_11652);
nand U12045 (N_12045,N_11817,N_11544);
nor U12046 (N_12046,N_11823,N_11990);
xnor U12047 (N_12047,N_11898,N_11836);
nand U12048 (N_12048,N_11682,N_11534);
or U12049 (N_12049,N_11654,N_11677);
nand U12050 (N_12050,N_11970,N_11828);
xnor U12051 (N_12051,N_11651,N_11542);
or U12052 (N_12052,N_11728,N_11646);
nand U12053 (N_12053,N_11533,N_11796);
nand U12054 (N_12054,N_11701,N_11614);
xnor U12055 (N_12055,N_11805,N_11717);
or U12056 (N_12056,N_11527,N_11516);
nand U12057 (N_12057,N_11824,N_11783);
nor U12058 (N_12058,N_11634,N_11963);
or U12059 (N_12059,N_11753,N_11875);
nand U12060 (N_12060,N_11872,N_11851);
xor U12061 (N_12061,N_11537,N_11562);
xor U12062 (N_12062,N_11799,N_11976);
nor U12063 (N_12063,N_11937,N_11601);
or U12064 (N_12064,N_11826,N_11867);
and U12065 (N_12065,N_11761,N_11548);
nor U12066 (N_12066,N_11920,N_11821);
and U12067 (N_12067,N_11727,N_11782);
or U12068 (N_12068,N_11797,N_11629);
xnor U12069 (N_12069,N_11865,N_11718);
nand U12070 (N_12070,N_11611,N_11762);
nand U12071 (N_12071,N_11733,N_11663);
nand U12072 (N_12072,N_11924,N_11632);
xnor U12073 (N_12073,N_11769,N_11819);
xor U12074 (N_12074,N_11669,N_11882);
nand U12075 (N_12075,N_11987,N_11641);
or U12076 (N_12076,N_11676,N_11503);
nor U12077 (N_12077,N_11879,N_11923);
xnor U12078 (N_12078,N_11758,N_11686);
xnor U12079 (N_12079,N_11543,N_11556);
or U12080 (N_12080,N_11656,N_11657);
xnor U12081 (N_12081,N_11943,N_11736);
nand U12082 (N_12082,N_11596,N_11655);
and U12083 (N_12083,N_11835,N_11584);
and U12084 (N_12084,N_11526,N_11606);
or U12085 (N_12085,N_11973,N_11863);
nor U12086 (N_12086,N_11771,N_11750);
or U12087 (N_12087,N_11893,N_11995);
xor U12088 (N_12088,N_11595,N_11810);
or U12089 (N_12089,N_11683,N_11748);
nor U12090 (N_12090,N_11941,N_11935);
xnor U12091 (N_12091,N_11884,N_11581);
xnor U12092 (N_12092,N_11928,N_11965);
xor U12093 (N_12093,N_11618,N_11820);
or U12094 (N_12094,N_11774,N_11784);
xor U12095 (N_12095,N_11557,N_11980);
or U12096 (N_12096,N_11768,N_11687);
or U12097 (N_12097,N_11789,N_11633);
xor U12098 (N_12098,N_11623,N_11684);
nand U12099 (N_12099,N_11904,N_11988);
xor U12100 (N_12100,N_11751,N_11752);
and U12101 (N_12101,N_11610,N_11779);
xnor U12102 (N_12102,N_11959,N_11644);
or U12103 (N_12103,N_11536,N_11952);
and U12104 (N_12104,N_11992,N_11658);
nor U12105 (N_12105,N_11692,N_11968);
nand U12106 (N_12106,N_11668,N_11800);
or U12107 (N_12107,N_11994,N_11594);
xor U12108 (N_12108,N_11615,N_11553);
nand U12109 (N_12109,N_11541,N_11529);
nor U12110 (N_12110,N_11699,N_11664);
xor U12111 (N_12111,N_11716,N_11532);
xnor U12112 (N_12112,N_11617,N_11812);
nor U12113 (N_12113,N_11808,N_11597);
nor U12114 (N_12114,N_11555,N_11791);
and U12115 (N_12115,N_11707,N_11960);
nand U12116 (N_12116,N_11837,N_11933);
nand U12117 (N_12117,N_11688,N_11585);
nand U12118 (N_12118,N_11661,N_11672);
nand U12119 (N_12119,N_11729,N_11983);
or U12120 (N_12120,N_11997,N_11638);
nor U12121 (N_12121,N_11739,N_11540);
and U12122 (N_12122,N_11807,N_11911);
nor U12123 (N_12123,N_11845,N_11860);
nand U12124 (N_12124,N_11730,N_11956);
nor U12125 (N_12125,N_11625,N_11874);
and U12126 (N_12126,N_11977,N_11841);
and U12127 (N_12127,N_11675,N_11723);
or U12128 (N_12128,N_11864,N_11743);
nand U12129 (N_12129,N_11785,N_11809);
and U12130 (N_12130,N_11619,N_11531);
xor U12131 (N_12131,N_11674,N_11680);
and U12132 (N_12132,N_11720,N_11856);
nor U12133 (N_12133,N_11915,N_11659);
xnor U12134 (N_12134,N_11693,N_11912);
nor U12135 (N_12135,N_11608,N_11520);
or U12136 (N_12136,N_11703,N_11563);
xnor U12137 (N_12137,N_11927,N_11545);
xor U12138 (N_12138,N_11901,N_11766);
or U12139 (N_12139,N_11514,N_11793);
and U12140 (N_12140,N_11605,N_11671);
and U12141 (N_12141,N_11786,N_11501);
or U12142 (N_12142,N_11588,N_11986);
nand U12143 (N_12143,N_11954,N_11706);
xor U12144 (N_12144,N_11978,N_11577);
or U12145 (N_12145,N_11709,N_11964);
nor U12146 (N_12146,N_11535,N_11936);
or U12147 (N_12147,N_11914,N_11673);
and U12148 (N_12148,N_11947,N_11613);
xor U12149 (N_12149,N_11929,N_11902);
or U12150 (N_12150,N_11877,N_11510);
nand U12151 (N_12151,N_11582,N_11685);
or U12152 (N_12152,N_11816,N_11759);
or U12153 (N_12153,N_11551,N_11846);
or U12154 (N_12154,N_11804,N_11910);
and U12155 (N_12155,N_11917,N_11578);
or U12156 (N_12156,N_11972,N_11993);
or U12157 (N_12157,N_11649,N_11982);
nor U12158 (N_12158,N_11559,N_11806);
xnor U12159 (N_12159,N_11907,N_11742);
xor U12160 (N_12160,N_11525,N_11887);
nor U12161 (N_12161,N_11694,N_11811);
nand U12162 (N_12162,N_11583,N_11580);
and U12163 (N_12163,N_11831,N_11519);
nand U12164 (N_12164,N_11848,N_11561);
or U12165 (N_12165,N_11896,N_11790);
nand U12166 (N_12166,N_11522,N_11958);
nand U12167 (N_12167,N_11918,N_11592);
nand U12168 (N_12168,N_11777,N_11852);
and U12169 (N_12169,N_11859,N_11511);
nor U12170 (N_12170,N_11825,N_11530);
xor U12171 (N_12171,N_11734,N_11776);
xor U12172 (N_12172,N_11552,N_11732);
nor U12173 (N_12173,N_11538,N_11949);
and U12174 (N_12174,N_11547,N_11622);
nand U12175 (N_12175,N_11985,N_11660);
and U12176 (N_12176,N_11981,N_11892);
and U12177 (N_12177,N_11833,N_11862);
xnor U12178 (N_12178,N_11938,N_11942);
or U12179 (N_12179,N_11568,N_11919);
xor U12180 (N_12180,N_11711,N_11741);
or U12181 (N_12181,N_11609,N_11621);
nand U12182 (N_12182,N_11991,N_11572);
nor U12183 (N_12183,N_11827,N_11574);
xnor U12184 (N_12184,N_11996,N_11500);
nand U12185 (N_12185,N_11853,N_11566);
nor U12186 (N_12186,N_11696,N_11869);
nor U12187 (N_12187,N_11829,N_11850);
nor U12188 (N_12188,N_11876,N_11726);
nor U12189 (N_12189,N_11616,N_11847);
nor U12190 (N_12190,N_11905,N_11818);
or U12191 (N_12191,N_11554,N_11974);
nor U12192 (N_12192,N_11897,N_11570);
or U12193 (N_12193,N_11528,N_11889);
nand U12194 (N_12194,N_11665,N_11512);
nand U12195 (N_12195,N_11813,N_11640);
xnor U12196 (N_12196,N_11868,N_11913);
xor U12197 (N_12197,N_11515,N_11903);
xnor U12198 (N_12198,N_11599,N_11506);
and U12199 (N_12199,N_11754,N_11539);
or U12200 (N_12200,N_11803,N_11971);
xnor U12201 (N_12201,N_11854,N_11950);
and U12202 (N_12202,N_11926,N_11695);
and U12203 (N_12203,N_11591,N_11934);
nand U12204 (N_12204,N_11722,N_11740);
xor U12205 (N_12205,N_11834,N_11931);
or U12206 (N_12206,N_11798,N_11744);
xnor U12207 (N_12207,N_11922,N_11814);
or U12208 (N_12208,N_11579,N_11648);
or U12209 (N_12209,N_11900,N_11839);
nor U12210 (N_12210,N_11691,N_11564);
or U12211 (N_12211,N_11822,N_11642);
xor U12212 (N_12212,N_11731,N_11637);
nand U12213 (N_12213,N_11681,N_11518);
nand U12214 (N_12214,N_11880,N_11628);
or U12215 (N_12215,N_11643,N_11906);
and U12216 (N_12216,N_11712,N_11607);
nand U12217 (N_12217,N_11815,N_11569);
nor U12218 (N_12218,N_11735,N_11702);
nand U12219 (N_12219,N_11830,N_11916);
nand U12220 (N_12220,N_11708,N_11746);
nand U12221 (N_12221,N_11961,N_11715);
nand U12222 (N_12222,N_11795,N_11721);
xor U12223 (N_12223,N_11770,N_11979);
nor U12224 (N_12224,N_11925,N_11967);
nand U12225 (N_12225,N_11794,N_11765);
nor U12226 (N_12226,N_11772,N_11946);
nor U12227 (N_12227,N_11921,N_11756);
nor U12228 (N_12228,N_11705,N_11792);
and U12229 (N_12229,N_11844,N_11612);
nor U12230 (N_12230,N_11571,N_11940);
xnor U12231 (N_12231,N_11944,N_11895);
nand U12232 (N_12232,N_11635,N_11573);
or U12233 (N_12233,N_11713,N_11890);
nor U12234 (N_12234,N_11507,N_11600);
nor U12235 (N_12235,N_11886,N_11576);
nor U12236 (N_12236,N_11502,N_11689);
nand U12237 (N_12237,N_11662,N_11873);
and U12238 (N_12238,N_11962,N_11738);
or U12239 (N_12239,N_11966,N_11870);
nor U12240 (N_12240,N_11843,N_11546);
nand U12241 (N_12241,N_11700,N_11647);
or U12242 (N_12242,N_11690,N_11939);
nor U12243 (N_12243,N_11505,N_11989);
and U12244 (N_12244,N_11909,N_11636);
xnor U12245 (N_12245,N_11589,N_11508);
xor U12246 (N_12246,N_11624,N_11509);
xor U12247 (N_12247,N_11857,N_11781);
or U12248 (N_12248,N_11984,N_11899);
or U12249 (N_12249,N_11719,N_11998);
or U12250 (N_12250,N_11923,N_11733);
nand U12251 (N_12251,N_11847,N_11585);
xnor U12252 (N_12252,N_11829,N_11806);
xor U12253 (N_12253,N_11656,N_11554);
nor U12254 (N_12254,N_11870,N_11783);
or U12255 (N_12255,N_11842,N_11543);
nand U12256 (N_12256,N_11590,N_11804);
nor U12257 (N_12257,N_11561,N_11930);
nand U12258 (N_12258,N_11880,N_11837);
nor U12259 (N_12259,N_11940,N_11991);
xor U12260 (N_12260,N_11845,N_11901);
and U12261 (N_12261,N_11571,N_11831);
and U12262 (N_12262,N_11661,N_11758);
and U12263 (N_12263,N_11605,N_11974);
xnor U12264 (N_12264,N_11500,N_11980);
or U12265 (N_12265,N_11665,N_11534);
and U12266 (N_12266,N_11598,N_11871);
or U12267 (N_12267,N_11714,N_11554);
nor U12268 (N_12268,N_11718,N_11860);
xor U12269 (N_12269,N_11758,N_11796);
nor U12270 (N_12270,N_11791,N_11842);
or U12271 (N_12271,N_11956,N_11562);
xnor U12272 (N_12272,N_11704,N_11594);
or U12273 (N_12273,N_11960,N_11593);
xor U12274 (N_12274,N_11924,N_11723);
nand U12275 (N_12275,N_11940,N_11999);
xor U12276 (N_12276,N_11998,N_11780);
nor U12277 (N_12277,N_11536,N_11571);
or U12278 (N_12278,N_11893,N_11940);
xnor U12279 (N_12279,N_11702,N_11937);
nor U12280 (N_12280,N_11515,N_11783);
xor U12281 (N_12281,N_11536,N_11605);
xor U12282 (N_12282,N_11561,N_11996);
nand U12283 (N_12283,N_11689,N_11847);
nor U12284 (N_12284,N_11782,N_11740);
nand U12285 (N_12285,N_11732,N_11996);
or U12286 (N_12286,N_11959,N_11859);
xnor U12287 (N_12287,N_11872,N_11500);
nor U12288 (N_12288,N_11827,N_11923);
nand U12289 (N_12289,N_11793,N_11667);
or U12290 (N_12290,N_11901,N_11799);
or U12291 (N_12291,N_11518,N_11944);
xor U12292 (N_12292,N_11717,N_11594);
and U12293 (N_12293,N_11948,N_11944);
nand U12294 (N_12294,N_11631,N_11997);
nand U12295 (N_12295,N_11843,N_11693);
and U12296 (N_12296,N_11914,N_11978);
nor U12297 (N_12297,N_11732,N_11704);
nor U12298 (N_12298,N_11750,N_11803);
nor U12299 (N_12299,N_11808,N_11957);
nor U12300 (N_12300,N_11744,N_11941);
nand U12301 (N_12301,N_11810,N_11538);
nand U12302 (N_12302,N_11623,N_11800);
nand U12303 (N_12303,N_11887,N_11924);
xor U12304 (N_12304,N_11844,N_11947);
or U12305 (N_12305,N_11823,N_11999);
nor U12306 (N_12306,N_11894,N_11644);
xor U12307 (N_12307,N_11606,N_11910);
nor U12308 (N_12308,N_11761,N_11876);
nand U12309 (N_12309,N_11874,N_11895);
or U12310 (N_12310,N_11527,N_11644);
or U12311 (N_12311,N_11762,N_11764);
and U12312 (N_12312,N_11606,N_11955);
or U12313 (N_12313,N_11745,N_11997);
and U12314 (N_12314,N_11590,N_11949);
or U12315 (N_12315,N_11989,N_11852);
nand U12316 (N_12316,N_11856,N_11773);
nand U12317 (N_12317,N_11740,N_11958);
nand U12318 (N_12318,N_11941,N_11618);
and U12319 (N_12319,N_11600,N_11574);
nand U12320 (N_12320,N_11944,N_11917);
nor U12321 (N_12321,N_11755,N_11591);
or U12322 (N_12322,N_11741,N_11915);
or U12323 (N_12323,N_11890,N_11720);
nor U12324 (N_12324,N_11768,N_11618);
or U12325 (N_12325,N_11842,N_11619);
nor U12326 (N_12326,N_11814,N_11586);
nor U12327 (N_12327,N_11785,N_11653);
nor U12328 (N_12328,N_11840,N_11555);
or U12329 (N_12329,N_11586,N_11924);
nand U12330 (N_12330,N_11900,N_11991);
nor U12331 (N_12331,N_11502,N_11886);
nand U12332 (N_12332,N_11770,N_11696);
and U12333 (N_12333,N_11967,N_11623);
nand U12334 (N_12334,N_11987,N_11948);
or U12335 (N_12335,N_11594,N_11543);
and U12336 (N_12336,N_11554,N_11988);
nor U12337 (N_12337,N_11781,N_11771);
nand U12338 (N_12338,N_11814,N_11714);
nor U12339 (N_12339,N_11685,N_11591);
nor U12340 (N_12340,N_11566,N_11738);
xnor U12341 (N_12341,N_11621,N_11695);
nor U12342 (N_12342,N_11557,N_11918);
and U12343 (N_12343,N_11694,N_11718);
nand U12344 (N_12344,N_11835,N_11812);
nand U12345 (N_12345,N_11792,N_11737);
or U12346 (N_12346,N_11900,N_11880);
nor U12347 (N_12347,N_11724,N_11574);
or U12348 (N_12348,N_11677,N_11681);
and U12349 (N_12349,N_11758,N_11920);
nor U12350 (N_12350,N_11908,N_11719);
or U12351 (N_12351,N_11612,N_11679);
xor U12352 (N_12352,N_11639,N_11706);
and U12353 (N_12353,N_11762,N_11621);
nor U12354 (N_12354,N_11971,N_11986);
xor U12355 (N_12355,N_11838,N_11717);
nor U12356 (N_12356,N_11910,N_11824);
xnor U12357 (N_12357,N_11574,N_11952);
nor U12358 (N_12358,N_11788,N_11701);
and U12359 (N_12359,N_11728,N_11836);
nor U12360 (N_12360,N_11874,N_11520);
nand U12361 (N_12361,N_11835,N_11644);
xor U12362 (N_12362,N_11976,N_11609);
xor U12363 (N_12363,N_11895,N_11667);
nand U12364 (N_12364,N_11780,N_11987);
and U12365 (N_12365,N_11635,N_11590);
or U12366 (N_12366,N_11931,N_11660);
nor U12367 (N_12367,N_11723,N_11528);
and U12368 (N_12368,N_11601,N_11897);
xor U12369 (N_12369,N_11955,N_11742);
nor U12370 (N_12370,N_11690,N_11874);
nor U12371 (N_12371,N_11648,N_11934);
and U12372 (N_12372,N_11906,N_11994);
nand U12373 (N_12373,N_11800,N_11517);
xor U12374 (N_12374,N_11712,N_11534);
xnor U12375 (N_12375,N_11966,N_11816);
nor U12376 (N_12376,N_11576,N_11625);
nand U12377 (N_12377,N_11944,N_11786);
and U12378 (N_12378,N_11934,N_11863);
nor U12379 (N_12379,N_11721,N_11778);
or U12380 (N_12380,N_11530,N_11689);
nor U12381 (N_12381,N_11706,N_11772);
xnor U12382 (N_12382,N_11809,N_11556);
or U12383 (N_12383,N_11802,N_11699);
or U12384 (N_12384,N_11719,N_11965);
nor U12385 (N_12385,N_11695,N_11804);
and U12386 (N_12386,N_11756,N_11533);
and U12387 (N_12387,N_11821,N_11876);
xnor U12388 (N_12388,N_11775,N_11850);
xor U12389 (N_12389,N_11836,N_11852);
nand U12390 (N_12390,N_11672,N_11947);
or U12391 (N_12391,N_11543,N_11629);
nor U12392 (N_12392,N_11904,N_11644);
nand U12393 (N_12393,N_11587,N_11504);
nand U12394 (N_12394,N_11911,N_11622);
xnor U12395 (N_12395,N_11655,N_11907);
nand U12396 (N_12396,N_11514,N_11928);
nor U12397 (N_12397,N_11896,N_11761);
nor U12398 (N_12398,N_11722,N_11531);
nor U12399 (N_12399,N_11726,N_11794);
nand U12400 (N_12400,N_11503,N_11878);
xor U12401 (N_12401,N_11889,N_11522);
or U12402 (N_12402,N_11861,N_11799);
nand U12403 (N_12403,N_11552,N_11995);
and U12404 (N_12404,N_11925,N_11563);
and U12405 (N_12405,N_11955,N_11762);
nand U12406 (N_12406,N_11513,N_11679);
nor U12407 (N_12407,N_11775,N_11674);
nor U12408 (N_12408,N_11604,N_11905);
or U12409 (N_12409,N_11897,N_11852);
nor U12410 (N_12410,N_11727,N_11623);
xnor U12411 (N_12411,N_11806,N_11758);
xnor U12412 (N_12412,N_11674,N_11734);
or U12413 (N_12413,N_11883,N_11952);
or U12414 (N_12414,N_11771,N_11896);
or U12415 (N_12415,N_11654,N_11693);
nand U12416 (N_12416,N_11923,N_11990);
xor U12417 (N_12417,N_11927,N_11921);
or U12418 (N_12418,N_11817,N_11848);
xor U12419 (N_12419,N_11712,N_11764);
nor U12420 (N_12420,N_11580,N_11585);
or U12421 (N_12421,N_11903,N_11665);
nor U12422 (N_12422,N_11616,N_11644);
nor U12423 (N_12423,N_11993,N_11754);
nand U12424 (N_12424,N_11573,N_11515);
or U12425 (N_12425,N_11682,N_11709);
or U12426 (N_12426,N_11611,N_11567);
nand U12427 (N_12427,N_11870,N_11587);
and U12428 (N_12428,N_11676,N_11512);
nand U12429 (N_12429,N_11517,N_11646);
and U12430 (N_12430,N_11550,N_11536);
xnor U12431 (N_12431,N_11986,N_11898);
nor U12432 (N_12432,N_11992,N_11610);
and U12433 (N_12433,N_11771,N_11543);
or U12434 (N_12434,N_11531,N_11707);
or U12435 (N_12435,N_11635,N_11520);
or U12436 (N_12436,N_11766,N_11693);
nor U12437 (N_12437,N_11572,N_11930);
nor U12438 (N_12438,N_11935,N_11552);
or U12439 (N_12439,N_11593,N_11645);
xnor U12440 (N_12440,N_11679,N_11566);
nor U12441 (N_12441,N_11844,N_11817);
nand U12442 (N_12442,N_11706,N_11717);
and U12443 (N_12443,N_11890,N_11517);
xor U12444 (N_12444,N_11520,N_11837);
nand U12445 (N_12445,N_11668,N_11872);
and U12446 (N_12446,N_11653,N_11510);
or U12447 (N_12447,N_11871,N_11980);
nor U12448 (N_12448,N_11951,N_11991);
nor U12449 (N_12449,N_11796,N_11766);
nand U12450 (N_12450,N_11684,N_11814);
and U12451 (N_12451,N_11998,N_11697);
or U12452 (N_12452,N_11685,N_11949);
nor U12453 (N_12453,N_11900,N_11847);
nor U12454 (N_12454,N_11587,N_11527);
nand U12455 (N_12455,N_11829,N_11773);
and U12456 (N_12456,N_11657,N_11564);
xnor U12457 (N_12457,N_11613,N_11635);
and U12458 (N_12458,N_11767,N_11624);
or U12459 (N_12459,N_11523,N_11912);
and U12460 (N_12460,N_11604,N_11992);
or U12461 (N_12461,N_11504,N_11939);
xnor U12462 (N_12462,N_11593,N_11789);
and U12463 (N_12463,N_11973,N_11837);
xor U12464 (N_12464,N_11887,N_11646);
nor U12465 (N_12465,N_11731,N_11932);
xor U12466 (N_12466,N_11986,N_11637);
or U12467 (N_12467,N_11689,N_11602);
nor U12468 (N_12468,N_11671,N_11802);
nand U12469 (N_12469,N_11812,N_11731);
nor U12470 (N_12470,N_11734,N_11787);
nand U12471 (N_12471,N_11592,N_11822);
or U12472 (N_12472,N_11591,N_11574);
or U12473 (N_12473,N_11761,N_11943);
nor U12474 (N_12474,N_11968,N_11888);
xnor U12475 (N_12475,N_11851,N_11806);
and U12476 (N_12476,N_11817,N_11980);
nand U12477 (N_12477,N_11513,N_11656);
nand U12478 (N_12478,N_11504,N_11933);
nand U12479 (N_12479,N_11931,N_11658);
or U12480 (N_12480,N_11519,N_11953);
nor U12481 (N_12481,N_11616,N_11722);
nor U12482 (N_12482,N_11835,N_11566);
or U12483 (N_12483,N_11843,N_11626);
nor U12484 (N_12484,N_11669,N_11934);
nor U12485 (N_12485,N_11832,N_11690);
nand U12486 (N_12486,N_11868,N_11852);
or U12487 (N_12487,N_11952,N_11656);
and U12488 (N_12488,N_11975,N_11596);
nor U12489 (N_12489,N_11945,N_11720);
nor U12490 (N_12490,N_11837,N_11698);
xor U12491 (N_12491,N_11593,N_11513);
xor U12492 (N_12492,N_11678,N_11941);
and U12493 (N_12493,N_11899,N_11780);
xnor U12494 (N_12494,N_11611,N_11899);
nor U12495 (N_12495,N_11625,N_11562);
or U12496 (N_12496,N_11512,N_11820);
nor U12497 (N_12497,N_11542,N_11932);
xnor U12498 (N_12498,N_11660,N_11723);
xor U12499 (N_12499,N_11654,N_11907);
xor U12500 (N_12500,N_12383,N_12046);
or U12501 (N_12501,N_12086,N_12217);
xnor U12502 (N_12502,N_12206,N_12095);
nor U12503 (N_12503,N_12278,N_12435);
or U12504 (N_12504,N_12471,N_12181);
and U12505 (N_12505,N_12223,N_12491);
and U12506 (N_12506,N_12088,N_12111);
nor U12507 (N_12507,N_12245,N_12405);
xor U12508 (N_12508,N_12215,N_12368);
nor U12509 (N_12509,N_12303,N_12320);
nor U12510 (N_12510,N_12065,N_12482);
or U12511 (N_12511,N_12304,N_12124);
and U12512 (N_12512,N_12269,N_12131);
nand U12513 (N_12513,N_12102,N_12361);
nand U12514 (N_12514,N_12209,N_12133);
xnor U12515 (N_12515,N_12387,N_12384);
or U12516 (N_12516,N_12317,N_12167);
or U12517 (N_12517,N_12324,N_12393);
xnor U12518 (N_12518,N_12319,N_12477);
nand U12519 (N_12519,N_12097,N_12479);
xnor U12520 (N_12520,N_12233,N_12262);
nand U12521 (N_12521,N_12195,N_12055);
and U12522 (N_12522,N_12173,N_12045);
nand U12523 (N_12523,N_12256,N_12483);
or U12524 (N_12524,N_12000,N_12196);
nor U12525 (N_12525,N_12313,N_12009);
or U12526 (N_12526,N_12467,N_12026);
nor U12527 (N_12527,N_12164,N_12335);
xnor U12528 (N_12528,N_12430,N_12035);
nor U12529 (N_12529,N_12087,N_12478);
xor U12530 (N_12530,N_12300,N_12421);
or U12531 (N_12531,N_12406,N_12083);
xor U12532 (N_12532,N_12386,N_12459);
xor U12533 (N_12533,N_12027,N_12194);
xor U12534 (N_12534,N_12487,N_12068);
and U12535 (N_12535,N_12450,N_12099);
xor U12536 (N_12536,N_12422,N_12100);
or U12537 (N_12537,N_12456,N_12161);
or U12538 (N_12538,N_12469,N_12307);
and U12539 (N_12539,N_12399,N_12006);
nor U12540 (N_12540,N_12080,N_12373);
xor U12541 (N_12541,N_12146,N_12123);
and U12542 (N_12542,N_12426,N_12486);
nor U12543 (N_12543,N_12150,N_12492);
nand U12544 (N_12544,N_12396,N_12163);
nand U12545 (N_12545,N_12473,N_12135);
nor U12546 (N_12546,N_12410,N_12170);
nor U12547 (N_12547,N_12231,N_12485);
nand U12548 (N_12548,N_12428,N_12371);
xnor U12549 (N_12549,N_12323,N_12263);
nor U12550 (N_12550,N_12416,N_12364);
or U12551 (N_12551,N_12214,N_12162);
nand U12552 (N_12552,N_12059,N_12367);
nor U12553 (N_12553,N_12295,N_12136);
nor U12554 (N_12554,N_12321,N_12011);
and U12555 (N_12555,N_12166,N_12172);
nand U12556 (N_12556,N_12415,N_12210);
nand U12557 (N_12557,N_12252,N_12454);
and U12558 (N_12558,N_12458,N_12293);
nor U12559 (N_12559,N_12061,N_12446);
nor U12560 (N_12560,N_12208,N_12365);
nor U12561 (N_12561,N_12104,N_12372);
nand U12562 (N_12562,N_12148,N_12126);
nand U12563 (N_12563,N_12407,N_12152);
nor U12564 (N_12564,N_12413,N_12344);
or U12565 (N_12565,N_12424,N_12075);
nor U12566 (N_12566,N_12230,N_12193);
and U12567 (N_12567,N_12178,N_12119);
or U12568 (N_12568,N_12191,N_12251);
nand U12569 (N_12569,N_12114,N_12240);
nor U12570 (N_12570,N_12211,N_12332);
or U12571 (N_12571,N_12468,N_12139);
or U12572 (N_12572,N_12184,N_12355);
and U12573 (N_12573,N_12460,N_12398);
xor U12574 (N_12574,N_12318,N_12484);
nand U12575 (N_12575,N_12499,N_12238);
xnor U12576 (N_12576,N_12154,N_12408);
and U12577 (N_12577,N_12089,N_12200);
or U12578 (N_12578,N_12334,N_12296);
xor U12579 (N_12579,N_12286,N_12069);
xor U12580 (N_12580,N_12040,N_12464);
nor U12581 (N_12581,N_12338,N_12457);
or U12582 (N_12582,N_12235,N_12056);
nor U12583 (N_12583,N_12310,N_12084);
and U12584 (N_12584,N_12369,N_12288);
xnor U12585 (N_12585,N_12187,N_12337);
or U12586 (N_12586,N_12264,N_12122);
xnor U12587 (N_12587,N_12349,N_12466);
and U12588 (N_12588,N_12322,N_12067);
and U12589 (N_12589,N_12107,N_12401);
xor U12590 (N_12590,N_12420,N_12047);
or U12591 (N_12591,N_12378,N_12397);
and U12592 (N_12592,N_12292,N_12077);
nand U12593 (N_12593,N_12297,N_12060);
nor U12594 (N_12594,N_12121,N_12140);
and U12595 (N_12595,N_12096,N_12168);
nor U12596 (N_12596,N_12429,N_12201);
and U12597 (N_12597,N_12352,N_12023);
and U12598 (N_12598,N_12388,N_12402);
and U12599 (N_12599,N_12325,N_12453);
xnor U12600 (N_12600,N_12205,N_12246);
or U12601 (N_12601,N_12409,N_12120);
nor U12602 (N_12602,N_12003,N_12366);
xnor U12603 (N_12603,N_12329,N_12129);
nand U12604 (N_12604,N_12073,N_12298);
nor U12605 (N_12605,N_12042,N_12203);
nor U12606 (N_12606,N_12132,N_12160);
xnor U12607 (N_12607,N_12273,N_12041);
nor U12608 (N_12608,N_12443,N_12177);
nand U12609 (N_12609,N_12391,N_12326);
xor U12610 (N_12610,N_12180,N_12182);
nor U12611 (N_12611,N_12390,N_12270);
nand U12612 (N_12612,N_12362,N_12036);
or U12613 (N_12613,N_12103,N_12495);
nor U12614 (N_12614,N_12227,N_12147);
nand U12615 (N_12615,N_12261,N_12091);
nor U12616 (N_12616,N_12171,N_12239);
nor U12617 (N_12617,N_12285,N_12071);
xor U12618 (N_12618,N_12336,N_12062);
or U12619 (N_12619,N_12439,N_12149);
and U12620 (N_12620,N_12145,N_12192);
xnor U12621 (N_12621,N_12185,N_12249);
nor U12622 (N_12622,N_12455,N_12382);
xor U12623 (N_12623,N_12019,N_12431);
xnor U12624 (N_12624,N_12440,N_12109);
and U12625 (N_12625,N_12012,N_12013);
and U12626 (N_12626,N_12277,N_12142);
nor U12627 (N_12627,N_12363,N_12275);
or U12628 (N_12628,N_12283,N_12445);
nand U12629 (N_12629,N_12225,N_12434);
xnor U12630 (N_12630,N_12034,N_12308);
or U12631 (N_12631,N_12353,N_12274);
nor U12632 (N_12632,N_12490,N_12280);
xnor U12633 (N_12633,N_12015,N_12221);
nand U12634 (N_12634,N_12279,N_12199);
nand U12635 (N_12635,N_12379,N_12465);
nand U12636 (N_12636,N_12494,N_12258);
and U12637 (N_12637,N_12299,N_12436);
and U12638 (N_12638,N_12289,N_12330);
nor U12639 (N_12639,N_12198,N_12052);
nor U12640 (N_12640,N_12057,N_12137);
nand U12641 (N_12641,N_12385,N_12389);
nor U12642 (N_12642,N_12017,N_12063);
and U12643 (N_12643,N_12400,N_12327);
and U12644 (N_12644,N_12462,N_12090);
nor U12645 (N_12645,N_12347,N_12476);
nor U12646 (N_12646,N_12081,N_12315);
nand U12647 (N_12647,N_12312,N_12255);
or U12648 (N_12648,N_12448,N_12309);
nand U12649 (N_12649,N_12333,N_12115);
nor U12650 (N_12650,N_12444,N_12475);
and U12651 (N_12651,N_12305,N_12447);
xor U12652 (N_12652,N_12417,N_12427);
and U12653 (N_12653,N_12425,N_12058);
or U12654 (N_12654,N_12449,N_12219);
and U12655 (N_12655,N_12116,N_12144);
xnor U12656 (N_12656,N_12064,N_12125);
nor U12657 (N_12657,N_12079,N_12271);
nand U12658 (N_12658,N_12282,N_12403);
or U12659 (N_12659,N_12496,N_12020);
nor U12660 (N_12660,N_12112,N_12244);
nand U12661 (N_12661,N_12302,N_12418);
xor U12662 (N_12662,N_12049,N_12250);
nor U12663 (N_12663,N_12498,N_12127);
xor U12664 (N_12664,N_12260,N_12392);
nand U12665 (N_12665,N_12374,N_12226);
or U12666 (N_12666,N_12480,N_12452);
or U12667 (N_12667,N_12357,N_12272);
and U12668 (N_12668,N_12105,N_12348);
nand U12669 (N_12669,N_12316,N_12207);
nand U12670 (N_12670,N_12204,N_12481);
or U12671 (N_12671,N_12281,N_12082);
or U12672 (N_12672,N_12029,N_12234);
or U12673 (N_12673,N_12039,N_12010);
and U12674 (N_12674,N_12222,N_12044);
and U12675 (N_12675,N_12007,N_12229);
nor U12676 (N_12676,N_12128,N_12380);
nand U12677 (N_12677,N_12016,N_12254);
nor U12678 (N_12678,N_12311,N_12346);
nand U12679 (N_12679,N_12257,N_12247);
or U12680 (N_12680,N_12018,N_12284);
and U12681 (N_12681,N_12008,N_12306);
nor U12682 (N_12682,N_12472,N_12241);
xnor U12683 (N_12683,N_12276,N_12159);
nand U12684 (N_12684,N_12339,N_12438);
nand U12685 (N_12685,N_12442,N_12404);
nand U12686 (N_12686,N_12359,N_12343);
nand U12687 (N_12687,N_12267,N_12268);
nor U12688 (N_12688,N_12224,N_12188);
or U12689 (N_12689,N_12101,N_12028);
or U12690 (N_12690,N_12394,N_12037);
nor U12691 (N_12691,N_12085,N_12213);
nor U12692 (N_12692,N_12113,N_12497);
or U12693 (N_12693,N_12048,N_12216);
xor U12694 (N_12694,N_12350,N_12053);
nand U12695 (N_12695,N_12423,N_12038);
xor U12696 (N_12696,N_12432,N_12354);
nor U12697 (N_12697,N_12176,N_12092);
and U12698 (N_12698,N_12025,N_12070);
nor U12699 (N_12699,N_12489,N_12461);
or U12700 (N_12700,N_12002,N_12138);
and U12701 (N_12701,N_12242,N_12074);
or U12702 (N_12702,N_12014,N_12381);
nand U12703 (N_12703,N_12232,N_12143);
and U12704 (N_12704,N_12179,N_12151);
and U12705 (N_12705,N_12220,N_12243);
nand U12706 (N_12706,N_12294,N_12021);
nor U12707 (N_12707,N_12377,N_12078);
xor U12708 (N_12708,N_12066,N_12441);
nand U12709 (N_12709,N_12345,N_12033);
xor U12710 (N_12710,N_12248,N_12054);
nand U12711 (N_12711,N_12165,N_12024);
xnor U12712 (N_12712,N_12004,N_12265);
xor U12713 (N_12713,N_12043,N_12118);
xor U12714 (N_12714,N_12470,N_12451);
xnor U12715 (N_12715,N_12331,N_12375);
or U12716 (N_12716,N_12157,N_12197);
nand U12717 (N_12717,N_12155,N_12395);
or U12718 (N_12718,N_12169,N_12094);
or U12719 (N_12719,N_12174,N_12287);
nor U12720 (N_12720,N_12360,N_12050);
nor U12721 (N_12721,N_12356,N_12175);
or U12722 (N_12722,N_12290,N_12493);
nand U12723 (N_12723,N_12051,N_12134);
xnor U12724 (N_12724,N_12259,N_12341);
or U12725 (N_12725,N_12032,N_12158);
xnor U12726 (N_12726,N_12253,N_12376);
nor U12727 (N_12727,N_12108,N_12106);
nand U12728 (N_12728,N_12212,N_12433);
or U12729 (N_12729,N_12340,N_12266);
nor U12730 (N_12730,N_12189,N_12412);
or U12731 (N_12731,N_12351,N_12370);
or U12732 (N_12732,N_12463,N_12328);
and U12733 (N_12733,N_12419,N_12130);
nor U12734 (N_12734,N_12183,N_12358);
nor U12735 (N_12735,N_12110,N_12031);
xor U12736 (N_12736,N_12291,N_12314);
xnor U12737 (N_12737,N_12156,N_12218);
nand U12738 (N_12738,N_12237,N_12411);
nand U12739 (N_12739,N_12202,N_12093);
and U12740 (N_12740,N_12414,N_12236);
and U12741 (N_12741,N_12098,N_12437);
and U12742 (N_12742,N_12186,N_12141);
nand U12743 (N_12743,N_12488,N_12474);
xnor U12744 (N_12744,N_12005,N_12342);
nand U12745 (N_12745,N_12228,N_12076);
and U12746 (N_12746,N_12022,N_12117);
or U12747 (N_12747,N_12030,N_12301);
and U12748 (N_12748,N_12072,N_12153);
xnor U12749 (N_12749,N_12190,N_12001);
or U12750 (N_12750,N_12471,N_12280);
nor U12751 (N_12751,N_12469,N_12084);
and U12752 (N_12752,N_12030,N_12297);
or U12753 (N_12753,N_12129,N_12396);
xor U12754 (N_12754,N_12101,N_12091);
nor U12755 (N_12755,N_12163,N_12123);
or U12756 (N_12756,N_12036,N_12350);
xor U12757 (N_12757,N_12471,N_12162);
nor U12758 (N_12758,N_12145,N_12024);
or U12759 (N_12759,N_12129,N_12332);
and U12760 (N_12760,N_12130,N_12224);
nor U12761 (N_12761,N_12380,N_12468);
xor U12762 (N_12762,N_12062,N_12198);
xnor U12763 (N_12763,N_12201,N_12278);
nor U12764 (N_12764,N_12219,N_12234);
xor U12765 (N_12765,N_12272,N_12432);
and U12766 (N_12766,N_12040,N_12367);
xor U12767 (N_12767,N_12031,N_12311);
xnor U12768 (N_12768,N_12407,N_12427);
nor U12769 (N_12769,N_12265,N_12440);
and U12770 (N_12770,N_12297,N_12459);
nor U12771 (N_12771,N_12135,N_12224);
nand U12772 (N_12772,N_12464,N_12296);
nor U12773 (N_12773,N_12477,N_12353);
and U12774 (N_12774,N_12316,N_12261);
xnor U12775 (N_12775,N_12024,N_12412);
nor U12776 (N_12776,N_12347,N_12080);
nor U12777 (N_12777,N_12087,N_12032);
or U12778 (N_12778,N_12329,N_12196);
xnor U12779 (N_12779,N_12392,N_12192);
and U12780 (N_12780,N_12026,N_12087);
or U12781 (N_12781,N_12327,N_12166);
or U12782 (N_12782,N_12049,N_12314);
or U12783 (N_12783,N_12337,N_12214);
xor U12784 (N_12784,N_12051,N_12021);
nor U12785 (N_12785,N_12124,N_12321);
xor U12786 (N_12786,N_12355,N_12241);
nor U12787 (N_12787,N_12200,N_12235);
xnor U12788 (N_12788,N_12197,N_12459);
or U12789 (N_12789,N_12363,N_12030);
nor U12790 (N_12790,N_12319,N_12251);
nor U12791 (N_12791,N_12097,N_12316);
nand U12792 (N_12792,N_12195,N_12051);
and U12793 (N_12793,N_12075,N_12218);
or U12794 (N_12794,N_12335,N_12285);
nor U12795 (N_12795,N_12481,N_12184);
xnor U12796 (N_12796,N_12332,N_12319);
nor U12797 (N_12797,N_12297,N_12027);
xnor U12798 (N_12798,N_12468,N_12423);
or U12799 (N_12799,N_12200,N_12250);
and U12800 (N_12800,N_12421,N_12022);
nand U12801 (N_12801,N_12256,N_12015);
nor U12802 (N_12802,N_12075,N_12040);
nand U12803 (N_12803,N_12456,N_12093);
nor U12804 (N_12804,N_12209,N_12285);
nand U12805 (N_12805,N_12034,N_12484);
nor U12806 (N_12806,N_12230,N_12377);
nor U12807 (N_12807,N_12336,N_12377);
or U12808 (N_12808,N_12079,N_12012);
and U12809 (N_12809,N_12111,N_12044);
or U12810 (N_12810,N_12239,N_12375);
or U12811 (N_12811,N_12125,N_12446);
or U12812 (N_12812,N_12499,N_12410);
nand U12813 (N_12813,N_12307,N_12149);
nand U12814 (N_12814,N_12316,N_12065);
nand U12815 (N_12815,N_12062,N_12097);
and U12816 (N_12816,N_12489,N_12497);
nor U12817 (N_12817,N_12472,N_12073);
and U12818 (N_12818,N_12101,N_12353);
xnor U12819 (N_12819,N_12082,N_12039);
nand U12820 (N_12820,N_12285,N_12404);
nor U12821 (N_12821,N_12388,N_12433);
and U12822 (N_12822,N_12187,N_12273);
nor U12823 (N_12823,N_12325,N_12345);
xnor U12824 (N_12824,N_12356,N_12251);
nand U12825 (N_12825,N_12120,N_12358);
or U12826 (N_12826,N_12083,N_12292);
nand U12827 (N_12827,N_12317,N_12443);
nor U12828 (N_12828,N_12270,N_12480);
xnor U12829 (N_12829,N_12322,N_12284);
and U12830 (N_12830,N_12315,N_12398);
xnor U12831 (N_12831,N_12372,N_12312);
and U12832 (N_12832,N_12083,N_12086);
and U12833 (N_12833,N_12039,N_12391);
nor U12834 (N_12834,N_12163,N_12161);
or U12835 (N_12835,N_12288,N_12467);
and U12836 (N_12836,N_12239,N_12140);
and U12837 (N_12837,N_12349,N_12402);
xnor U12838 (N_12838,N_12455,N_12283);
nand U12839 (N_12839,N_12201,N_12289);
nor U12840 (N_12840,N_12487,N_12085);
nand U12841 (N_12841,N_12077,N_12256);
xor U12842 (N_12842,N_12411,N_12431);
and U12843 (N_12843,N_12089,N_12496);
nor U12844 (N_12844,N_12108,N_12385);
xor U12845 (N_12845,N_12297,N_12296);
xor U12846 (N_12846,N_12005,N_12129);
nand U12847 (N_12847,N_12394,N_12499);
nor U12848 (N_12848,N_12444,N_12155);
nand U12849 (N_12849,N_12192,N_12443);
and U12850 (N_12850,N_12423,N_12339);
nand U12851 (N_12851,N_12403,N_12091);
nand U12852 (N_12852,N_12400,N_12485);
xnor U12853 (N_12853,N_12199,N_12027);
nand U12854 (N_12854,N_12434,N_12080);
nor U12855 (N_12855,N_12126,N_12195);
xnor U12856 (N_12856,N_12105,N_12162);
nor U12857 (N_12857,N_12275,N_12303);
xnor U12858 (N_12858,N_12399,N_12491);
nand U12859 (N_12859,N_12388,N_12220);
or U12860 (N_12860,N_12158,N_12440);
and U12861 (N_12861,N_12288,N_12304);
nor U12862 (N_12862,N_12116,N_12074);
nand U12863 (N_12863,N_12481,N_12009);
or U12864 (N_12864,N_12358,N_12415);
nor U12865 (N_12865,N_12137,N_12369);
nor U12866 (N_12866,N_12495,N_12108);
and U12867 (N_12867,N_12316,N_12449);
nand U12868 (N_12868,N_12228,N_12404);
or U12869 (N_12869,N_12169,N_12471);
and U12870 (N_12870,N_12477,N_12438);
nor U12871 (N_12871,N_12380,N_12442);
or U12872 (N_12872,N_12134,N_12370);
or U12873 (N_12873,N_12147,N_12231);
and U12874 (N_12874,N_12141,N_12316);
and U12875 (N_12875,N_12211,N_12377);
nand U12876 (N_12876,N_12472,N_12280);
and U12877 (N_12877,N_12151,N_12342);
xnor U12878 (N_12878,N_12313,N_12429);
nand U12879 (N_12879,N_12423,N_12175);
nor U12880 (N_12880,N_12228,N_12306);
xnor U12881 (N_12881,N_12409,N_12098);
and U12882 (N_12882,N_12142,N_12358);
and U12883 (N_12883,N_12133,N_12063);
xnor U12884 (N_12884,N_12028,N_12477);
and U12885 (N_12885,N_12372,N_12337);
xor U12886 (N_12886,N_12229,N_12188);
xor U12887 (N_12887,N_12012,N_12431);
nor U12888 (N_12888,N_12138,N_12402);
nand U12889 (N_12889,N_12025,N_12191);
xnor U12890 (N_12890,N_12422,N_12029);
and U12891 (N_12891,N_12430,N_12234);
nand U12892 (N_12892,N_12437,N_12094);
xnor U12893 (N_12893,N_12183,N_12273);
xor U12894 (N_12894,N_12414,N_12024);
and U12895 (N_12895,N_12218,N_12423);
nand U12896 (N_12896,N_12109,N_12238);
xor U12897 (N_12897,N_12114,N_12484);
nand U12898 (N_12898,N_12262,N_12277);
nand U12899 (N_12899,N_12489,N_12057);
nand U12900 (N_12900,N_12163,N_12055);
nor U12901 (N_12901,N_12092,N_12204);
xor U12902 (N_12902,N_12096,N_12364);
xor U12903 (N_12903,N_12078,N_12350);
nand U12904 (N_12904,N_12227,N_12216);
nor U12905 (N_12905,N_12480,N_12417);
xnor U12906 (N_12906,N_12196,N_12222);
and U12907 (N_12907,N_12234,N_12287);
nand U12908 (N_12908,N_12117,N_12213);
and U12909 (N_12909,N_12404,N_12170);
or U12910 (N_12910,N_12446,N_12318);
xnor U12911 (N_12911,N_12328,N_12487);
or U12912 (N_12912,N_12279,N_12043);
xnor U12913 (N_12913,N_12347,N_12127);
nand U12914 (N_12914,N_12455,N_12029);
nor U12915 (N_12915,N_12356,N_12184);
xnor U12916 (N_12916,N_12336,N_12476);
or U12917 (N_12917,N_12161,N_12108);
nand U12918 (N_12918,N_12135,N_12191);
nand U12919 (N_12919,N_12463,N_12367);
nor U12920 (N_12920,N_12380,N_12006);
and U12921 (N_12921,N_12136,N_12348);
nand U12922 (N_12922,N_12153,N_12340);
xor U12923 (N_12923,N_12085,N_12230);
and U12924 (N_12924,N_12369,N_12075);
nand U12925 (N_12925,N_12483,N_12303);
xnor U12926 (N_12926,N_12203,N_12233);
or U12927 (N_12927,N_12308,N_12070);
and U12928 (N_12928,N_12234,N_12238);
xnor U12929 (N_12929,N_12279,N_12432);
nor U12930 (N_12930,N_12172,N_12448);
or U12931 (N_12931,N_12432,N_12182);
nor U12932 (N_12932,N_12123,N_12407);
nor U12933 (N_12933,N_12329,N_12109);
nor U12934 (N_12934,N_12460,N_12070);
nand U12935 (N_12935,N_12142,N_12354);
nor U12936 (N_12936,N_12493,N_12057);
and U12937 (N_12937,N_12056,N_12432);
nor U12938 (N_12938,N_12045,N_12238);
nand U12939 (N_12939,N_12395,N_12261);
and U12940 (N_12940,N_12013,N_12174);
nand U12941 (N_12941,N_12153,N_12325);
and U12942 (N_12942,N_12132,N_12163);
nor U12943 (N_12943,N_12173,N_12016);
and U12944 (N_12944,N_12277,N_12294);
nor U12945 (N_12945,N_12395,N_12275);
nor U12946 (N_12946,N_12178,N_12057);
or U12947 (N_12947,N_12088,N_12106);
nand U12948 (N_12948,N_12259,N_12133);
nor U12949 (N_12949,N_12229,N_12343);
or U12950 (N_12950,N_12352,N_12406);
and U12951 (N_12951,N_12197,N_12137);
and U12952 (N_12952,N_12224,N_12063);
nand U12953 (N_12953,N_12290,N_12380);
xnor U12954 (N_12954,N_12371,N_12334);
and U12955 (N_12955,N_12425,N_12459);
or U12956 (N_12956,N_12478,N_12221);
xor U12957 (N_12957,N_12297,N_12086);
xor U12958 (N_12958,N_12032,N_12384);
or U12959 (N_12959,N_12366,N_12006);
or U12960 (N_12960,N_12020,N_12179);
xnor U12961 (N_12961,N_12439,N_12072);
nand U12962 (N_12962,N_12393,N_12151);
xor U12963 (N_12963,N_12187,N_12493);
xor U12964 (N_12964,N_12243,N_12298);
or U12965 (N_12965,N_12041,N_12127);
or U12966 (N_12966,N_12219,N_12325);
xnor U12967 (N_12967,N_12108,N_12363);
xor U12968 (N_12968,N_12226,N_12015);
nor U12969 (N_12969,N_12237,N_12257);
or U12970 (N_12970,N_12256,N_12331);
nand U12971 (N_12971,N_12007,N_12196);
xnor U12972 (N_12972,N_12229,N_12428);
xor U12973 (N_12973,N_12234,N_12167);
and U12974 (N_12974,N_12342,N_12455);
nor U12975 (N_12975,N_12368,N_12405);
nor U12976 (N_12976,N_12080,N_12439);
and U12977 (N_12977,N_12032,N_12187);
or U12978 (N_12978,N_12120,N_12465);
nor U12979 (N_12979,N_12369,N_12385);
nor U12980 (N_12980,N_12373,N_12116);
and U12981 (N_12981,N_12246,N_12319);
or U12982 (N_12982,N_12043,N_12119);
xor U12983 (N_12983,N_12213,N_12256);
xor U12984 (N_12984,N_12014,N_12265);
or U12985 (N_12985,N_12162,N_12190);
and U12986 (N_12986,N_12026,N_12206);
xnor U12987 (N_12987,N_12027,N_12164);
and U12988 (N_12988,N_12306,N_12478);
or U12989 (N_12989,N_12442,N_12156);
xor U12990 (N_12990,N_12107,N_12283);
and U12991 (N_12991,N_12107,N_12115);
and U12992 (N_12992,N_12407,N_12069);
and U12993 (N_12993,N_12173,N_12200);
and U12994 (N_12994,N_12461,N_12354);
and U12995 (N_12995,N_12173,N_12100);
xnor U12996 (N_12996,N_12355,N_12248);
xnor U12997 (N_12997,N_12328,N_12442);
nand U12998 (N_12998,N_12148,N_12447);
or U12999 (N_12999,N_12345,N_12304);
or U13000 (N_13000,N_12802,N_12648);
and U13001 (N_13001,N_12930,N_12841);
xnor U13002 (N_13002,N_12625,N_12753);
or U13003 (N_13003,N_12966,N_12565);
or U13004 (N_13004,N_12993,N_12917);
nand U13005 (N_13005,N_12830,N_12618);
nand U13006 (N_13006,N_12752,N_12867);
xor U13007 (N_13007,N_12956,N_12513);
or U13008 (N_13008,N_12738,N_12939);
or U13009 (N_13009,N_12835,N_12736);
nand U13010 (N_13010,N_12673,N_12554);
and U13011 (N_13011,N_12793,N_12903);
or U13012 (N_13012,N_12622,N_12872);
or U13013 (N_13013,N_12571,N_12636);
nand U13014 (N_13014,N_12574,N_12711);
xnor U13015 (N_13015,N_12696,N_12539);
and U13016 (N_13016,N_12984,N_12986);
and U13017 (N_13017,N_12613,N_12931);
xnor U13018 (N_13018,N_12656,N_12639);
or U13019 (N_13019,N_12954,N_12932);
nor U13020 (N_13020,N_12786,N_12681);
xnor U13021 (N_13021,N_12628,N_12935);
nor U13022 (N_13022,N_12808,N_12923);
xor U13023 (N_13023,N_12694,N_12688);
and U13024 (N_13024,N_12972,N_12858);
and U13025 (N_13025,N_12739,N_12607);
nor U13026 (N_13026,N_12719,N_12703);
nand U13027 (N_13027,N_12655,N_12937);
or U13028 (N_13028,N_12627,N_12896);
or U13029 (N_13029,N_12838,N_12992);
and U13030 (N_13030,N_12723,N_12644);
or U13031 (N_13031,N_12887,N_12970);
nand U13032 (N_13032,N_12927,N_12947);
nand U13033 (N_13033,N_12654,N_12633);
or U13034 (N_13034,N_12647,N_12891);
and U13035 (N_13035,N_12596,N_12997);
or U13036 (N_13036,N_12682,N_12505);
nand U13037 (N_13037,N_12806,N_12729);
and U13038 (N_13038,N_12536,N_12785);
nor U13039 (N_13039,N_12781,N_12704);
xnor U13040 (N_13040,N_12632,N_12812);
nor U13041 (N_13041,N_12726,N_12518);
xor U13042 (N_13042,N_12934,N_12717);
nand U13043 (N_13043,N_12591,N_12826);
and U13044 (N_13044,N_12965,N_12669);
nand U13045 (N_13045,N_12832,N_12905);
xnor U13046 (N_13046,N_12816,N_12801);
xnor U13047 (N_13047,N_12900,N_12728);
nor U13048 (N_13048,N_12698,N_12991);
nand U13049 (N_13049,N_12573,N_12883);
or U13050 (N_13050,N_12908,N_12646);
and U13051 (N_13051,N_12549,N_12784);
nor U13052 (N_13052,N_12585,N_12843);
and U13053 (N_13053,N_12674,N_12779);
nor U13054 (N_13054,N_12778,N_12760);
nand U13055 (N_13055,N_12665,N_12770);
nand U13056 (N_13056,N_12584,N_12515);
xor U13057 (N_13057,N_12548,N_12706);
or U13058 (N_13058,N_12678,N_12857);
xor U13059 (N_13059,N_12777,N_12910);
nand U13060 (N_13060,N_12963,N_12718);
nand U13061 (N_13061,N_12895,N_12837);
or U13062 (N_13062,N_12996,N_12512);
and U13063 (N_13063,N_12767,N_12823);
and U13064 (N_13064,N_12960,N_12790);
xor U13065 (N_13065,N_12948,N_12886);
or U13066 (N_13066,N_12980,N_12873);
nor U13067 (N_13067,N_12707,N_12995);
xnor U13068 (N_13068,N_12720,N_12773);
and U13069 (N_13069,N_12897,N_12868);
nor U13070 (N_13070,N_12922,N_12672);
nor U13071 (N_13071,N_12985,N_12564);
and U13072 (N_13072,N_12893,N_12615);
nand U13073 (N_13073,N_12904,N_12533);
or U13074 (N_13074,N_12982,N_12683);
nand U13075 (N_13075,N_12977,N_12881);
or U13076 (N_13076,N_12884,N_12504);
nor U13077 (N_13077,N_12503,N_12761);
xnor U13078 (N_13078,N_12606,N_12671);
and U13079 (N_13079,N_12730,N_12799);
nand U13080 (N_13080,N_12560,N_12815);
or U13081 (N_13081,N_12611,N_12999);
nand U13082 (N_13082,N_12880,N_12936);
or U13083 (N_13083,N_12556,N_12814);
nor U13084 (N_13084,N_12701,N_12747);
and U13085 (N_13085,N_12994,N_12545);
and U13086 (N_13086,N_12551,N_12700);
nor U13087 (N_13087,N_12959,N_12710);
and U13088 (N_13088,N_12938,N_12661);
nand U13089 (N_13089,N_12553,N_12679);
xor U13090 (N_13090,N_12949,N_12530);
or U13091 (N_13091,N_12612,N_12740);
nand U13092 (N_13092,N_12769,N_12928);
or U13093 (N_13093,N_12863,N_12563);
and U13094 (N_13094,N_12501,N_12609);
nand U13095 (N_13095,N_12820,N_12940);
xor U13096 (N_13096,N_12919,N_12697);
or U13097 (N_13097,N_12750,N_12663);
or U13098 (N_13098,N_12692,N_12525);
xor U13099 (N_13099,N_12676,N_12805);
and U13100 (N_13100,N_12875,N_12541);
xnor U13101 (N_13101,N_12955,N_12526);
nand U13102 (N_13102,N_12798,N_12668);
nor U13103 (N_13103,N_12540,N_12732);
nor U13104 (N_13104,N_12978,N_12855);
nand U13105 (N_13105,N_12929,N_12918);
and U13106 (N_13106,N_12637,N_12942);
or U13107 (N_13107,N_12580,N_12754);
nor U13108 (N_13108,N_12594,N_12831);
nor U13109 (N_13109,N_12925,N_12755);
and U13110 (N_13110,N_12856,N_12521);
xnor U13111 (N_13111,N_12537,N_12776);
nor U13112 (N_13112,N_12522,N_12677);
and U13113 (N_13113,N_12791,N_12666);
or U13114 (N_13114,N_12662,N_12667);
or U13115 (N_13115,N_12762,N_12593);
and U13116 (N_13116,N_12557,N_12691);
nand U13117 (N_13117,N_12527,N_12902);
nand U13118 (N_13118,N_12705,N_12950);
xor U13119 (N_13119,N_12714,N_12976);
xor U13120 (N_13120,N_12507,N_12601);
xnor U13121 (N_13121,N_12913,N_12829);
nor U13122 (N_13122,N_12699,N_12825);
nor U13123 (N_13123,N_12854,N_12953);
nand U13124 (N_13124,N_12828,N_12734);
nor U13125 (N_13125,N_12589,N_12568);
nand U13126 (N_13126,N_12869,N_12810);
and U13127 (N_13127,N_12797,N_12890);
or U13128 (N_13128,N_12559,N_12708);
or U13129 (N_13129,N_12968,N_12821);
xor U13130 (N_13130,N_12653,N_12975);
nor U13131 (N_13131,N_12532,N_12592);
nor U13132 (N_13132,N_12725,N_12836);
xor U13133 (N_13133,N_12642,N_12765);
or U13134 (N_13134,N_12787,N_12885);
xor U13135 (N_13135,N_12610,N_12840);
and U13136 (N_13136,N_12619,N_12794);
or U13137 (N_13137,N_12689,N_12864);
and U13138 (N_13138,N_12690,N_12620);
nand U13139 (N_13139,N_12638,N_12933);
nand U13140 (N_13140,N_12575,N_12743);
nand U13141 (N_13141,N_12749,N_12795);
nand U13142 (N_13142,N_12952,N_12624);
nand U13143 (N_13143,N_12882,N_12614);
nor U13144 (N_13144,N_12983,N_12684);
nor U13145 (N_13145,N_12561,N_12626);
and U13146 (N_13146,N_12608,N_12783);
and U13147 (N_13147,N_12898,N_12715);
and U13148 (N_13148,N_12531,N_12722);
and U13149 (N_13149,N_12889,N_12675);
xnor U13150 (N_13150,N_12879,N_12538);
or U13151 (N_13151,N_12617,N_12578);
and U13152 (N_13152,N_12604,N_12981);
and U13153 (N_13153,N_12848,N_12788);
or U13154 (N_13154,N_12988,N_12969);
or U13155 (N_13155,N_12542,N_12543);
and U13156 (N_13156,N_12870,N_12915);
nor U13157 (N_13157,N_12724,N_12866);
or U13158 (N_13158,N_12772,N_12660);
nor U13159 (N_13159,N_12766,N_12780);
or U13160 (N_13160,N_12861,N_12758);
and U13161 (N_13161,N_12789,N_12957);
xnor U13162 (N_13162,N_12641,N_12894);
nor U13163 (N_13163,N_12588,N_12631);
and U13164 (N_13164,N_12876,N_12813);
or U13165 (N_13165,N_12586,N_12595);
nand U13166 (N_13166,N_12817,N_12800);
nand U13167 (N_13167,N_12603,N_12599);
xnor U13168 (N_13168,N_12524,N_12774);
and U13169 (N_13169,N_12845,N_12844);
xor U13170 (N_13170,N_12598,N_12756);
or U13171 (N_13171,N_12558,N_12500);
nand U13172 (N_13172,N_12569,N_12746);
xor U13173 (N_13173,N_12693,N_12721);
xor U13174 (N_13174,N_12748,N_12892);
xnor U13175 (N_13175,N_12664,N_12842);
and U13176 (N_13176,N_12967,N_12818);
or U13177 (N_13177,N_12634,N_12712);
xor U13178 (N_13178,N_12519,N_12916);
nand U13179 (N_13179,N_12579,N_12782);
xnor U13180 (N_13180,N_12745,N_12643);
nand U13181 (N_13181,N_12834,N_12649);
and U13182 (N_13182,N_12751,N_12888);
or U13183 (N_13183,N_12912,N_12964);
or U13184 (N_13184,N_12713,N_12909);
nand U13185 (N_13185,N_12878,N_12846);
xnor U13186 (N_13186,N_12901,N_12582);
or U13187 (N_13187,N_12944,N_12852);
and U13188 (N_13188,N_12796,N_12853);
nor U13189 (N_13189,N_12597,N_12506);
and U13190 (N_13190,N_12602,N_12635);
nor U13191 (N_13191,N_12695,N_12943);
xor U13192 (N_13192,N_12502,N_12528);
nand U13193 (N_13193,N_12979,N_12973);
nor U13194 (N_13194,N_12517,N_12827);
nor U13195 (N_13195,N_12514,N_12529);
or U13196 (N_13196,N_12733,N_12998);
xnor U13197 (N_13197,N_12651,N_12847);
or U13198 (N_13198,N_12576,N_12792);
nand U13199 (N_13199,N_12581,N_12680);
xor U13200 (N_13200,N_12971,N_12907);
xor U13201 (N_13201,N_12851,N_12562);
nand U13202 (N_13202,N_12811,N_12871);
nand U13203 (N_13203,N_12946,N_12990);
nand U13204 (N_13204,N_12819,N_12865);
and U13205 (N_13205,N_12621,N_12763);
or U13206 (N_13206,N_12824,N_12658);
and U13207 (N_13207,N_12555,N_12616);
nand U13208 (N_13208,N_12544,N_12659);
and U13209 (N_13209,N_12546,N_12630);
and U13210 (N_13210,N_12583,N_12716);
xor U13211 (N_13211,N_12640,N_12906);
nand U13212 (N_13212,N_12516,N_12727);
and U13213 (N_13213,N_12987,N_12652);
nor U13214 (N_13214,N_12657,N_12804);
nor U13215 (N_13215,N_12803,N_12687);
nand U13216 (N_13216,N_12702,N_12862);
nand U13217 (N_13217,N_12914,N_12771);
nand U13218 (N_13218,N_12709,N_12961);
and U13219 (N_13219,N_12764,N_12552);
or U13220 (N_13220,N_12570,N_12850);
nor U13221 (N_13221,N_12744,N_12511);
or U13222 (N_13222,N_12520,N_12775);
nand U13223 (N_13223,N_12566,N_12742);
or U13224 (N_13224,N_12833,N_12509);
and U13225 (N_13225,N_12590,N_12577);
nor U13226 (N_13226,N_12523,N_12629);
nand U13227 (N_13227,N_12534,N_12550);
nand U13228 (N_13228,N_12757,N_12650);
nor U13229 (N_13229,N_12962,N_12510);
nand U13230 (N_13230,N_12759,N_12859);
nor U13231 (N_13231,N_12768,N_12874);
nand U13232 (N_13232,N_12839,N_12547);
nor U13233 (N_13233,N_12572,N_12924);
and U13234 (N_13234,N_12741,N_12809);
nor U13235 (N_13235,N_12600,N_12567);
and U13236 (N_13236,N_12535,N_12941);
xor U13237 (N_13237,N_12958,N_12645);
or U13238 (N_13238,N_12974,N_12508);
nand U13239 (N_13239,N_12686,N_12926);
nor U13240 (N_13240,N_12587,N_12899);
xor U13241 (N_13241,N_12877,N_12685);
or U13242 (N_13242,N_12911,N_12849);
and U13243 (N_13243,N_12989,N_12737);
and U13244 (N_13244,N_12860,N_12735);
nor U13245 (N_13245,N_12921,N_12951);
nand U13246 (N_13246,N_12670,N_12920);
xnor U13247 (N_13247,N_12623,N_12945);
nor U13248 (N_13248,N_12807,N_12731);
nor U13249 (N_13249,N_12605,N_12822);
and U13250 (N_13250,N_12588,N_12698);
xnor U13251 (N_13251,N_12868,N_12816);
nor U13252 (N_13252,N_12687,N_12633);
nand U13253 (N_13253,N_12898,N_12886);
xnor U13254 (N_13254,N_12908,N_12774);
nor U13255 (N_13255,N_12876,N_12758);
or U13256 (N_13256,N_12571,N_12939);
nor U13257 (N_13257,N_12579,N_12643);
and U13258 (N_13258,N_12682,N_12544);
and U13259 (N_13259,N_12716,N_12641);
xor U13260 (N_13260,N_12712,N_12618);
xnor U13261 (N_13261,N_12801,N_12856);
nand U13262 (N_13262,N_12559,N_12960);
nor U13263 (N_13263,N_12593,N_12597);
nor U13264 (N_13264,N_12965,N_12835);
nor U13265 (N_13265,N_12719,N_12843);
and U13266 (N_13266,N_12508,N_12998);
or U13267 (N_13267,N_12581,N_12935);
or U13268 (N_13268,N_12594,N_12837);
nand U13269 (N_13269,N_12786,N_12654);
or U13270 (N_13270,N_12575,N_12776);
nor U13271 (N_13271,N_12864,N_12678);
xnor U13272 (N_13272,N_12987,N_12810);
or U13273 (N_13273,N_12608,N_12897);
nor U13274 (N_13274,N_12785,N_12819);
and U13275 (N_13275,N_12564,N_12581);
nor U13276 (N_13276,N_12655,N_12921);
xor U13277 (N_13277,N_12678,N_12978);
xnor U13278 (N_13278,N_12882,N_12644);
nand U13279 (N_13279,N_12793,N_12778);
nand U13280 (N_13280,N_12787,N_12775);
nor U13281 (N_13281,N_12500,N_12952);
or U13282 (N_13282,N_12506,N_12598);
nor U13283 (N_13283,N_12684,N_12903);
or U13284 (N_13284,N_12888,N_12665);
nor U13285 (N_13285,N_12768,N_12511);
nor U13286 (N_13286,N_12696,N_12995);
nor U13287 (N_13287,N_12828,N_12519);
or U13288 (N_13288,N_12845,N_12853);
nor U13289 (N_13289,N_12897,N_12701);
xor U13290 (N_13290,N_12851,N_12848);
nand U13291 (N_13291,N_12826,N_12597);
nor U13292 (N_13292,N_12639,N_12633);
nor U13293 (N_13293,N_12964,N_12588);
and U13294 (N_13294,N_12774,N_12789);
xnor U13295 (N_13295,N_12710,N_12998);
xnor U13296 (N_13296,N_12750,N_12811);
and U13297 (N_13297,N_12683,N_12527);
nor U13298 (N_13298,N_12723,N_12645);
or U13299 (N_13299,N_12935,N_12999);
nor U13300 (N_13300,N_12631,N_12594);
nor U13301 (N_13301,N_12898,N_12521);
or U13302 (N_13302,N_12576,N_12538);
or U13303 (N_13303,N_12954,N_12814);
nor U13304 (N_13304,N_12719,N_12866);
nand U13305 (N_13305,N_12551,N_12968);
or U13306 (N_13306,N_12640,N_12769);
and U13307 (N_13307,N_12669,N_12619);
nand U13308 (N_13308,N_12829,N_12784);
or U13309 (N_13309,N_12744,N_12607);
nor U13310 (N_13310,N_12856,N_12845);
or U13311 (N_13311,N_12562,N_12720);
xnor U13312 (N_13312,N_12507,N_12801);
xor U13313 (N_13313,N_12849,N_12603);
nor U13314 (N_13314,N_12666,N_12653);
xor U13315 (N_13315,N_12568,N_12756);
and U13316 (N_13316,N_12726,N_12962);
nand U13317 (N_13317,N_12526,N_12541);
nor U13318 (N_13318,N_12539,N_12622);
or U13319 (N_13319,N_12770,N_12515);
nand U13320 (N_13320,N_12655,N_12595);
or U13321 (N_13321,N_12821,N_12862);
nand U13322 (N_13322,N_12660,N_12788);
nand U13323 (N_13323,N_12816,N_12624);
or U13324 (N_13324,N_12756,N_12525);
nand U13325 (N_13325,N_12950,N_12902);
nor U13326 (N_13326,N_12987,N_12892);
xnor U13327 (N_13327,N_12608,N_12843);
nand U13328 (N_13328,N_12988,N_12800);
nor U13329 (N_13329,N_12721,N_12744);
xnor U13330 (N_13330,N_12940,N_12626);
or U13331 (N_13331,N_12820,N_12639);
and U13332 (N_13332,N_12917,N_12949);
nor U13333 (N_13333,N_12510,N_12545);
and U13334 (N_13334,N_12748,N_12844);
xor U13335 (N_13335,N_12725,N_12910);
xor U13336 (N_13336,N_12959,N_12942);
nor U13337 (N_13337,N_12508,N_12986);
or U13338 (N_13338,N_12680,N_12969);
nand U13339 (N_13339,N_12598,N_12709);
nand U13340 (N_13340,N_12659,N_12723);
xor U13341 (N_13341,N_12773,N_12594);
nand U13342 (N_13342,N_12524,N_12659);
nand U13343 (N_13343,N_12780,N_12867);
nand U13344 (N_13344,N_12798,N_12619);
xor U13345 (N_13345,N_12783,N_12672);
nor U13346 (N_13346,N_12581,N_12597);
nand U13347 (N_13347,N_12921,N_12679);
and U13348 (N_13348,N_12909,N_12733);
or U13349 (N_13349,N_12588,N_12644);
and U13350 (N_13350,N_12846,N_12736);
nand U13351 (N_13351,N_12769,N_12983);
and U13352 (N_13352,N_12744,N_12655);
and U13353 (N_13353,N_12991,N_12930);
nor U13354 (N_13354,N_12591,N_12817);
nand U13355 (N_13355,N_12597,N_12773);
or U13356 (N_13356,N_12926,N_12746);
nor U13357 (N_13357,N_12761,N_12828);
or U13358 (N_13358,N_12945,N_12671);
nor U13359 (N_13359,N_12777,N_12916);
and U13360 (N_13360,N_12683,N_12619);
and U13361 (N_13361,N_12553,N_12657);
and U13362 (N_13362,N_12759,N_12690);
xor U13363 (N_13363,N_12978,N_12663);
and U13364 (N_13364,N_12656,N_12602);
nor U13365 (N_13365,N_12734,N_12590);
nor U13366 (N_13366,N_12803,N_12517);
and U13367 (N_13367,N_12825,N_12598);
xor U13368 (N_13368,N_12726,N_12500);
nor U13369 (N_13369,N_12834,N_12980);
xnor U13370 (N_13370,N_12779,N_12550);
nor U13371 (N_13371,N_12668,N_12915);
xor U13372 (N_13372,N_12740,N_12974);
and U13373 (N_13373,N_12780,N_12834);
nand U13374 (N_13374,N_12991,N_12584);
xnor U13375 (N_13375,N_12871,N_12606);
nor U13376 (N_13376,N_12779,N_12576);
nor U13377 (N_13377,N_12913,N_12881);
xor U13378 (N_13378,N_12999,N_12735);
or U13379 (N_13379,N_12509,N_12944);
and U13380 (N_13380,N_12552,N_12966);
xnor U13381 (N_13381,N_12717,N_12743);
nor U13382 (N_13382,N_12664,N_12539);
xnor U13383 (N_13383,N_12741,N_12667);
nand U13384 (N_13384,N_12865,N_12591);
and U13385 (N_13385,N_12777,N_12574);
or U13386 (N_13386,N_12765,N_12874);
or U13387 (N_13387,N_12619,N_12665);
nand U13388 (N_13388,N_12612,N_12938);
or U13389 (N_13389,N_12955,N_12974);
xnor U13390 (N_13390,N_12917,N_12567);
nand U13391 (N_13391,N_12535,N_12886);
nand U13392 (N_13392,N_12772,N_12786);
nand U13393 (N_13393,N_12882,N_12951);
xor U13394 (N_13394,N_12873,N_12763);
xnor U13395 (N_13395,N_12598,N_12828);
or U13396 (N_13396,N_12502,N_12623);
and U13397 (N_13397,N_12588,N_12558);
and U13398 (N_13398,N_12554,N_12992);
and U13399 (N_13399,N_12715,N_12524);
or U13400 (N_13400,N_12760,N_12672);
or U13401 (N_13401,N_12899,N_12841);
and U13402 (N_13402,N_12625,N_12562);
nand U13403 (N_13403,N_12990,N_12686);
and U13404 (N_13404,N_12717,N_12696);
xor U13405 (N_13405,N_12665,N_12980);
nand U13406 (N_13406,N_12575,N_12586);
and U13407 (N_13407,N_12808,N_12595);
or U13408 (N_13408,N_12598,N_12645);
nor U13409 (N_13409,N_12875,N_12914);
and U13410 (N_13410,N_12985,N_12881);
nor U13411 (N_13411,N_12645,N_12693);
and U13412 (N_13412,N_12671,N_12952);
and U13413 (N_13413,N_12761,N_12820);
xnor U13414 (N_13414,N_12892,N_12797);
or U13415 (N_13415,N_12928,N_12529);
and U13416 (N_13416,N_12688,N_12547);
or U13417 (N_13417,N_12791,N_12998);
xnor U13418 (N_13418,N_12814,N_12696);
nand U13419 (N_13419,N_12930,N_12917);
nand U13420 (N_13420,N_12571,N_12603);
and U13421 (N_13421,N_12534,N_12504);
and U13422 (N_13422,N_12930,N_12578);
nand U13423 (N_13423,N_12768,N_12579);
xor U13424 (N_13424,N_12588,N_12984);
or U13425 (N_13425,N_12860,N_12820);
and U13426 (N_13426,N_12930,N_12640);
nor U13427 (N_13427,N_12624,N_12976);
xor U13428 (N_13428,N_12710,N_12672);
and U13429 (N_13429,N_12676,N_12806);
or U13430 (N_13430,N_12928,N_12584);
nand U13431 (N_13431,N_12867,N_12879);
nand U13432 (N_13432,N_12787,N_12723);
nand U13433 (N_13433,N_12758,N_12598);
or U13434 (N_13434,N_12630,N_12619);
nor U13435 (N_13435,N_12697,N_12973);
nor U13436 (N_13436,N_12801,N_12948);
xnor U13437 (N_13437,N_12552,N_12557);
or U13438 (N_13438,N_12875,N_12967);
and U13439 (N_13439,N_12626,N_12725);
nand U13440 (N_13440,N_12872,N_12778);
or U13441 (N_13441,N_12901,N_12601);
and U13442 (N_13442,N_12630,N_12542);
nand U13443 (N_13443,N_12532,N_12522);
xnor U13444 (N_13444,N_12984,N_12823);
nor U13445 (N_13445,N_12580,N_12927);
xor U13446 (N_13446,N_12652,N_12567);
or U13447 (N_13447,N_12860,N_12672);
xor U13448 (N_13448,N_12840,N_12748);
nand U13449 (N_13449,N_12565,N_12979);
nor U13450 (N_13450,N_12584,N_12500);
nand U13451 (N_13451,N_12917,N_12676);
and U13452 (N_13452,N_12924,N_12816);
xnor U13453 (N_13453,N_12806,N_12507);
or U13454 (N_13454,N_12789,N_12924);
xnor U13455 (N_13455,N_12824,N_12605);
nand U13456 (N_13456,N_12633,N_12728);
or U13457 (N_13457,N_12604,N_12999);
or U13458 (N_13458,N_12514,N_12988);
and U13459 (N_13459,N_12871,N_12689);
nand U13460 (N_13460,N_12760,N_12544);
and U13461 (N_13461,N_12741,N_12736);
xnor U13462 (N_13462,N_12909,N_12591);
and U13463 (N_13463,N_12552,N_12927);
nor U13464 (N_13464,N_12677,N_12784);
xnor U13465 (N_13465,N_12533,N_12519);
nand U13466 (N_13466,N_12664,N_12815);
and U13467 (N_13467,N_12798,N_12790);
nor U13468 (N_13468,N_12839,N_12503);
nor U13469 (N_13469,N_12766,N_12946);
xnor U13470 (N_13470,N_12514,N_12972);
nor U13471 (N_13471,N_12855,N_12646);
nor U13472 (N_13472,N_12571,N_12851);
nor U13473 (N_13473,N_12618,N_12946);
nor U13474 (N_13474,N_12636,N_12559);
nand U13475 (N_13475,N_12903,N_12889);
or U13476 (N_13476,N_12982,N_12693);
nand U13477 (N_13477,N_12772,N_12877);
nand U13478 (N_13478,N_12954,N_12502);
and U13479 (N_13479,N_12757,N_12864);
xnor U13480 (N_13480,N_12722,N_12547);
and U13481 (N_13481,N_12918,N_12815);
or U13482 (N_13482,N_12903,N_12625);
xor U13483 (N_13483,N_12622,N_12713);
xor U13484 (N_13484,N_12562,N_12931);
nor U13485 (N_13485,N_12795,N_12938);
and U13486 (N_13486,N_12783,N_12580);
nand U13487 (N_13487,N_12617,N_12999);
nor U13488 (N_13488,N_12615,N_12879);
and U13489 (N_13489,N_12663,N_12787);
nand U13490 (N_13490,N_12952,N_12868);
and U13491 (N_13491,N_12816,N_12948);
and U13492 (N_13492,N_12650,N_12763);
xnor U13493 (N_13493,N_12587,N_12938);
xor U13494 (N_13494,N_12838,N_12881);
xnor U13495 (N_13495,N_12890,N_12840);
nand U13496 (N_13496,N_12997,N_12597);
nand U13497 (N_13497,N_12501,N_12533);
nand U13498 (N_13498,N_12509,N_12565);
nand U13499 (N_13499,N_12528,N_12967);
and U13500 (N_13500,N_13309,N_13178);
xnor U13501 (N_13501,N_13156,N_13470);
nor U13502 (N_13502,N_13194,N_13247);
xor U13503 (N_13503,N_13191,N_13270);
or U13504 (N_13504,N_13232,N_13184);
or U13505 (N_13505,N_13196,N_13289);
xor U13506 (N_13506,N_13255,N_13003);
nor U13507 (N_13507,N_13324,N_13080);
nand U13508 (N_13508,N_13084,N_13154);
or U13509 (N_13509,N_13418,N_13095);
and U13510 (N_13510,N_13248,N_13085);
nand U13511 (N_13511,N_13376,N_13395);
xor U13512 (N_13512,N_13261,N_13441);
or U13513 (N_13513,N_13391,N_13164);
and U13514 (N_13514,N_13299,N_13158);
and U13515 (N_13515,N_13268,N_13139);
xor U13516 (N_13516,N_13235,N_13282);
xor U13517 (N_13517,N_13153,N_13367);
nand U13518 (N_13518,N_13373,N_13471);
and U13519 (N_13519,N_13416,N_13474);
and U13520 (N_13520,N_13362,N_13325);
xnor U13521 (N_13521,N_13203,N_13072);
xor U13522 (N_13522,N_13183,N_13461);
xnor U13523 (N_13523,N_13252,N_13071);
xnor U13524 (N_13524,N_13216,N_13348);
and U13525 (N_13525,N_13163,N_13368);
nand U13526 (N_13526,N_13382,N_13206);
and U13527 (N_13527,N_13166,N_13244);
nor U13528 (N_13528,N_13132,N_13228);
xor U13529 (N_13529,N_13039,N_13408);
or U13530 (N_13530,N_13176,N_13210);
nor U13531 (N_13531,N_13375,N_13338);
xnor U13532 (N_13532,N_13077,N_13295);
or U13533 (N_13533,N_13221,N_13093);
and U13534 (N_13534,N_13073,N_13300);
nor U13535 (N_13535,N_13025,N_13259);
nor U13536 (N_13536,N_13353,N_13466);
or U13537 (N_13537,N_13207,N_13243);
and U13538 (N_13538,N_13406,N_13114);
nand U13539 (N_13539,N_13401,N_13017);
xnor U13540 (N_13540,N_13070,N_13274);
nand U13541 (N_13541,N_13251,N_13069);
xnor U13542 (N_13542,N_13028,N_13054);
nand U13543 (N_13543,N_13396,N_13415);
and U13544 (N_13544,N_13107,N_13349);
or U13545 (N_13545,N_13143,N_13242);
nand U13546 (N_13546,N_13460,N_13030);
nand U13547 (N_13547,N_13287,N_13465);
xor U13548 (N_13548,N_13257,N_13056);
nand U13549 (N_13549,N_13222,N_13266);
nor U13550 (N_13550,N_13313,N_13004);
and U13551 (N_13551,N_13102,N_13245);
nor U13552 (N_13552,N_13220,N_13212);
nor U13553 (N_13553,N_13205,N_13484);
nor U13554 (N_13554,N_13439,N_13438);
xnor U13555 (N_13555,N_13403,N_13144);
and U13556 (N_13556,N_13010,N_13451);
nor U13557 (N_13557,N_13202,N_13480);
or U13558 (N_13558,N_13468,N_13001);
or U13559 (N_13559,N_13481,N_13078);
nor U13560 (N_13560,N_13414,N_13038);
and U13561 (N_13561,N_13286,N_13253);
nand U13562 (N_13562,N_13435,N_13464);
xor U13563 (N_13563,N_13197,N_13098);
and U13564 (N_13564,N_13423,N_13061);
nor U13565 (N_13565,N_13174,N_13113);
nand U13566 (N_13566,N_13490,N_13452);
nand U13567 (N_13567,N_13173,N_13074);
xor U13568 (N_13568,N_13089,N_13058);
xor U13569 (N_13569,N_13249,N_13021);
and U13570 (N_13570,N_13083,N_13260);
xor U13571 (N_13571,N_13246,N_13473);
nand U13572 (N_13572,N_13112,N_13230);
or U13573 (N_13573,N_13281,N_13227);
and U13574 (N_13574,N_13055,N_13298);
or U13575 (N_13575,N_13312,N_13379);
and U13576 (N_13576,N_13090,N_13135);
and U13577 (N_13577,N_13350,N_13137);
xnor U13578 (N_13578,N_13442,N_13020);
xnor U13579 (N_13579,N_13326,N_13491);
xor U13580 (N_13580,N_13272,N_13131);
xnor U13581 (N_13581,N_13489,N_13434);
xor U13582 (N_13582,N_13226,N_13343);
nand U13583 (N_13583,N_13192,N_13002);
and U13584 (N_13584,N_13366,N_13063);
nor U13585 (N_13585,N_13273,N_13024);
and U13586 (N_13586,N_13467,N_13447);
nand U13587 (N_13587,N_13427,N_13472);
and U13588 (N_13588,N_13327,N_13340);
and U13589 (N_13589,N_13339,N_13317);
nor U13590 (N_13590,N_13162,N_13456);
and U13591 (N_13591,N_13284,N_13032);
nand U13592 (N_13592,N_13407,N_13271);
xnor U13593 (N_13593,N_13128,N_13181);
xor U13594 (N_13594,N_13123,N_13487);
and U13595 (N_13595,N_13404,N_13269);
xnor U13596 (N_13596,N_13378,N_13031);
nor U13597 (N_13597,N_13359,N_13386);
and U13598 (N_13598,N_13400,N_13041);
or U13599 (N_13599,N_13431,N_13385);
nor U13600 (N_13600,N_13397,N_13081);
or U13601 (N_13601,N_13110,N_13262);
and U13602 (N_13602,N_13046,N_13458);
xor U13603 (N_13603,N_13351,N_13015);
and U13604 (N_13604,N_13433,N_13417);
nor U13605 (N_13605,N_13355,N_13424);
and U13606 (N_13606,N_13006,N_13172);
nand U13607 (N_13607,N_13053,N_13319);
and U13608 (N_13608,N_13280,N_13315);
and U13609 (N_13609,N_13167,N_13236);
nand U13610 (N_13610,N_13231,N_13264);
nand U13611 (N_13611,N_13168,N_13322);
or U13612 (N_13612,N_13432,N_13067);
and U13613 (N_13613,N_13399,N_13088);
and U13614 (N_13614,N_13023,N_13288);
and U13615 (N_13615,N_13377,N_13492);
or U13616 (N_13616,N_13180,N_13494);
nor U13617 (N_13617,N_13482,N_13405);
nand U13618 (N_13618,N_13008,N_13250);
nand U13619 (N_13619,N_13170,N_13346);
xnor U13620 (N_13620,N_13354,N_13169);
and U13621 (N_13621,N_13263,N_13372);
nand U13622 (N_13622,N_13337,N_13239);
nand U13623 (N_13623,N_13329,N_13332);
xor U13624 (N_13624,N_13022,N_13219);
xnor U13625 (N_13625,N_13277,N_13450);
and U13626 (N_13626,N_13064,N_13496);
or U13627 (N_13627,N_13308,N_13459);
and U13628 (N_13628,N_13483,N_13142);
and U13629 (N_13629,N_13103,N_13215);
or U13630 (N_13630,N_13240,N_13224);
nand U13631 (N_13631,N_13402,N_13106);
and U13632 (N_13632,N_13443,N_13237);
and U13633 (N_13633,N_13384,N_13422);
nor U13634 (N_13634,N_13426,N_13097);
nand U13635 (N_13635,N_13087,N_13413);
xnor U13636 (N_13636,N_13225,N_13394);
or U13637 (N_13637,N_13410,N_13291);
and U13638 (N_13638,N_13146,N_13347);
xor U13639 (N_13639,N_13233,N_13218);
or U13640 (N_13640,N_13420,N_13486);
or U13641 (N_13641,N_13119,N_13182);
xnor U13642 (N_13642,N_13276,N_13209);
and U13643 (N_13643,N_13043,N_13303);
or U13644 (N_13644,N_13152,N_13436);
xor U13645 (N_13645,N_13305,N_13149);
nor U13646 (N_13646,N_13013,N_13136);
or U13647 (N_13647,N_13296,N_13454);
nor U13648 (N_13648,N_13429,N_13120);
or U13649 (N_13649,N_13175,N_13374);
and U13650 (N_13650,N_13201,N_13334);
nand U13651 (N_13651,N_13425,N_13390);
and U13652 (N_13652,N_13499,N_13306);
and U13653 (N_13653,N_13371,N_13393);
and U13654 (N_13654,N_13094,N_13099);
and U13655 (N_13655,N_13241,N_13488);
and U13656 (N_13656,N_13117,N_13051);
and U13657 (N_13657,N_13147,N_13057);
nand U13658 (N_13658,N_13141,N_13133);
xnor U13659 (N_13659,N_13159,N_13370);
or U13660 (N_13660,N_13485,N_13014);
nand U13661 (N_13661,N_13333,N_13336);
and U13662 (N_13662,N_13040,N_13050);
nor U13663 (N_13663,N_13437,N_13344);
nor U13664 (N_13664,N_13208,N_13389);
xor U13665 (N_13665,N_13285,N_13108);
or U13666 (N_13666,N_13294,N_13320);
nor U13667 (N_13667,N_13138,N_13316);
nand U13668 (N_13668,N_13392,N_13462);
or U13669 (N_13669,N_13318,N_13195);
nand U13670 (N_13670,N_13211,N_13047);
nor U13671 (N_13671,N_13495,N_13331);
nor U13672 (N_13672,N_13140,N_13186);
nand U13673 (N_13673,N_13200,N_13311);
xor U13674 (N_13674,N_13335,N_13412);
nor U13675 (N_13675,N_13189,N_13477);
nand U13676 (N_13676,N_13027,N_13160);
and U13677 (N_13677,N_13304,N_13035);
xor U13678 (N_13678,N_13357,N_13005);
or U13679 (N_13679,N_13387,N_13104);
nor U13680 (N_13680,N_13301,N_13364);
xnor U13681 (N_13681,N_13079,N_13217);
or U13682 (N_13682,N_13042,N_13165);
or U13683 (N_13683,N_13341,N_13121);
nand U13684 (N_13684,N_13048,N_13440);
or U13685 (N_13685,N_13044,N_13115);
xor U13686 (N_13686,N_13428,N_13129);
and U13687 (N_13687,N_13049,N_13234);
nand U13688 (N_13688,N_13185,N_13475);
nand U13689 (N_13689,N_13265,N_13292);
xor U13690 (N_13690,N_13029,N_13100);
and U13691 (N_13691,N_13111,N_13118);
or U13692 (N_13692,N_13016,N_13302);
nor U13693 (N_13693,N_13122,N_13125);
nand U13694 (N_13694,N_13190,N_13290);
nor U13695 (N_13695,N_13062,N_13009);
nor U13696 (N_13696,N_13076,N_13254);
nand U13697 (N_13697,N_13199,N_13476);
nand U13698 (N_13698,N_13096,N_13469);
xnor U13699 (N_13699,N_13369,N_13238);
or U13700 (N_13700,N_13297,N_13150);
nor U13701 (N_13701,N_13321,N_13279);
or U13702 (N_13702,N_13161,N_13068);
xnor U13703 (N_13703,N_13398,N_13179);
and U13704 (N_13704,N_13026,N_13036);
nor U13705 (N_13705,N_13453,N_13409);
nand U13706 (N_13706,N_13307,N_13479);
xor U13707 (N_13707,N_13019,N_13000);
nand U13708 (N_13708,N_13109,N_13330);
xnor U13709 (N_13709,N_13478,N_13449);
and U13710 (N_13710,N_13360,N_13342);
nand U13711 (N_13711,N_13198,N_13092);
nor U13712 (N_13712,N_13223,N_13145);
and U13713 (N_13713,N_13445,N_13011);
or U13714 (N_13714,N_13086,N_13157);
xnor U13715 (N_13715,N_13105,N_13059);
and U13716 (N_13716,N_13034,N_13381);
xor U13717 (N_13717,N_13012,N_13116);
nor U13718 (N_13718,N_13323,N_13388);
nor U13719 (N_13719,N_13148,N_13411);
nand U13720 (N_13720,N_13421,N_13124);
xor U13721 (N_13721,N_13126,N_13018);
and U13722 (N_13722,N_13075,N_13091);
and U13723 (N_13723,N_13258,N_13497);
or U13724 (N_13724,N_13363,N_13033);
nor U13725 (N_13725,N_13463,N_13127);
or U13726 (N_13726,N_13204,N_13293);
xnor U13727 (N_13727,N_13151,N_13134);
xor U13728 (N_13728,N_13187,N_13155);
nor U13729 (N_13729,N_13358,N_13213);
or U13730 (N_13730,N_13345,N_13101);
nor U13731 (N_13731,N_13446,N_13060);
and U13732 (N_13732,N_13007,N_13498);
xnor U13733 (N_13733,N_13052,N_13082);
and U13734 (N_13734,N_13066,N_13352);
and U13735 (N_13735,N_13310,N_13214);
and U13736 (N_13736,N_13229,N_13193);
nor U13737 (N_13737,N_13419,N_13448);
nand U13738 (N_13738,N_13130,N_13037);
nand U13739 (N_13739,N_13188,N_13328);
nor U13740 (N_13740,N_13457,N_13278);
nand U13741 (N_13741,N_13177,N_13430);
and U13742 (N_13742,N_13045,N_13356);
xor U13743 (N_13743,N_13380,N_13455);
xor U13744 (N_13744,N_13383,N_13361);
nor U13745 (N_13745,N_13493,N_13444);
xnor U13746 (N_13746,N_13365,N_13314);
xor U13747 (N_13747,N_13283,N_13267);
nor U13748 (N_13748,N_13065,N_13171);
xor U13749 (N_13749,N_13275,N_13256);
or U13750 (N_13750,N_13068,N_13040);
nand U13751 (N_13751,N_13497,N_13318);
and U13752 (N_13752,N_13391,N_13483);
nand U13753 (N_13753,N_13025,N_13053);
nand U13754 (N_13754,N_13370,N_13389);
and U13755 (N_13755,N_13063,N_13221);
xor U13756 (N_13756,N_13006,N_13133);
nand U13757 (N_13757,N_13319,N_13234);
or U13758 (N_13758,N_13282,N_13396);
xor U13759 (N_13759,N_13111,N_13122);
or U13760 (N_13760,N_13300,N_13038);
nand U13761 (N_13761,N_13453,N_13080);
or U13762 (N_13762,N_13284,N_13271);
nor U13763 (N_13763,N_13459,N_13202);
xnor U13764 (N_13764,N_13373,N_13429);
nand U13765 (N_13765,N_13179,N_13407);
xnor U13766 (N_13766,N_13013,N_13015);
nand U13767 (N_13767,N_13143,N_13094);
nand U13768 (N_13768,N_13032,N_13425);
nand U13769 (N_13769,N_13086,N_13301);
nand U13770 (N_13770,N_13485,N_13106);
nor U13771 (N_13771,N_13070,N_13383);
nand U13772 (N_13772,N_13418,N_13243);
or U13773 (N_13773,N_13023,N_13445);
or U13774 (N_13774,N_13225,N_13480);
nand U13775 (N_13775,N_13352,N_13327);
and U13776 (N_13776,N_13295,N_13345);
or U13777 (N_13777,N_13191,N_13355);
xor U13778 (N_13778,N_13032,N_13012);
nor U13779 (N_13779,N_13163,N_13010);
nand U13780 (N_13780,N_13039,N_13212);
nor U13781 (N_13781,N_13138,N_13307);
or U13782 (N_13782,N_13027,N_13236);
nor U13783 (N_13783,N_13045,N_13327);
xnor U13784 (N_13784,N_13128,N_13046);
and U13785 (N_13785,N_13056,N_13304);
and U13786 (N_13786,N_13060,N_13285);
nand U13787 (N_13787,N_13101,N_13011);
xnor U13788 (N_13788,N_13424,N_13444);
or U13789 (N_13789,N_13266,N_13109);
xor U13790 (N_13790,N_13205,N_13474);
and U13791 (N_13791,N_13308,N_13093);
and U13792 (N_13792,N_13134,N_13076);
nand U13793 (N_13793,N_13323,N_13449);
nor U13794 (N_13794,N_13208,N_13443);
and U13795 (N_13795,N_13115,N_13365);
or U13796 (N_13796,N_13213,N_13144);
and U13797 (N_13797,N_13485,N_13256);
and U13798 (N_13798,N_13246,N_13472);
nor U13799 (N_13799,N_13106,N_13039);
or U13800 (N_13800,N_13197,N_13175);
nor U13801 (N_13801,N_13379,N_13167);
nand U13802 (N_13802,N_13032,N_13262);
nand U13803 (N_13803,N_13449,N_13167);
or U13804 (N_13804,N_13153,N_13159);
xor U13805 (N_13805,N_13196,N_13468);
or U13806 (N_13806,N_13091,N_13179);
xnor U13807 (N_13807,N_13479,N_13196);
or U13808 (N_13808,N_13164,N_13082);
or U13809 (N_13809,N_13176,N_13311);
nand U13810 (N_13810,N_13022,N_13159);
or U13811 (N_13811,N_13382,N_13420);
xnor U13812 (N_13812,N_13444,N_13003);
and U13813 (N_13813,N_13259,N_13155);
nor U13814 (N_13814,N_13326,N_13244);
xor U13815 (N_13815,N_13248,N_13064);
and U13816 (N_13816,N_13437,N_13268);
and U13817 (N_13817,N_13314,N_13264);
nor U13818 (N_13818,N_13036,N_13063);
and U13819 (N_13819,N_13084,N_13264);
nand U13820 (N_13820,N_13126,N_13243);
or U13821 (N_13821,N_13405,N_13495);
nand U13822 (N_13822,N_13387,N_13312);
xnor U13823 (N_13823,N_13275,N_13269);
and U13824 (N_13824,N_13402,N_13328);
nor U13825 (N_13825,N_13390,N_13245);
or U13826 (N_13826,N_13244,N_13223);
or U13827 (N_13827,N_13210,N_13054);
nor U13828 (N_13828,N_13021,N_13369);
nor U13829 (N_13829,N_13464,N_13223);
nand U13830 (N_13830,N_13196,N_13202);
and U13831 (N_13831,N_13225,N_13242);
xor U13832 (N_13832,N_13081,N_13330);
or U13833 (N_13833,N_13432,N_13282);
nor U13834 (N_13834,N_13192,N_13437);
or U13835 (N_13835,N_13342,N_13133);
nand U13836 (N_13836,N_13249,N_13477);
xor U13837 (N_13837,N_13269,N_13478);
or U13838 (N_13838,N_13393,N_13180);
or U13839 (N_13839,N_13325,N_13286);
and U13840 (N_13840,N_13216,N_13152);
nor U13841 (N_13841,N_13203,N_13224);
nor U13842 (N_13842,N_13405,N_13041);
nor U13843 (N_13843,N_13174,N_13232);
xnor U13844 (N_13844,N_13241,N_13458);
or U13845 (N_13845,N_13180,N_13382);
xnor U13846 (N_13846,N_13398,N_13049);
nor U13847 (N_13847,N_13124,N_13319);
nor U13848 (N_13848,N_13141,N_13050);
xnor U13849 (N_13849,N_13166,N_13160);
nand U13850 (N_13850,N_13251,N_13280);
and U13851 (N_13851,N_13010,N_13249);
nor U13852 (N_13852,N_13140,N_13187);
xnor U13853 (N_13853,N_13294,N_13353);
and U13854 (N_13854,N_13494,N_13348);
nand U13855 (N_13855,N_13419,N_13057);
and U13856 (N_13856,N_13443,N_13316);
nand U13857 (N_13857,N_13085,N_13226);
and U13858 (N_13858,N_13361,N_13007);
and U13859 (N_13859,N_13017,N_13215);
nand U13860 (N_13860,N_13194,N_13225);
nor U13861 (N_13861,N_13134,N_13206);
nor U13862 (N_13862,N_13211,N_13239);
nand U13863 (N_13863,N_13494,N_13366);
nand U13864 (N_13864,N_13051,N_13159);
and U13865 (N_13865,N_13149,N_13050);
nand U13866 (N_13866,N_13043,N_13414);
xor U13867 (N_13867,N_13344,N_13253);
or U13868 (N_13868,N_13158,N_13395);
or U13869 (N_13869,N_13122,N_13081);
nor U13870 (N_13870,N_13401,N_13199);
nor U13871 (N_13871,N_13237,N_13330);
nand U13872 (N_13872,N_13216,N_13365);
xnor U13873 (N_13873,N_13206,N_13424);
nor U13874 (N_13874,N_13189,N_13361);
nand U13875 (N_13875,N_13388,N_13313);
and U13876 (N_13876,N_13396,N_13311);
or U13877 (N_13877,N_13169,N_13164);
nor U13878 (N_13878,N_13105,N_13474);
or U13879 (N_13879,N_13409,N_13197);
and U13880 (N_13880,N_13449,N_13401);
and U13881 (N_13881,N_13403,N_13228);
or U13882 (N_13882,N_13334,N_13065);
or U13883 (N_13883,N_13208,N_13203);
or U13884 (N_13884,N_13115,N_13298);
or U13885 (N_13885,N_13228,N_13163);
nand U13886 (N_13886,N_13107,N_13194);
nor U13887 (N_13887,N_13089,N_13464);
xnor U13888 (N_13888,N_13083,N_13273);
and U13889 (N_13889,N_13263,N_13287);
or U13890 (N_13890,N_13409,N_13460);
or U13891 (N_13891,N_13197,N_13318);
and U13892 (N_13892,N_13259,N_13325);
nand U13893 (N_13893,N_13459,N_13338);
xor U13894 (N_13894,N_13092,N_13378);
and U13895 (N_13895,N_13069,N_13343);
or U13896 (N_13896,N_13452,N_13423);
xnor U13897 (N_13897,N_13094,N_13080);
nor U13898 (N_13898,N_13128,N_13398);
nor U13899 (N_13899,N_13064,N_13451);
and U13900 (N_13900,N_13256,N_13199);
nand U13901 (N_13901,N_13390,N_13123);
or U13902 (N_13902,N_13329,N_13157);
nand U13903 (N_13903,N_13392,N_13464);
nand U13904 (N_13904,N_13388,N_13436);
or U13905 (N_13905,N_13120,N_13478);
xor U13906 (N_13906,N_13323,N_13418);
or U13907 (N_13907,N_13445,N_13343);
xor U13908 (N_13908,N_13153,N_13446);
nor U13909 (N_13909,N_13163,N_13292);
nand U13910 (N_13910,N_13032,N_13102);
or U13911 (N_13911,N_13383,N_13481);
and U13912 (N_13912,N_13361,N_13417);
xnor U13913 (N_13913,N_13197,N_13228);
or U13914 (N_13914,N_13312,N_13485);
and U13915 (N_13915,N_13407,N_13216);
and U13916 (N_13916,N_13079,N_13418);
and U13917 (N_13917,N_13210,N_13211);
xor U13918 (N_13918,N_13125,N_13492);
and U13919 (N_13919,N_13310,N_13147);
nor U13920 (N_13920,N_13457,N_13034);
nand U13921 (N_13921,N_13111,N_13008);
or U13922 (N_13922,N_13271,N_13246);
nand U13923 (N_13923,N_13064,N_13459);
xnor U13924 (N_13924,N_13281,N_13194);
nand U13925 (N_13925,N_13460,N_13070);
nor U13926 (N_13926,N_13097,N_13043);
and U13927 (N_13927,N_13222,N_13379);
nor U13928 (N_13928,N_13090,N_13271);
nor U13929 (N_13929,N_13289,N_13205);
xnor U13930 (N_13930,N_13126,N_13408);
xnor U13931 (N_13931,N_13329,N_13076);
nor U13932 (N_13932,N_13384,N_13142);
xor U13933 (N_13933,N_13037,N_13410);
nand U13934 (N_13934,N_13258,N_13324);
xnor U13935 (N_13935,N_13000,N_13404);
nor U13936 (N_13936,N_13241,N_13097);
or U13937 (N_13937,N_13396,N_13316);
nor U13938 (N_13938,N_13203,N_13087);
nor U13939 (N_13939,N_13088,N_13080);
xnor U13940 (N_13940,N_13490,N_13361);
xnor U13941 (N_13941,N_13324,N_13019);
nand U13942 (N_13942,N_13295,N_13440);
nand U13943 (N_13943,N_13004,N_13026);
and U13944 (N_13944,N_13178,N_13060);
nand U13945 (N_13945,N_13069,N_13341);
nor U13946 (N_13946,N_13010,N_13303);
and U13947 (N_13947,N_13072,N_13317);
and U13948 (N_13948,N_13406,N_13416);
and U13949 (N_13949,N_13072,N_13331);
nand U13950 (N_13950,N_13289,N_13369);
or U13951 (N_13951,N_13015,N_13331);
or U13952 (N_13952,N_13253,N_13016);
nand U13953 (N_13953,N_13380,N_13322);
and U13954 (N_13954,N_13050,N_13177);
nand U13955 (N_13955,N_13111,N_13178);
and U13956 (N_13956,N_13129,N_13133);
nand U13957 (N_13957,N_13028,N_13178);
nor U13958 (N_13958,N_13048,N_13460);
nor U13959 (N_13959,N_13484,N_13085);
or U13960 (N_13960,N_13235,N_13074);
and U13961 (N_13961,N_13033,N_13415);
nand U13962 (N_13962,N_13349,N_13425);
nor U13963 (N_13963,N_13414,N_13008);
xnor U13964 (N_13964,N_13282,N_13406);
nor U13965 (N_13965,N_13428,N_13185);
nor U13966 (N_13966,N_13339,N_13204);
or U13967 (N_13967,N_13043,N_13281);
nand U13968 (N_13968,N_13054,N_13268);
and U13969 (N_13969,N_13252,N_13365);
nor U13970 (N_13970,N_13304,N_13010);
nor U13971 (N_13971,N_13337,N_13055);
nand U13972 (N_13972,N_13374,N_13015);
nand U13973 (N_13973,N_13184,N_13381);
and U13974 (N_13974,N_13110,N_13282);
xor U13975 (N_13975,N_13285,N_13047);
or U13976 (N_13976,N_13145,N_13071);
xor U13977 (N_13977,N_13077,N_13473);
xnor U13978 (N_13978,N_13164,N_13378);
and U13979 (N_13979,N_13300,N_13333);
and U13980 (N_13980,N_13281,N_13335);
nor U13981 (N_13981,N_13298,N_13209);
nor U13982 (N_13982,N_13138,N_13429);
xnor U13983 (N_13983,N_13152,N_13229);
or U13984 (N_13984,N_13207,N_13121);
or U13985 (N_13985,N_13353,N_13482);
and U13986 (N_13986,N_13426,N_13320);
xnor U13987 (N_13987,N_13142,N_13229);
and U13988 (N_13988,N_13353,N_13197);
or U13989 (N_13989,N_13322,N_13144);
or U13990 (N_13990,N_13314,N_13282);
nor U13991 (N_13991,N_13438,N_13481);
nand U13992 (N_13992,N_13427,N_13038);
nor U13993 (N_13993,N_13361,N_13240);
and U13994 (N_13994,N_13184,N_13257);
xor U13995 (N_13995,N_13367,N_13245);
or U13996 (N_13996,N_13215,N_13436);
or U13997 (N_13997,N_13289,N_13297);
nand U13998 (N_13998,N_13144,N_13038);
or U13999 (N_13999,N_13435,N_13027);
nand U14000 (N_14000,N_13796,N_13521);
or U14001 (N_14001,N_13986,N_13906);
nand U14002 (N_14002,N_13612,N_13572);
xnor U14003 (N_14003,N_13916,N_13504);
nand U14004 (N_14004,N_13748,N_13896);
or U14005 (N_14005,N_13712,N_13539);
xnor U14006 (N_14006,N_13802,N_13506);
and U14007 (N_14007,N_13611,N_13700);
nand U14008 (N_14008,N_13727,N_13540);
and U14009 (N_14009,N_13651,N_13541);
xnor U14010 (N_14010,N_13656,N_13733);
nor U14011 (N_14011,N_13621,N_13744);
or U14012 (N_14012,N_13983,N_13790);
and U14013 (N_14013,N_13674,N_13884);
or U14014 (N_14014,N_13514,N_13838);
xnor U14015 (N_14015,N_13616,N_13509);
xnor U14016 (N_14016,N_13633,N_13515);
nand U14017 (N_14017,N_13822,N_13669);
and U14018 (N_14018,N_13556,N_13771);
or U14019 (N_14019,N_13930,N_13565);
xor U14020 (N_14020,N_13809,N_13649);
and U14021 (N_14021,N_13927,N_13879);
or U14022 (N_14022,N_13530,N_13694);
xor U14023 (N_14023,N_13936,N_13566);
and U14024 (N_14024,N_13682,N_13797);
xnor U14025 (N_14025,N_13898,N_13500);
nor U14026 (N_14026,N_13569,N_13555);
and U14027 (N_14027,N_13726,N_13816);
and U14028 (N_14028,N_13581,N_13586);
xor U14029 (N_14029,N_13736,N_13827);
xnor U14030 (N_14030,N_13720,N_13824);
or U14031 (N_14031,N_13971,N_13761);
nor U14032 (N_14032,N_13803,N_13928);
and U14033 (N_14033,N_13585,N_13654);
and U14034 (N_14034,N_13794,N_13676);
or U14035 (N_14035,N_13534,N_13538);
xor U14036 (N_14036,N_13766,N_13661);
or U14037 (N_14037,N_13878,N_13917);
and U14038 (N_14038,N_13683,N_13759);
xor U14039 (N_14039,N_13647,N_13954);
nand U14040 (N_14040,N_13704,N_13834);
nor U14041 (N_14041,N_13687,N_13776);
nand U14042 (N_14042,N_13889,N_13897);
nor U14043 (N_14043,N_13644,N_13801);
nand U14044 (N_14044,N_13812,N_13597);
and U14045 (N_14045,N_13778,N_13558);
or U14046 (N_14046,N_13642,N_13531);
nor U14047 (N_14047,N_13529,N_13552);
and U14048 (N_14048,N_13602,N_13937);
nand U14049 (N_14049,N_13839,N_13547);
nand U14050 (N_14050,N_13899,N_13598);
nand U14051 (N_14051,N_13945,N_13672);
xnor U14052 (N_14052,N_13909,N_13628);
or U14053 (N_14053,N_13607,N_13730);
nand U14054 (N_14054,N_13833,N_13901);
nand U14055 (N_14055,N_13503,N_13814);
or U14056 (N_14056,N_13970,N_13645);
or U14057 (N_14057,N_13888,N_13703);
xnor U14058 (N_14058,N_13636,N_13883);
xnor U14059 (N_14059,N_13717,N_13979);
nor U14060 (N_14060,N_13624,N_13934);
or U14061 (N_14061,N_13872,N_13867);
nand U14062 (N_14062,N_13855,N_13543);
nor U14063 (N_14063,N_13958,N_13873);
and U14064 (N_14064,N_13606,N_13957);
and U14065 (N_14065,N_13882,N_13892);
and U14066 (N_14066,N_13886,N_13707);
and U14067 (N_14067,N_13603,N_13973);
nor U14068 (N_14068,N_13863,N_13955);
xor U14069 (N_14069,N_13593,N_13559);
nand U14070 (N_14070,N_13537,N_13815);
xor U14071 (N_14071,N_13743,N_13548);
nor U14072 (N_14072,N_13574,N_13871);
nor U14073 (N_14073,N_13938,N_13792);
xnor U14074 (N_14074,N_13508,N_13974);
and U14075 (N_14075,N_13750,N_13856);
nor U14076 (N_14076,N_13610,N_13620);
or U14077 (N_14077,N_13943,N_13763);
xnor U14078 (N_14078,N_13595,N_13829);
nor U14079 (N_14079,N_13751,N_13915);
nand U14080 (N_14080,N_13632,N_13741);
xnor U14081 (N_14081,N_13671,N_13578);
nor U14082 (N_14082,N_13890,N_13705);
nor U14083 (N_14083,N_13653,N_13977);
nand U14084 (N_14084,N_13623,N_13989);
nor U14085 (N_14085,N_13918,N_13735);
or U14086 (N_14086,N_13791,N_13788);
nor U14087 (N_14087,N_13895,N_13859);
or U14088 (N_14088,N_13601,N_13903);
or U14089 (N_14089,N_13501,N_13599);
and U14090 (N_14090,N_13525,N_13630);
xnor U14091 (N_14091,N_13512,N_13900);
nand U14092 (N_14092,N_13625,N_13577);
nor U14093 (N_14093,N_13613,N_13589);
nor U14094 (N_14094,N_13535,N_13667);
nand U14095 (N_14095,N_13846,N_13554);
or U14096 (N_14096,N_13617,N_13520);
and U14097 (N_14097,N_13995,N_13688);
nand U14098 (N_14098,N_13887,N_13770);
nand U14099 (N_14099,N_13946,N_13841);
or U14100 (N_14100,N_13874,N_13907);
nand U14101 (N_14101,N_13587,N_13960);
nand U14102 (N_14102,N_13695,N_13505);
xnor U14103 (N_14103,N_13951,N_13686);
nand U14104 (N_14104,N_13680,N_13817);
and U14105 (N_14105,N_13935,N_13780);
and U14106 (N_14106,N_13622,N_13522);
and U14107 (N_14107,N_13831,N_13532);
xor U14108 (N_14108,N_13590,N_13865);
and U14109 (N_14109,N_13724,N_13755);
and U14110 (N_14110,N_13904,N_13737);
and U14111 (N_14111,N_13584,N_13518);
nor U14112 (N_14112,N_13965,N_13708);
nand U14113 (N_14113,N_13968,N_13911);
nand U14114 (N_14114,N_13706,N_13742);
xor U14115 (N_14115,N_13562,N_13697);
nand U14116 (N_14116,N_13963,N_13605);
and U14117 (N_14117,N_13575,N_13825);
nor U14118 (N_14118,N_13710,N_13773);
and U14119 (N_14119,N_13905,N_13826);
nor U14120 (N_14120,N_13752,N_13837);
nor U14121 (N_14121,N_13699,N_13787);
nor U14122 (N_14122,N_13964,N_13681);
xnor U14123 (N_14123,N_13866,N_13711);
and U14124 (N_14124,N_13894,N_13808);
xnor U14125 (N_14125,N_13967,N_13725);
or U14126 (N_14126,N_13852,N_13910);
xor U14127 (N_14127,N_13600,N_13570);
xor U14128 (N_14128,N_13768,N_13640);
or U14129 (N_14129,N_13746,N_13563);
nand U14130 (N_14130,N_13926,N_13657);
and U14131 (N_14131,N_13939,N_13975);
and U14132 (N_14132,N_13805,N_13952);
nand U14133 (N_14133,N_13764,N_13774);
xor U14134 (N_14134,N_13848,N_13713);
xnor U14135 (N_14135,N_13721,N_13594);
nand U14136 (N_14136,N_13627,N_13519);
nor U14137 (N_14137,N_13580,N_13550);
nor U14138 (N_14138,N_13881,N_13648);
and U14139 (N_14139,N_13953,N_13643);
nor U14140 (N_14140,N_13658,N_13772);
and U14141 (N_14141,N_13853,N_13948);
and U14142 (N_14142,N_13678,N_13925);
nor U14143 (N_14143,N_13782,N_13567);
and U14144 (N_14144,N_13984,N_13760);
nand U14145 (N_14145,N_13641,N_13722);
or U14146 (N_14146,N_13844,N_13779);
and U14147 (N_14147,N_13561,N_13840);
and U14148 (N_14148,N_13850,N_13893);
or U14149 (N_14149,N_13847,N_13868);
nor U14150 (N_14150,N_13675,N_13777);
or U14151 (N_14151,N_13545,N_13691);
xnor U14152 (N_14152,N_13511,N_13858);
and U14153 (N_14153,N_13614,N_13637);
and U14154 (N_14154,N_13969,N_13997);
xor U14155 (N_14155,N_13758,N_13823);
xnor U14156 (N_14156,N_13663,N_13854);
nand U14157 (N_14157,N_13789,N_13698);
xnor U14158 (N_14158,N_13956,N_13571);
xor U14159 (N_14159,N_13877,N_13998);
or U14160 (N_14160,N_13806,N_13551);
xnor U14161 (N_14161,N_13832,N_13655);
nand U14162 (N_14162,N_13738,N_13857);
and U14163 (N_14163,N_13626,N_13944);
xnor U14164 (N_14164,N_13679,N_13830);
nor U14165 (N_14165,N_13582,N_13861);
xnor U14166 (N_14166,N_13793,N_13573);
nor U14167 (N_14167,N_13576,N_13608);
nand U14168 (N_14168,N_13769,N_13502);
and U14169 (N_14169,N_13604,N_13664);
nor U14170 (N_14170,N_13875,N_13731);
or U14171 (N_14171,N_13560,N_13673);
nand U14172 (N_14172,N_13591,N_13966);
xor U14173 (N_14173,N_13931,N_13950);
xnor U14174 (N_14174,N_13942,N_13544);
nand U14175 (N_14175,N_13821,N_13811);
and U14176 (N_14176,N_13709,N_13804);
nor U14177 (N_14177,N_13835,N_13959);
xor U14178 (N_14178,N_13920,N_13949);
nand U14179 (N_14179,N_13976,N_13729);
or U14180 (N_14180,N_13813,N_13988);
xnor U14181 (N_14181,N_13836,N_13728);
nand U14182 (N_14182,N_13919,N_13528);
nand U14183 (N_14183,N_13756,N_13798);
nand U14184 (N_14184,N_13516,N_13659);
and U14185 (N_14185,N_13740,N_13762);
or U14186 (N_14186,N_13991,N_13715);
and U14187 (N_14187,N_13799,N_13629);
xor U14188 (N_14188,N_13513,N_13961);
or U14189 (N_14189,N_13851,N_13526);
nor U14190 (N_14190,N_13922,N_13891);
xor U14191 (N_14191,N_13870,N_13639);
and U14192 (N_14192,N_13785,N_13818);
or U14193 (N_14193,N_13747,N_13842);
nand U14194 (N_14194,N_13786,N_13908);
nor U14195 (N_14195,N_13860,N_13781);
nor U14196 (N_14196,N_13869,N_13523);
or U14197 (N_14197,N_13596,N_13993);
and U14198 (N_14198,N_13723,N_13757);
or U14199 (N_14199,N_13734,N_13783);
nand U14200 (N_14200,N_13862,N_13684);
and U14201 (N_14201,N_13940,N_13885);
nand U14202 (N_14202,N_13981,N_13533);
nor U14203 (N_14203,N_13527,N_13739);
nor U14204 (N_14204,N_13690,N_13843);
nand U14205 (N_14205,N_13996,N_13696);
and U14206 (N_14206,N_13987,N_13564);
nand U14207 (N_14207,N_13646,N_13619);
nor U14208 (N_14208,N_13828,N_13921);
xnor U14209 (N_14209,N_13719,N_13716);
nand U14210 (N_14210,N_13666,N_13615);
nor U14211 (N_14211,N_13932,N_13849);
nand U14212 (N_14212,N_13800,N_13701);
or U14213 (N_14213,N_13767,N_13933);
or U14214 (N_14214,N_13912,N_13702);
xor U14215 (N_14215,N_13864,N_13665);
or U14216 (N_14216,N_13994,N_13784);
nand U14217 (N_14217,N_13553,N_13810);
and U14218 (N_14218,N_13689,N_13765);
nand U14219 (N_14219,N_13807,N_13753);
xnor U14220 (N_14220,N_13923,N_13982);
and U14221 (N_14221,N_13978,N_13999);
nand U14222 (N_14222,N_13517,N_13913);
and U14223 (N_14223,N_13510,N_13660);
or U14224 (N_14224,N_13631,N_13652);
and U14225 (N_14225,N_13588,N_13549);
or U14226 (N_14226,N_13557,N_13670);
xor U14227 (N_14227,N_13775,N_13880);
nand U14228 (N_14228,N_13579,N_13714);
nor U14229 (N_14229,N_13745,N_13754);
nand U14230 (N_14230,N_13990,N_13924);
nor U14231 (N_14231,N_13876,N_13568);
or U14232 (N_14232,N_13583,N_13662);
nor U14233 (N_14233,N_13592,N_13718);
nand U14234 (N_14234,N_13929,N_13902);
or U14235 (N_14235,N_13546,N_13638);
and U14236 (N_14236,N_13941,N_13985);
xnor U14237 (N_14237,N_13685,N_13692);
or U14238 (N_14238,N_13992,N_13635);
or U14239 (N_14239,N_13972,N_13524);
nand U14240 (N_14240,N_13962,N_13634);
and U14241 (N_14241,N_13693,N_13820);
nor U14242 (N_14242,N_13914,N_13845);
nand U14243 (N_14243,N_13732,N_13947);
nor U14244 (N_14244,N_13609,N_13795);
nand U14245 (N_14245,N_13650,N_13542);
or U14246 (N_14246,N_13677,N_13819);
or U14247 (N_14247,N_13749,N_13536);
or U14248 (N_14248,N_13980,N_13618);
nor U14249 (N_14249,N_13507,N_13668);
nand U14250 (N_14250,N_13674,N_13723);
nor U14251 (N_14251,N_13809,N_13898);
and U14252 (N_14252,N_13843,N_13754);
nand U14253 (N_14253,N_13990,N_13748);
xnor U14254 (N_14254,N_13990,N_13914);
nor U14255 (N_14255,N_13778,N_13633);
or U14256 (N_14256,N_13704,N_13972);
nor U14257 (N_14257,N_13515,N_13530);
xnor U14258 (N_14258,N_13758,N_13704);
nand U14259 (N_14259,N_13685,N_13901);
nand U14260 (N_14260,N_13989,N_13613);
nor U14261 (N_14261,N_13601,N_13558);
nor U14262 (N_14262,N_13865,N_13974);
or U14263 (N_14263,N_13626,N_13710);
and U14264 (N_14264,N_13874,N_13825);
nand U14265 (N_14265,N_13554,N_13505);
xor U14266 (N_14266,N_13899,N_13678);
and U14267 (N_14267,N_13870,N_13937);
xnor U14268 (N_14268,N_13807,N_13895);
nor U14269 (N_14269,N_13620,N_13513);
and U14270 (N_14270,N_13952,N_13710);
nand U14271 (N_14271,N_13781,N_13596);
or U14272 (N_14272,N_13818,N_13538);
nand U14273 (N_14273,N_13986,N_13587);
xnor U14274 (N_14274,N_13530,N_13872);
or U14275 (N_14275,N_13724,N_13637);
and U14276 (N_14276,N_13570,N_13968);
nor U14277 (N_14277,N_13652,N_13683);
nand U14278 (N_14278,N_13726,N_13849);
or U14279 (N_14279,N_13901,N_13823);
nor U14280 (N_14280,N_13894,N_13520);
nor U14281 (N_14281,N_13616,N_13878);
or U14282 (N_14282,N_13594,N_13712);
nand U14283 (N_14283,N_13811,N_13660);
xnor U14284 (N_14284,N_13544,N_13881);
nand U14285 (N_14285,N_13990,N_13544);
nor U14286 (N_14286,N_13980,N_13579);
and U14287 (N_14287,N_13541,N_13703);
nand U14288 (N_14288,N_13873,N_13766);
and U14289 (N_14289,N_13590,N_13928);
and U14290 (N_14290,N_13598,N_13651);
nor U14291 (N_14291,N_13944,N_13884);
or U14292 (N_14292,N_13836,N_13924);
and U14293 (N_14293,N_13754,N_13899);
nand U14294 (N_14294,N_13887,N_13809);
and U14295 (N_14295,N_13757,N_13789);
xor U14296 (N_14296,N_13703,N_13982);
or U14297 (N_14297,N_13552,N_13940);
or U14298 (N_14298,N_13988,N_13982);
and U14299 (N_14299,N_13883,N_13537);
and U14300 (N_14300,N_13568,N_13731);
or U14301 (N_14301,N_13715,N_13701);
nand U14302 (N_14302,N_13686,N_13708);
nor U14303 (N_14303,N_13613,N_13711);
or U14304 (N_14304,N_13789,N_13592);
xnor U14305 (N_14305,N_13864,N_13577);
and U14306 (N_14306,N_13796,N_13642);
or U14307 (N_14307,N_13550,N_13745);
and U14308 (N_14308,N_13779,N_13941);
xnor U14309 (N_14309,N_13926,N_13754);
xor U14310 (N_14310,N_13863,N_13708);
and U14311 (N_14311,N_13916,N_13645);
xnor U14312 (N_14312,N_13947,N_13887);
xnor U14313 (N_14313,N_13576,N_13862);
nand U14314 (N_14314,N_13798,N_13801);
xnor U14315 (N_14315,N_13710,N_13555);
or U14316 (N_14316,N_13559,N_13943);
or U14317 (N_14317,N_13847,N_13694);
or U14318 (N_14318,N_13685,N_13547);
xnor U14319 (N_14319,N_13831,N_13828);
nand U14320 (N_14320,N_13843,N_13857);
xnor U14321 (N_14321,N_13868,N_13798);
and U14322 (N_14322,N_13708,N_13670);
or U14323 (N_14323,N_13887,N_13824);
nor U14324 (N_14324,N_13730,N_13510);
nand U14325 (N_14325,N_13625,N_13652);
xor U14326 (N_14326,N_13904,N_13741);
nand U14327 (N_14327,N_13720,N_13583);
xor U14328 (N_14328,N_13878,N_13961);
or U14329 (N_14329,N_13634,N_13890);
nand U14330 (N_14330,N_13821,N_13893);
or U14331 (N_14331,N_13706,N_13584);
nor U14332 (N_14332,N_13972,N_13720);
nor U14333 (N_14333,N_13780,N_13816);
and U14334 (N_14334,N_13847,N_13633);
xnor U14335 (N_14335,N_13930,N_13588);
and U14336 (N_14336,N_13977,N_13699);
nand U14337 (N_14337,N_13774,N_13885);
nand U14338 (N_14338,N_13988,N_13586);
or U14339 (N_14339,N_13913,N_13945);
nor U14340 (N_14340,N_13546,N_13652);
and U14341 (N_14341,N_13658,N_13640);
nor U14342 (N_14342,N_13514,N_13708);
xnor U14343 (N_14343,N_13638,N_13567);
or U14344 (N_14344,N_13834,N_13891);
and U14345 (N_14345,N_13629,N_13923);
nor U14346 (N_14346,N_13856,N_13503);
or U14347 (N_14347,N_13594,N_13593);
nor U14348 (N_14348,N_13626,N_13981);
xnor U14349 (N_14349,N_13871,N_13553);
and U14350 (N_14350,N_13690,N_13735);
nand U14351 (N_14351,N_13554,N_13956);
xnor U14352 (N_14352,N_13929,N_13641);
and U14353 (N_14353,N_13677,N_13872);
nor U14354 (N_14354,N_13519,N_13566);
and U14355 (N_14355,N_13716,N_13772);
and U14356 (N_14356,N_13670,N_13675);
xor U14357 (N_14357,N_13865,N_13981);
or U14358 (N_14358,N_13805,N_13842);
nand U14359 (N_14359,N_13943,N_13501);
nand U14360 (N_14360,N_13790,N_13978);
and U14361 (N_14361,N_13973,N_13806);
nor U14362 (N_14362,N_13647,N_13823);
nor U14363 (N_14363,N_13711,N_13919);
nand U14364 (N_14364,N_13871,N_13653);
xnor U14365 (N_14365,N_13694,N_13610);
or U14366 (N_14366,N_13880,N_13945);
xnor U14367 (N_14367,N_13625,N_13607);
xnor U14368 (N_14368,N_13794,N_13677);
xor U14369 (N_14369,N_13755,N_13722);
nand U14370 (N_14370,N_13710,N_13968);
nand U14371 (N_14371,N_13791,N_13922);
nand U14372 (N_14372,N_13702,N_13987);
xor U14373 (N_14373,N_13761,N_13707);
xor U14374 (N_14374,N_13615,N_13805);
or U14375 (N_14375,N_13934,N_13518);
nor U14376 (N_14376,N_13820,N_13859);
xnor U14377 (N_14377,N_13568,N_13993);
nand U14378 (N_14378,N_13687,N_13553);
nor U14379 (N_14379,N_13631,N_13778);
nor U14380 (N_14380,N_13931,N_13619);
xor U14381 (N_14381,N_13718,N_13724);
nor U14382 (N_14382,N_13666,N_13596);
xor U14383 (N_14383,N_13534,N_13648);
or U14384 (N_14384,N_13851,N_13548);
or U14385 (N_14385,N_13875,N_13868);
nor U14386 (N_14386,N_13676,N_13740);
nor U14387 (N_14387,N_13654,N_13653);
and U14388 (N_14388,N_13839,N_13822);
xor U14389 (N_14389,N_13979,N_13899);
xnor U14390 (N_14390,N_13733,N_13662);
and U14391 (N_14391,N_13899,N_13617);
nand U14392 (N_14392,N_13836,N_13884);
xor U14393 (N_14393,N_13829,N_13918);
nor U14394 (N_14394,N_13680,N_13514);
nor U14395 (N_14395,N_13569,N_13934);
nor U14396 (N_14396,N_13949,N_13674);
and U14397 (N_14397,N_13770,N_13732);
xor U14398 (N_14398,N_13760,N_13520);
nor U14399 (N_14399,N_13607,N_13876);
nand U14400 (N_14400,N_13724,N_13824);
or U14401 (N_14401,N_13985,N_13532);
nor U14402 (N_14402,N_13762,N_13684);
nand U14403 (N_14403,N_13688,N_13937);
nor U14404 (N_14404,N_13754,N_13750);
or U14405 (N_14405,N_13603,N_13577);
nand U14406 (N_14406,N_13980,N_13615);
or U14407 (N_14407,N_13857,N_13654);
nand U14408 (N_14408,N_13550,N_13637);
and U14409 (N_14409,N_13541,N_13965);
xnor U14410 (N_14410,N_13644,N_13800);
nor U14411 (N_14411,N_13526,N_13855);
and U14412 (N_14412,N_13916,N_13508);
nand U14413 (N_14413,N_13961,N_13699);
or U14414 (N_14414,N_13864,N_13796);
xnor U14415 (N_14415,N_13613,N_13574);
xnor U14416 (N_14416,N_13679,N_13896);
and U14417 (N_14417,N_13610,N_13568);
or U14418 (N_14418,N_13583,N_13547);
nor U14419 (N_14419,N_13591,N_13983);
nor U14420 (N_14420,N_13759,N_13894);
xor U14421 (N_14421,N_13506,N_13598);
nor U14422 (N_14422,N_13670,N_13640);
nand U14423 (N_14423,N_13884,N_13621);
xnor U14424 (N_14424,N_13984,N_13987);
nand U14425 (N_14425,N_13658,N_13672);
xnor U14426 (N_14426,N_13928,N_13904);
xor U14427 (N_14427,N_13974,N_13778);
or U14428 (N_14428,N_13673,N_13512);
and U14429 (N_14429,N_13998,N_13771);
nand U14430 (N_14430,N_13911,N_13912);
and U14431 (N_14431,N_13904,N_13596);
nand U14432 (N_14432,N_13680,N_13952);
xnor U14433 (N_14433,N_13567,N_13843);
nor U14434 (N_14434,N_13856,N_13627);
nand U14435 (N_14435,N_13749,N_13835);
xnor U14436 (N_14436,N_13628,N_13739);
nor U14437 (N_14437,N_13918,N_13720);
nor U14438 (N_14438,N_13690,N_13630);
nand U14439 (N_14439,N_13798,N_13637);
xnor U14440 (N_14440,N_13691,N_13917);
xnor U14441 (N_14441,N_13681,N_13615);
xnor U14442 (N_14442,N_13988,N_13809);
xnor U14443 (N_14443,N_13854,N_13544);
nand U14444 (N_14444,N_13600,N_13758);
and U14445 (N_14445,N_13591,N_13542);
nor U14446 (N_14446,N_13792,N_13588);
and U14447 (N_14447,N_13677,N_13795);
nor U14448 (N_14448,N_13609,N_13685);
nor U14449 (N_14449,N_13728,N_13801);
xnor U14450 (N_14450,N_13822,N_13962);
nor U14451 (N_14451,N_13793,N_13687);
nor U14452 (N_14452,N_13754,N_13888);
xnor U14453 (N_14453,N_13908,N_13929);
nor U14454 (N_14454,N_13699,N_13998);
nand U14455 (N_14455,N_13515,N_13796);
and U14456 (N_14456,N_13588,N_13893);
nand U14457 (N_14457,N_13735,N_13891);
or U14458 (N_14458,N_13787,N_13682);
xnor U14459 (N_14459,N_13560,N_13978);
or U14460 (N_14460,N_13821,N_13732);
xor U14461 (N_14461,N_13685,N_13775);
xnor U14462 (N_14462,N_13599,N_13678);
or U14463 (N_14463,N_13652,N_13501);
nor U14464 (N_14464,N_13681,N_13730);
or U14465 (N_14465,N_13634,N_13582);
nor U14466 (N_14466,N_13799,N_13886);
xnor U14467 (N_14467,N_13612,N_13911);
or U14468 (N_14468,N_13960,N_13861);
xnor U14469 (N_14469,N_13610,N_13614);
or U14470 (N_14470,N_13759,N_13797);
or U14471 (N_14471,N_13698,N_13827);
and U14472 (N_14472,N_13855,N_13732);
nand U14473 (N_14473,N_13506,N_13747);
and U14474 (N_14474,N_13771,N_13620);
or U14475 (N_14475,N_13630,N_13946);
or U14476 (N_14476,N_13570,N_13892);
nand U14477 (N_14477,N_13506,N_13604);
xor U14478 (N_14478,N_13578,N_13768);
and U14479 (N_14479,N_13695,N_13902);
nand U14480 (N_14480,N_13542,N_13586);
and U14481 (N_14481,N_13706,N_13691);
nor U14482 (N_14482,N_13514,N_13982);
nor U14483 (N_14483,N_13532,N_13541);
or U14484 (N_14484,N_13636,N_13761);
xor U14485 (N_14485,N_13543,N_13551);
and U14486 (N_14486,N_13739,N_13646);
nand U14487 (N_14487,N_13520,N_13739);
and U14488 (N_14488,N_13954,N_13507);
nand U14489 (N_14489,N_13814,N_13870);
xnor U14490 (N_14490,N_13669,N_13842);
xnor U14491 (N_14491,N_13792,N_13524);
nand U14492 (N_14492,N_13826,N_13662);
xor U14493 (N_14493,N_13836,N_13860);
nand U14494 (N_14494,N_13918,N_13805);
nor U14495 (N_14495,N_13733,N_13513);
or U14496 (N_14496,N_13626,N_13903);
and U14497 (N_14497,N_13665,N_13560);
and U14498 (N_14498,N_13953,N_13660);
or U14499 (N_14499,N_13560,N_13864);
and U14500 (N_14500,N_14068,N_14347);
nand U14501 (N_14501,N_14120,N_14007);
and U14502 (N_14502,N_14059,N_14144);
xnor U14503 (N_14503,N_14153,N_14360);
and U14504 (N_14504,N_14037,N_14205);
nor U14505 (N_14505,N_14168,N_14338);
nor U14506 (N_14506,N_14266,N_14417);
xor U14507 (N_14507,N_14036,N_14203);
and U14508 (N_14508,N_14455,N_14175);
and U14509 (N_14509,N_14420,N_14199);
nor U14510 (N_14510,N_14478,N_14270);
xor U14511 (N_14511,N_14336,N_14453);
xnor U14512 (N_14512,N_14089,N_14469);
and U14513 (N_14513,N_14082,N_14458);
xnor U14514 (N_14514,N_14450,N_14404);
and U14515 (N_14515,N_14191,N_14471);
xnor U14516 (N_14516,N_14373,N_14066);
nor U14517 (N_14517,N_14479,N_14167);
and U14518 (N_14518,N_14158,N_14031);
xor U14519 (N_14519,N_14047,N_14343);
xnor U14520 (N_14520,N_14442,N_14311);
nor U14521 (N_14521,N_14043,N_14254);
or U14522 (N_14522,N_14058,N_14359);
or U14523 (N_14523,N_14474,N_14314);
nand U14524 (N_14524,N_14171,N_14088);
nand U14525 (N_14525,N_14257,N_14333);
xor U14526 (N_14526,N_14095,N_14014);
nand U14527 (N_14527,N_14204,N_14081);
nor U14528 (N_14528,N_14448,N_14462);
nand U14529 (N_14529,N_14444,N_14402);
and U14530 (N_14530,N_14273,N_14030);
nand U14531 (N_14531,N_14432,N_14316);
and U14532 (N_14532,N_14488,N_14102);
xor U14533 (N_14533,N_14134,N_14433);
nor U14534 (N_14534,N_14487,N_14123);
nor U14535 (N_14535,N_14370,N_14372);
nor U14536 (N_14536,N_14287,N_14354);
nand U14537 (N_14537,N_14419,N_14159);
nand U14538 (N_14538,N_14012,N_14140);
xor U14539 (N_14539,N_14213,N_14284);
xnor U14540 (N_14540,N_14434,N_14376);
xnor U14541 (N_14541,N_14309,N_14077);
or U14542 (N_14542,N_14172,N_14313);
nor U14543 (N_14543,N_14422,N_14391);
and U14544 (N_14544,N_14210,N_14356);
xnor U14545 (N_14545,N_14407,N_14228);
or U14546 (N_14546,N_14119,N_14242);
nor U14547 (N_14547,N_14253,N_14006);
nor U14548 (N_14548,N_14099,N_14364);
and U14549 (N_14549,N_14033,N_14476);
and U14550 (N_14550,N_14292,N_14108);
nor U14551 (N_14551,N_14497,N_14499);
and U14552 (N_14552,N_14352,N_14018);
nand U14553 (N_14553,N_14465,N_14100);
or U14554 (N_14554,N_14184,N_14250);
or U14555 (N_14555,N_14070,N_14435);
xor U14556 (N_14556,N_14481,N_14430);
and U14557 (N_14557,N_14492,N_14276);
or U14558 (N_14558,N_14247,N_14240);
and U14559 (N_14559,N_14281,N_14048);
xor U14560 (N_14560,N_14148,N_14357);
xnor U14561 (N_14561,N_14016,N_14482);
or U14562 (N_14562,N_14054,N_14489);
nand U14563 (N_14563,N_14177,N_14325);
nor U14564 (N_14564,N_14132,N_14264);
xor U14565 (N_14565,N_14207,N_14441);
xnor U14566 (N_14566,N_14121,N_14387);
and U14567 (N_14567,N_14446,N_14383);
and U14568 (N_14568,N_14003,N_14115);
or U14569 (N_14569,N_14398,N_14439);
or U14570 (N_14570,N_14396,N_14261);
or U14571 (N_14571,N_14377,N_14187);
and U14572 (N_14572,N_14447,N_14085);
nor U14573 (N_14573,N_14348,N_14290);
and U14574 (N_14574,N_14278,N_14063);
or U14575 (N_14575,N_14258,N_14227);
or U14576 (N_14576,N_14353,N_14368);
xor U14577 (N_14577,N_14091,N_14234);
and U14578 (N_14578,N_14301,N_14463);
nand U14579 (N_14579,N_14229,N_14445);
xor U14580 (N_14580,N_14457,N_14295);
nand U14581 (N_14581,N_14004,N_14157);
or U14582 (N_14582,N_14023,N_14274);
and U14583 (N_14583,N_14180,N_14154);
xor U14584 (N_14584,N_14306,N_14375);
nor U14585 (N_14585,N_14028,N_14071);
nor U14586 (N_14586,N_14239,N_14015);
nand U14587 (N_14587,N_14366,N_14209);
and U14588 (N_14588,N_14032,N_14389);
nand U14589 (N_14589,N_14045,N_14092);
and U14590 (N_14590,N_14285,N_14268);
nor U14591 (N_14591,N_14416,N_14223);
nor U14592 (N_14592,N_14466,N_14019);
nor U14593 (N_14593,N_14449,N_14294);
xnor U14594 (N_14594,N_14190,N_14367);
and U14595 (N_14595,N_14124,N_14055);
nand U14596 (N_14596,N_14262,N_14189);
nand U14597 (N_14597,N_14183,N_14103);
nand U14598 (N_14598,N_14110,N_14118);
nor U14599 (N_14599,N_14219,N_14069);
and U14600 (N_14600,N_14025,N_14141);
nor U14601 (N_14601,N_14206,N_14020);
nand U14602 (N_14602,N_14073,N_14112);
nand U14603 (N_14603,N_14414,N_14395);
nor U14604 (N_14604,N_14271,N_14378);
or U14605 (N_14605,N_14026,N_14302);
nand U14606 (N_14606,N_14310,N_14039);
and U14607 (N_14607,N_14221,N_14040);
xor U14608 (N_14608,N_14405,N_14472);
nor U14609 (N_14609,N_14490,N_14361);
nor U14610 (N_14610,N_14215,N_14300);
nor U14611 (N_14611,N_14374,N_14320);
and U14612 (N_14612,N_14315,N_14297);
nand U14613 (N_14613,N_14098,N_14044);
or U14614 (N_14614,N_14238,N_14052);
or U14615 (N_14615,N_14339,N_14452);
nor U14616 (N_14616,N_14113,N_14001);
and U14617 (N_14617,N_14265,N_14362);
nor U14618 (N_14618,N_14437,N_14243);
or U14619 (N_14619,N_14161,N_14116);
or U14620 (N_14620,N_14256,N_14351);
nand U14621 (N_14621,N_14096,N_14222);
and U14622 (N_14622,N_14379,N_14371);
nand U14623 (N_14623,N_14399,N_14321);
and U14624 (N_14624,N_14277,N_14185);
nor U14625 (N_14625,N_14076,N_14079);
nor U14626 (N_14626,N_14329,N_14067);
xor U14627 (N_14627,N_14291,N_14000);
and U14628 (N_14628,N_14304,N_14241);
xnor U14629 (N_14629,N_14393,N_14461);
and U14630 (N_14630,N_14224,N_14400);
and U14631 (N_14631,N_14440,N_14217);
and U14632 (N_14632,N_14438,N_14473);
nor U14633 (N_14633,N_14041,N_14226);
nand U14634 (N_14634,N_14104,N_14129);
and U14635 (N_14635,N_14057,N_14260);
or U14636 (N_14636,N_14220,N_14388);
nand U14637 (N_14637,N_14214,N_14498);
nor U14638 (N_14638,N_14431,N_14334);
and U14639 (N_14639,N_14384,N_14010);
or U14640 (N_14640,N_14236,N_14299);
nand U14641 (N_14641,N_14021,N_14174);
nand U14642 (N_14642,N_14078,N_14186);
nand U14643 (N_14643,N_14401,N_14008);
nand U14644 (N_14644,N_14332,N_14415);
nand U14645 (N_14645,N_14225,N_14111);
nand U14646 (N_14646,N_14249,N_14188);
nand U14647 (N_14647,N_14145,N_14412);
nand U14648 (N_14648,N_14024,N_14410);
nand U14649 (N_14649,N_14013,N_14164);
nor U14650 (N_14650,N_14114,N_14346);
nor U14651 (N_14651,N_14151,N_14232);
nand U14652 (N_14652,N_14197,N_14344);
and U14653 (N_14653,N_14170,N_14074);
or U14654 (N_14654,N_14051,N_14283);
nand U14655 (N_14655,N_14193,N_14105);
xnor U14656 (N_14656,N_14293,N_14208);
nor U14657 (N_14657,N_14459,N_14097);
or U14658 (N_14658,N_14252,N_14195);
or U14659 (N_14659,N_14212,N_14272);
nor U14660 (N_14660,N_14486,N_14147);
or U14661 (N_14661,N_14328,N_14251);
nand U14662 (N_14662,N_14005,N_14392);
nand U14663 (N_14663,N_14211,N_14194);
xnor U14664 (N_14664,N_14470,N_14156);
nor U14665 (N_14665,N_14075,N_14382);
nand U14666 (N_14666,N_14495,N_14303);
or U14667 (N_14667,N_14122,N_14056);
xor U14668 (N_14668,N_14341,N_14418);
nor U14669 (N_14669,N_14327,N_14307);
nand U14670 (N_14670,N_14200,N_14323);
xor U14671 (N_14671,N_14046,N_14084);
nor U14672 (N_14672,N_14324,N_14155);
nor U14673 (N_14673,N_14049,N_14162);
nand U14674 (N_14674,N_14259,N_14308);
nor U14675 (N_14675,N_14429,N_14083);
and U14676 (N_14676,N_14425,N_14286);
nand U14677 (N_14677,N_14173,N_14143);
nand U14678 (N_14678,N_14133,N_14086);
xor U14679 (N_14679,N_14178,N_14318);
or U14680 (N_14680,N_14386,N_14305);
nand U14681 (N_14681,N_14355,N_14279);
and U14682 (N_14682,N_14468,N_14390);
nor U14683 (N_14683,N_14142,N_14101);
nand U14684 (N_14684,N_14369,N_14165);
nor U14685 (N_14685,N_14131,N_14050);
or U14686 (N_14686,N_14350,N_14423);
nor U14687 (N_14687,N_14233,N_14288);
nand U14688 (N_14688,N_14218,N_14093);
nand U14689 (N_14689,N_14107,N_14484);
or U14690 (N_14690,N_14380,N_14087);
nand U14691 (N_14691,N_14330,N_14125);
nor U14692 (N_14692,N_14009,N_14060);
nor U14693 (N_14693,N_14248,N_14267);
xor U14694 (N_14694,N_14342,N_14460);
and U14695 (N_14695,N_14176,N_14080);
or U14696 (N_14696,N_14034,N_14496);
and U14697 (N_14697,N_14427,N_14160);
nand U14698 (N_14698,N_14017,N_14246);
and U14699 (N_14699,N_14331,N_14454);
nor U14700 (N_14700,N_14263,N_14201);
or U14701 (N_14701,N_14062,N_14231);
nand U14702 (N_14702,N_14152,N_14094);
and U14703 (N_14703,N_14467,N_14117);
nand U14704 (N_14704,N_14319,N_14042);
nor U14705 (N_14705,N_14179,N_14149);
xor U14706 (N_14706,N_14138,N_14282);
nand U14707 (N_14707,N_14406,N_14136);
and U14708 (N_14708,N_14485,N_14029);
nand U14709 (N_14709,N_14477,N_14163);
nand U14710 (N_14710,N_14491,N_14109);
nor U14711 (N_14711,N_14358,N_14245);
nor U14712 (N_14712,N_14192,N_14451);
or U14713 (N_14713,N_14061,N_14397);
or U14714 (N_14714,N_14135,N_14426);
xor U14715 (N_14715,N_14230,N_14072);
xor U14716 (N_14716,N_14475,N_14106);
and U14717 (N_14717,N_14337,N_14408);
and U14718 (N_14718,N_14322,N_14411);
or U14719 (N_14719,N_14443,N_14182);
nand U14720 (N_14720,N_14127,N_14169);
and U14721 (N_14721,N_14464,N_14064);
and U14722 (N_14722,N_14137,N_14493);
xor U14723 (N_14723,N_14166,N_14002);
or U14724 (N_14724,N_14022,N_14413);
nor U14725 (N_14725,N_14053,N_14421);
nor U14726 (N_14726,N_14146,N_14483);
nand U14727 (N_14727,N_14428,N_14345);
xnor U14728 (N_14728,N_14296,N_14235);
nand U14729 (N_14729,N_14385,N_14424);
xor U14730 (N_14730,N_14035,N_14065);
nand U14731 (N_14731,N_14381,N_14403);
nand U14732 (N_14732,N_14038,N_14196);
or U14733 (N_14733,N_14128,N_14340);
nor U14734 (N_14734,N_14275,N_14494);
and U14735 (N_14735,N_14280,N_14216);
nor U14736 (N_14736,N_14409,N_14150);
or U14737 (N_14737,N_14326,N_14090);
and U14738 (N_14738,N_14456,N_14298);
or U14739 (N_14739,N_14198,N_14011);
nand U14740 (N_14740,N_14349,N_14181);
and U14741 (N_14741,N_14027,N_14335);
nand U14742 (N_14742,N_14365,N_14480);
and U14743 (N_14743,N_14317,N_14312);
or U14744 (N_14744,N_14126,N_14202);
nand U14745 (N_14745,N_14255,N_14363);
nor U14746 (N_14746,N_14130,N_14436);
nor U14747 (N_14747,N_14289,N_14269);
nor U14748 (N_14748,N_14244,N_14237);
nand U14749 (N_14749,N_14139,N_14394);
or U14750 (N_14750,N_14479,N_14395);
nand U14751 (N_14751,N_14075,N_14047);
nor U14752 (N_14752,N_14308,N_14294);
or U14753 (N_14753,N_14467,N_14112);
or U14754 (N_14754,N_14286,N_14196);
and U14755 (N_14755,N_14031,N_14174);
or U14756 (N_14756,N_14431,N_14167);
nor U14757 (N_14757,N_14237,N_14192);
nand U14758 (N_14758,N_14394,N_14360);
xnor U14759 (N_14759,N_14003,N_14466);
or U14760 (N_14760,N_14006,N_14393);
or U14761 (N_14761,N_14236,N_14259);
and U14762 (N_14762,N_14497,N_14192);
or U14763 (N_14763,N_14301,N_14106);
nand U14764 (N_14764,N_14326,N_14444);
or U14765 (N_14765,N_14387,N_14486);
nor U14766 (N_14766,N_14335,N_14285);
nand U14767 (N_14767,N_14412,N_14212);
and U14768 (N_14768,N_14108,N_14277);
or U14769 (N_14769,N_14293,N_14127);
or U14770 (N_14770,N_14161,N_14233);
or U14771 (N_14771,N_14074,N_14234);
xor U14772 (N_14772,N_14408,N_14437);
and U14773 (N_14773,N_14181,N_14463);
or U14774 (N_14774,N_14155,N_14387);
nand U14775 (N_14775,N_14183,N_14274);
nand U14776 (N_14776,N_14046,N_14137);
nor U14777 (N_14777,N_14368,N_14207);
nand U14778 (N_14778,N_14194,N_14364);
nand U14779 (N_14779,N_14098,N_14001);
xnor U14780 (N_14780,N_14157,N_14246);
xnor U14781 (N_14781,N_14416,N_14071);
nor U14782 (N_14782,N_14152,N_14111);
nand U14783 (N_14783,N_14446,N_14195);
nand U14784 (N_14784,N_14315,N_14248);
or U14785 (N_14785,N_14447,N_14483);
nor U14786 (N_14786,N_14030,N_14077);
xor U14787 (N_14787,N_14366,N_14389);
and U14788 (N_14788,N_14404,N_14393);
and U14789 (N_14789,N_14115,N_14470);
xor U14790 (N_14790,N_14186,N_14350);
nor U14791 (N_14791,N_14408,N_14094);
and U14792 (N_14792,N_14328,N_14120);
or U14793 (N_14793,N_14087,N_14154);
nor U14794 (N_14794,N_14477,N_14324);
nand U14795 (N_14795,N_14123,N_14071);
xnor U14796 (N_14796,N_14232,N_14108);
or U14797 (N_14797,N_14250,N_14364);
nand U14798 (N_14798,N_14394,N_14148);
or U14799 (N_14799,N_14366,N_14120);
nor U14800 (N_14800,N_14144,N_14363);
and U14801 (N_14801,N_14352,N_14368);
or U14802 (N_14802,N_14472,N_14074);
or U14803 (N_14803,N_14190,N_14086);
nor U14804 (N_14804,N_14060,N_14260);
nor U14805 (N_14805,N_14386,N_14416);
or U14806 (N_14806,N_14291,N_14322);
or U14807 (N_14807,N_14223,N_14430);
xor U14808 (N_14808,N_14261,N_14440);
xnor U14809 (N_14809,N_14221,N_14061);
nand U14810 (N_14810,N_14272,N_14454);
and U14811 (N_14811,N_14111,N_14075);
xor U14812 (N_14812,N_14010,N_14262);
nor U14813 (N_14813,N_14385,N_14301);
nand U14814 (N_14814,N_14158,N_14299);
nor U14815 (N_14815,N_14380,N_14497);
xnor U14816 (N_14816,N_14471,N_14325);
and U14817 (N_14817,N_14484,N_14407);
or U14818 (N_14818,N_14145,N_14448);
nand U14819 (N_14819,N_14430,N_14140);
xor U14820 (N_14820,N_14311,N_14455);
nor U14821 (N_14821,N_14308,N_14330);
and U14822 (N_14822,N_14172,N_14378);
nor U14823 (N_14823,N_14251,N_14205);
xor U14824 (N_14824,N_14376,N_14080);
and U14825 (N_14825,N_14497,N_14285);
nand U14826 (N_14826,N_14445,N_14465);
xnor U14827 (N_14827,N_14438,N_14311);
or U14828 (N_14828,N_14492,N_14216);
and U14829 (N_14829,N_14043,N_14058);
or U14830 (N_14830,N_14164,N_14159);
nand U14831 (N_14831,N_14165,N_14166);
and U14832 (N_14832,N_14190,N_14098);
nand U14833 (N_14833,N_14415,N_14004);
and U14834 (N_14834,N_14131,N_14492);
and U14835 (N_14835,N_14000,N_14374);
nand U14836 (N_14836,N_14173,N_14380);
and U14837 (N_14837,N_14230,N_14148);
or U14838 (N_14838,N_14264,N_14162);
or U14839 (N_14839,N_14228,N_14398);
nand U14840 (N_14840,N_14040,N_14106);
or U14841 (N_14841,N_14316,N_14373);
nor U14842 (N_14842,N_14189,N_14279);
or U14843 (N_14843,N_14256,N_14002);
nor U14844 (N_14844,N_14166,N_14490);
nor U14845 (N_14845,N_14474,N_14370);
nand U14846 (N_14846,N_14242,N_14261);
xor U14847 (N_14847,N_14072,N_14169);
xor U14848 (N_14848,N_14029,N_14259);
nor U14849 (N_14849,N_14098,N_14474);
or U14850 (N_14850,N_14209,N_14382);
nor U14851 (N_14851,N_14246,N_14311);
and U14852 (N_14852,N_14123,N_14489);
xor U14853 (N_14853,N_14358,N_14247);
xnor U14854 (N_14854,N_14487,N_14214);
xor U14855 (N_14855,N_14381,N_14108);
xnor U14856 (N_14856,N_14446,N_14088);
or U14857 (N_14857,N_14472,N_14200);
and U14858 (N_14858,N_14359,N_14336);
nand U14859 (N_14859,N_14073,N_14480);
xnor U14860 (N_14860,N_14252,N_14396);
xor U14861 (N_14861,N_14352,N_14196);
xnor U14862 (N_14862,N_14074,N_14069);
and U14863 (N_14863,N_14007,N_14308);
nor U14864 (N_14864,N_14079,N_14212);
or U14865 (N_14865,N_14264,N_14161);
nand U14866 (N_14866,N_14259,N_14458);
or U14867 (N_14867,N_14071,N_14181);
or U14868 (N_14868,N_14407,N_14262);
nand U14869 (N_14869,N_14376,N_14166);
nand U14870 (N_14870,N_14343,N_14259);
nand U14871 (N_14871,N_14310,N_14419);
xor U14872 (N_14872,N_14092,N_14050);
xor U14873 (N_14873,N_14170,N_14285);
and U14874 (N_14874,N_14414,N_14061);
and U14875 (N_14875,N_14379,N_14007);
and U14876 (N_14876,N_14330,N_14397);
or U14877 (N_14877,N_14259,N_14382);
and U14878 (N_14878,N_14472,N_14492);
or U14879 (N_14879,N_14066,N_14069);
nand U14880 (N_14880,N_14111,N_14088);
or U14881 (N_14881,N_14448,N_14150);
or U14882 (N_14882,N_14419,N_14083);
or U14883 (N_14883,N_14068,N_14376);
nand U14884 (N_14884,N_14402,N_14346);
and U14885 (N_14885,N_14307,N_14044);
or U14886 (N_14886,N_14021,N_14340);
xor U14887 (N_14887,N_14412,N_14391);
nand U14888 (N_14888,N_14031,N_14136);
and U14889 (N_14889,N_14237,N_14248);
nor U14890 (N_14890,N_14339,N_14236);
nor U14891 (N_14891,N_14453,N_14128);
xnor U14892 (N_14892,N_14118,N_14286);
xnor U14893 (N_14893,N_14342,N_14309);
and U14894 (N_14894,N_14405,N_14413);
or U14895 (N_14895,N_14279,N_14499);
and U14896 (N_14896,N_14462,N_14217);
and U14897 (N_14897,N_14495,N_14463);
nand U14898 (N_14898,N_14205,N_14239);
and U14899 (N_14899,N_14355,N_14367);
nor U14900 (N_14900,N_14442,N_14386);
nor U14901 (N_14901,N_14320,N_14078);
nand U14902 (N_14902,N_14200,N_14487);
xnor U14903 (N_14903,N_14267,N_14495);
and U14904 (N_14904,N_14159,N_14371);
and U14905 (N_14905,N_14327,N_14170);
or U14906 (N_14906,N_14027,N_14074);
nand U14907 (N_14907,N_14487,N_14206);
xor U14908 (N_14908,N_14419,N_14210);
or U14909 (N_14909,N_14488,N_14249);
nand U14910 (N_14910,N_14128,N_14144);
nand U14911 (N_14911,N_14179,N_14176);
xnor U14912 (N_14912,N_14238,N_14407);
nand U14913 (N_14913,N_14254,N_14133);
nor U14914 (N_14914,N_14178,N_14466);
nor U14915 (N_14915,N_14430,N_14270);
nand U14916 (N_14916,N_14144,N_14279);
nand U14917 (N_14917,N_14466,N_14266);
nand U14918 (N_14918,N_14199,N_14337);
and U14919 (N_14919,N_14235,N_14481);
xor U14920 (N_14920,N_14390,N_14491);
xnor U14921 (N_14921,N_14399,N_14394);
xor U14922 (N_14922,N_14456,N_14209);
and U14923 (N_14923,N_14366,N_14065);
xor U14924 (N_14924,N_14089,N_14439);
xor U14925 (N_14925,N_14277,N_14011);
nand U14926 (N_14926,N_14227,N_14485);
nor U14927 (N_14927,N_14182,N_14069);
or U14928 (N_14928,N_14061,N_14287);
and U14929 (N_14929,N_14289,N_14277);
or U14930 (N_14930,N_14255,N_14150);
nor U14931 (N_14931,N_14288,N_14024);
or U14932 (N_14932,N_14023,N_14186);
xor U14933 (N_14933,N_14427,N_14134);
and U14934 (N_14934,N_14424,N_14059);
xor U14935 (N_14935,N_14102,N_14114);
and U14936 (N_14936,N_14381,N_14241);
and U14937 (N_14937,N_14378,N_14451);
nor U14938 (N_14938,N_14216,N_14266);
and U14939 (N_14939,N_14233,N_14176);
nor U14940 (N_14940,N_14017,N_14327);
or U14941 (N_14941,N_14098,N_14232);
and U14942 (N_14942,N_14442,N_14301);
and U14943 (N_14943,N_14121,N_14327);
and U14944 (N_14944,N_14197,N_14229);
and U14945 (N_14945,N_14049,N_14372);
nand U14946 (N_14946,N_14371,N_14116);
nand U14947 (N_14947,N_14392,N_14242);
xor U14948 (N_14948,N_14240,N_14211);
nand U14949 (N_14949,N_14259,N_14063);
nand U14950 (N_14950,N_14428,N_14336);
xor U14951 (N_14951,N_14049,N_14045);
nor U14952 (N_14952,N_14140,N_14071);
and U14953 (N_14953,N_14263,N_14151);
and U14954 (N_14954,N_14194,N_14083);
and U14955 (N_14955,N_14463,N_14433);
xor U14956 (N_14956,N_14218,N_14278);
nor U14957 (N_14957,N_14310,N_14114);
xor U14958 (N_14958,N_14352,N_14460);
and U14959 (N_14959,N_14467,N_14305);
or U14960 (N_14960,N_14370,N_14055);
nor U14961 (N_14961,N_14298,N_14153);
nand U14962 (N_14962,N_14002,N_14346);
or U14963 (N_14963,N_14433,N_14368);
xor U14964 (N_14964,N_14395,N_14107);
xor U14965 (N_14965,N_14451,N_14113);
xor U14966 (N_14966,N_14209,N_14428);
nor U14967 (N_14967,N_14064,N_14152);
or U14968 (N_14968,N_14043,N_14461);
or U14969 (N_14969,N_14137,N_14413);
nand U14970 (N_14970,N_14122,N_14389);
or U14971 (N_14971,N_14069,N_14416);
or U14972 (N_14972,N_14077,N_14459);
or U14973 (N_14973,N_14354,N_14338);
and U14974 (N_14974,N_14113,N_14121);
and U14975 (N_14975,N_14324,N_14060);
nand U14976 (N_14976,N_14084,N_14022);
nand U14977 (N_14977,N_14498,N_14145);
xnor U14978 (N_14978,N_14016,N_14440);
and U14979 (N_14979,N_14394,N_14107);
xor U14980 (N_14980,N_14369,N_14328);
nand U14981 (N_14981,N_14116,N_14111);
xnor U14982 (N_14982,N_14435,N_14426);
nor U14983 (N_14983,N_14375,N_14059);
nand U14984 (N_14984,N_14466,N_14126);
or U14985 (N_14985,N_14148,N_14262);
and U14986 (N_14986,N_14436,N_14154);
nor U14987 (N_14987,N_14362,N_14283);
and U14988 (N_14988,N_14322,N_14428);
nor U14989 (N_14989,N_14272,N_14276);
xnor U14990 (N_14990,N_14189,N_14106);
nand U14991 (N_14991,N_14385,N_14225);
or U14992 (N_14992,N_14317,N_14009);
nand U14993 (N_14993,N_14173,N_14485);
nand U14994 (N_14994,N_14256,N_14280);
or U14995 (N_14995,N_14382,N_14079);
nand U14996 (N_14996,N_14442,N_14215);
and U14997 (N_14997,N_14430,N_14412);
nor U14998 (N_14998,N_14103,N_14442);
nor U14999 (N_14999,N_14386,N_14014);
or U15000 (N_15000,N_14539,N_14534);
nor U15001 (N_15001,N_14797,N_14576);
or U15002 (N_15002,N_14923,N_14617);
nand U15003 (N_15003,N_14513,N_14888);
and U15004 (N_15004,N_14804,N_14932);
or U15005 (N_15005,N_14670,N_14502);
nand U15006 (N_15006,N_14922,N_14725);
nor U15007 (N_15007,N_14986,N_14575);
or U15008 (N_15008,N_14963,N_14755);
xnor U15009 (N_15009,N_14500,N_14561);
and U15010 (N_15010,N_14763,N_14876);
nor U15011 (N_15011,N_14880,N_14759);
or U15012 (N_15012,N_14529,N_14770);
or U15013 (N_15013,N_14998,N_14895);
and U15014 (N_15014,N_14659,N_14852);
nor U15015 (N_15015,N_14785,N_14811);
xnor U15016 (N_15016,N_14819,N_14648);
and U15017 (N_15017,N_14574,N_14959);
nand U15018 (N_15018,N_14765,N_14739);
xnor U15019 (N_15019,N_14704,N_14847);
or U15020 (N_15020,N_14691,N_14597);
or U15021 (N_15021,N_14610,N_14793);
xnor U15022 (N_15022,N_14622,N_14948);
nand U15023 (N_15023,N_14593,N_14536);
and U15024 (N_15024,N_14666,N_14857);
nor U15025 (N_15025,N_14911,N_14612);
and U15026 (N_15026,N_14885,N_14631);
nand U15027 (N_15027,N_14916,N_14958);
nor U15028 (N_15028,N_14594,N_14680);
nand U15029 (N_15029,N_14766,N_14938);
or U15030 (N_15030,N_14525,N_14578);
or U15031 (N_15031,N_14787,N_14689);
xor U15032 (N_15032,N_14940,N_14969);
or U15033 (N_15033,N_14786,N_14915);
nand U15034 (N_15034,N_14508,N_14868);
and U15035 (N_15035,N_14736,N_14873);
or U15036 (N_15036,N_14867,N_14552);
or U15037 (N_15037,N_14961,N_14834);
nor U15038 (N_15038,N_14846,N_14606);
xnor U15039 (N_15039,N_14562,N_14646);
nor U15040 (N_15040,N_14935,N_14853);
nor U15041 (N_15041,N_14924,N_14907);
and U15042 (N_15042,N_14828,N_14690);
and U15043 (N_15043,N_14727,N_14798);
and U15044 (N_15044,N_14845,N_14750);
xor U15045 (N_15045,N_14545,N_14544);
nand U15046 (N_15046,N_14625,N_14627);
or U15047 (N_15047,N_14843,N_14955);
and U15048 (N_15048,N_14554,N_14548);
and U15049 (N_15049,N_14814,N_14863);
and U15050 (N_15050,N_14564,N_14501);
nand U15051 (N_15051,N_14897,N_14975);
xnor U15052 (N_15052,N_14609,N_14920);
nand U15053 (N_15053,N_14607,N_14862);
or U15054 (N_15054,N_14592,N_14683);
or U15055 (N_15055,N_14778,N_14864);
nor U15056 (N_15056,N_14957,N_14790);
xor U15057 (N_15057,N_14926,N_14737);
nor U15058 (N_15058,N_14717,N_14914);
xor U15059 (N_15059,N_14818,N_14912);
nor U15060 (N_15060,N_14875,N_14726);
nand U15061 (N_15061,N_14568,N_14692);
or U15062 (N_15062,N_14524,N_14638);
and U15063 (N_15063,N_14619,N_14655);
nand U15064 (N_15064,N_14710,N_14767);
nand U15065 (N_15065,N_14591,N_14604);
xnor U15066 (N_15066,N_14669,N_14700);
nor U15067 (N_15067,N_14516,N_14694);
nor U15068 (N_15068,N_14891,N_14728);
and U15069 (N_15069,N_14647,N_14799);
xnor U15070 (N_15070,N_14849,N_14719);
or U15071 (N_15071,N_14774,N_14553);
or U15072 (N_15072,N_14526,N_14898);
or U15073 (N_15073,N_14510,N_14679);
and U15074 (N_15074,N_14662,N_14972);
nand U15075 (N_15075,N_14893,N_14599);
or U15076 (N_15076,N_14964,N_14733);
or U15077 (N_15077,N_14543,N_14577);
nand U15078 (N_15078,N_14702,N_14688);
or U15079 (N_15079,N_14663,N_14974);
nor U15080 (N_15080,N_14829,N_14987);
nor U15081 (N_15081,N_14514,N_14760);
xnor U15082 (N_15082,N_14518,N_14716);
nand U15083 (N_15083,N_14677,N_14933);
nor U15084 (N_15084,N_14980,N_14632);
nand U15085 (N_15085,N_14644,N_14567);
nor U15086 (N_15086,N_14678,N_14565);
or U15087 (N_15087,N_14628,N_14626);
nor U15088 (N_15088,N_14832,N_14573);
nor U15089 (N_15089,N_14754,N_14503);
nor U15090 (N_15090,N_14533,N_14855);
xor U15091 (N_15091,N_14676,N_14571);
nand U15092 (N_15092,N_14584,N_14990);
and U15093 (N_15093,N_14674,N_14996);
nand U15094 (N_15094,N_14640,N_14944);
nor U15095 (N_15095,N_14967,N_14758);
nor U15096 (N_15096,N_14721,N_14901);
xor U15097 (N_15097,N_14656,N_14921);
or U15098 (N_15098,N_14781,N_14848);
xnor U15099 (N_15099,N_14634,N_14950);
or U15100 (N_15100,N_14751,N_14879);
and U15101 (N_15101,N_14796,N_14817);
nor U15102 (N_15102,N_14805,N_14742);
or U15103 (N_15103,N_14587,N_14757);
nor U15104 (N_15104,N_14989,N_14773);
and U15105 (N_15105,N_14635,N_14777);
nand U15106 (N_15106,N_14673,N_14572);
and U15107 (N_15107,N_14801,N_14771);
nor U15108 (N_15108,N_14546,N_14899);
xor U15109 (N_15109,N_14951,N_14511);
nand U15110 (N_15110,N_14675,N_14650);
nor U15111 (N_15111,N_14512,N_14822);
or U15112 (N_15112,N_14639,N_14743);
and U15113 (N_15113,N_14858,N_14839);
nand U15114 (N_15114,N_14782,N_14703);
nand U15115 (N_15115,N_14715,N_14837);
or U15116 (N_15116,N_14841,N_14976);
and U15117 (N_15117,N_14658,N_14555);
nand U15118 (N_15118,N_14913,N_14515);
xnor U15119 (N_15119,N_14722,N_14667);
nor U15120 (N_15120,N_14874,N_14827);
xnor U15121 (N_15121,N_14842,N_14713);
or U15122 (N_15122,N_14551,N_14586);
nor U15123 (N_15123,N_14971,N_14535);
xor U15124 (N_15124,N_14791,N_14992);
xor U15125 (N_15125,N_14560,N_14633);
xnor U15126 (N_15126,N_14783,N_14825);
xor U15127 (N_15127,N_14746,N_14865);
nor U15128 (N_15128,N_14910,N_14854);
nor U15129 (N_15129,N_14982,N_14960);
or U15130 (N_15130,N_14735,N_14894);
or U15131 (N_15131,N_14823,N_14869);
and U15132 (N_15132,N_14711,N_14517);
xor U15133 (N_15133,N_14657,N_14753);
and U15134 (N_15134,N_14954,N_14589);
or U15135 (N_15135,N_14764,N_14952);
or U15136 (N_15136,N_14686,N_14820);
nor U15137 (N_15137,N_14664,N_14671);
nand U15138 (N_15138,N_14831,N_14844);
xnor U15139 (N_15139,N_14979,N_14541);
xnor U15140 (N_15140,N_14630,N_14557);
and U15141 (N_15141,N_14925,N_14707);
nor U15142 (N_15142,N_14613,N_14918);
nand U15143 (N_15143,N_14614,N_14549);
xnor U15144 (N_15144,N_14984,N_14883);
and U15145 (N_15145,N_14927,N_14946);
nand U15146 (N_15146,N_14917,N_14570);
nand U15147 (N_15147,N_14537,N_14596);
or U15148 (N_15148,N_14652,N_14772);
and U15149 (N_15149,N_14813,N_14520);
or U15150 (N_15150,N_14642,N_14697);
nand U15151 (N_15151,N_14569,N_14623);
xor U15152 (N_15152,N_14929,N_14705);
xnor U15153 (N_15153,N_14977,N_14890);
nor U15154 (N_15154,N_14540,N_14824);
and U15155 (N_15155,N_14991,N_14838);
or U15156 (N_15156,N_14882,N_14878);
and U15157 (N_15157,N_14809,N_14579);
nand U15158 (N_15158,N_14800,N_14653);
and U15159 (N_15159,N_14872,N_14601);
xnor U15160 (N_15160,N_14660,N_14744);
nand U15161 (N_15161,N_14902,N_14611);
and U15162 (N_15162,N_14507,N_14840);
and U15163 (N_15163,N_14775,N_14695);
nor U15164 (N_15164,N_14509,N_14956);
and U15165 (N_15165,N_14608,N_14931);
nor U15166 (N_15166,N_14745,N_14881);
nor U15167 (N_15167,N_14877,N_14884);
nand U15168 (N_15168,N_14906,N_14618);
nor U15169 (N_15169,N_14649,N_14706);
or U15170 (N_15170,N_14637,N_14965);
xor U15171 (N_15171,N_14966,N_14600);
nand U15172 (N_15172,N_14768,N_14731);
xnor U15173 (N_15173,N_14860,N_14833);
nand U15174 (N_15174,N_14693,N_14896);
and U15175 (N_15175,N_14522,N_14826);
or U15176 (N_15176,N_14523,N_14563);
xnor U15177 (N_15177,N_14581,N_14714);
nor U15178 (N_15178,N_14740,N_14761);
and U15179 (N_15179,N_14661,N_14682);
or U15180 (N_15180,N_14803,N_14550);
nand U15181 (N_15181,N_14780,N_14530);
and U15182 (N_15182,N_14784,N_14821);
or U15183 (N_15183,N_14684,N_14668);
nor U15184 (N_15184,N_14978,N_14590);
and U15185 (N_15185,N_14851,N_14995);
nor U15186 (N_15186,N_14943,N_14724);
nor U15187 (N_15187,N_14506,N_14905);
nor U15188 (N_15188,N_14732,N_14580);
and U15189 (N_15189,N_14730,N_14605);
and U15190 (N_15190,N_14741,N_14701);
and U15191 (N_15191,N_14542,N_14887);
nor U15192 (N_15192,N_14687,N_14947);
nand U15193 (N_15193,N_14930,N_14808);
and U15194 (N_15194,N_14504,N_14538);
or U15195 (N_15195,N_14696,N_14624);
xor U15196 (N_15196,N_14531,N_14685);
xnor U15197 (N_15197,N_14934,N_14962);
or U15198 (N_15198,N_14942,N_14861);
and U15199 (N_15199,N_14908,N_14997);
and U15200 (N_15200,N_14866,N_14900);
nand U15201 (N_15201,N_14672,N_14709);
nor U15202 (N_15202,N_14532,N_14810);
and U15203 (N_15203,N_14598,N_14681);
nor U15204 (N_15204,N_14892,N_14723);
nor U15205 (N_15205,N_14953,N_14643);
nand U15206 (N_15206,N_14651,N_14889);
xnor U15207 (N_15207,N_14558,N_14812);
nor U15208 (N_15208,N_14527,N_14973);
xor U15209 (N_15209,N_14999,N_14788);
and U15210 (N_15210,N_14939,N_14779);
or U15211 (N_15211,N_14936,N_14985);
or U15212 (N_15212,N_14871,N_14665);
nand U15213 (N_15213,N_14699,N_14856);
xnor U15214 (N_15214,N_14928,N_14830);
nand U15215 (N_15215,N_14835,N_14582);
nor U15216 (N_15216,N_14993,N_14983);
nand U15217 (N_15217,N_14749,N_14792);
nand U15218 (N_15218,N_14968,N_14904);
xor U15219 (N_15219,N_14615,N_14949);
or U15220 (N_15220,N_14718,N_14595);
or U15221 (N_15221,N_14945,N_14603);
or U15222 (N_15222,N_14528,N_14886);
nor U15223 (N_15223,N_14519,N_14836);
or U15224 (N_15224,N_14970,N_14981);
and U15225 (N_15225,N_14641,N_14566);
xnor U15226 (N_15226,N_14698,N_14620);
and U15227 (N_15227,N_14602,N_14521);
xnor U15228 (N_15228,N_14756,N_14769);
and U15229 (N_15229,N_14616,N_14729);
or U15230 (N_15230,N_14816,N_14815);
nor U15231 (N_15231,N_14988,N_14941);
xnor U15232 (N_15232,N_14629,N_14583);
nor U15233 (N_15233,N_14794,N_14909);
or U15234 (N_15234,N_14734,N_14547);
and U15235 (N_15235,N_14645,N_14795);
xnor U15236 (N_15236,N_14802,N_14559);
xor U15237 (N_15237,N_14654,N_14870);
xnor U15238 (N_15238,N_14994,N_14903);
xnor U15239 (N_15239,N_14708,N_14738);
and U15240 (N_15240,N_14789,N_14621);
nor U15241 (N_15241,N_14807,N_14747);
nor U15242 (N_15242,N_14752,N_14859);
nand U15243 (N_15243,N_14748,N_14636);
or U15244 (N_15244,N_14712,N_14556);
or U15245 (N_15245,N_14850,N_14720);
xnor U15246 (N_15246,N_14505,N_14588);
nor U15247 (N_15247,N_14776,N_14937);
xor U15248 (N_15248,N_14585,N_14806);
or U15249 (N_15249,N_14919,N_14762);
nand U15250 (N_15250,N_14889,N_14766);
xor U15251 (N_15251,N_14600,N_14630);
nand U15252 (N_15252,N_14677,N_14668);
nor U15253 (N_15253,N_14681,N_14672);
nor U15254 (N_15254,N_14719,N_14958);
and U15255 (N_15255,N_14518,N_14899);
nor U15256 (N_15256,N_14864,N_14902);
nor U15257 (N_15257,N_14629,N_14567);
nand U15258 (N_15258,N_14821,N_14569);
nor U15259 (N_15259,N_14912,N_14508);
and U15260 (N_15260,N_14788,N_14507);
and U15261 (N_15261,N_14555,N_14503);
nand U15262 (N_15262,N_14941,N_14963);
nand U15263 (N_15263,N_14990,N_14764);
or U15264 (N_15264,N_14519,N_14984);
nor U15265 (N_15265,N_14945,N_14881);
or U15266 (N_15266,N_14953,N_14937);
or U15267 (N_15267,N_14834,N_14892);
and U15268 (N_15268,N_14523,N_14693);
or U15269 (N_15269,N_14559,N_14841);
and U15270 (N_15270,N_14629,N_14612);
or U15271 (N_15271,N_14569,N_14596);
xnor U15272 (N_15272,N_14724,N_14843);
xor U15273 (N_15273,N_14667,N_14599);
xnor U15274 (N_15274,N_14858,N_14910);
nor U15275 (N_15275,N_14883,N_14587);
nand U15276 (N_15276,N_14746,N_14893);
nor U15277 (N_15277,N_14861,N_14580);
and U15278 (N_15278,N_14772,N_14842);
and U15279 (N_15279,N_14694,N_14925);
nand U15280 (N_15280,N_14673,N_14919);
nor U15281 (N_15281,N_14502,N_14800);
nand U15282 (N_15282,N_14610,N_14967);
nand U15283 (N_15283,N_14768,N_14880);
nand U15284 (N_15284,N_14686,N_14569);
and U15285 (N_15285,N_14779,N_14662);
or U15286 (N_15286,N_14900,N_14771);
or U15287 (N_15287,N_14648,N_14927);
or U15288 (N_15288,N_14884,N_14913);
and U15289 (N_15289,N_14849,N_14953);
nor U15290 (N_15290,N_14894,N_14848);
nand U15291 (N_15291,N_14891,N_14536);
xnor U15292 (N_15292,N_14945,N_14894);
nor U15293 (N_15293,N_14544,N_14855);
xor U15294 (N_15294,N_14839,N_14661);
or U15295 (N_15295,N_14751,N_14601);
nand U15296 (N_15296,N_14922,N_14908);
nand U15297 (N_15297,N_14683,N_14785);
nor U15298 (N_15298,N_14830,N_14879);
and U15299 (N_15299,N_14729,N_14999);
and U15300 (N_15300,N_14841,N_14887);
or U15301 (N_15301,N_14995,N_14935);
or U15302 (N_15302,N_14946,N_14788);
nor U15303 (N_15303,N_14970,N_14677);
and U15304 (N_15304,N_14637,N_14984);
or U15305 (N_15305,N_14928,N_14606);
or U15306 (N_15306,N_14959,N_14902);
and U15307 (N_15307,N_14715,N_14609);
or U15308 (N_15308,N_14759,N_14946);
xor U15309 (N_15309,N_14785,N_14810);
nand U15310 (N_15310,N_14826,N_14998);
nor U15311 (N_15311,N_14865,N_14936);
nand U15312 (N_15312,N_14997,N_14775);
nand U15313 (N_15313,N_14792,N_14928);
xor U15314 (N_15314,N_14945,N_14877);
or U15315 (N_15315,N_14673,N_14969);
and U15316 (N_15316,N_14936,N_14903);
nor U15317 (N_15317,N_14551,N_14721);
nor U15318 (N_15318,N_14773,N_14645);
nor U15319 (N_15319,N_14836,N_14817);
nand U15320 (N_15320,N_14746,N_14566);
or U15321 (N_15321,N_14777,N_14796);
xnor U15322 (N_15322,N_14905,N_14777);
nand U15323 (N_15323,N_14920,N_14597);
xor U15324 (N_15324,N_14744,N_14608);
and U15325 (N_15325,N_14821,N_14777);
xnor U15326 (N_15326,N_14741,N_14910);
nor U15327 (N_15327,N_14831,N_14503);
or U15328 (N_15328,N_14642,N_14519);
nor U15329 (N_15329,N_14690,N_14751);
nand U15330 (N_15330,N_14881,N_14693);
nand U15331 (N_15331,N_14968,N_14845);
xor U15332 (N_15332,N_14512,N_14642);
xnor U15333 (N_15333,N_14977,N_14987);
nor U15334 (N_15334,N_14800,N_14593);
nor U15335 (N_15335,N_14626,N_14669);
and U15336 (N_15336,N_14904,N_14818);
nor U15337 (N_15337,N_14832,N_14921);
nor U15338 (N_15338,N_14556,N_14564);
and U15339 (N_15339,N_14781,N_14785);
nor U15340 (N_15340,N_14862,N_14993);
or U15341 (N_15341,N_14693,N_14732);
nor U15342 (N_15342,N_14956,N_14592);
nand U15343 (N_15343,N_14842,N_14970);
nand U15344 (N_15344,N_14580,N_14695);
and U15345 (N_15345,N_14776,N_14818);
or U15346 (N_15346,N_14541,N_14831);
and U15347 (N_15347,N_14745,N_14577);
or U15348 (N_15348,N_14742,N_14555);
nand U15349 (N_15349,N_14952,N_14910);
and U15350 (N_15350,N_14515,N_14645);
nand U15351 (N_15351,N_14792,N_14530);
nor U15352 (N_15352,N_14521,N_14656);
nand U15353 (N_15353,N_14575,N_14515);
xnor U15354 (N_15354,N_14974,N_14737);
nand U15355 (N_15355,N_14730,N_14532);
or U15356 (N_15356,N_14796,N_14531);
nor U15357 (N_15357,N_14844,N_14864);
or U15358 (N_15358,N_14554,N_14787);
and U15359 (N_15359,N_14845,N_14976);
nor U15360 (N_15360,N_14866,N_14893);
xnor U15361 (N_15361,N_14846,N_14570);
nor U15362 (N_15362,N_14861,N_14817);
nor U15363 (N_15363,N_14962,N_14578);
and U15364 (N_15364,N_14770,N_14735);
nand U15365 (N_15365,N_14595,N_14979);
xnor U15366 (N_15366,N_14700,N_14653);
nand U15367 (N_15367,N_14612,N_14922);
or U15368 (N_15368,N_14865,N_14980);
or U15369 (N_15369,N_14750,N_14808);
nand U15370 (N_15370,N_14992,N_14766);
nand U15371 (N_15371,N_14694,N_14615);
nor U15372 (N_15372,N_14860,N_14999);
xor U15373 (N_15373,N_14580,N_14667);
nand U15374 (N_15374,N_14858,N_14694);
xor U15375 (N_15375,N_14898,N_14646);
and U15376 (N_15376,N_14777,N_14548);
or U15377 (N_15377,N_14839,N_14688);
or U15378 (N_15378,N_14761,N_14728);
xor U15379 (N_15379,N_14649,N_14835);
and U15380 (N_15380,N_14809,N_14533);
and U15381 (N_15381,N_14577,N_14578);
nand U15382 (N_15382,N_14772,N_14735);
and U15383 (N_15383,N_14625,N_14721);
xor U15384 (N_15384,N_14764,N_14978);
or U15385 (N_15385,N_14595,N_14705);
and U15386 (N_15386,N_14635,N_14620);
and U15387 (N_15387,N_14580,N_14705);
nand U15388 (N_15388,N_14888,N_14830);
nor U15389 (N_15389,N_14647,N_14901);
nor U15390 (N_15390,N_14931,N_14933);
nor U15391 (N_15391,N_14650,N_14920);
nor U15392 (N_15392,N_14946,N_14646);
nand U15393 (N_15393,N_14834,N_14532);
nand U15394 (N_15394,N_14828,N_14929);
nor U15395 (N_15395,N_14775,N_14834);
and U15396 (N_15396,N_14870,N_14788);
or U15397 (N_15397,N_14915,N_14651);
and U15398 (N_15398,N_14881,N_14716);
nand U15399 (N_15399,N_14500,N_14991);
or U15400 (N_15400,N_14785,N_14637);
or U15401 (N_15401,N_14628,N_14971);
xnor U15402 (N_15402,N_14937,N_14556);
nand U15403 (N_15403,N_14578,N_14716);
xor U15404 (N_15404,N_14705,N_14877);
nor U15405 (N_15405,N_14816,N_14728);
xor U15406 (N_15406,N_14941,N_14947);
nor U15407 (N_15407,N_14710,N_14548);
and U15408 (N_15408,N_14950,N_14967);
xnor U15409 (N_15409,N_14795,N_14573);
nor U15410 (N_15410,N_14790,N_14950);
xnor U15411 (N_15411,N_14777,N_14746);
xor U15412 (N_15412,N_14753,N_14789);
xnor U15413 (N_15413,N_14629,N_14517);
xnor U15414 (N_15414,N_14884,N_14692);
or U15415 (N_15415,N_14534,N_14804);
and U15416 (N_15416,N_14973,N_14910);
nor U15417 (N_15417,N_14608,N_14518);
and U15418 (N_15418,N_14968,N_14811);
xor U15419 (N_15419,N_14831,N_14951);
and U15420 (N_15420,N_14642,N_14841);
and U15421 (N_15421,N_14987,N_14860);
nor U15422 (N_15422,N_14514,N_14831);
and U15423 (N_15423,N_14943,N_14504);
xor U15424 (N_15424,N_14558,N_14538);
nor U15425 (N_15425,N_14541,N_14766);
nand U15426 (N_15426,N_14651,N_14624);
nor U15427 (N_15427,N_14823,N_14879);
xnor U15428 (N_15428,N_14756,N_14791);
nand U15429 (N_15429,N_14785,N_14551);
and U15430 (N_15430,N_14842,N_14923);
xnor U15431 (N_15431,N_14518,N_14788);
xnor U15432 (N_15432,N_14685,N_14940);
and U15433 (N_15433,N_14700,N_14969);
xnor U15434 (N_15434,N_14785,N_14853);
nor U15435 (N_15435,N_14985,N_14759);
and U15436 (N_15436,N_14585,N_14740);
xor U15437 (N_15437,N_14518,N_14712);
and U15438 (N_15438,N_14958,N_14524);
xor U15439 (N_15439,N_14975,N_14891);
xor U15440 (N_15440,N_14856,N_14968);
nor U15441 (N_15441,N_14896,N_14919);
and U15442 (N_15442,N_14517,N_14654);
nor U15443 (N_15443,N_14589,N_14786);
nand U15444 (N_15444,N_14630,N_14595);
or U15445 (N_15445,N_14906,N_14922);
and U15446 (N_15446,N_14729,N_14747);
nand U15447 (N_15447,N_14547,N_14501);
nor U15448 (N_15448,N_14822,N_14652);
xor U15449 (N_15449,N_14667,N_14608);
xnor U15450 (N_15450,N_14632,N_14567);
or U15451 (N_15451,N_14847,N_14862);
xor U15452 (N_15452,N_14933,N_14984);
and U15453 (N_15453,N_14537,N_14801);
xor U15454 (N_15454,N_14718,N_14584);
xnor U15455 (N_15455,N_14863,N_14568);
xnor U15456 (N_15456,N_14869,N_14736);
nand U15457 (N_15457,N_14811,N_14658);
and U15458 (N_15458,N_14527,N_14962);
or U15459 (N_15459,N_14595,N_14917);
nor U15460 (N_15460,N_14743,N_14526);
and U15461 (N_15461,N_14513,N_14751);
nor U15462 (N_15462,N_14658,N_14829);
nand U15463 (N_15463,N_14821,N_14735);
xnor U15464 (N_15464,N_14909,N_14718);
nand U15465 (N_15465,N_14723,N_14635);
nor U15466 (N_15466,N_14762,N_14932);
xor U15467 (N_15467,N_14647,N_14800);
or U15468 (N_15468,N_14859,N_14937);
nor U15469 (N_15469,N_14563,N_14848);
nand U15470 (N_15470,N_14896,N_14928);
nand U15471 (N_15471,N_14581,N_14636);
nand U15472 (N_15472,N_14864,N_14934);
xor U15473 (N_15473,N_14541,N_14697);
nor U15474 (N_15474,N_14667,N_14963);
xnor U15475 (N_15475,N_14807,N_14831);
nand U15476 (N_15476,N_14673,N_14566);
or U15477 (N_15477,N_14643,N_14853);
nand U15478 (N_15478,N_14859,N_14652);
nand U15479 (N_15479,N_14820,N_14601);
nor U15480 (N_15480,N_14582,N_14500);
nand U15481 (N_15481,N_14632,N_14818);
nand U15482 (N_15482,N_14548,N_14534);
nor U15483 (N_15483,N_14762,N_14561);
nor U15484 (N_15484,N_14816,N_14569);
nand U15485 (N_15485,N_14573,N_14593);
or U15486 (N_15486,N_14823,N_14994);
nor U15487 (N_15487,N_14772,N_14873);
or U15488 (N_15488,N_14638,N_14687);
and U15489 (N_15489,N_14809,N_14699);
or U15490 (N_15490,N_14887,N_14698);
xor U15491 (N_15491,N_14503,N_14614);
and U15492 (N_15492,N_14903,N_14864);
and U15493 (N_15493,N_14553,N_14819);
xnor U15494 (N_15494,N_14810,N_14816);
or U15495 (N_15495,N_14878,N_14640);
xor U15496 (N_15496,N_14624,N_14833);
or U15497 (N_15497,N_14810,N_14939);
xnor U15498 (N_15498,N_14806,N_14595);
nor U15499 (N_15499,N_14870,N_14847);
and U15500 (N_15500,N_15176,N_15384);
or U15501 (N_15501,N_15391,N_15070);
or U15502 (N_15502,N_15257,N_15405);
nand U15503 (N_15503,N_15228,N_15169);
nor U15504 (N_15504,N_15040,N_15146);
and U15505 (N_15505,N_15322,N_15382);
nand U15506 (N_15506,N_15251,N_15101);
nor U15507 (N_15507,N_15227,N_15387);
and U15508 (N_15508,N_15219,N_15300);
xor U15509 (N_15509,N_15184,N_15107);
xor U15510 (N_15510,N_15483,N_15167);
and U15511 (N_15511,N_15465,N_15256);
nand U15512 (N_15512,N_15094,N_15296);
xor U15513 (N_15513,N_15435,N_15341);
and U15514 (N_15514,N_15074,N_15024);
and U15515 (N_15515,N_15314,N_15245);
and U15516 (N_15516,N_15099,N_15374);
xor U15517 (N_15517,N_15434,N_15447);
and U15518 (N_15518,N_15338,N_15208);
and U15519 (N_15519,N_15444,N_15021);
xor U15520 (N_15520,N_15223,N_15105);
or U15521 (N_15521,N_15480,N_15095);
and U15522 (N_15522,N_15351,N_15274);
nor U15523 (N_15523,N_15306,N_15285);
xnor U15524 (N_15524,N_15267,N_15014);
nand U15525 (N_15525,N_15232,N_15453);
or U15526 (N_15526,N_15344,N_15038);
xnor U15527 (N_15527,N_15001,N_15211);
nor U15528 (N_15528,N_15277,N_15017);
nand U15529 (N_15529,N_15468,N_15416);
nand U15530 (N_15530,N_15034,N_15467);
nor U15531 (N_15531,N_15181,N_15250);
or U15532 (N_15532,N_15477,N_15497);
nor U15533 (N_15533,N_15226,N_15240);
xor U15534 (N_15534,N_15361,N_15195);
and U15535 (N_15535,N_15152,N_15090);
nand U15536 (N_15536,N_15263,N_15178);
or U15537 (N_15537,N_15421,N_15114);
nor U15538 (N_15538,N_15022,N_15424);
or U15539 (N_15539,N_15136,N_15316);
and U15540 (N_15540,N_15495,N_15264);
or U15541 (N_15541,N_15119,N_15047);
nor U15542 (N_15542,N_15403,N_15102);
nand U15543 (N_15543,N_15057,N_15259);
xor U15544 (N_15544,N_15145,N_15253);
xnor U15545 (N_15545,N_15224,N_15419);
xnor U15546 (N_15546,N_15270,N_15089);
nand U15547 (N_15547,N_15269,N_15121);
or U15548 (N_15548,N_15205,N_15364);
nand U15549 (N_15549,N_15078,N_15108);
or U15550 (N_15550,N_15430,N_15396);
nand U15551 (N_15551,N_15427,N_15097);
or U15552 (N_15552,N_15323,N_15206);
nand U15553 (N_15553,N_15473,N_15451);
nand U15554 (N_15554,N_15182,N_15423);
xor U15555 (N_15555,N_15366,N_15392);
and U15556 (N_15556,N_15254,N_15059);
or U15557 (N_15557,N_15312,N_15428);
or U15558 (N_15558,N_15415,N_15018);
xor U15559 (N_15559,N_15360,N_15383);
nor U15560 (N_15560,N_15093,N_15393);
nand U15561 (N_15561,N_15013,N_15476);
or U15562 (N_15562,N_15440,N_15303);
nor U15563 (N_15563,N_15048,N_15032);
and U15564 (N_15564,N_15412,N_15455);
nor U15565 (N_15565,N_15369,N_15413);
nand U15566 (N_15566,N_15156,N_15484);
or U15567 (N_15567,N_15050,N_15062);
xnor U15568 (N_15568,N_15190,N_15437);
or U15569 (N_15569,N_15456,N_15071);
nor U15570 (N_15570,N_15137,N_15399);
xnor U15571 (N_15571,N_15088,N_15160);
and U15572 (N_15572,N_15326,N_15367);
nand U15573 (N_15573,N_15112,N_15357);
xnor U15574 (N_15574,N_15164,N_15124);
xor U15575 (N_15575,N_15493,N_15289);
and U15576 (N_15576,N_15087,N_15340);
nand U15577 (N_15577,N_15450,N_15066);
or U15578 (N_15578,N_15307,N_15129);
nor U15579 (N_15579,N_15148,N_15298);
nand U15580 (N_15580,N_15449,N_15273);
nand U15581 (N_15581,N_15370,N_15487);
nor U15582 (N_15582,N_15420,N_15331);
xor U15583 (N_15583,N_15149,N_15309);
and U15584 (N_15584,N_15464,N_15459);
nor U15585 (N_15585,N_15131,N_15337);
and U15586 (N_15586,N_15045,N_15194);
nand U15587 (N_15587,N_15216,N_15239);
xor U15588 (N_15588,N_15359,N_15162);
nand U15589 (N_15589,N_15371,N_15261);
and U15590 (N_15590,N_15073,N_15400);
or U15591 (N_15591,N_15068,N_15395);
and U15592 (N_15592,N_15054,N_15422);
and U15593 (N_15593,N_15317,N_15083);
xnor U15594 (N_15594,N_15457,N_15011);
and U15595 (N_15595,N_15470,N_15436);
and U15596 (N_15596,N_15386,N_15329);
nor U15597 (N_15597,N_15486,N_15446);
and U15598 (N_15598,N_15220,N_15246);
and U15599 (N_15599,N_15077,N_15026);
nor U15600 (N_15600,N_15002,N_15321);
nor U15601 (N_15601,N_15212,N_15202);
or U15602 (N_15602,N_15043,N_15174);
xor U15603 (N_15603,N_15004,N_15474);
and U15604 (N_15604,N_15033,N_15041);
nor U15605 (N_15605,N_15260,N_15282);
xnor U15606 (N_15606,N_15499,N_15439);
or U15607 (N_15607,N_15117,N_15110);
nor U15608 (N_15608,N_15368,N_15354);
xnor U15609 (N_15609,N_15081,N_15381);
and U15610 (N_15610,N_15111,N_15086);
nor U15611 (N_15611,N_15198,N_15471);
xor U15612 (N_15612,N_15469,N_15299);
or U15613 (N_15613,N_15172,N_15379);
xor U15614 (N_15614,N_15333,N_15376);
and U15615 (N_15615,N_15179,N_15200);
xnor U15616 (N_15616,N_15452,N_15291);
and U15617 (N_15617,N_15052,N_15063);
nor U15618 (N_15618,N_15482,N_15204);
xor U15619 (N_15619,N_15377,N_15330);
or U15620 (N_15620,N_15056,N_15494);
nand U15621 (N_15621,N_15166,N_15460);
nand U15622 (N_15622,N_15217,N_15290);
xnor U15623 (N_15623,N_15003,N_15236);
and U15624 (N_15624,N_15008,N_15157);
nor U15625 (N_15625,N_15397,N_15142);
or U15626 (N_15626,N_15143,N_15007);
xnor U15627 (N_15627,N_15346,N_15044);
nor U15628 (N_15628,N_15127,N_15170);
and U15629 (N_15629,N_15378,N_15414);
xnor U15630 (N_15630,N_15229,N_15147);
xor U15631 (N_15631,N_15362,N_15139);
nand U15632 (N_15632,N_15012,N_15265);
nor U15633 (N_15633,N_15278,N_15272);
xor U15634 (N_15634,N_15356,N_15027);
nor U15635 (N_15635,N_15103,N_15431);
xor U15636 (N_15636,N_15492,N_15308);
nand U15637 (N_15637,N_15418,N_15025);
nand U15638 (N_15638,N_15130,N_15275);
xnor U15639 (N_15639,N_15132,N_15214);
and U15640 (N_15640,N_15417,N_15177);
xnor U15641 (N_15641,N_15292,N_15429);
nor U15642 (N_15642,N_15019,N_15100);
nor U15643 (N_15643,N_15201,N_15342);
or U15644 (N_15644,N_15046,N_15029);
xor U15645 (N_15645,N_15475,N_15363);
xor U15646 (N_15646,N_15140,N_15225);
or U15647 (N_15647,N_15458,N_15247);
nand U15648 (N_15648,N_15173,N_15442);
or U15649 (N_15649,N_15055,N_15203);
or U15650 (N_15650,N_15138,N_15061);
nor U15651 (N_15651,N_15092,N_15113);
nand U15652 (N_15652,N_15485,N_15481);
and U15653 (N_15653,N_15000,N_15060);
nor U15654 (N_15654,N_15080,N_15283);
and U15655 (N_15655,N_15398,N_15293);
nand U15656 (N_15656,N_15268,N_15249);
xnor U15657 (N_15657,N_15065,N_15281);
and U15658 (N_15658,N_15058,N_15334);
or U15659 (N_15659,N_15401,N_15238);
xnor U15660 (N_15660,N_15009,N_15318);
nand U15661 (N_15661,N_15037,N_15325);
or U15662 (N_15662,N_15158,N_15276);
or U15663 (N_15663,N_15154,N_15258);
nand U15664 (N_15664,N_15118,N_15310);
nor U15665 (N_15665,N_15410,N_15091);
or U15666 (N_15666,N_15496,N_15248);
nand U15667 (N_15667,N_15295,N_15096);
and U15668 (N_15668,N_15463,N_15339);
nor U15669 (N_15669,N_15355,N_15472);
nor U15670 (N_15670,N_15163,N_15175);
nand U15671 (N_15671,N_15049,N_15301);
or U15672 (N_15672,N_15235,N_15133);
xnor U15673 (N_15673,N_15213,N_15031);
or U15674 (N_15674,N_15144,N_15262);
and U15675 (N_15675,N_15336,N_15005);
or U15676 (N_15676,N_15030,N_15425);
nor U15677 (N_15677,N_15454,N_15388);
nor U15678 (N_15678,N_15462,N_15255);
and U15679 (N_15679,N_15284,N_15327);
or U15680 (N_15680,N_15150,N_15151);
or U15681 (N_15681,N_15209,N_15441);
nor U15682 (N_15682,N_15188,N_15319);
nand U15683 (N_15683,N_15016,N_15404);
nor U15684 (N_15684,N_15443,N_15015);
nand U15685 (N_15685,N_15324,N_15234);
nor U15686 (N_15686,N_15116,N_15155);
nand U15687 (N_15687,N_15141,N_15478);
xor U15688 (N_15688,N_15104,N_15115);
nand U15689 (N_15689,N_15237,N_15320);
or U15690 (N_15690,N_15406,N_15006);
nand U15691 (N_15691,N_15222,N_15122);
xor U15692 (N_15692,N_15328,N_15286);
nor U15693 (N_15693,N_15279,N_15039);
and U15694 (N_15694,N_15199,N_15168);
and U15695 (N_15695,N_15353,N_15023);
nand U15696 (N_15696,N_15385,N_15294);
and U15697 (N_15697,N_15488,N_15304);
nand U15698 (N_15698,N_15243,N_15347);
xor U15699 (N_15699,N_15067,N_15305);
nand U15700 (N_15700,N_15221,N_15171);
or U15701 (N_15701,N_15409,N_15372);
and U15702 (N_15702,N_15271,N_15051);
xor U15703 (N_15703,N_15010,N_15332);
nor U15704 (N_15704,N_15389,N_15180);
nand U15705 (N_15705,N_15438,N_15123);
or U15706 (N_15706,N_15280,N_15135);
nor U15707 (N_15707,N_15394,N_15231);
nand U15708 (N_15708,N_15244,N_15215);
nor U15709 (N_15709,N_15466,N_15287);
nand U15710 (N_15710,N_15373,N_15218);
and U15711 (N_15711,N_15426,N_15109);
or U15712 (N_15712,N_15076,N_15375);
and U15713 (N_15713,N_15266,N_15432);
or U15714 (N_15714,N_15230,N_15069);
nand U15715 (N_15715,N_15185,N_15183);
nand U15716 (N_15716,N_15082,N_15407);
xor U15717 (N_15717,N_15348,N_15197);
nand U15718 (N_15718,N_15128,N_15036);
or U15719 (N_15719,N_15350,N_15120);
or U15720 (N_15720,N_15159,N_15315);
nor U15721 (N_15721,N_15084,N_15134);
and U15722 (N_15722,N_15064,N_15498);
nand U15723 (N_15723,N_15075,N_15489);
and U15724 (N_15724,N_15358,N_15402);
nand U15725 (N_15725,N_15491,N_15313);
nand U15726 (N_15726,N_15490,N_15380);
and U15727 (N_15727,N_15153,N_15411);
nand U15728 (N_15728,N_15311,N_15233);
nand U15729 (N_15729,N_15297,N_15165);
nand U15730 (N_15730,N_15161,N_15365);
and U15731 (N_15731,N_15252,N_15098);
and U15732 (N_15732,N_15352,N_15448);
or U15733 (N_15733,N_15193,N_15079);
nor U15734 (N_15734,N_15479,N_15186);
or U15735 (N_15735,N_15349,N_15210);
nor U15736 (N_15736,N_15242,N_15053);
or U15737 (N_15737,N_15028,N_15192);
or U15738 (N_15738,N_15241,N_15335);
xnor U15739 (N_15739,N_15020,N_15035);
nand U15740 (N_15740,N_15106,N_15302);
or U15741 (N_15741,N_15345,N_15288);
and U15742 (N_15742,N_15461,N_15072);
nor U15743 (N_15743,N_15408,N_15126);
nand U15744 (N_15744,N_15125,N_15207);
xnor U15745 (N_15745,N_15390,N_15433);
and U15746 (N_15746,N_15189,N_15187);
nor U15747 (N_15747,N_15445,N_15196);
or U15748 (N_15748,N_15042,N_15085);
or U15749 (N_15749,N_15343,N_15191);
and U15750 (N_15750,N_15054,N_15236);
xnor U15751 (N_15751,N_15270,N_15112);
and U15752 (N_15752,N_15272,N_15119);
nand U15753 (N_15753,N_15332,N_15047);
nand U15754 (N_15754,N_15340,N_15371);
xor U15755 (N_15755,N_15314,N_15101);
or U15756 (N_15756,N_15303,N_15213);
or U15757 (N_15757,N_15391,N_15468);
or U15758 (N_15758,N_15414,N_15445);
nand U15759 (N_15759,N_15130,N_15367);
and U15760 (N_15760,N_15016,N_15434);
nor U15761 (N_15761,N_15331,N_15346);
nor U15762 (N_15762,N_15471,N_15325);
or U15763 (N_15763,N_15062,N_15302);
nand U15764 (N_15764,N_15148,N_15401);
nand U15765 (N_15765,N_15290,N_15468);
or U15766 (N_15766,N_15365,N_15293);
nor U15767 (N_15767,N_15289,N_15328);
and U15768 (N_15768,N_15468,N_15464);
nor U15769 (N_15769,N_15460,N_15031);
nand U15770 (N_15770,N_15094,N_15374);
or U15771 (N_15771,N_15344,N_15234);
and U15772 (N_15772,N_15116,N_15050);
nor U15773 (N_15773,N_15080,N_15268);
nor U15774 (N_15774,N_15461,N_15367);
and U15775 (N_15775,N_15264,N_15103);
or U15776 (N_15776,N_15484,N_15008);
and U15777 (N_15777,N_15456,N_15013);
xor U15778 (N_15778,N_15037,N_15108);
or U15779 (N_15779,N_15272,N_15143);
nand U15780 (N_15780,N_15041,N_15042);
nor U15781 (N_15781,N_15366,N_15136);
nand U15782 (N_15782,N_15383,N_15283);
nand U15783 (N_15783,N_15471,N_15070);
or U15784 (N_15784,N_15349,N_15327);
xor U15785 (N_15785,N_15202,N_15104);
nand U15786 (N_15786,N_15479,N_15177);
nand U15787 (N_15787,N_15167,N_15017);
nand U15788 (N_15788,N_15278,N_15320);
and U15789 (N_15789,N_15153,N_15341);
nand U15790 (N_15790,N_15453,N_15221);
nand U15791 (N_15791,N_15109,N_15206);
nor U15792 (N_15792,N_15077,N_15211);
and U15793 (N_15793,N_15288,N_15354);
and U15794 (N_15794,N_15311,N_15430);
and U15795 (N_15795,N_15123,N_15138);
xor U15796 (N_15796,N_15184,N_15029);
xnor U15797 (N_15797,N_15345,N_15023);
xnor U15798 (N_15798,N_15362,N_15203);
nand U15799 (N_15799,N_15016,N_15290);
xor U15800 (N_15800,N_15100,N_15464);
xnor U15801 (N_15801,N_15103,N_15311);
nand U15802 (N_15802,N_15034,N_15475);
and U15803 (N_15803,N_15144,N_15165);
nand U15804 (N_15804,N_15267,N_15005);
nand U15805 (N_15805,N_15387,N_15241);
xor U15806 (N_15806,N_15010,N_15080);
nand U15807 (N_15807,N_15150,N_15075);
and U15808 (N_15808,N_15126,N_15372);
or U15809 (N_15809,N_15085,N_15218);
nor U15810 (N_15810,N_15408,N_15248);
nand U15811 (N_15811,N_15004,N_15332);
xor U15812 (N_15812,N_15476,N_15068);
or U15813 (N_15813,N_15241,N_15008);
nor U15814 (N_15814,N_15025,N_15468);
or U15815 (N_15815,N_15295,N_15139);
nand U15816 (N_15816,N_15168,N_15094);
nand U15817 (N_15817,N_15447,N_15015);
nor U15818 (N_15818,N_15047,N_15029);
nand U15819 (N_15819,N_15407,N_15498);
xnor U15820 (N_15820,N_15286,N_15297);
nand U15821 (N_15821,N_15282,N_15397);
or U15822 (N_15822,N_15042,N_15324);
and U15823 (N_15823,N_15178,N_15494);
nand U15824 (N_15824,N_15368,N_15321);
nor U15825 (N_15825,N_15248,N_15349);
nor U15826 (N_15826,N_15115,N_15161);
and U15827 (N_15827,N_15076,N_15028);
nor U15828 (N_15828,N_15138,N_15093);
nand U15829 (N_15829,N_15458,N_15321);
and U15830 (N_15830,N_15350,N_15060);
or U15831 (N_15831,N_15047,N_15489);
and U15832 (N_15832,N_15307,N_15047);
nor U15833 (N_15833,N_15403,N_15096);
nand U15834 (N_15834,N_15074,N_15350);
xor U15835 (N_15835,N_15240,N_15225);
and U15836 (N_15836,N_15335,N_15161);
nand U15837 (N_15837,N_15065,N_15153);
nor U15838 (N_15838,N_15356,N_15017);
nor U15839 (N_15839,N_15169,N_15066);
nor U15840 (N_15840,N_15078,N_15005);
nor U15841 (N_15841,N_15436,N_15046);
and U15842 (N_15842,N_15389,N_15446);
or U15843 (N_15843,N_15397,N_15466);
or U15844 (N_15844,N_15260,N_15114);
and U15845 (N_15845,N_15323,N_15342);
and U15846 (N_15846,N_15424,N_15133);
or U15847 (N_15847,N_15017,N_15212);
nand U15848 (N_15848,N_15465,N_15270);
xor U15849 (N_15849,N_15238,N_15060);
and U15850 (N_15850,N_15374,N_15308);
or U15851 (N_15851,N_15255,N_15141);
and U15852 (N_15852,N_15431,N_15417);
xor U15853 (N_15853,N_15229,N_15242);
xnor U15854 (N_15854,N_15452,N_15309);
or U15855 (N_15855,N_15107,N_15419);
or U15856 (N_15856,N_15383,N_15419);
and U15857 (N_15857,N_15328,N_15445);
xnor U15858 (N_15858,N_15151,N_15274);
nor U15859 (N_15859,N_15321,N_15084);
nor U15860 (N_15860,N_15105,N_15309);
nand U15861 (N_15861,N_15402,N_15311);
nand U15862 (N_15862,N_15411,N_15198);
nand U15863 (N_15863,N_15315,N_15474);
or U15864 (N_15864,N_15086,N_15104);
or U15865 (N_15865,N_15155,N_15370);
and U15866 (N_15866,N_15372,N_15353);
or U15867 (N_15867,N_15348,N_15167);
nand U15868 (N_15868,N_15282,N_15362);
nand U15869 (N_15869,N_15096,N_15492);
nor U15870 (N_15870,N_15268,N_15315);
or U15871 (N_15871,N_15192,N_15108);
nand U15872 (N_15872,N_15039,N_15188);
nand U15873 (N_15873,N_15079,N_15452);
or U15874 (N_15874,N_15221,N_15050);
xnor U15875 (N_15875,N_15069,N_15036);
xor U15876 (N_15876,N_15120,N_15016);
nor U15877 (N_15877,N_15267,N_15259);
and U15878 (N_15878,N_15474,N_15047);
nor U15879 (N_15879,N_15490,N_15358);
and U15880 (N_15880,N_15458,N_15274);
nand U15881 (N_15881,N_15200,N_15355);
and U15882 (N_15882,N_15432,N_15041);
nand U15883 (N_15883,N_15437,N_15413);
nor U15884 (N_15884,N_15258,N_15128);
and U15885 (N_15885,N_15150,N_15360);
xnor U15886 (N_15886,N_15303,N_15461);
nand U15887 (N_15887,N_15121,N_15032);
xor U15888 (N_15888,N_15377,N_15075);
nor U15889 (N_15889,N_15293,N_15022);
and U15890 (N_15890,N_15129,N_15050);
and U15891 (N_15891,N_15392,N_15484);
or U15892 (N_15892,N_15281,N_15260);
and U15893 (N_15893,N_15237,N_15147);
nand U15894 (N_15894,N_15102,N_15055);
and U15895 (N_15895,N_15035,N_15297);
xor U15896 (N_15896,N_15383,N_15224);
and U15897 (N_15897,N_15019,N_15239);
nor U15898 (N_15898,N_15220,N_15318);
xnor U15899 (N_15899,N_15188,N_15339);
nand U15900 (N_15900,N_15465,N_15301);
or U15901 (N_15901,N_15415,N_15492);
xnor U15902 (N_15902,N_15197,N_15101);
or U15903 (N_15903,N_15103,N_15057);
and U15904 (N_15904,N_15165,N_15008);
nor U15905 (N_15905,N_15493,N_15229);
nand U15906 (N_15906,N_15197,N_15064);
nand U15907 (N_15907,N_15037,N_15210);
xnor U15908 (N_15908,N_15205,N_15110);
xor U15909 (N_15909,N_15459,N_15356);
or U15910 (N_15910,N_15235,N_15111);
or U15911 (N_15911,N_15088,N_15068);
xor U15912 (N_15912,N_15245,N_15017);
nand U15913 (N_15913,N_15053,N_15496);
nand U15914 (N_15914,N_15199,N_15420);
xnor U15915 (N_15915,N_15144,N_15423);
nor U15916 (N_15916,N_15030,N_15238);
xnor U15917 (N_15917,N_15445,N_15385);
xnor U15918 (N_15918,N_15146,N_15251);
or U15919 (N_15919,N_15220,N_15170);
nand U15920 (N_15920,N_15334,N_15128);
xnor U15921 (N_15921,N_15214,N_15215);
or U15922 (N_15922,N_15231,N_15430);
nor U15923 (N_15923,N_15114,N_15332);
and U15924 (N_15924,N_15160,N_15092);
nor U15925 (N_15925,N_15087,N_15193);
nand U15926 (N_15926,N_15193,N_15396);
and U15927 (N_15927,N_15245,N_15263);
xnor U15928 (N_15928,N_15162,N_15056);
or U15929 (N_15929,N_15299,N_15480);
nand U15930 (N_15930,N_15457,N_15024);
nor U15931 (N_15931,N_15485,N_15472);
and U15932 (N_15932,N_15033,N_15472);
nand U15933 (N_15933,N_15276,N_15378);
or U15934 (N_15934,N_15377,N_15219);
nor U15935 (N_15935,N_15348,N_15367);
or U15936 (N_15936,N_15212,N_15267);
nand U15937 (N_15937,N_15045,N_15364);
or U15938 (N_15938,N_15131,N_15360);
nor U15939 (N_15939,N_15184,N_15373);
or U15940 (N_15940,N_15486,N_15011);
nor U15941 (N_15941,N_15256,N_15011);
nor U15942 (N_15942,N_15399,N_15445);
xnor U15943 (N_15943,N_15481,N_15324);
nor U15944 (N_15944,N_15267,N_15450);
nor U15945 (N_15945,N_15153,N_15247);
and U15946 (N_15946,N_15386,N_15170);
and U15947 (N_15947,N_15176,N_15119);
nand U15948 (N_15948,N_15450,N_15375);
xnor U15949 (N_15949,N_15392,N_15190);
nor U15950 (N_15950,N_15339,N_15136);
nor U15951 (N_15951,N_15075,N_15282);
nor U15952 (N_15952,N_15255,N_15077);
and U15953 (N_15953,N_15304,N_15254);
nand U15954 (N_15954,N_15237,N_15229);
xor U15955 (N_15955,N_15105,N_15000);
xnor U15956 (N_15956,N_15058,N_15309);
or U15957 (N_15957,N_15485,N_15339);
nor U15958 (N_15958,N_15473,N_15297);
nor U15959 (N_15959,N_15266,N_15386);
nor U15960 (N_15960,N_15004,N_15271);
nand U15961 (N_15961,N_15429,N_15370);
nor U15962 (N_15962,N_15096,N_15304);
nor U15963 (N_15963,N_15051,N_15171);
xor U15964 (N_15964,N_15378,N_15069);
and U15965 (N_15965,N_15058,N_15359);
nor U15966 (N_15966,N_15165,N_15226);
nor U15967 (N_15967,N_15457,N_15235);
or U15968 (N_15968,N_15232,N_15252);
nand U15969 (N_15969,N_15334,N_15187);
nor U15970 (N_15970,N_15223,N_15314);
nand U15971 (N_15971,N_15282,N_15453);
xor U15972 (N_15972,N_15212,N_15255);
or U15973 (N_15973,N_15235,N_15237);
nor U15974 (N_15974,N_15272,N_15355);
nand U15975 (N_15975,N_15316,N_15033);
nand U15976 (N_15976,N_15357,N_15467);
nand U15977 (N_15977,N_15321,N_15455);
nor U15978 (N_15978,N_15217,N_15307);
nand U15979 (N_15979,N_15072,N_15121);
xnor U15980 (N_15980,N_15273,N_15412);
xor U15981 (N_15981,N_15029,N_15180);
and U15982 (N_15982,N_15483,N_15123);
xnor U15983 (N_15983,N_15492,N_15344);
nor U15984 (N_15984,N_15149,N_15112);
xor U15985 (N_15985,N_15081,N_15426);
nand U15986 (N_15986,N_15493,N_15093);
and U15987 (N_15987,N_15188,N_15086);
xor U15988 (N_15988,N_15261,N_15127);
and U15989 (N_15989,N_15273,N_15458);
nor U15990 (N_15990,N_15039,N_15124);
xnor U15991 (N_15991,N_15408,N_15002);
and U15992 (N_15992,N_15294,N_15447);
and U15993 (N_15993,N_15240,N_15360);
or U15994 (N_15994,N_15325,N_15287);
nor U15995 (N_15995,N_15244,N_15423);
xor U15996 (N_15996,N_15489,N_15049);
nand U15997 (N_15997,N_15392,N_15193);
nand U15998 (N_15998,N_15330,N_15442);
nand U15999 (N_15999,N_15395,N_15492);
and U16000 (N_16000,N_15833,N_15944);
nor U16001 (N_16001,N_15821,N_15684);
xor U16002 (N_16002,N_15705,N_15646);
nand U16003 (N_16003,N_15767,N_15527);
xnor U16004 (N_16004,N_15538,N_15945);
nor U16005 (N_16005,N_15597,N_15605);
and U16006 (N_16006,N_15976,N_15642);
nand U16007 (N_16007,N_15774,N_15588);
nand U16008 (N_16008,N_15972,N_15730);
xnor U16009 (N_16009,N_15969,N_15932);
or U16010 (N_16010,N_15926,N_15675);
xnor U16011 (N_16011,N_15952,N_15554);
or U16012 (N_16012,N_15671,N_15780);
and U16013 (N_16013,N_15814,N_15792);
xor U16014 (N_16014,N_15744,N_15974);
xnor U16015 (N_16015,N_15580,N_15513);
xnor U16016 (N_16016,N_15759,N_15865);
or U16017 (N_16017,N_15719,N_15817);
nand U16018 (N_16018,N_15530,N_15748);
and U16019 (N_16019,N_15989,N_15739);
nor U16020 (N_16020,N_15870,N_15914);
nor U16021 (N_16021,N_15656,N_15828);
nand U16022 (N_16022,N_15815,N_15502);
or U16023 (N_16023,N_15956,N_15900);
nand U16024 (N_16024,N_15555,N_15832);
xor U16025 (N_16025,N_15922,N_15604);
and U16026 (N_16026,N_15583,N_15633);
xor U16027 (N_16027,N_15856,N_15764);
and U16028 (N_16028,N_15677,N_15954);
xnor U16029 (N_16029,N_15716,N_15570);
nor U16030 (N_16030,N_15717,N_15875);
nor U16031 (N_16031,N_15881,N_15876);
and U16032 (N_16032,N_15806,N_15840);
and U16033 (N_16033,N_15779,N_15561);
and U16034 (N_16034,N_15718,N_15590);
nand U16035 (N_16035,N_15754,N_15579);
or U16036 (N_16036,N_15586,N_15853);
xnor U16037 (N_16037,N_15746,N_15635);
xnor U16038 (N_16038,N_15740,N_15596);
nor U16039 (N_16039,N_15645,N_15621);
nor U16040 (N_16040,N_15843,N_15686);
and U16041 (N_16041,N_15618,N_15712);
or U16042 (N_16042,N_15894,N_15564);
and U16043 (N_16043,N_15988,N_15623);
nor U16044 (N_16044,N_15528,N_15902);
xor U16045 (N_16045,N_15504,N_15690);
and U16046 (N_16046,N_15882,N_15884);
and U16047 (N_16047,N_15785,N_15743);
xor U16048 (N_16048,N_15795,N_15598);
and U16049 (N_16049,N_15631,N_15542);
xnor U16050 (N_16050,N_15593,N_15575);
and U16051 (N_16051,N_15903,N_15763);
or U16052 (N_16052,N_15729,N_15786);
nor U16053 (N_16053,N_15951,N_15638);
nor U16054 (N_16054,N_15626,N_15727);
xnor U16055 (N_16055,N_15994,N_15898);
xnor U16056 (N_16056,N_15658,N_15906);
or U16057 (N_16057,N_15724,N_15640);
or U16058 (N_16058,N_15868,N_15861);
xor U16059 (N_16059,N_15693,N_15560);
nor U16060 (N_16060,N_15711,N_15602);
nand U16061 (N_16061,N_15851,N_15966);
or U16062 (N_16062,N_15948,N_15526);
nand U16063 (N_16063,N_15973,N_15760);
and U16064 (N_16064,N_15960,N_15608);
xor U16065 (N_16065,N_15909,N_15939);
or U16066 (N_16066,N_15582,N_15837);
xor U16067 (N_16067,N_15933,N_15812);
nor U16068 (N_16068,N_15920,N_15563);
and U16069 (N_16069,N_15797,N_15857);
xnor U16070 (N_16070,N_15811,N_15664);
or U16071 (N_16071,N_15572,N_15747);
or U16072 (N_16072,N_15508,N_15609);
xnor U16073 (N_16073,N_15999,N_15663);
nor U16074 (N_16074,N_15681,N_15819);
nand U16075 (N_16075,N_15889,N_15521);
or U16076 (N_16076,N_15991,N_15592);
nor U16077 (N_16077,N_15942,N_15629);
nand U16078 (N_16078,N_15810,N_15659);
or U16079 (N_16079,N_15577,N_15987);
and U16080 (N_16080,N_15917,N_15761);
nor U16081 (N_16081,N_15784,N_15878);
nor U16082 (N_16082,N_15678,N_15835);
or U16083 (N_16083,N_15568,N_15616);
or U16084 (N_16084,N_15726,N_15807);
or U16085 (N_16085,N_15982,N_15808);
xnor U16086 (N_16086,N_15818,N_15888);
or U16087 (N_16087,N_15573,N_15802);
xnor U16088 (N_16088,N_15611,N_15632);
nand U16089 (N_16089,N_15648,N_15787);
nor U16090 (N_16090,N_15581,N_15736);
and U16091 (N_16091,N_15524,N_15995);
nor U16092 (N_16092,N_15970,N_15587);
or U16093 (N_16093,N_15644,N_15546);
xor U16094 (N_16094,N_15829,N_15692);
xor U16095 (N_16095,N_15978,N_15858);
or U16096 (N_16096,N_15866,N_15507);
and U16097 (N_16097,N_15556,N_15643);
xor U16098 (N_16098,N_15937,N_15517);
and U16099 (N_16099,N_15533,N_15585);
or U16100 (N_16100,N_15733,N_15963);
or U16101 (N_16101,N_15698,N_15790);
nand U16102 (N_16102,N_15836,N_15531);
nor U16103 (N_16103,N_15850,N_15691);
xor U16104 (N_16104,N_15919,N_15669);
and U16105 (N_16105,N_15599,N_15839);
nand U16106 (N_16106,N_15890,N_15725);
nor U16107 (N_16107,N_15694,N_15607);
nor U16108 (N_16108,N_15591,N_15750);
xor U16109 (N_16109,N_15891,N_15957);
nand U16110 (N_16110,N_15755,N_15905);
or U16111 (N_16111,N_15911,N_15673);
xnor U16112 (N_16112,N_15990,N_15799);
xnor U16113 (N_16113,N_15916,N_15789);
or U16114 (N_16114,N_15996,N_15578);
or U16115 (N_16115,N_15804,N_15619);
xor U16116 (N_16116,N_15877,N_15612);
or U16117 (N_16117,N_15674,N_15523);
and U16118 (N_16118,N_15895,N_15627);
or U16119 (N_16119,N_15864,N_15688);
and U16120 (N_16120,N_15834,N_15672);
or U16121 (N_16121,N_15859,N_15636);
nand U16122 (N_16122,N_15749,N_15732);
xor U16123 (N_16123,N_15964,N_15938);
and U16124 (N_16124,N_15738,N_15641);
or U16125 (N_16125,N_15845,N_15901);
or U16126 (N_16126,N_15953,N_15869);
nor U16127 (N_16127,N_15628,N_15863);
xnor U16128 (N_16128,N_15514,N_15552);
nand U16129 (N_16129,N_15852,N_15775);
or U16130 (N_16130,N_15997,N_15661);
and U16131 (N_16131,N_15981,N_15512);
nand U16132 (N_16132,N_15701,N_15772);
xnor U16133 (N_16133,N_15562,N_15867);
nor U16134 (N_16134,N_15910,N_15915);
and U16135 (N_16135,N_15522,N_15505);
nor U16136 (N_16136,N_15846,N_15699);
xor U16137 (N_16137,N_15715,N_15549);
or U16138 (N_16138,N_15501,N_15624);
nor U16139 (N_16139,N_15689,N_15924);
nand U16140 (N_16140,N_15687,N_15929);
xnor U16141 (N_16141,N_15768,N_15620);
nor U16142 (N_16142,N_15883,N_15637);
nand U16143 (N_16143,N_15566,N_15601);
and U16144 (N_16144,N_15551,N_15830);
xor U16145 (N_16145,N_15510,N_15913);
xnor U16146 (N_16146,N_15565,N_15820);
and U16147 (N_16147,N_15855,N_15907);
and U16148 (N_16148,N_15660,N_15662);
and U16149 (N_16149,N_15928,N_15930);
xnor U16150 (N_16150,N_15992,N_15742);
and U16151 (N_16151,N_15547,N_15935);
or U16152 (N_16152,N_15751,N_15516);
nor U16153 (N_16153,N_15921,N_15847);
xor U16154 (N_16154,N_15803,N_15961);
or U16155 (N_16155,N_15553,N_15844);
nor U16156 (N_16156,N_15842,N_15927);
or U16157 (N_16157,N_15872,N_15793);
xnor U16158 (N_16158,N_15816,N_15777);
nor U16159 (N_16159,N_15685,N_15762);
and U16160 (N_16160,N_15827,N_15946);
nor U16161 (N_16161,N_15943,N_15649);
xnor U16162 (N_16162,N_15657,N_15756);
or U16163 (N_16163,N_15918,N_15569);
nand U16164 (N_16164,N_15571,N_15770);
or U16165 (N_16165,N_15511,N_15600);
xor U16166 (N_16166,N_15652,N_15899);
nand U16167 (N_16167,N_15515,N_15520);
and U16168 (N_16168,N_15540,N_15539);
xor U16169 (N_16169,N_15809,N_15731);
and U16170 (N_16170,N_15791,N_15979);
or U16171 (N_16171,N_15603,N_15695);
or U16172 (N_16172,N_15838,N_15848);
nor U16173 (N_16173,N_15653,N_15558);
nand U16174 (N_16174,N_15529,N_15634);
or U16175 (N_16175,N_15950,N_15545);
xnor U16176 (N_16176,N_15841,N_15670);
nand U16177 (N_16177,N_15782,N_15766);
nand U16178 (N_16178,N_15977,N_15610);
or U16179 (N_16179,N_15798,N_15548);
and U16180 (N_16180,N_15765,N_15896);
and U16181 (N_16181,N_15860,N_15541);
nand U16182 (N_16182,N_15544,N_15783);
nor U16183 (N_16183,N_15959,N_15500);
or U16184 (N_16184,N_15885,N_15874);
and U16185 (N_16185,N_15525,N_15776);
and U16186 (N_16186,N_15745,N_15697);
and U16187 (N_16187,N_15655,N_15532);
and U16188 (N_16188,N_15639,N_15589);
and U16189 (N_16189,N_15503,N_15615);
nand U16190 (N_16190,N_15702,N_15788);
nand U16191 (N_16191,N_15947,N_15936);
and U16192 (N_16192,N_15617,N_15824);
nand U16193 (N_16193,N_15826,N_15622);
nor U16194 (N_16194,N_15993,N_15757);
nand U16195 (N_16195,N_15703,N_15506);
or U16196 (N_16196,N_15796,N_15752);
nor U16197 (N_16197,N_15949,N_15892);
xor U16198 (N_16198,N_15904,N_15614);
or U16199 (N_16199,N_15714,N_15737);
nor U16200 (N_16200,N_15594,N_15567);
nor U16201 (N_16201,N_15721,N_15535);
nor U16202 (N_16202,N_15706,N_15801);
xnor U16203 (N_16203,N_15720,N_15536);
nand U16204 (N_16204,N_15606,N_15965);
nor U16205 (N_16205,N_15537,N_15543);
or U16206 (N_16206,N_15975,N_15758);
nand U16207 (N_16207,N_15651,N_15519);
nand U16208 (N_16208,N_15931,N_15955);
and U16209 (N_16209,N_15668,N_15584);
nor U16210 (N_16210,N_15813,N_15576);
nor U16211 (N_16211,N_15985,N_15962);
nand U16212 (N_16212,N_15704,N_15849);
xnor U16213 (N_16213,N_15823,N_15958);
or U16214 (N_16214,N_15940,N_15822);
nand U16215 (N_16215,N_15613,N_15912);
and U16216 (N_16216,N_15700,N_15980);
nor U16217 (N_16217,N_15871,N_15696);
nand U16218 (N_16218,N_15778,N_15908);
nand U16219 (N_16219,N_15873,N_15534);
nand U16220 (N_16220,N_15923,N_15707);
xor U16221 (N_16221,N_15771,N_15934);
or U16222 (N_16222,N_15831,N_15879);
and U16223 (N_16223,N_15680,N_15887);
or U16224 (N_16224,N_15984,N_15509);
xor U16225 (N_16225,N_15773,N_15968);
and U16226 (N_16226,N_15557,N_15781);
nand U16227 (N_16227,N_15825,N_15666);
or U16228 (N_16228,N_15800,N_15971);
nor U16229 (N_16229,N_15998,N_15654);
nand U16230 (N_16230,N_15983,N_15880);
xor U16231 (N_16231,N_15794,N_15713);
and U16232 (N_16232,N_15886,N_15862);
and U16233 (N_16233,N_15518,N_15676);
and U16234 (N_16234,N_15574,N_15650);
or U16235 (N_16235,N_15559,N_15667);
or U16236 (N_16236,N_15682,N_15741);
nor U16237 (N_16237,N_15854,N_15679);
and U16238 (N_16238,N_15967,N_15665);
nor U16239 (N_16239,N_15897,N_15550);
xnor U16240 (N_16240,N_15708,N_15986);
and U16241 (N_16241,N_15709,N_15722);
or U16242 (N_16242,N_15734,N_15941);
nand U16243 (N_16243,N_15735,N_15710);
nor U16244 (N_16244,N_15753,N_15723);
nor U16245 (N_16245,N_15625,N_15630);
xnor U16246 (N_16246,N_15893,N_15805);
nor U16247 (N_16247,N_15728,N_15595);
xor U16248 (N_16248,N_15647,N_15769);
or U16249 (N_16249,N_15683,N_15925);
and U16250 (N_16250,N_15784,N_15855);
xor U16251 (N_16251,N_15547,N_15766);
nand U16252 (N_16252,N_15745,N_15663);
or U16253 (N_16253,N_15532,N_15672);
nand U16254 (N_16254,N_15814,N_15919);
xor U16255 (N_16255,N_15593,N_15854);
nor U16256 (N_16256,N_15707,N_15699);
and U16257 (N_16257,N_15967,N_15730);
xor U16258 (N_16258,N_15555,N_15858);
nand U16259 (N_16259,N_15608,N_15883);
nand U16260 (N_16260,N_15504,N_15658);
and U16261 (N_16261,N_15787,N_15778);
or U16262 (N_16262,N_15631,N_15831);
and U16263 (N_16263,N_15526,N_15586);
nor U16264 (N_16264,N_15966,N_15724);
nor U16265 (N_16265,N_15963,N_15578);
nor U16266 (N_16266,N_15539,N_15993);
and U16267 (N_16267,N_15676,N_15611);
xnor U16268 (N_16268,N_15997,N_15923);
xor U16269 (N_16269,N_15717,N_15863);
xor U16270 (N_16270,N_15748,N_15526);
nor U16271 (N_16271,N_15795,N_15700);
or U16272 (N_16272,N_15629,N_15948);
or U16273 (N_16273,N_15945,N_15701);
nor U16274 (N_16274,N_15735,N_15570);
and U16275 (N_16275,N_15979,N_15779);
and U16276 (N_16276,N_15684,N_15712);
nand U16277 (N_16277,N_15738,N_15797);
nor U16278 (N_16278,N_15703,N_15975);
xor U16279 (N_16279,N_15771,N_15785);
nor U16280 (N_16280,N_15523,N_15822);
and U16281 (N_16281,N_15750,N_15803);
or U16282 (N_16282,N_15610,N_15811);
nor U16283 (N_16283,N_15548,N_15911);
nor U16284 (N_16284,N_15998,N_15771);
or U16285 (N_16285,N_15510,N_15724);
nor U16286 (N_16286,N_15757,N_15658);
nand U16287 (N_16287,N_15646,N_15701);
xnor U16288 (N_16288,N_15956,N_15882);
and U16289 (N_16289,N_15630,N_15729);
or U16290 (N_16290,N_15999,N_15594);
or U16291 (N_16291,N_15665,N_15620);
nand U16292 (N_16292,N_15573,N_15842);
or U16293 (N_16293,N_15529,N_15652);
nand U16294 (N_16294,N_15692,N_15685);
and U16295 (N_16295,N_15830,N_15836);
xor U16296 (N_16296,N_15904,N_15977);
xor U16297 (N_16297,N_15792,N_15949);
or U16298 (N_16298,N_15762,N_15676);
nand U16299 (N_16299,N_15546,N_15778);
and U16300 (N_16300,N_15987,N_15983);
and U16301 (N_16301,N_15948,N_15936);
or U16302 (N_16302,N_15589,N_15852);
and U16303 (N_16303,N_15915,N_15567);
and U16304 (N_16304,N_15679,N_15678);
and U16305 (N_16305,N_15641,N_15940);
xor U16306 (N_16306,N_15592,N_15998);
or U16307 (N_16307,N_15798,N_15912);
and U16308 (N_16308,N_15939,N_15740);
xnor U16309 (N_16309,N_15659,N_15807);
nor U16310 (N_16310,N_15748,N_15939);
nand U16311 (N_16311,N_15908,N_15689);
nand U16312 (N_16312,N_15571,N_15643);
xnor U16313 (N_16313,N_15840,N_15887);
or U16314 (N_16314,N_15872,N_15885);
and U16315 (N_16315,N_15804,N_15668);
nand U16316 (N_16316,N_15774,N_15699);
nand U16317 (N_16317,N_15632,N_15889);
nor U16318 (N_16318,N_15897,N_15914);
or U16319 (N_16319,N_15627,N_15823);
xor U16320 (N_16320,N_15552,N_15638);
nand U16321 (N_16321,N_15600,N_15970);
and U16322 (N_16322,N_15946,N_15786);
nand U16323 (N_16323,N_15670,N_15678);
nand U16324 (N_16324,N_15553,N_15667);
or U16325 (N_16325,N_15818,N_15616);
nand U16326 (N_16326,N_15502,N_15576);
nor U16327 (N_16327,N_15980,N_15594);
xnor U16328 (N_16328,N_15681,N_15594);
xor U16329 (N_16329,N_15915,N_15969);
nor U16330 (N_16330,N_15662,N_15937);
or U16331 (N_16331,N_15503,N_15973);
or U16332 (N_16332,N_15993,N_15540);
nand U16333 (N_16333,N_15952,N_15532);
nor U16334 (N_16334,N_15517,N_15865);
nor U16335 (N_16335,N_15533,N_15589);
and U16336 (N_16336,N_15545,N_15607);
xor U16337 (N_16337,N_15565,N_15728);
xnor U16338 (N_16338,N_15852,N_15550);
nor U16339 (N_16339,N_15850,N_15504);
nor U16340 (N_16340,N_15606,N_15763);
nor U16341 (N_16341,N_15932,N_15596);
nand U16342 (N_16342,N_15985,N_15871);
and U16343 (N_16343,N_15784,N_15608);
nor U16344 (N_16344,N_15501,N_15867);
nor U16345 (N_16345,N_15664,N_15868);
or U16346 (N_16346,N_15544,N_15646);
and U16347 (N_16347,N_15563,N_15989);
xor U16348 (N_16348,N_15820,N_15787);
xor U16349 (N_16349,N_15785,N_15504);
nand U16350 (N_16350,N_15651,N_15994);
or U16351 (N_16351,N_15577,N_15854);
nor U16352 (N_16352,N_15570,N_15793);
and U16353 (N_16353,N_15547,N_15650);
xor U16354 (N_16354,N_15845,N_15518);
xor U16355 (N_16355,N_15713,N_15989);
nor U16356 (N_16356,N_15884,N_15906);
nand U16357 (N_16357,N_15833,N_15548);
or U16358 (N_16358,N_15544,N_15702);
or U16359 (N_16359,N_15743,N_15923);
nand U16360 (N_16360,N_15739,N_15855);
xor U16361 (N_16361,N_15941,N_15722);
nor U16362 (N_16362,N_15774,N_15614);
or U16363 (N_16363,N_15828,N_15781);
nand U16364 (N_16364,N_15559,N_15870);
nor U16365 (N_16365,N_15762,N_15787);
and U16366 (N_16366,N_15946,N_15854);
xor U16367 (N_16367,N_15537,N_15525);
or U16368 (N_16368,N_15728,N_15536);
or U16369 (N_16369,N_15623,N_15549);
nand U16370 (N_16370,N_15640,N_15829);
nor U16371 (N_16371,N_15948,N_15787);
nand U16372 (N_16372,N_15856,N_15713);
nor U16373 (N_16373,N_15880,N_15628);
nor U16374 (N_16374,N_15922,N_15816);
nand U16375 (N_16375,N_15793,N_15605);
and U16376 (N_16376,N_15788,N_15933);
xnor U16377 (N_16377,N_15735,N_15707);
xnor U16378 (N_16378,N_15718,N_15932);
xnor U16379 (N_16379,N_15802,N_15544);
nor U16380 (N_16380,N_15859,N_15516);
and U16381 (N_16381,N_15519,N_15631);
or U16382 (N_16382,N_15842,N_15740);
nor U16383 (N_16383,N_15866,N_15696);
and U16384 (N_16384,N_15693,N_15944);
nand U16385 (N_16385,N_15504,N_15800);
or U16386 (N_16386,N_15934,N_15780);
xnor U16387 (N_16387,N_15579,N_15900);
nand U16388 (N_16388,N_15701,N_15655);
nand U16389 (N_16389,N_15939,N_15989);
nor U16390 (N_16390,N_15657,N_15895);
nor U16391 (N_16391,N_15825,N_15646);
or U16392 (N_16392,N_15823,N_15755);
or U16393 (N_16393,N_15803,N_15576);
or U16394 (N_16394,N_15875,N_15932);
and U16395 (N_16395,N_15526,N_15528);
or U16396 (N_16396,N_15589,N_15814);
or U16397 (N_16397,N_15997,N_15864);
and U16398 (N_16398,N_15617,N_15860);
or U16399 (N_16399,N_15954,N_15977);
or U16400 (N_16400,N_15866,N_15682);
and U16401 (N_16401,N_15611,N_15997);
and U16402 (N_16402,N_15800,N_15821);
or U16403 (N_16403,N_15855,N_15989);
and U16404 (N_16404,N_15885,N_15521);
and U16405 (N_16405,N_15793,N_15850);
and U16406 (N_16406,N_15702,N_15615);
nor U16407 (N_16407,N_15963,N_15696);
xnor U16408 (N_16408,N_15577,N_15751);
or U16409 (N_16409,N_15513,N_15880);
xnor U16410 (N_16410,N_15562,N_15794);
and U16411 (N_16411,N_15840,N_15626);
nand U16412 (N_16412,N_15678,N_15910);
nand U16413 (N_16413,N_15561,N_15857);
xor U16414 (N_16414,N_15658,N_15532);
or U16415 (N_16415,N_15849,N_15678);
xor U16416 (N_16416,N_15697,N_15746);
nor U16417 (N_16417,N_15837,N_15983);
or U16418 (N_16418,N_15793,N_15784);
and U16419 (N_16419,N_15876,N_15935);
xnor U16420 (N_16420,N_15917,N_15800);
nand U16421 (N_16421,N_15746,N_15503);
or U16422 (N_16422,N_15512,N_15746);
or U16423 (N_16423,N_15845,N_15698);
xor U16424 (N_16424,N_15647,N_15842);
and U16425 (N_16425,N_15580,N_15584);
and U16426 (N_16426,N_15748,N_15830);
nor U16427 (N_16427,N_15859,N_15978);
or U16428 (N_16428,N_15540,N_15729);
and U16429 (N_16429,N_15616,N_15525);
and U16430 (N_16430,N_15865,N_15628);
and U16431 (N_16431,N_15854,N_15521);
and U16432 (N_16432,N_15733,N_15857);
or U16433 (N_16433,N_15796,N_15647);
nor U16434 (N_16434,N_15716,N_15953);
and U16435 (N_16435,N_15743,N_15841);
or U16436 (N_16436,N_15611,N_15980);
xnor U16437 (N_16437,N_15803,N_15797);
nor U16438 (N_16438,N_15981,N_15843);
and U16439 (N_16439,N_15623,N_15934);
and U16440 (N_16440,N_15536,N_15564);
xnor U16441 (N_16441,N_15751,N_15590);
nand U16442 (N_16442,N_15810,N_15548);
nor U16443 (N_16443,N_15806,N_15607);
and U16444 (N_16444,N_15552,N_15691);
xnor U16445 (N_16445,N_15614,N_15965);
and U16446 (N_16446,N_15723,N_15552);
and U16447 (N_16447,N_15692,N_15857);
and U16448 (N_16448,N_15947,N_15554);
or U16449 (N_16449,N_15732,N_15944);
nand U16450 (N_16450,N_15904,N_15599);
or U16451 (N_16451,N_15770,N_15851);
or U16452 (N_16452,N_15727,N_15573);
xor U16453 (N_16453,N_15827,N_15627);
xnor U16454 (N_16454,N_15525,N_15882);
or U16455 (N_16455,N_15729,N_15877);
nand U16456 (N_16456,N_15664,N_15869);
nor U16457 (N_16457,N_15895,N_15587);
nor U16458 (N_16458,N_15961,N_15566);
nor U16459 (N_16459,N_15512,N_15957);
or U16460 (N_16460,N_15571,N_15975);
and U16461 (N_16461,N_15878,N_15779);
or U16462 (N_16462,N_15909,N_15579);
or U16463 (N_16463,N_15566,N_15537);
and U16464 (N_16464,N_15548,N_15787);
and U16465 (N_16465,N_15939,N_15544);
or U16466 (N_16466,N_15973,N_15898);
or U16467 (N_16467,N_15646,N_15813);
and U16468 (N_16468,N_15869,N_15978);
xnor U16469 (N_16469,N_15953,N_15862);
xor U16470 (N_16470,N_15971,N_15797);
and U16471 (N_16471,N_15585,N_15551);
or U16472 (N_16472,N_15599,N_15743);
or U16473 (N_16473,N_15781,N_15733);
nor U16474 (N_16474,N_15518,N_15930);
and U16475 (N_16475,N_15629,N_15756);
nand U16476 (N_16476,N_15677,N_15894);
or U16477 (N_16477,N_15877,N_15835);
or U16478 (N_16478,N_15517,N_15537);
or U16479 (N_16479,N_15963,N_15743);
nor U16480 (N_16480,N_15692,N_15876);
xnor U16481 (N_16481,N_15766,N_15512);
and U16482 (N_16482,N_15973,N_15507);
nand U16483 (N_16483,N_15605,N_15884);
and U16484 (N_16484,N_15788,N_15668);
xor U16485 (N_16485,N_15955,N_15858);
or U16486 (N_16486,N_15756,N_15806);
xnor U16487 (N_16487,N_15751,N_15688);
and U16488 (N_16488,N_15574,N_15663);
nor U16489 (N_16489,N_15978,N_15707);
xnor U16490 (N_16490,N_15994,N_15988);
nand U16491 (N_16491,N_15777,N_15618);
or U16492 (N_16492,N_15906,N_15660);
or U16493 (N_16493,N_15804,N_15743);
nand U16494 (N_16494,N_15837,N_15779);
nand U16495 (N_16495,N_15600,N_15549);
and U16496 (N_16496,N_15689,N_15562);
nor U16497 (N_16497,N_15774,N_15778);
or U16498 (N_16498,N_15660,N_15877);
nor U16499 (N_16499,N_15719,N_15730);
and U16500 (N_16500,N_16205,N_16440);
and U16501 (N_16501,N_16178,N_16073);
or U16502 (N_16502,N_16299,N_16447);
nand U16503 (N_16503,N_16272,N_16431);
xnor U16504 (N_16504,N_16010,N_16059);
nand U16505 (N_16505,N_16462,N_16354);
or U16506 (N_16506,N_16048,N_16244);
or U16507 (N_16507,N_16441,N_16115);
and U16508 (N_16508,N_16335,N_16193);
nand U16509 (N_16509,N_16327,N_16082);
nand U16510 (N_16510,N_16255,N_16152);
xor U16511 (N_16511,N_16035,N_16287);
or U16512 (N_16512,N_16127,N_16045);
and U16513 (N_16513,N_16364,N_16175);
nand U16514 (N_16514,N_16375,N_16294);
nand U16515 (N_16515,N_16003,N_16459);
nand U16516 (N_16516,N_16376,N_16492);
nand U16517 (N_16517,N_16147,N_16305);
nand U16518 (N_16518,N_16382,N_16164);
xnor U16519 (N_16519,N_16187,N_16460);
and U16520 (N_16520,N_16151,N_16015);
nor U16521 (N_16521,N_16249,N_16261);
nor U16522 (N_16522,N_16209,N_16320);
and U16523 (N_16523,N_16143,N_16225);
nand U16524 (N_16524,N_16300,N_16068);
xnor U16525 (N_16525,N_16090,N_16475);
or U16526 (N_16526,N_16271,N_16367);
and U16527 (N_16527,N_16269,N_16153);
and U16528 (N_16528,N_16442,N_16438);
nor U16529 (N_16529,N_16464,N_16408);
nor U16530 (N_16530,N_16061,N_16423);
nor U16531 (N_16531,N_16257,N_16030);
and U16532 (N_16532,N_16302,N_16121);
and U16533 (N_16533,N_16312,N_16072);
xnor U16534 (N_16534,N_16331,N_16124);
and U16535 (N_16535,N_16432,N_16325);
or U16536 (N_16536,N_16465,N_16201);
or U16537 (N_16537,N_16337,N_16065);
nor U16538 (N_16538,N_16208,N_16400);
nor U16539 (N_16539,N_16322,N_16087);
nand U16540 (N_16540,N_16052,N_16393);
and U16541 (N_16541,N_16234,N_16498);
nor U16542 (N_16542,N_16185,N_16230);
nor U16543 (N_16543,N_16350,N_16424);
or U16544 (N_16544,N_16319,N_16406);
nand U16545 (N_16545,N_16425,N_16278);
nor U16546 (N_16546,N_16142,N_16493);
xnor U16547 (N_16547,N_16069,N_16222);
xor U16548 (N_16548,N_16101,N_16081);
xor U16549 (N_16549,N_16495,N_16414);
nor U16550 (N_16550,N_16398,N_16445);
and U16551 (N_16551,N_16231,N_16140);
xnor U16552 (N_16552,N_16169,N_16444);
nand U16553 (N_16553,N_16085,N_16245);
xnor U16554 (N_16554,N_16025,N_16119);
and U16555 (N_16555,N_16077,N_16292);
nor U16556 (N_16556,N_16372,N_16144);
xnor U16557 (N_16557,N_16088,N_16353);
nand U16558 (N_16558,N_16053,N_16387);
nand U16559 (N_16559,N_16499,N_16186);
or U16560 (N_16560,N_16226,N_16420);
and U16561 (N_16561,N_16135,N_16026);
nor U16562 (N_16562,N_16282,N_16395);
nor U16563 (N_16563,N_16397,N_16456);
nand U16564 (N_16564,N_16416,N_16166);
xnor U16565 (N_16565,N_16307,N_16428);
xor U16566 (N_16566,N_16288,N_16276);
xor U16567 (N_16567,N_16062,N_16358);
nand U16568 (N_16568,N_16289,N_16012);
or U16569 (N_16569,N_16404,N_16401);
nor U16570 (N_16570,N_16363,N_16032);
and U16571 (N_16571,N_16345,N_16277);
nand U16572 (N_16572,N_16008,N_16157);
nand U16573 (N_16573,N_16033,N_16324);
xor U16574 (N_16574,N_16366,N_16311);
and U16575 (N_16575,N_16283,N_16041);
nand U16576 (N_16576,N_16471,N_16227);
xnor U16577 (N_16577,N_16336,N_16391);
xnor U16578 (N_16578,N_16125,N_16197);
xnor U16579 (N_16579,N_16089,N_16238);
nor U16580 (N_16580,N_16494,N_16468);
or U16581 (N_16581,N_16159,N_16100);
nand U16582 (N_16582,N_16021,N_16128);
xor U16583 (N_16583,N_16383,N_16267);
and U16584 (N_16584,N_16285,N_16176);
xor U16585 (N_16585,N_16449,N_16196);
nand U16586 (N_16586,N_16242,N_16403);
xor U16587 (N_16587,N_16040,N_16343);
nand U16588 (N_16588,N_16338,N_16023);
nor U16589 (N_16589,N_16229,N_16361);
and U16590 (N_16590,N_16374,N_16083);
and U16591 (N_16591,N_16020,N_16031);
and U16592 (N_16592,N_16339,N_16241);
nand U16593 (N_16593,N_16123,N_16098);
and U16594 (N_16594,N_16239,N_16019);
nand U16595 (N_16595,N_16351,N_16480);
or U16596 (N_16596,N_16388,N_16407);
and U16597 (N_16597,N_16007,N_16000);
or U16598 (N_16598,N_16247,N_16349);
nand U16599 (N_16599,N_16473,N_16221);
xnor U16600 (N_16600,N_16111,N_16070);
and U16601 (N_16601,N_16352,N_16160);
nand U16602 (N_16602,N_16156,N_16155);
and U16603 (N_16603,N_16038,N_16108);
or U16604 (N_16604,N_16434,N_16315);
nand U16605 (N_16605,N_16126,N_16248);
nand U16606 (N_16606,N_16369,N_16092);
or U16607 (N_16607,N_16483,N_16443);
nand U16608 (N_16608,N_16355,N_16190);
xnor U16609 (N_16609,N_16146,N_16120);
or U16610 (N_16610,N_16304,N_16470);
or U16611 (N_16611,N_16419,N_16290);
xor U16612 (N_16612,N_16411,N_16392);
nand U16613 (N_16613,N_16162,N_16298);
and U16614 (N_16614,N_16017,N_16344);
nand U16615 (N_16615,N_16154,N_16265);
xnor U16616 (N_16616,N_16268,N_16028);
xor U16617 (N_16617,N_16340,N_16009);
or U16618 (N_16618,N_16105,N_16079);
nand U16619 (N_16619,N_16433,N_16198);
xor U16620 (N_16620,N_16472,N_16066);
nand U16621 (N_16621,N_16297,N_16212);
and U16622 (N_16622,N_16384,N_16368);
and U16623 (N_16623,N_16084,N_16006);
nor U16624 (N_16624,N_16183,N_16301);
nand U16625 (N_16625,N_16262,N_16145);
or U16626 (N_16626,N_16415,N_16273);
xor U16627 (N_16627,N_16005,N_16477);
nor U16628 (N_16628,N_16341,N_16426);
nor U16629 (N_16629,N_16260,N_16256);
nand U16630 (N_16630,N_16463,N_16488);
xnor U16631 (N_16631,N_16099,N_16455);
nor U16632 (N_16632,N_16056,N_16394);
and U16633 (N_16633,N_16218,N_16210);
nor U16634 (N_16634,N_16200,N_16043);
or U16635 (N_16635,N_16252,N_16094);
or U16636 (N_16636,N_16150,N_16024);
nand U16637 (N_16637,N_16001,N_16286);
xnor U16638 (N_16638,N_16075,N_16485);
and U16639 (N_16639,N_16203,N_16129);
nand U16640 (N_16640,N_16047,N_16138);
and U16641 (N_16641,N_16096,N_16170);
xnor U16642 (N_16642,N_16022,N_16211);
nor U16643 (N_16643,N_16109,N_16356);
nor U16644 (N_16644,N_16293,N_16148);
nor U16645 (N_16645,N_16114,N_16250);
or U16646 (N_16646,N_16274,N_16359);
nand U16647 (N_16647,N_16107,N_16491);
or U16648 (N_16648,N_16004,N_16131);
nand U16649 (N_16649,N_16189,N_16371);
nor U16650 (N_16650,N_16132,N_16313);
nand U16651 (N_16651,N_16191,N_16281);
or U16652 (N_16652,N_16163,N_16466);
or U16653 (N_16653,N_16046,N_16042);
or U16654 (N_16654,N_16417,N_16049);
xor U16655 (N_16655,N_16064,N_16430);
xnor U16656 (N_16656,N_16452,N_16013);
or U16657 (N_16657,N_16333,N_16215);
nand U16658 (N_16658,N_16116,N_16214);
or U16659 (N_16659,N_16165,N_16410);
and U16660 (N_16660,N_16018,N_16217);
and U16661 (N_16661,N_16037,N_16027);
xor U16662 (N_16662,N_16034,N_16332);
and U16663 (N_16663,N_16095,N_16450);
and U16664 (N_16664,N_16490,N_16122);
or U16665 (N_16665,N_16323,N_16439);
xnor U16666 (N_16666,N_16029,N_16204);
and U16667 (N_16667,N_16451,N_16213);
and U16668 (N_16668,N_16264,N_16318);
xnor U16669 (N_16669,N_16233,N_16243);
nor U16670 (N_16670,N_16103,N_16251);
xnor U16671 (N_16671,N_16291,N_16326);
xnor U16672 (N_16672,N_16448,N_16457);
and U16673 (N_16673,N_16334,N_16117);
nand U16674 (N_16674,N_16453,N_16235);
xor U16675 (N_16675,N_16346,N_16469);
nand U16676 (N_16676,N_16259,N_16435);
and U16677 (N_16677,N_16220,N_16192);
or U16678 (N_16678,N_16014,N_16295);
xnor U16679 (N_16679,N_16474,N_16489);
xor U16680 (N_16680,N_16482,N_16275);
nor U16681 (N_16681,N_16476,N_16362);
nor U16682 (N_16682,N_16418,N_16380);
xor U16683 (N_16683,N_16232,N_16130);
and U16684 (N_16684,N_16303,N_16481);
nand U16685 (N_16685,N_16429,N_16314);
nand U16686 (N_16686,N_16427,N_16389);
nand U16687 (N_16687,N_16102,N_16078);
or U16688 (N_16688,N_16342,N_16051);
xnor U16689 (N_16689,N_16060,N_16044);
xnor U16690 (N_16690,N_16076,N_16202);
nand U16691 (N_16691,N_16199,N_16219);
and U16692 (N_16692,N_16036,N_16136);
nand U16693 (N_16693,N_16478,N_16421);
nand U16694 (N_16694,N_16437,N_16195);
or U16695 (N_16695,N_16174,N_16496);
nand U16696 (N_16696,N_16284,N_16236);
and U16697 (N_16697,N_16321,N_16308);
and U16698 (N_16698,N_16497,N_16039);
xnor U16699 (N_16699,N_16172,N_16263);
nor U16700 (N_16700,N_16378,N_16412);
nand U16701 (N_16701,N_16309,N_16379);
nor U16702 (N_16702,N_16158,N_16347);
and U16703 (N_16703,N_16373,N_16370);
nand U16704 (N_16704,N_16106,N_16055);
or U16705 (N_16705,N_16484,N_16011);
and U16706 (N_16706,N_16184,N_16137);
or U16707 (N_16707,N_16306,N_16134);
xor U16708 (N_16708,N_16173,N_16310);
nor U16709 (N_16709,N_16330,N_16167);
and U16710 (N_16710,N_16206,N_16016);
nand U16711 (N_16711,N_16074,N_16458);
nor U16712 (N_16712,N_16405,N_16002);
or U16713 (N_16713,N_16086,N_16317);
nor U16714 (N_16714,N_16118,N_16254);
and U16715 (N_16715,N_16058,N_16253);
nand U16716 (N_16716,N_16228,N_16181);
nor U16717 (N_16717,N_16357,N_16180);
nor U16718 (N_16718,N_16385,N_16402);
and U16719 (N_16719,N_16246,N_16329);
or U16720 (N_16720,N_16133,N_16179);
nor U16721 (N_16721,N_16194,N_16461);
nand U16722 (N_16722,N_16091,N_16381);
or U16723 (N_16723,N_16396,N_16360);
or U16724 (N_16724,N_16258,N_16177);
xor U16725 (N_16725,N_16054,N_16348);
xor U16726 (N_16726,N_16139,N_16168);
xnor U16727 (N_16727,N_16270,N_16207);
nand U16728 (N_16728,N_16182,N_16454);
and U16729 (N_16729,N_16390,N_16266);
nand U16730 (N_16730,N_16328,N_16188);
or U16731 (N_16731,N_16071,N_16436);
and U16732 (N_16732,N_16467,N_16067);
nor U16733 (N_16733,N_16141,N_16093);
or U16734 (N_16734,N_16413,N_16104);
nand U16735 (N_16735,N_16171,N_16479);
xor U16736 (N_16736,N_16237,N_16097);
or U16737 (N_16737,N_16446,N_16422);
nand U16738 (N_16738,N_16112,N_16063);
and U16739 (N_16739,N_16296,N_16223);
nor U16740 (N_16740,N_16224,N_16161);
xnor U16741 (N_16741,N_16080,N_16377);
xor U16742 (N_16742,N_16486,N_16280);
xor U16743 (N_16743,N_16399,N_16386);
nand U16744 (N_16744,N_16365,N_16050);
nand U16745 (N_16745,N_16149,N_16316);
or U16746 (N_16746,N_16409,N_16279);
or U16747 (N_16747,N_16240,N_16110);
and U16748 (N_16748,N_16216,N_16113);
xor U16749 (N_16749,N_16487,N_16057);
nand U16750 (N_16750,N_16181,N_16436);
nor U16751 (N_16751,N_16306,N_16372);
xor U16752 (N_16752,N_16312,N_16005);
nor U16753 (N_16753,N_16495,N_16147);
or U16754 (N_16754,N_16440,N_16413);
nor U16755 (N_16755,N_16212,N_16371);
and U16756 (N_16756,N_16467,N_16116);
nor U16757 (N_16757,N_16333,N_16377);
xor U16758 (N_16758,N_16231,N_16092);
or U16759 (N_16759,N_16451,N_16445);
nand U16760 (N_16760,N_16295,N_16090);
xnor U16761 (N_16761,N_16407,N_16125);
nor U16762 (N_16762,N_16202,N_16302);
nand U16763 (N_16763,N_16235,N_16103);
nor U16764 (N_16764,N_16249,N_16378);
nor U16765 (N_16765,N_16259,N_16241);
and U16766 (N_16766,N_16256,N_16125);
xnor U16767 (N_16767,N_16438,N_16121);
or U16768 (N_16768,N_16310,N_16153);
and U16769 (N_16769,N_16119,N_16291);
nand U16770 (N_16770,N_16408,N_16434);
xor U16771 (N_16771,N_16160,N_16137);
nand U16772 (N_16772,N_16049,N_16235);
nor U16773 (N_16773,N_16162,N_16239);
and U16774 (N_16774,N_16340,N_16238);
or U16775 (N_16775,N_16049,N_16357);
and U16776 (N_16776,N_16421,N_16180);
or U16777 (N_16777,N_16313,N_16459);
nand U16778 (N_16778,N_16393,N_16215);
or U16779 (N_16779,N_16357,N_16255);
nor U16780 (N_16780,N_16046,N_16381);
or U16781 (N_16781,N_16250,N_16362);
and U16782 (N_16782,N_16497,N_16259);
nand U16783 (N_16783,N_16227,N_16194);
nor U16784 (N_16784,N_16477,N_16474);
nor U16785 (N_16785,N_16146,N_16494);
or U16786 (N_16786,N_16476,N_16240);
nand U16787 (N_16787,N_16134,N_16457);
and U16788 (N_16788,N_16199,N_16245);
and U16789 (N_16789,N_16019,N_16459);
xor U16790 (N_16790,N_16372,N_16106);
and U16791 (N_16791,N_16288,N_16370);
nor U16792 (N_16792,N_16410,N_16444);
or U16793 (N_16793,N_16416,N_16443);
xnor U16794 (N_16794,N_16011,N_16290);
or U16795 (N_16795,N_16410,N_16384);
nand U16796 (N_16796,N_16212,N_16258);
nor U16797 (N_16797,N_16102,N_16125);
xor U16798 (N_16798,N_16357,N_16187);
or U16799 (N_16799,N_16239,N_16128);
nand U16800 (N_16800,N_16231,N_16113);
xor U16801 (N_16801,N_16421,N_16034);
nor U16802 (N_16802,N_16133,N_16025);
nand U16803 (N_16803,N_16290,N_16116);
and U16804 (N_16804,N_16318,N_16224);
and U16805 (N_16805,N_16108,N_16403);
nand U16806 (N_16806,N_16240,N_16222);
and U16807 (N_16807,N_16405,N_16256);
or U16808 (N_16808,N_16373,N_16456);
xor U16809 (N_16809,N_16294,N_16150);
nor U16810 (N_16810,N_16038,N_16046);
nand U16811 (N_16811,N_16094,N_16247);
or U16812 (N_16812,N_16090,N_16411);
and U16813 (N_16813,N_16179,N_16409);
xnor U16814 (N_16814,N_16375,N_16139);
and U16815 (N_16815,N_16187,N_16168);
nor U16816 (N_16816,N_16215,N_16459);
nor U16817 (N_16817,N_16098,N_16358);
xor U16818 (N_16818,N_16398,N_16081);
or U16819 (N_16819,N_16458,N_16255);
and U16820 (N_16820,N_16335,N_16436);
nand U16821 (N_16821,N_16363,N_16325);
xnor U16822 (N_16822,N_16049,N_16023);
and U16823 (N_16823,N_16364,N_16334);
xnor U16824 (N_16824,N_16075,N_16397);
nor U16825 (N_16825,N_16375,N_16402);
nand U16826 (N_16826,N_16027,N_16051);
or U16827 (N_16827,N_16310,N_16160);
xnor U16828 (N_16828,N_16188,N_16468);
or U16829 (N_16829,N_16449,N_16068);
nand U16830 (N_16830,N_16472,N_16114);
or U16831 (N_16831,N_16087,N_16488);
xnor U16832 (N_16832,N_16277,N_16211);
xor U16833 (N_16833,N_16433,N_16415);
and U16834 (N_16834,N_16099,N_16283);
or U16835 (N_16835,N_16455,N_16435);
xnor U16836 (N_16836,N_16060,N_16495);
xnor U16837 (N_16837,N_16165,N_16376);
nor U16838 (N_16838,N_16432,N_16173);
nand U16839 (N_16839,N_16238,N_16431);
and U16840 (N_16840,N_16078,N_16408);
or U16841 (N_16841,N_16359,N_16455);
or U16842 (N_16842,N_16045,N_16244);
xor U16843 (N_16843,N_16025,N_16094);
nor U16844 (N_16844,N_16247,N_16006);
nand U16845 (N_16845,N_16479,N_16226);
nor U16846 (N_16846,N_16310,N_16252);
and U16847 (N_16847,N_16145,N_16389);
or U16848 (N_16848,N_16025,N_16248);
nand U16849 (N_16849,N_16453,N_16310);
nor U16850 (N_16850,N_16352,N_16487);
nand U16851 (N_16851,N_16016,N_16196);
nand U16852 (N_16852,N_16464,N_16017);
and U16853 (N_16853,N_16358,N_16353);
or U16854 (N_16854,N_16035,N_16433);
and U16855 (N_16855,N_16398,N_16233);
nand U16856 (N_16856,N_16096,N_16123);
nand U16857 (N_16857,N_16086,N_16456);
or U16858 (N_16858,N_16152,N_16184);
and U16859 (N_16859,N_16195,N_16052);
or U16860 (N_16860,N_16163,N_16006);
or U16861 (N_16861,N_16432,N_16060);
nor U16862 (N_16862,N_16273,N_16055);
or U16863 (N_16863,N_16175,N_16014);
and U16864 (N_16864,N_16002,N_16279);
or U16865 (N_16865,N_16005,N_16037);
and U16866 (N_16866,N_16078,N_16375);
or U16867 (N_16867,N_16152,N_16032);
nand U16868 (N_16868,N_16389,N_16445);
nand U16869 (N_16869,N_16146,N_16045);
or U16870 (N_16870,N_16031,N_16444);
or U16871 (N_16871,N_16216,N_16015);
xnor U16872 (N_16872,N_16135,N_16043);
nand U16873 (N_16873,N_16496,N_16077);
and U16874 (N_16874,N_16042,N_16144);
nor U16875 (N_16875,N_16053,N_16229);
nor U16876 (N_16876,N_16098,N_16254);
nand U16877 (N_16877,N_16123,N_16298);
nor U16878 (N_16878,N_16462,N_16294);
and U16879 (N_16879,N_16498,N_16280);
or U16880 (N_16880,N_16094,N_16113);
or U16881 (N_16881,N_16394,N_16203);
or U16882 (N_16882,N_16482,N_16047);
and U16883 (N_16883,N_16082,N_16218);
nor U16884 (N_16884,N_16147,N_16030);
xnor U16885 (N_16885,N_16183,N_16171);
nand U16886 (N_16886,N_16308,N_16414);
or U16887 (N_16887,N_16246,N_16380);
xor U16888 (N_16888,N_16056,N_16223);
nor U16889 (N_16889,N_16083,N_16396);
xor U16890 (N_16890,N_16279,N_16376);
nor U16891 (N_16891,N_16155,N_16474);
and U16892 (N_16892,N_16462,N_16211);
and U16893 (N_16893,N_16023,N_16446);
nor U16894 (N_16894,N_16406,N_16093);
nand U16895 (N_16895,N_16293,N_16225);
xnor U16896 (N_16896,N_16437,N_16048);
nor U16897 (N_16897,N_16332,N_16235);
nor U16898 (N_16898,N_16208,N_16369);
nor U16899 (N_16899,N_16444,N_16285);
and U16900 (N_16900,N_16374,N_16159);
xnor U16901 (N_16901,N_16091,N_16350);
and U16902 (N_16902,N_16479,N_16112);
and U16903 (N_16903,N_16498,N_16053);
or U16904 (N_16904,N_16468,N_16112);
nand U16905 (N_16905,N_16285,N_16073);
and U16906 (N_16906,N_16296,N_16036);
nor U16907 (N_16907,N_16266,N_16056);
nor U16908 (N_16908,N_16058,N_16459);
xnor U16909 (N_16909,N_16132,N_16499);
nand U16910 (N_16910,N_16078,N_16452);
nand U16911 (N_16911,N_16032,N_16165);
and U16912 (N_16912,N_16018,N_16384);
or U16913 (N_16913,N_16092,N_16488);
xnor U16914 (N_16914,N_16236,N_16430);
nand U16915 (N_16915,N_16412,N_16397);
or U16916 (N_16916,N_16406,N_16463);
xor U16917 (N_16917,N_16355,N_16345);
or U16918 (N_16918,N_16294,N_16432);
nand U16919 (N_16919,N_16140,N_16321);
and U16920 (N_16920,N_16014,N_16120);
nor U16921 (N_16921,N_16346,N_16371);
and U16922 (N_16922,N_16108,N_16288);
nor U16923 (N_16923,N_16277,N_16386);
nand U16924 (N_16924,N_16254,N_16161);
and U16925 (N_16925,N_16380,N_16252);
or U16926 (N_16926,N_16158,N_16180);
nor U16927 (N_16927,N_16484,N_16022);
nand U16928 (N_16928,N_16469,N_16331);
xnor U16929 (N_16929,N_16068,N_16253);
xnor U16930 (N_16930,N_16301,N_16460);
or U16931 (N_16931,N_16173,N_16269);
xnor U16932 (N_16932,N_16355,N_16149);
nand U16933 (N_16933,N_16456,N_16327);
and U16934 (N_16934,N_16174,N_16061);
and U16935 (N_16935,N_16109,N_16097);
nand U16936 (N_16936,N_16210,N_16097);
and U16937 (N_16937,N_16393,N_16367);
nor U16938 (N_16938,N_16144,N_16202);
nor U16939 (N_16939,N_16089,N_16301);
nor U16940 (N_16940,N_16243,N_16224);
nor U16941 (N_16941,N_16171,N_16008);
xor U16942 (N_16942,N_16297,N_16097);
xnor U16943 (N_16943,N_16327,N_16438);
nor U16944 (N_16944,N_16454,N_16370);
or U16945 (N_16945,N_16241,N_16018);
xnor U16946 (N_16946,N_16011,N_16470);
and U16947 (N_16947,N_16187,N_16294);
and U16948 (N_16948,N_16138,N_16171);
xnor U16949 (N_16949,N_16392,N_16079);
and U16950 (N_16950,N_16348,N_16017);
xnor U16951 (N_16951,N_16398,N_16469);
nand U16952 (N_16952,N_16490,N_16211);
nand U16953 (N_16953,N_16014,N_16376);
nand U16954 (N_16954,N_16231,N_16340);
xnor U16955 (N_16955,N_16463,N_16069);
and U16956 (N_16956,N_16085,N_16233);
or U16957 (N_16957,N_16498,N_16397);
nor U16958 (N_16958,N_16255,N_16481);
and U16959 (N_16959,N_16207,N_16223);
or U16960 (N_16960,N_16214,N_16451);
nand U16961 (N_16961,N_16171,N_16021);
nor U16962 (N_16962,N_16436,N_16209);
or U16963 (N_16963,N_16032,N_16017);
or U16964 (N_16964,N_16423,N_16480);
or U16965 (N_16965,N_16174,N_16449);
or U16966 (N_16966,N_16091,N_16171);
xor U16967 (N_16967,N_16037,N_16225);
nor U16968 (N_16968,N_16196,N_16375);
nand U16969 (N_16969,N_16334,N_16062);
xnor U16970 (N_16970,N_16409,N_16050);
nand U16971 (N_16971,N_16008,N_16046);
and U16972 (N_16972,N_16460,N_16282);
or U16973 (N_16973,N_16413,N_16155);
xor U16974 (N_16974,N_16345,N_16270);
nor U16975 (N_16975,N_16281,N_16393);
or U16976 (N_16976,N_16093,N_16106);
nor U16977 (N_16977,N_16453,N_16116);
or U16978 (N_16978,N_16170,N_16432);
nor U16979 (N_16979,N_16208,N_16374);
nor U16980 (N_16980,N_16466,N_16496);
and U16981 (N_16981,N_16179,N_16369);
xnor U16982 (N_16982,N_16195,N_16090);
nor U16983 (N_16983,N_16450,N_16005);
nor U16984 (N_16984,N_16352,N_16099);
nand U16985 (N_16985,N_16147,N_16362);
nor U16986 (N_16986,N_16428,N_16017);
nor U16987 (N_16987,N_16161,N_16368);
xor U16988 (N_16988,N_16288,N_16147);
or U16989 (N_16989,N_16101,N_16274);
or U16990 (N_16990,N_16413,N_16062);
or U16991 (N_16991,N_16465,N_16119);
or U16992 (N_16992,N_16049,N_16153);
and U16993 (N_16993,N_16063,N_16231);
or U16994 (N_16994,N_16353,N_16032);
nor U16995 (N_16995,N_16066,N_16261);
nor U16996 (N_16996,N_16306,N_16102);
and U16997 (N_16997,N_16032,N_16064);
xor U16998 (N_16998,N_16191,N_16363);
xnor U16999 (N_16999,N_16301,N_16373);
or U17000 (N_17000,N_16727,N_16969);
nand U17001 (N_17001,N_16803,N_16936);
nand U17002 (N_17002,N_16733,N_16909);
xor U17003 (N_17003,N_16543,N_16514);
xnor U17004 (N_17004,N_16724,N_16694);
xnor U17005 (N_17005,N_16524,N_16855);
nor U17006 (N_17006,N_16538,N_16691);
or U17007 (N_17007,N_16789,N_16632);
xnor U17008 (N_17008,N_16534,N_16555);
or U17009 (N_17009,N_16625,N_16525);
xor U17010 (N_17010,N_16857,N_16847);
nand U17011 (N_17011,N_16908,N_16834);
nor U17012 (N_17012,N_16946,N_16942);
or U17013 (N_17013,N_16790,N_16948);
nor U17014 (N_17014,N_16673,N_16622);
nor U17015 (N_17015,N_16949,N_16983);
nor U17016 (N_17016,N_16672,N_16626);
xnor U17017 (N_17017,N_16843,N_16648);
and U17018 (N_17018,N_16647,N_16777);
nand U17019 (N_17019,N_16878,N_16655);
and U17020 (N_17020,N_16831,N_16561);
xor U17021 (N_17021,N_16886,N_16980);
nor U17022 (N_17022,N_16928,N_16917);
or U17023 (N_17023,N_16558,N_16897);
or U17024 (N_17024,N_16863,N_16771);
or U17025 (N_17025,N_16877,N_16984);
nor U17026 (N_17026,N_16978,N_16574);
or U17027 (N_17027,N_16992,N_16546);
or U17028 (N_17028,N_16669,N_16660);
or U17029 (N_17029,N_16624,N_16504);
nor U17030 (N_17030,N_16628,N_16519);
xnor U17031 (N_17031,N_16792,N_16810);
xnor U17032 (N_17032,N_16697,N_16554);
nor U17033 (N_17033,N_16541,N_16545);
and U17034 (N_17034,N_16720,N_16702);
xnor U17035 (N_17035,N_16904,N_16664);
and U17036 (N_17036,N_16607,N_16767);
nor U17037 (N_17037,N_16522,N_16850);
nor U17038 (N_17038,N_16744,N_16993);
xor U17039 (N_17039,N_16586,N_16570);
nand U17040 (N_17040,N_16851,N_16910);
xor U17041 (N_17041,N_16921,N_16703);
or U17042 (N_17042,N_16700,N_16927);
and U17043 (N_17043,N_16696,N_16950);
nor U17044 (N_17044,N_16520,N_16838);
nor U17045 (N_17045,N_16802,N_16595);
nor U17046 (N_17046,N_16516,N_16846);
nor U17047 (N_17047,N_16941,N_16723);
nand U17048 (N_17048,N_16788,N_16666);
xor U17049 (N_17049,N_16571,N_16807);
nor U17050 (N_17050,N_16704,N_16606);
nor U17051 (N_17051,N_16630,N_16532);
nor U17052 (N_17052,N_16508,N_16935);
xor U17053 (N_17053,N_16797,N_16615);
or U17054 (N_17054,N_16619,N_16536);
or U17055 (N_17055,N_16825,N_16583);
nand U17056 (N_17056,N_16675,N_16912);
or U17057 (N_17057,N_16743,N_16649);
or U17058 (N_17058,N_16753,N_16565);
or U17059 (N_17059,N_16568,N_16506);
nand U17060 (N_17060,N_16816,N_16715);
and U17061 (N_17061,N_16533,N_16730);
and U17062 (N_17062,N_16799,N_16903);
nor U17063 (N_17063,N_16572,N_16501);
nand U17064 (N_17064,N_16828,N_16783);
nor U17065 (N_17065,N_16631,N_16888);
nand U17066 (N_17066,N_16830,N_16526);
xnor U17067 (N_17067,N_16662,N_16502);
and U17068 (N_17068,N_16968,N_16894);
and U17069 (N_17069,N_16965,N_16820);
nor U17070 (N_17070,N_16684,N_16940);
nor U17071 (N_17071,N_16865,N_16605);
or U17072 (N_17072,N_16922,N_16937);
nand U17073 (N_17073,N_16891,N_16915);
nand U17074 (N_17074,N_16805,N_16852);
nor U17075 (N_17075,N_16542,N_16885);
nand U17076 (N_17076,N_16592,N_16701);
nand U17077 (N_17077,N_16889,N_16837);
or U17078 (N_17078,N_16769,N_16550);
xor U17079 (N_17079,N_16804,N_16994);
and U17080 (N_17080,N_16713,N_16573);
or U17081 (N_17081,N_16944,N_16613);
xnor U17082 (N_17082,N_16657,N_16785);
nand U17083 (N_17083,N_16609,N_16587);
nor U17084 (N_17084,N_16787,N_16761);
nor U17085 (N_17085,N_16966,N_16644);
nor U17086 (N_17086,N_16832,N_16902);
or U17087 (N_17087,N_16557,N_16989);
or U17088 (N_17088,N_16779,N_16801);
xor U17089 (N_17089,N_16869,N_16862);
xor U17090 (N_17090,N_16784,N_16896);
nor U17091 (N_17091,N_16641,N_16589);
or U17092 (N_17092,N_16836,N_16822);
and U17093 (N_17093,N_16640,N_16719);
nand U17094 (N_17094,N_16745,N_16637);
and U17095 (N_17095,N_16798,N_16566);
and U17096 (N_17096,N_16859,N_16699);
nand U17097 (N_17097,N_16659,N_16521);
xor U17098 (N_17098,N_16668,N_16650);
and U17099 (N_17099,N_16695,N_16796);
nor U17100 (N_17100,N_16551,N_16868);
xor U17101 (N_17101,N_16653,N_16602);
and U17102 (N_17102,N_16617,N_16663);
xor U17103 (N_17103,N_16887,N_16782);
nand U17104 (N_17104,N_16812,N_16982);
nand U17105 (N_17105,N_16867,N_16890);
and U17106 (N_17106,N_16527,N_16560);
or U17107 (N_17107,N_16575,N_16898);
nand U17108 (N_17108,N_16594,N_16945);
xnor U17109 (N_17109,N_16848,N_16698);
or U17110 (N_17110,N_16665,N_16651);
xor U17111 (N_17111,N_16577,N_16518);
nor U17112 (N_17112,N_16755,N_16814);
xnor U17113 (N_17113,N_16567,N_16770);
nor U17114 (N_17114,N_16997,N_16593);
and U17115 (N_17115,N_16576,N_16710);
nor U17116 (N_17116,N_16731,N_16823);
and U17117 (N_17117,N_16809,N_16718);
xnor U17118 (N_17118,N_16584,N_16866);
xnor U17119 (N_17119,N_16582,N_16732);
and U17120 (N_17120,N_16870,N_16629);
and U17121 (N_17121,N_16773,N_16728);
and U17122 (N_17122,N_16692,N_16706);
or U17123 (N_17123,N_16547,N_16974);
xor U17124 (N_17124,N_16725,N_16549);
nand U17125 (N_17125,N_16633,N_16975);
and U17126 (N_17126,N_16634,N_16849);
xor U17127 (N_17127,N_16930,N_16858);
or U17128 (N_17128,N_16958,N_16599);
or U17129 (N_17129,N_16776,N_16774);
nand U17130 (N_17130,N_16539,N_16986);
and U17131 (N_17131,N_16537,N_16712);
and U17132 (N_17132,N_16750,N_16962);
and U17133 (N_17133,N_16711,N_16620);
or U17134 (N_17134,N_16924,N_16709);
nand U17135 (N_17135,N_16772,N_16726);
and U17136 (N_17136,N_16509,N_16970);
and U17137 (N_17137,N_16998,N_16841);
nand U17138 (N_17138,N_16678,N_16597);
and U17139 (N_17139,N_16562,N_16786);
xor U17140 (N_17140,N_16614,N_16717);
nor U17141 (N_17141,N_16690,N_16923);
and U17142 (N_17142,N_16737,N_16736);
nor U17143 (N_17143,N_16929,N_16907);
nor U17144 (N_17144,N_16680,N_16623);
nand U17145 (N_17145,N_16611,N_16919);
nand U17146 (N_17146,N_16938,N_16860);
nor U17147 (N_17147,N_16754,N_16528);
nor U17148 (N_17148,N_16742,N_16729);
nor U17149 (N_17149,N_16747,N_16515);
or U17150 (N_17150,N_16676,N_16839);
nor U17151 (N_17151,N_16705,N_16734);
and U17152 (N_17152,N_16811,N_16735);
xnor U17153 (N_17153,N_16708,N_16916);
or U17154 (N_17154,N_16876,N_16616);
nor U17155 (N_17155,N_16685,N_16960);
and U17156 (N_17156,N_16740,N_16645);
xor U17157 (N_17157,N_16580,N_16591);
nand U17158 (N_17158,N_16642,N_16748);
xor U17159 (N_17159,N_16564,N_16901);
xor U17160 (N_17160,N_16842,N_16996);
and U17161 (N_17161,N_16531,N_16953);
or U17162 (N_17162,N_16768,N_16559);
xnor U17163 (N_17163,N_16920,N_16529);
or U17164 (N_17164,N_16905,N_16791);
nand U17165 (N_17165,N_16618,N_16636);
nor U17166 (N_17166,N_16925,N_16864);
nand U17167 (N_17167,N_16893,N_16967);
xor U17168 (N_17168,N_16721,N_16505);
nor U17169 (N_17169,N_16513,N_16535);
nand U17170 (N_17170,N_16511,N_16815);
or U17171 (N_17171,N_16933,N_16598);
nor U17172 (N_17172,N_16979,N_16510);
xor U17173 (N_17173,N_16507,N_16835);
nand U17174 (N_17174,N_16741,N_16914);
or U17175 (N_17175,N_16687,N_16739);
nor U17176 (N_17176,N_16961,N_16872);
nand U17177 (N_17177,N_16523,N_16714);
nor U17178 (N_17178,N_16795,N_16627);
or U17179 (N_17179,N_16621,N_16818);
and U17180 (N_17180,N_16827,N_16759);
or U17181 (N_17181,N_16590,N_16646);
nor U17182 (N_17182,N_16899,N_16661);
and U17183 (N_17183,N_16579,N_16840);
nand U17184 (N_17184,N_16985,N_16656);
or U17185 (N_17185,N_16977,N_16638);
xor U17186 (N_17186,N_16861,N_16756);
nand U17187 (N_17187,N_16871,N_16987);
or U17188 (N_17188,N_16856,N_16544);
and U17189 (N_17189,N_16749,N_16794);
nand U17190 (N_17190,N_16512,N_16947);
or U17191 (N_17191,N_16988,N_16931);
and U17192 (N_17192,N_16826,N_16503);
or U17193 (N_17193,N_16563,N_16879);
nor U17194 (N_17194,N_16758,N_16596);
nand U17195 (N_17195,N_16604,N_16762);
nor U17196 (N_17196,N_16873,N_16681);
nand U17197 (N_17197,N_16610,N_16757);
and U17198 (N_17198,N_16845,N_16517);
or U17199 (N_17199,N_16667,N_16926);
xnor U17200 (N_17200,N_16722,N_16934);
xor U17201 (N_17201,N_16778,N_16658);
or U17202 (N_17202,N_16781,N_16682);
nand U17203 (N_17203,N_16635,N_16746);
or U17204 (N_17204,N_16652,N_16763);
or U17205 (N_17205,N_16957,N_16892);
or U17206 (N_17206,N_16603,N_16500);
nor U17207 (N_17207,N_16766,N_16883);
or U17208 (N_17208,N_16693,N_16707);
xnor U17209 (N_17209,N_16800,N_16874);
nor U17210 (N_17210,N_16601,N_16973);
nor U17211 (N_17211,N_16751,N_16530);
xnor U17212 (N_17212,N_16793,N_16963);
or U17213 (N_17213,N_16854,N_16581);
and U17214 (N_17214,N_16760,N_16990);
xnor U17215 (N_17215,N_16808,N_16951);
and U17216 (N_17216,N_16677,N_16671);
xnor U17217 (N_17217,N_16643,N_16943);
or U17218 (N_17218,N_16954,N_16556);
xnor U17219 (N_17219,N_16670,N_16780);
or U17220 (N_17220,N_16578,N_16964);
or U17221 (N_17221,N_16829,N_16600);
or U17222 (N_17222,N_16833,N_16884);
and U17223 (N_17223,N_16853,N_16552);
xnor U17224 (N_17224,N_16553,N_16738);
or U17225 (N_17225,N_16683,N_16585);
or U17226 (N_17226,N_16881,N_16806);
and U17227 (N_17227,N_16752,N_16686);
nor U17228 (N_17228,N_16608,N_16895);
nor U17229 (N_17229,N_16918,N_16821);
nand U17230 (N_17230,N_16959,N_16540);
nand U17231 (N_17231,N_16976,N_16639);
nor U17232 (N_17232,N_16882,N_16972);
or U17233 (N_17233,N_16939,N_16679);
or U17234 (N_17234,N_16995,N_16654);
and U17235 (N_17235,N_16932,N_16764);
or U17236 (N_17236,N_16900,N_16991);
and U17237 (N_17237,N_16971,N_16875);
xor U17238 (N_17238,N_16999,N_16913);
or U17239 (N_17239,N_16981,N_16765);
or U17240 (N_17240,N_16775,N_16612);
xor U17241 (N_17241,N_16911,N_16569);
nand U17242 (N_17242,N_16688,N_16674);
or U17243 (N_17243,N_16955,N_16817);
or U17244 (N_17244,N_16588,N_16906);
nor U17245 (N_17245,N_16819,N_16952);
nand U17246 (N_17246,N_16844,N_16716);
nand U17247 (N_17247,N_16824,N_16956);
or U17248 (N_17248,N_16880,N_16689);
nand U17249 (N_17249,N_16548,N_16813);
or U17250 (N_17250,N_16812,N_16581);
or U17251 (N_17251,N_16506,N_16552);
or U17252 (N_17252,N_16862,N_16509);
or U17253 (N_17253,N_16919,N_16552);
and U17254 (N_17254,N_16776,N_16729);
and U17255 (N_17255,N_16809,N_16652);
or U17256 (N_17256,N_16734,N_16716);
xor U17257 (N_17257,N_16667,N_16800);
nand U17258 (N_17258,N_16635,N_16808);
and U17259 (N_17259,N_16557,N_16613);
and U17260 (N_17260,N_16605,N_16968);
xor U17261 (N_17261,N_16710,N_16859);
and U17262 (N_17262,N_16667,N_16966);
and U17263 (N_17263,N_16658,N_16825);
nand U17264 (N_17264,N_16527,N_16803);
nand U17265 (N_17265,N_16672,N_16900);
xnor U17266 (N_17266,N_16612,N_16717);
nor U17267 (N_17267,N_16784,N_16653);
nand U17268 (N_17268,N_16886,N_16604);
nor U17269 (N_17269,N_16989,N_16990);
nor U17270 (N_17270,N_16641,N_16711);
xnor U17271 (N_17271,N_16908,N_16571);
or U17272 (N_17272,N_16961,N_16642);
xor U17273 (N_17273,N_16528,N_16785);
and U17274 (N_17274,N_16623,N_16537);
xor U17275 (N_17275,N_16975,N_16992);
or U17276 (N_17276,N_16524,N_16832);
nand U17277 (N_17277,N_16929,N_16867);
xor U17278 (N_17278,N_16969,N_16628);
xnor U17279 (N_17279,N_16761,N_16542);
and U17280 (N_17280,N_16813,N_16779);
or U17281 (N_17281,N_16748,N_16501);
nand U17282 (N_17282,N_16764,N_16633);
or U17283 (N_17283,N_16771,N_16567);
nand U17284 (N_17284,N_16736,N_16602);
and U17285 (N_17285,N_16729,N_16862);
xnor U17286 (N_17286,N_16623,N_16575);
nor U17287 (N_17287,N_16574,N_16742);
or U17288 (N_17288,N_16743,N_16827);
nor U17289 (N_17289,N_16502,N_16893);
or U17290 (N_17290,N_16885,N_16670);
nor U17291 (N_17291,N_16507,N_16779);
xor U17292 (N_17292,N_16681,N_16819);
nand U17293 (N_17293,N_16630,N_16563);
nand U17294 (N_17294,N_16567,N_16723);
nor U17295 (N_17295,N_16646,N_16508);
xor U17296 (N_17296,N_16759,N_16691);
or U17297 (N_17297,N_16801,N_16897);
xnor U17298 (N_17298,N_16668,N_16914);
and U17299 (N_17299,N_16731,N_16809);
xor U17300 (N_17300,N_16560,N_16518);
and U17301 (N_17301,N_16681,N_16634);
or U17302 (N_17302,N_16952,N_16523);
or U17303 (N_17303,N_16697,N_16656);
nor U17304 (N_17304,N_16641,N_16570);
and U17305 (N_17305,N_16825,N_16990);
or U17306 (N_17306,N_16528,N_16579);
or U17307 (N_17307,N_16715,N_16894);
xor U17308 (N_17308,N_16919,N_16594);
nand U17309 (N_17309,N_16886,N_16656);
xor U17310 (N_17310,N_16895,N_16788);
nor U17311 (N_17311,N_16855,N_16923);
or U17312 (N_17312,N_16886,N_16984);
or U17313 (N_17313,N_16562,N_16946);
nand U17314 (N_17314,N_16603,N_16640);
and U17315 (N_17315,N_16748,N_16880);
nand U17316 (N_17316,N_16965,N_16551);
xor U17317 (N_17317,N_16879,N_16659);
nor U17318 (N_17318,N_16624,N_16704);
nor U17319 (N_17319,N_16664,N_16580);
xnor U17320 (N_17320,N_16924,N_16754);
xnor U17321 (N_17321,N_16588,N_16942);
or U17322 (N_17322,N_16929,N_16528);
nand U17323 (N_17323,N_16531,N_16759);
or U17324 (N_17324,N_16790,N_16839);
nand U17325 (N_17325,N_16740,N_16675);
nand U17326 (N_17326,N_16938,N_16782);
xnor U17327 (N_17327,N_16987,N_16875);
nand U17328 (N_17328,N_16780,N_16504);
nor U17329 (N_17329,N_16888,N_16654);
xor U17330 (N_17330,N_16945,N_16643);
nor U17331 (N_17331,N_16883,N_16585);
xnor U17332 (N_17332,N_16777,N_16718);
nor U17333 (N_17333,N_16738,N_16628);
nand U17334 (N_17334,N_16936,N_16940);
nand U17335 (N_17335,N_16767,N_16638);
nor U17336 (N_17336,N_16995,N_16722);
or U17337 (N_17337,N_16714,N_16759);
and U17338 (N_17338,N_16722,N_16976);
or U17339 (N_17339,N_16832,N_16852);
nor U17340 (N_17340,N_16531,N_16550);
nand U17341 (N_17341,N_16614,N_16704);
or U17342 (N_17342,N_16615,N_16620);
nand U17343 (N_17343,N_16718,N_16636);
xnor U17344 (N_17344,N_16759,N_16939);
nand U17345 (N_17345,N_16545,N_16730);
or U17346 (N_17346,N_16534,N_16675);
or U17347 (N_17347,N_16516,N_16552);
nor U17348 (N_17348,N_16658,N_16767);
and U17349 (N_17349,N_16867,N_16562);
nand U17350 (N_17350,N_16532,N_16889);
or U17351 (N_17351,N_16958,N_16861);
nor U17352 (N_17352,N_16746,N_16991);
nand U17353 (N_17353,N_16773,N_16915);
or U17354 (N_17354,N_16955,N_16811);
and U17355 (N_17355,N_16817,N_16634);
nand U17356 (N_17356,N_16581,N_16511);
nor U17357 (N_17357,N_16644,N_16909);
xor U17358 (N_17358,N_16972,N_16941);
or U17359 (N_17359,N_16718,N_16899);
nor U17360 (N_17360,N_16541,N_16862);
xor U17361 (N_17361,N_16756,N_16731);
nand U17362 (N_17362,N_16556,N_16704);
or U17363 (N_17363,N_16758,N_16852);
nor U17364 (N_17364,N_16981,N_16620);
nor U17365 (N_17365,N_16750,N_16660);
or U17366 (N_17366,N_16684,N_16667);
and U17367 (N_17367,N_16765,N_16940);
or U17368 (N_17368,N_16674,N_16877);
and U17369 (N_17369,N_16644,N_16938);
xnor U17370 (N_17370,N_16801,N_16893);
nor U17371 (N_17371,N_16903,N_16539);
and U17372 (N_17372,N_16630,N_16633);
nand U17373 (N_17373,N_16818,N_16722);
nand U17374 (N_17374,N_16960,N_16505);
nor U17375 (N_17375,N_16736,N_16754);
nand U17376 (N_17376,N_16507,N_16637);
or U17377 (N_17377,N_16751,N_16519);
nand U17378 (N_17378,N_16874,N_16582);
or U17379 (N_17379,N_16573,N_16675);
nand U17380 (N_17380,N_16874,N_16782);
nand U17381 (N_17381,N_16686,N_16865);
nor U17382 (N_17382,N_16704,N_16866);
and U17383 (N_17383,N_16867,N_16966);
xor U17384 (N_17384,N_16782,N_16978);
nand U17385 (N_17385,N_16707,N_16734);
nand U17386 (N_17386,N_16863,N_16526);
nor U17387 (N_17387,N_16610,N_16918);
nand U17388 (N_17388,N_16714,N_16858);
nand U17389 (N_17389,N_16675,N_16977);
nand U17390 (N_17390,N_16893,N_16561);
and U17391 (N_17391,N_16565,N_16750);
xnor U17392 (N_17392,N_16530,N_16799);
nand U17393 (N_17393,N_16618,N_16819);
nor U17394 (N_17394,N_16587,N_16696);
nor U17395 (N_17395,N_16915,N_16862);
nand U17396 (N_17396,N_16686,N_16569);
and U17397 (N_17397,N_16808,N_16728);
nand U17398 (N_17398,N_16735,N_16657);
xnor U17399 (N_17399,N_16682,N_16507);
xnor U17400 (N_17400,N_16794,N_16970);
nand U17401 (N_17401,N_16754,N_16902);
and U17402 (N_17402,N_16563,N_16935);
nor U17403 (N_17403,N_16853,N_16544);
nor U17404 (N_17404,N_16923,N_16792);
nor U17405 (N_17405,N_16908,N_16530);
nor U17406 (N_17406,N_16538,N_16745);
or U17407 (N_17407,N_16781,N_16956);
nand U17408 (N_17408,N_16978,N_16669);
or U17409 (N_17409,N_16613,N_16668);
nor U17410 (N_17410,N_16589,N_16580);
or U17411 (N_17411,N_16971,N_16831);
or U17412 (N_17412,N_16880,N_16944);
nor U17413 (N_17413,N_16776,N_16865);
and U17414 (N_17414,N_16809,N_16997);
or U17415 (N_17415,N_16862,N_16986);
and U17416 (N_17416,N_16559,N_16618);
nand U17417 (N_17417,N_16894,N_16936);
xnor U17418 (N_17418,N_16878,N_16836);
nand U17419 (N_17419,N_16676,N_16824);
xor U17420 (N_17420,N_16870,N_16687);
xnor U17421 (N_17421,N_16965,N_16593);
xor U17422 (N_17422,N_16894,N_16944);
nand U17423 (N_17423,N_16663,N_16652);
or U17424 (N_17424,N_16962,N_16883);
and U17425 (N_17425,N_16726,N_16854);
nand U17426 (N_17426,N_16593,N_16678);
xnor U17427 (N_17427,N_16872,N_16825);
or U17428 (N_17428,N_16960,N_16596);
and U17429 (N_17429,N_16985,N_16617);
or U17430 (N_17430,N_16862,N_16837);
and U17431 (N_17431,N_16601,N_16776);
or U17432 (N_17432,N_16784,N_16599);
nor U17433 (N_17433,N_16749,N_16605);
xnor U17434 (N_17434,N_16575,N_16650);
xor U17435 (N_17435,N_16560,N_16638);
xnor U17436 (N_17436,N_16502,N_16695);
and U17437 (N_17437,N_16922,N_16736);
and U17438 (N_17438,N_16528,N_16509);
or U17439 (N_17439,N_16540,N_16946);
or U17440 (N_17440,N_16504,N_16667);
nor U17441 (N_17441,N_16734,N_16929);
or U17442 (N_17442,N_16853,N_16795);
xor U17443 (N_17443,N_16905,N_16884);
xnor U17444 (N_17444,N_16528,N_16947);
xnor U17445 (N_17445,N_16784,N_16862);
nand U17446 (N_17446,N_16630,N_16819);
nor U17447 (N_17447,N_16748,N_16640);
nand U17448 (N_17448,N_16636,N_16866);
or U17449 (N_17449,N_16696,N_16801);
and U17450 (N_17450,N_16912,N_16890);
xor U17451 (N_17451,N_16873,N_16705);
nand U17452 (N_17452,N_16636,N_16557);
nor U17453 (N_17453,N_16945,N_16887);
nor U17454 (N_17454,N_16992,N_16955);
and U17455 (N_17455,N_16949,N_16801);
or U17456 (N_17456,N_16798,N_16986);
nor U17457 (N_17457,N_16917,N_16907);
nor U17458 (N_17458,N_16919,N_16534);
and U17459 (N_17459,N_16785,N_16926);
and U17460 (N_17460,N_16747,N_16507);
or U17461 (N_17461,N_16769,N_16611);
and U17462 (N_17462,N_16660,N_16513);
nor U17463 (N_17463,N_16770,N_16681);
or U17464 (N_17464,N_16563,N_16577);
and U17465 (N_17465,N_16914,N_16543);
nand U17466 (N_17466,N_16951,N_16790);
and U17467 (N_17467,N_16828,N_16605);
and U17468 (N_17468,N_16760,N_16919);
xnor U17469 (N_17469,N_16995,N_16904);
nor U17470 (N_17470,N_16597,N_16986);
and U17471 (N_17471,N_16743,N_16794);
xor U17472 (N_17472,N_16576,N_16823);
nor U17473 (N_17473,N_16886,N_16759);
xnor U17474 (N_17474,N_16559,N_16736);
xor U17475 (N_17475,N_16936,N_16596);
xnor U17476 (N_17476,N_16595,N_16916);
nand U17477 (N_17477,N_16663,N_16743);
nand U17478 (N_17478,N_16741,N_16673);
and U17479 (N_17479,N_16744,N_16996);
and U17480 (N_17480,N_16861,N_16842);
or U17481 (N_17481,N_16726,N_16847);
nand U17482 (N_17482,N_16662,N_16712);
nand U17483 (N_17483,N_16796,N_16810);
nand U17484 (N_17484,N_16794,N_16736);
nor U17485 (N_17485,N_16889,N_16609);
xor U17486 (N_17486,N_16746,N_16930);
and U17487 (N_17487,N_16815,N_16807);
nor U17488 (N_17488,N_16782,N_16975);
or U17489 (N_17489,N_16796,N_16827);
or U17490 (N_17490,N_16587,N_16520);
nor U17491 (N_17491,N_16719,N_16953);
or U17492 (N_17492,N_16721,N_16563);
xor U17493 (N_17493,N_16658,N_16652);
nor U17494 (N_17494,N_16577,N_16544);
or U17495 (N_17495,N_16715,N_16627);
xor U17496 (N_17496,N_16952,N_16654);
xor U17497 (N_17497,N_16517,N_16564);
or U17498 (N_17498,N_16849,N_16589);
and U17499 (N_17499,N_16642,N_16876);
and U17500 (N_17500,N_17101,N_17059);
or U17501 (N_17501,N_17133,N_17477);
nor U17502 (N_17502,N_17333,N_17453);
nand U17503 (N_17503,N_17200,N_17265);
nand U17504 (N_17504,N_17423,N_17237);
nor U17505 (N_17505,N_17252,N_17000);
xnor U17506 (N_17506,N_17148,N_17212);
nor U17507 (N_17507,N_17343,N_17066);
or U17508 (N_17508,N_17466,N_17422);
nand U17509 (N_17509,N_17224,N_17073);
nand U17510 (N_17510,N_17206,N_17313);
nor U17511 (N_17511,N_17419,N_17410);
nor U17512 (N_17512,N_17281,N_17289);
or U17513 (N_17513,N_17007,N_17069);
nor U17514 (N_17514,N_17068,N_17050);
xor U17515 (N_17515,N_17219,N_17121);
nand U17516 (N_17516,N_17296,N_17338);
nand U17517 (N_17517,N_17149,N_17418);
and U17518 (N_17518,N_17468,N_17352);
xor U17519 (N_17519,N_17063,N_17027);
nand U17520 (N_17520,N_17037,N_17258);
and U17521 (N_17521,N_17361,N_17303);
or U17522 (N_17522,N_17354,N_17010);
or U17523 (N_17523,N_17432,N_17260);
xnor U17524 (N_17524,N_17385,N_17062);
or U17525 (N_17525,N_17482,N_17285);
nor U17526 (N_17526,N_17401,N_17249);
or U17527 (N_17527,N_17056,N_17012);
nand U17528 (N_17528,N_17328,N_17194);
xor U17529 (N_17529,N_17132,N_17127);
nand U17530 (N_17530,N_17025,N_17225);
or U17531 (N_17531,N_17198,N_17039);
nor U17532 (N_17532,N_17091,N_17368);
or U17533 (N_17533,N_17088,N_17040);
or U17534 (N_17534,N_17118,N_17465);
nand U17535 (N_17535,N_17264,N_17229);
or U17536 (N_17536,N_17145,N_17072);
nand U17537 (N_17537,N_17452,N_17388);
nor U17538 (N_17538,N_17254,N_17028);
nand U17539 (N_17539,N_17097,N_17160);
and U17540 (N_17540,N_17332,N_17446);
nand U17541 (N_17541,N_17309,N_17142);
and U17542 (N_17542,N_17112,N_17382);
xor U17543 (N_17543,N_17394,N_17403);
and U17544 (N_17544,N_17483,N_17263);
and U17545 (N_17545,N_17287,N_17307);
nand U17546 (N_17546,N_17234,N_17030);
nand U17547 (N_17547,N_17045,N_17034);
and U17548 (N_17548,N_17353,N_17440);
nand U17549 (N_17549,N_17146,N_17284);
xnor U17550 (N_17550,N_17412,N_17359);
and U17551 (N_17551,N_17201,N_17444);
nor U17552 (N_17552,N_17086,N_17499);
and U17553 (N_17553,N_17397,N_17250);
nor U17554 (N_17554,N_17277,N_17203);
and U17555 (N_17555,N_17192,N_17116);
or U17556 (N_17556,N_17496,N_17235);
or U17557 (N_17557,N_17035,N_17020);
or U17558 (N_17558,N_17367,N_17271);
nor U17559 (N_17559,N_17016,N_17084);
xor U17560 (N_17560,N_17227,N_17002);
nor U17561 (N_17561,N_17436,N_17438);
and U17562 (N_17562,N_17255,N_17318);
nor U17563 (N_17563,N_17075,N_17378);
nand U17564 (N_17564,N_17341,N_17408);
and U17565 (N_17565,N_17288,N_17240);
or U17566 (N_17566,N_17302,N_17449);
nand U17567 (N_17567,N_17129,N_17492);
and U17568 (N_17568,N_17104,N_17464);
nand U17569 (N_17569,N_17349,N_17162);
xnor U17570 (N_17570,N_17498,N_17126);
or U17571 (N_17571,N_17373,N_17488);
xor U17572 (N_17572,N_17082,N_17380);
nand U17573 (N_17573,N_17166,N_17369);
and U17574 (N_17574,N_17154,N_17305);
and U17575 (N_17575,N_17413,N_17023);
or U17576 (N_17576,N_17014,N_17430);
or U17577 (N_17577,N_17135,N_17003);
nand U17578 (N_17578,N_17360,N_17304);
or U17579 (N_17579,N_17321,N_17090);
nand U17580 (N_17580,N_17467,N_17013);
nand U17581 (N_17581,N_17077,N_17085);
or U17582 (N_17582,N_17024,N_17152);
and U17583 (N_17583,N_17099,N_17017);
or U17584 (N_17584,N_17136,N_17243);
nor U17585 (N_17585,N_17437,N_17124);
or U17586 (N_17586,N_17119,N_17167);
xor U17587 (N_17587,N_17141,N_17331);
and U17588 (N_17588,N_17241,N_17424);
nor U17589 (N_17589,N_17386,N_17336);
or U17590 (N_17590,N_17163,N_17159);
and U17591 (N_17591,N_17290,N_17251);
nand U17592 (N_17592,N_17402,N_17270);
nor U17593 (N_17593,N_17046,N_17448);
nor U17594 (N_17594,N_17355,N_17026);
and U17595 (N_17595,N_17247,N_17215);
and U17596 (N_17596,N_17151,N_17473);
and U17597 (N_17597,N_17130,N_17348);
nor U17598 (N_17598,N_17187,N_17295);
or U17599 (N_17599,N_17393,N_17398);
xor U17600 (N_17600,N_17409,N_17174);
nand U17601 (N_17601,N_17233,N_17186);
and U17602 (N_17602,N_17087,N_17497);
nand U17603 (N_17603,N_17232,N_17370);
nand U17604 (N_17604,N_17274,N_17070);
nand U17605 (N_17605,N_17414,N_17098);
xor U17606 (N_17606,N_17376,N_17122);
nand U17607 (N_17607,N_17214,N_17218);
xnor U17608 (N_17608,N_17381,N_17029);
nor U17609 (N_17609,N_17058,N_17479);
nor U17610 (N_17610,N_17404,N_17207);
xnor U17611 (N_17611,N_17351,N_17399);
and U17612 (N_17612,N_17458,N_17415);
and U17613 (N_17613,N_17036,N_17257);
nand U17614 (N_17614,N_17253,N_17245);
xnor U17615 (N_17615,N_17226,N_17317);
and U17616 (N_17616,N_17366,N_17079);
and U17617 (N_17617,N_17078,N_17442);
or U17618 (N_17618,N_17182,N_17044);
or U17619 (N_17619,N_17161,N_17334);
or U17620 (N_17620,N_17076,N_17048);
xor U17621 (N_17621,N_17322,N_17259);
nor U17622 (N_17622,N_17139,N_17469);
and U17623 (N_17623,N_17278,N_17276);
or U17624 (N_17624,N_17481,N_17327);
or U17625 (N_17625,N_17049,N_17093);
xnor U17626 (N_17626,N_17391,N_17312);
nand U17627 (N_17627,N_17096,N_17495);
or U17628 (N_17628,N_17291,N_17137);
nor U17629 (N_17629,N_17282,N_17364);
and U17630 (N_17630,N_17392,N_17463);
or U17631 (N_17631,N_17443,N_17319);
and U17632 (N_17632,N_17365,N_17065);
and U17633 (N_17633,N_17205,N_17306);
nor U17634 (N_17634,N_17406,N_17131);
xnor U17635 (N_17635,N_17294,N_17197);
or U17636 (N_17636,N_17164,N_17390);
and U17637 (N_17637,N_17177,N_17363);
xnor U17638 (N_17638,N_17478,N_17342);
and U17639 (N_17639,N_17293,N_17202);
nand U17640 (N_17640,N_17396,N_17326);
nand U17641 (N_17641,N_17196,N_17178);
and U17642 (N_17642,N_17387,N_17221);
or U17643 (N_17643,N_17081,N_17032);
xor U17644 (N_17644,N_17143,N_17213);
or U17645 (N_17645,N_17439,N_17494);
xnor U17646 (N_17646,N_17374,N_17314);
nand U17647 (N_17647,N_17171,N_17019);
and U17648 (N_17648,N_17457,N_17009);
and U17649 (N_17649,N_17067,N_17324);
or U17650 (N_17650,N_17301,N_17286);
xor U17651 (N_17651,N_17450,N_17199);
nor U17652 (N_17652,N_17184,N_17421);
and U17653 (N_17653,N_17176,N_17346);
or U17654 (N_17654,N_17471,N_17375);
and U17655 (N_17655,N_17231,N_17242);
nor U17656 (N_17656,N_17022,N_17470);
and U17657 (N_17657,N_17134,N_17300);
xor U17658 (N_17658,N_17005,N_17111);
xor U17659 (N_17659,N_17001,N_17474);
nor U17660 (N_17660,N_17172,N_17055);
and U17661 (N_17661,N_17433,N_17292);
or U17662 (N_17662,N_17004,N_17445);
xnor U17663 (N_17663,N_17175,N_17060);
and U17664 (N_17664,N_17114,N_17180);
xnor U17665 (N_17665,N_17230,N_17357);
and U17666 (N_17666,N_17041,N_17475);
nor U17667 (N_17667,N_17083,N_17095);
nand U17668 (N_17668,N_17211,N_17246);
nor U17669 (N_17669,N_17427,N_17074);
and U17670 (N_17670,N_17108,N_17429);
nand U17671 (N_17671,N_17447,N_17435);
xnor U17672 (N_17672,N_17185,N_17311);
nand U17673 (N_17673,N_17384,N_17047);
or U17674 (N_17674,N_17248,N_17189);
and U17675 (N_17675,N_17476,N_17279);
nand U17676 (N_17676,N_17372,N_17490);
or U17677 (N_17677,N_17209,N_17157);
or U17678 (N_17678,N_17428,N_17280);
and U17679 (N_17679,N_17238,N_17094);
or U17680 (N_17680,N_17244,N_17299);
and U17681 (N_17681,N_17472,N_17434);
nand U17682 (N_17682,N_17109,N_17191);
nor U17683 (N_17683,N_17011,N_17165);
or U17684 (N_17684,N_17018,N_17308);
and U17685 (N_17685,N_17183,N_17115);
nor U17686 (N_17686,N_17272,N_17275);
nand U17687 (N_17687,N_17223,N_17273);
or U17688 (N_17688,N_17451,N_17092);
xnor U17689 (N_17689,N_17057,N_17316);
and U17690 (N_17690,N_17400,N_17195);
nor U17691 (N_17691,N_17340,N_17485);
xnor U17692 (N_17692,N_17217,N_17015);
or U17693 (N_17693,N_17416,N_17347);
xnor U17694 (N_17694,N_17426,N_17460);
nand U17695 (N_17695,N_17283,N_17325);
and U17696 (N_17696,N_17236,N_17008);
nor U17697 (N_17697,N_17123,N_17220);
or U17698 (N_17698,N_17155,N_17459);
xor U17699 (N_17699,N_17089,N_17106);
and U17700 (N_17700,N_17486,N_17051);
nand U17701 (N_17701,N_17038,N_17033);
nor U17702 (N_17702,N_17125,N_17345);
and U17703 (N_17703,N_17169,N_17407);
and U17704 (N_17704,N_17168,N_17480);
or U17705 (N_17705,N_17128,N_17193);
xor U17706 (N_17706,N_17021,N_17042);
nand U17707 (N_17707,N_17454,N_17239);
or U17708 (N_17708,N_17350,N_17204);
nor U17709 (N_17709,N_17054,N_17190);
xor U17710 (N_17710,N_17102,N_17487);
or U17711 (N_17711,N_17188,N_17140);
or U17712 (N_17712,N_17031,N_17071);
nand U17713 (N_17713,N_17344,N_17491);
xor U17714 (N_17714,N_17179,N_17268);
nand U17715 (N_17715,N_17310,N_17120);
nand U17716 (N_17716,N_17377,N_17358);
xnor U17717 (N_17717,N_17107,N_17425);
nor U17718 (N_17718,N_17337,N_17150);
nor U17719 (N_17719,N_17383,N_17228);
or U17720 (N_17720,N_17256,N_17103);
and U17721 (N_17721,N_17323,N_17262);
and U17722 (N_17722,N_17456,N_17297);
and U17723 (N_17723,N_17329,N_17420);
nor U17724 (N_17724,N_17170,N_17105);
nor U17725 (N_17725,N_17315,N_17261);
or U17726 (N_17726,N_17389,N_17153);
xor U17727 (N_17727,N_17100,N_17493);
or U17728 (N_17728,N_17222,N_17356);
and U17729 (N_17729,N_17489,N_17441);
xnor U17730 (N_17730,N_17064,N_17462);
xor U17731 (N_17731,N_17144,N_17267);
or U17732 (N_17732,N_17117,N_17006);
and U17733 (N_17733,N_17080,N_17147);
or U17734 (N_17734,N_17043,N_17216);
and U17735 (N_17735,N_17113,N_17320);
xnor U17736 (N_17736,N_17379,N_17181);
xnor U17737 (N_17737,N_17411,N_17210);
or U17738 (N_17738,N_17208,N_17484);
or U17739 (N_17739,N_17053,N_17339);
nand U17740 (N_17740,N_17395,N_17330);
nand U17741 (N_17741,N_17173,N_17461);
nand U17742 (N_17742,N_17371,N_17061);
nand U17743 (N_17743,N_17417,N_17455);
or U17744 (N_17744,N_17110,N_17052);
or U17745 (N_17745,N_17269,N_17405);
or U17746 (N_17746,N_17266,N_17156);
nor U17747 (N_17747,N_17138,N_17335);
and U17748 (N_17748,N_17298,N_17158);
or U17749 (N_17749,N_17362,N_17431);
nand U17750 (N_17750,N_17236,N_17155);
and U17751 (N_17751,N_17053,N_17480);
nor U17752 (N_17752,N_17325,N_17367);
and U17753 (N_17753,N_17193,N_17046);
nand U17754 (N_17754,N_17180,N_17238);
or U17755 (N_17755,N_17145,N_17150);
nand U17756 (N_17756,N_17020,N_17477);
nand U17757 (N_17757,N_17285,N_17082);
or U17758 (N_17758,N_17418,N_17168);
nor U17759 (N_17759,N_17105,N_17371);
and U17760 (N_17760,N_17299,N_17227);
xnor U17761 (N_17761,N_17475,N_17338);
nand U17762 (N_17762,N_17183,N_17381);
or U17763 (N_17763,N_17346,N_17314);
and U17764 (N_17764,N_17375,N_17477);
xor U17765 (N_17765,N_17180,N_17073);
and U17766 (N_17766,N_17463,N_17017);
and U17767 (N_17767,N_17467,N_17223);
nand U17768 (N_17768,N_17482,N_17352);
nand U17769 (N_17769,N_17203,N_17428);
nand U17770 (N_17770,N_17287,N_17175);
nand U17771 (N_17771,N_17155,N_17378);
or U17772 (N_17772,N_17057,N_17097);
nor U17773 (N_17773,N_17132,N_17194);
and U17774 (N_17774,N_17416,N_17420);
or U17775 (N_17775,N_17340,N_17491);
or U17776 (N_17776,N_17327,N_17403);
and U17777 (N_17777,N_17278,N_17254);
nor U17778 (N_17778,N_17097,N_17061);
nand U17779 (N_17779,N_17322,N_17343);
xnor U17780 (N_17780,N_17086,N_17468);
or U17781 (N_17781,N_17099,N_17253);
or U17782 (N_17782,N_17183,N_17199);
nor U17783 (N_17783,N_17163,N_17199);
xor U17784 (N_17784,N_17215,N_17071);
xnor U17785 (N_17785,N_17327,N_17224);
and U17786 (N_17786,N_17235,N_17312);
and U17787 (N_17787,N_17105,N_17020);
xor U17788 (N_17788,N_17243,N_17266);
and U17789 (N_17789,N_17165,N_17254);
nand U17790 (N_17790,N_17190,N_17091);
xor U17791 (N_17791,N_17430,N_17290);
nor U17792 (N_17792,N_17431,N_17230);
or U17793 (N_17793,N_17348,N_17145);
or U17794 (N_17794,N_17380,N_17214);
nor U17795 (N_17795,N_17368,N_17395);
xor U17796 (N_17796,N_17250,N_17080);
nor U17797 (N_17797,N_17224,N_17196);
and U17798 (N_17798,N_17343,N_17236);
and U17799 (N_17799,N_17291,N_17464);
and U17800 (N_17800,N_17281,N_17159);
and U17801 (N_17801,N_17242,N_17086);
xnor U17802 (N_17802,N_17287,N_17339);
and U17803 (N_17803,N_17315,N_17388);
xnor U17804 (N_17804,N_17498,N_17133);
xor U17805 (N_17805,N_17159,N_17415);
xnor U17806 (N_17806,N_17095,N_17076);
nand U17807 (N_17807,N_17371,N_17359);
nor U17808 (N_17808,N_17101,N_17350);
and U17809 (N_17809,N_17480,N_17148);
nor U17810 (N_17810,N_17059,N_17073);
and U17811 (N_17811,N_17048,N_17169);
or U17812 (N_17812,N_17192,N_17319);
nand U17813 (N_17813,N_17360,N_17288);
nand U17814 (N_17814,N_17306,N_17299);
nor U17815 (N_17815,N_17498,N_17187);
or U17816 (N_17816,N_17117,N_17141);
and U17817 (N_17817,N_17320,N_17176);
xnor U17818 (N_17818,N_17479,N_17147);
nand U17819 (N_17819,N_17449,N_17345);
or U17820 (N_17820,N_17273,N_17414);
nand U17821 (N_17821,N_17348,N_17223);
nand U17822 (N_17822,N_17211,N_17063);
nor U17823 (N_17823,N_17061,N_17426);
xor U17824 (N_17824,N_17064,N_17463);
nand U17825 (N_17825,N_17301,N_17386);
or U17826 (N_17826,N_17228,N_17330);
and U17827 (N_17827,N_17033,N_17203);
xnor U17828 (N_17828,N_17243,N_17373);
xnor U17829 (N_17829,N_17470,N_17293);
nor U17830 (N_17830,N_17017,N_17220);
nand U17831 (N_17831,N_17230,N_17471);
xnor U17832 (N_17832,N_17414,N_17269);
nor U17833 (N_17833,N_17214,N_17328);
nand U17834 (N_17834,N_17371,N_17071);
nor U17835 (N_17835,N_17264,N_17051);
xor U17836 (N_17836,N_17268,N_17061);
and U17837 (N_17837,N_17312,N_17441);
and U17838 (N_17838,N_17429,N_17431);
and U17839 (N_17839,N_17293,N_17187);
and U17840 (N_17840,N_17356,N_17487);
nor U17841 (N_17841,N_17087,N_17444);
nor U17842 (N_17842,N_17198,N_17055);
nor U17843 (N_17843,N_17176,N_17163);
xnor U17844 (N_17844,N_17333,N_17430);
nor U17845 (N_17845,N_17013,N_17287);
and U17846 (N_17846,N_17106,N_17393);
nor U17847 (N_17847,N_17420,N_17336);
and U17848 (N_17848,N_17366,N_17416);
nand U17849 (N_17849,N_17326,N_17040);
xor U17850 (N_17850,N_17445,N_17163);
or U17851 (N_17851,N_17082,N_17078);
nand U17852 (N_17852,N_17159,N_17324);
xor U17853 (N_17853,N_17138,N_17420);
xnor U17854 (N_17854,N_17074,N_17075);
and U17855 (N_17855,N_17000,N_17360);
nor U17856 (N_17856,N_17305,N_17429);
nand U17857 (N_17857,N_17493,N_17337);
xor U17858 (N_17858,N_17340,N_17134);
nand U17859 (N_17859,N_17193,N_17059);
xnor U17860 (N_17860,N_17173,N_17330);
nand U17861 (N_17861,N_17022,N_17192);
nor U17862 (N_17862,N_17139,N_17045);
nor U17863 (N_17863,N_17243,N_17128);
or U17864 (N_17864,N_17315,N_17174);
xnor U17865 (N_17865,N_17218,N_17469);
xnor U17866 (N_17866,N_17449,N_17070);
and U17867 (N_17867,N_17213,N_17403);
nor U17868 (N_17868,N_17115,N_17326);
nand U17869 (N_17869,N_17141,N_17020);
nor U17870 (N_17870,N_17481,N_17204);
nand U17871 (N_17871,N_17389,N_17492);
nor U17872 (N_17872,N_17303,N_17040);
nand U17873 (N_17873,N_17274,N_17072);
xnor U17874 (N_17874,N_17266,N_17265);
or U17875 (N_17875,N_17462,N_17366);
nor U17876 (N_17876,N_17236,N_17266);
and U17877 (N_17877,N_17191,N_17052);
nand U17878 (N_17878,N_17329,N_17353);
nand U17879 (N_17879,N_17021,N_17337);
nor U17880 (N_17880,N_17268,N_17109);
or U17881 (N_17881,N_17485,N_17123);
xnor U17882 (N_17882,N_17498,N_17124);
and U17883 (N_17883,N_17251,N_17065);
nand U17884 (N_17884,N_17043,N_17334);
and U17885 (N_17885,N_17218,N_17338);
and U17886 (N_17886,N_17303,N_17420);
or U17887 (N_17887,N_17101,N_17131);
nor U17888 (N_17888,N_17286,N_17107);
xor U17889 (N_17889,N_17371,N_17337);
and U17890 (N_17890,N_17171,N_17139);
or U17891 (N_17891,N_17082,N_17468);
or U17892 (N_17892,N_17338,N_17415);
and U17893 (N_17893,N_17234,N_17154);
nor U17894 (N_17894,N_17186,N_17085);
nand U17895 (N_17895,N_17255,N_17268);
nor U17896 (N_17896,N_17258,N_17341);
nor U17897 (N_17897,N_17038,N_17277);
nand U17898 (N_17898,N_17166,N_17308);
or U17899 (N_17899,N_17302,N_17062);
or U17900 (N_17900,N_17127,N_17164);
and U17901 (N_17901,N_17300,N_17084);
nor U17902 (N_17902,N_17315,N_17416);
xor U17903 (N_17903,N_17068,N_17220);
and U17904 (N_17904,N_17343,N_17239);
or U17905 (N_17905,N_17348,N_17456);
nand U17906 (N_17906,N_17489,N_17052);
and U17907 (N_17907,N_17477,N_17347);
xnor U17908 (N_17908,N_17168,N_17332);
nand U17909 (N_17909,N_17117,N_17452);
nand U17910 (N_17910,N_17062,N_17050);
and U17911 (N_17911,N_17188,N_17334);
and U17912 (N_17912,N_17233,N_17255);
or U17913 (N_17913,N_17084,N_17349);
nand U17914 (N_17914,N_17111,N_17175);
nand U17915 (N_17915,N_17319,N_17015);
nor U17916 (N_17916,N_17307,N_17282);
xnor U17917 (N_17917,N_17134,N_17150);
nor U17918 (N_17918,N_17081,N_17111);
and U17919 (N_17919,N_17306,N_17148);
or U17920 (N_17920,N_17113,N_17152);
xor U17921 (N_17921,N_17294,N_17331);
nor U17922 (N_17922,N_17026,N_17289);
nor U17923 (N_17923,N_17481,N_17350);
nand U17924 (N_17924,N_17084,N_17037);
and U17925 (N_17925,N_17302,N_17194);
xor U17926 (N_17926,N_17301,N_17300);
xor U17927 (N_17927,N_17083,N_17332);
and U17928 (N_17928,N_17408,N_17311);
or U17929 (N_17929,N_17047,N_17479);
xor U17930 (N_17930,N_17361,N_17013);
and U17931 (N_17931,N_17379,N_17288);
nand U17932 (N_17932,N_17293,N_17235);
nor U17933 (N_17933,N_17478,N_17162);
or U17934 (N_17934,N_17056,N_17447);
xor U17935 (N_17935,N_17229,N_17182);
nor U17936 (N_17936,N_17399,N_17466);
nor U17937 (N_17937,N_17065,N_17087);
nor U17938 (N_17938,N_17255,N_17426);
or U17939 (N_17939,N_17086,N_17440);
or U17940 (N_17940,N_17016,N_17316);
nand U17941 (N_17941,N_17016,N_17381);
or U17942 (N_17942,N_17102,N_17469);
and U17943 (N_17943,N_17445,N_17124);
and U17944 (N_17944,N_17456,N_17133);
xnor U17945 (N_17945,N_17094,N_17164);
xor U17946 (N_17946,N_17447,N_17362);
or U17947 (N_17947,N_17415,N_17477);
nand U17948 (N_17948,N_17316,N_17023);
and U17949 (N_17949,N_17353,N_17143);
and U17950 (N_17950,N_17345,N_17309);
nand U17951 (N_17951,N_17115,N_17232);
and U17952 (N_17952,N_17294,N_17417);
and U17953 (N_17953,N_17088,N_17279);
xor U17954 (N_17954,N_17450,N_17312);
or U17955 (N_17955,N_17162,N_17128);
nand U17956 (N_17956,N_17131,N_17413);
nor U17957 (N_17957,N_17067,N_17355);
or U17958 (N_17958,N_17368,N_17479);
xnor U17959 (N_17959,N_17374,N_17048);
and U17960 (N_17960,N_17265,N_17261);
or U17961 (N_17961,N_17220,N_17124);
xnor U17962 (N_17962,N_17001,N_17034);
xnor U17963 (N_17963,N_17231,N_17351);
nand U17964 (N_17964,N_17479,N_17324);
nand U17965 (N_17965,N_17353,N_17221);
nand U17966 (N_17966,N_17146,N_17202);
nor U17967 (N_17967,N_17116,N_17485);
nor U17968 (N_17968,N_17437,N_17138);
or U17969 (N_17969,N_17164,N_17258);
nand U17970 (N_17970,N_17017,N_17268);
and U17971 (N_17971,N_17140,N_17227);
nor U17972 (N_17972,N_17250,N_17187);
or U17973 (N_17973,N_17395,N_17431);
xor U17974 (N_17974,N_17086,N_17239);
or U17975 (N_17975,N_17214,N_17034);
xnor U17976 (N_17976,N_17095,N_17257);
xnor U17977 (N_17977,N_17279,N_17055);
xor U17978 (N_17978,N_17174,N_17319);
or U17979 (N_17979,N_17477,N_17085);
nor U17980 (N_17980,N_17105,N_17225);
or U17981 (N_17981,N_17002,N_17199);
nor U17982 (N_17982,N_17235,N_17339);
or U17983 (N_17983,N_17233,N_17470);
nor U17984 (N_17984,N_17092,N_17272);
nor U17985 (N_17985,N_17139,N_17069);
nand U17986 (N_17986,N_17091,N_17240);
nor U17987 (N_17987,N_17139,N_17134);
or U17988 (N_17988,N_17089,N_17190);
nor U17989 (N_17989,N_17494,N_17218);
or U17990 (N_17990,N_17311,N_17074);
and U17991 (N_17991,N_17317,N_17275);
xnor U17992 (N_17992,N_17411,N_17198);
xor U17993 (N_17993,N_17324,N_17217);
nand U17994 (N_17994,N_17029,N_17097);
xnor U17995 (N_17995,N_17161,N_17232);
xnor U17996 (N_17996,N_17382,N_17245);
and U17997 (N_17997,N_17219,N_17206);
xor U17998 (N_17998,N_17285,N_17316);
or U17999 (N_17999,N_17255,N_17481);
xor U18000 (N_18000,N_17736,N_17541);
or U18001 (N_18001,N_17554,N_17869);
xor U18002 (N_18002,N_17596,N_17862);
xor U18003 (N_18003,N_17966,N_17840);
or U18004 (N_18004,N_17581,N_17572);
or U18005 (N_18005,N_17659,N_17500);
nand U18006 (N_18006,N_17597,N_17786);
or U18007 (N_18007,N_17922,N_17986);
nor U18008 (N_18008,N_17912,N_17880);
xnor U18009 (N_18009,N_17956,N_17672);
and U18010 (N_18010,N_17645,N_17867);
and U18011 (N_18011,N_17531,N_17997);
xor U18012 (N_18012,N_17741,N_17951);
and U18013 (N_18013,N_17651,N_17982);
or U18014 (N_18014,N_17923,N_17522);
or U18015 (N_18015,N_17953,N_17977);
and U18016 (N_18016,N_17802,N_17657);
xnor U18017 (N_18017,N_17706,N_17715);
nand U18018 (N_18018,N_17954,N_17726);
nor U18019 (N_18019,N_17910,N_17969);
and U18020 (N_18020,N_17944,N_17996);
nor U18021 (N_18021,N_17720,N_17760);
nor U18022 (N_18022,N_17902,N_17762);
nor U18023 (N_18023,N_17767,N_17559);
nor U18024 (N_18024,N_17794,N_17945);
xor U18025 (N_18025,N_17989,N_17864);
xor U18026 (N_18026,N_17872,N_17918);
nand U18027 (N_18027,N_17623,N_17777);
or U18028 (N_18028,N_17805,N_17856);
xnor U18029 (N_18029,N_17782,N_17682);
nor U18030 (N_18030,N_17789,N_17851);
nand U18031 (N_18031,N_17564,N_17661);
nor U18032 (N_18032,N_17974,N_17981);
nand U18033 (N_18033,N_17671,N_17666);
or U18034 (N_18034,N_17928,N_17825);
xnor U18035 (N_18035,N_17523,N_17933);
and U18036 (N_18036,N_17943,N_17545);
nand U18037 (N_18037,N_17549,N_17538);
and U18038 (N_18038,N_17506,N_17568);
nand U18039 (N_18039,N_17937,N_17703);
or U18040 (N_18040,N_17861,N_17926);
nor U18041 (N_18041,N_17868,N_17664);
xnor U18042 (N_18042,N_17900,N_17562);
nor U18043 (N_18043,N_17758,N_17759);
xnor U18044 (N_18044,N_17935,N_17587);
nand U18045 (N_18045,N_17779,N_17719);
xnor U18046 (N_18046,N_17740,N_17739);
xnor U18047 (N_18047,N_17853,N_17775);
or U18048 (N_18048,N_17924,N_17738);
or U18049 (N_18049,N_17624,N_17622);
xnor U18050 (N_18050,N_17774,N_17536);
nand U18051 (N_18051,N_17705,N_17504);
nand U18052 (N_18052,N_17772,N_17567);
and U18053 (N_18053,N_17848,N_17887);
nand U18054 (N_18054,N_17746,N_17668);
and U18055 (N_18055,N_17617,N_17785);
or U18056 (N_18056,N_17612,N_17898);
xor U18057 (N_18057,N_17631,N_17971);
nand U18058 (N_18058,N_17566,N_17803);
or U18059 (N_18059,N_17710,N_17896);
xnor U18060 (N_18060,N_17917,N_17921);
xor U18061 (N_18061,N_17532,N_17535);
and U18062 (N_18062,N_17580,N_17806);
nor U18063 (N_18063,N_17721,N_17801);
or U18064 (N_18064,N_17808,N_17525);
nor U18065 (N_18065,N_17750,N_17993);
nand U18066 (N_18066,N_17984,N_17905);
xnor U18067 (N_18067,N_17938,N_17914);
nor U18068 (N_18068,N_17609,N_17569);
nor U18069 (N_18069,N_17708,N_17698);
nand U18070 (N_18070,N_17968,N_17714);
nand U18071 (N_18071,N_17503,N_17979);
nor U18072 (N_18072,N_17618,N_17611);
xnor U18073 (N_18073,N_17595,N_17990);
or U18074 (N_18074,N_17748,N_17857);
nor U18075 (N_18075,N_17925,N_17734);
and U18076 (N_18076,N_17859,N_17790);
and U18077 (N_18077,N_17565,N_17826);
xor U18078 (N_18078,N_17553,N_17930);
nor U18079 (N_18079,N_17970,N_17787);
or U18080 (N_18080,N_17879,N_17874);
nor U18081 (N_18081,N_17598,N_17819);
and U18082 (N_18082,N_17662,N_17636);
xor U18083 (N_18083,N_17891,N_17828);
or U18084 (N_18084,N_17831,N_17843);
xor U18085 (N_18085,N_17585,N_17836);
and U18086 (N_18086,N_17793,N_17780);
and U18087 (N_18087,N_17627,N_17892);
nand U18088 (N_18088,N_17508,N_17512);
nor U18089 (N_18089,N_17730,N_17605);
and U18090 (N_18090,N_17599,N_17792);
nor U18091 (N_18091,N_17501,N_17854);
nor U18092 (N_18092,N_17886,N_17834);
or U18093 (N_18093,N_17707,N_17547);
and U18094 (N_18094,N_17696,N_17528);
and U18095 (N_18095,N_17517,N_17621);
nand U18096 (N_18096,N_17781,N_17578);
and U18097 (N_18097,N_17791,N_17600);
or U18098 (N_18098,N_17514,N_17766);
nand U18099 (N_18099,N_17976,N_17995);
nor U18100 (N_18100,N_17871,N_17718);
and U18101 (N_18101,N_17711,N_17509);
nor U18102 (N_18102,N_17634,N_17798);
nand U18103 (N_18103,N_17589,N_17709);
xnor U18104 (N_18104,N_17692,N_17510);
and U18105 (N_18105,N_17804,N_17911);
and U18106 (N_18106,N_17560,N_17888);
or U18107 (N_18107,N_17638,N_17588);
xnor U18108 (N_18108,N_17811,N_17965);
and U18109 (N_18109,N_17906,N_17593);
nand U18110 (N_18110,N_17717,N_17908);
and U18111 (N_18111,N_17521,N_17749);
and U18112 (N_18112,N_17815,N_17899);
and U18113 (N_18113,N_17702,N_17768);
xor U18114 (N_18114,N_17783,N_17642);
nor U18115 (N_18115,N_17959,N_17812);
or U18116 (N_18116,N_17530,N_17576);
nor U18117 (N_18117,N_17680,N_17903);
or U18118 (N_18118,N_17778,N_17881);
or U18119 (N_18119,N_17684,N_17909);
or U18120 (N_18120,N_17690,N_17629);
and U18121 (N_18121,N_17543,N_17747);
and U18122 (N_18122,N_17570,N_17687);
nor U18123 (N_18123,N_17556,N_17765);
nand U18124 (N_18124,N_17901,N_17643);
nor U18125 (N_18125,N_17763,N_17919);
or U18126 (N_18126,N_17630,N_17941);
and U18127 (N_18127,N_17653,N_17849);
nand U18128 (N_18128,N_17950,N_17628);
xnor U18129 (N_18129,N_17654,N_17992);
xnor U18130 (N_18130,N_17890,N_17732);
xor U18131 (N_18131,N_17655,N_17674);
and U18132 (N_18132,N_17827,N_17870);
nor U18133 (N_18133,N_17975,N_17894);
nor U18134 (N_18134,N_17579,N_17942);
nand U18135 (N_18135,N_17863,N_17962);
nand U18136 (N_18136,N_17809,N_17877);
or U18137 (N_18137,N_17967,N_17797);
xnor U18138 (N_18138,N_17603,N_17728);
or U18139 (N_18139,N_17987,N_17876);
nor U18140 (N_18140,N_17841,N_17694);
or U18141 (N_18141,N_17625,N_17934);
and U18142 (N_18142,N_17733,N_17561);
or U18143 (N_18143,N_17582,N_17816);
or U18144 (N_18144,N_17725,N_17632);
or U18145 (N_18145,N_17907,N_17520);
and U18146 (N_18146,N_17606,N_17800);
or U18147 (N_18147,N_17776,N_17675);
and U18148 (N_18148,N_17855,N_17614);
and U18149 (N_18149,N_17745,N_17552);
or U18150 (N_18150,N_17729,N_17681);
nand U18151 (N_18151,N_17546,N_17704);
nor U18152 (N_18152,N_17640,N_17770);
xnor U18153 (N_18153,N_17991,N_17590);
and U18154 (N_18154,N_17665,N_17577);
and U18155 (N_18155,N_17650,N_17737);
or U18156 (N_18156,N_17515,N_17586);
or U18157 (N_18157,N_17940,N_17865);
and U18158 (N_18158,N_17539,N_17847);
nand U18159 (N_18159,N_17754,N_17573);
xnor U18160 (N_18160,N_17727,N_17511);
nand U18161 (N_18161,N_17833,N_17689);
or U18162 (N_18162,N_17616,N_17821);
nor U18163 (N_18163,N_17761,N_17663);
nand U18164 (N_18164,N_17529,N_17829);
and U18165 (N_18165,N_17883,N_17931);
and U18166 (N_18166,N_17858,N_17527);
and U18167 (N_18167,N_17755,N_17507);
and U18168 (N_18168,N_17571,N_17574);
or U18169 (N_18169,N_17895,N_17752);
nor U18170 (N_18170,N_17756,N_17686);
or U18171 (N_18171,N_17673,N_17505);
or U18172 (N_18172,N_17832,N_17677);
or U18173 (N_18173,N_17540,N_17592);
and U18174 (N_18174,N_17866,N_17700);
and U18175 (N_18175,N_17626,N_17646);
nand U18176 (N_18176,N_17742,N_17980);
nand U18177 (N_18177,N_17830,N_17813);
nor U18178 (N_18178,N_17929,N_17695);
nor U18179 (N_18179,N_17658,N_17839);
nor U18180 (N_18180,N_17722,N_17648);
or U18181 (N_18181,N_17607,N_17913);
nand U18182 (N_18182,N_17619,N_17875);
or U18183 (N_18183,N_17660,N_17985);
and U18184 (N_18184,N_17608,N_17927);
nand U18185 (N_18185,N_17939,N_17807);
nand U18186 (N_18186,N_17519,N_17788);
nor U18187 (N_18187,N_17731,N_17563);
and U18188 (N_18188,N_17583,N_17795);
and U18189 (N_18189,N_17988,N_17701);
nor U18190 (N_18190,N_17610,N_17757);
and U18191 (N_18191,N_17688,N_17822);
or U18192 (N_18192,N_17947,N_17835);
nand U18193 (N_18193,N_17667,N_17724);
nor U18194 (N_18194,N_17946,N_17670);
nand U18195 (N_18195,N_17649,N_17973);
nor U18196 (N_18196,N_17915,N_17591);
xor U18197 (N_18197,N_17542,N_17961);
nand U18198 (N_18198,N_17647,N_17999);
nor U18199 (N_18199,N_17963,N_17697);
nand U18200 (N_18200,N_17916,N_17955);
and U18201 (N_18201,N_17920,N_17893);
xnor U18202 (N_18202,N_17544,N_17693);
and U18203 (N_18203,N_17769,N_17604);
and U18204 (N_18204,N_17824,N_17817);
xnor U18205 (N_18205,N_17964,N_17852);
or U18206 (N_18206,N_17818,N_17678);
nor U18207 (N_18207,N_17524,N_17601);
and U18208 (N_18208,N_17602,N_17846);
nor U18209 (N_18209,N_17949,N_17735);
or U18210 (N_18210,N_17635,N_17723);
or U18211 (N_18211,N_17936,N_17958);
and U18212 (N_18212,N_17972,N_17526);
nor U18213 (N_18213,N_17837,N_17613);
nor U18214 (N_18214,N_17998,N_17620);
xnor U18215 (N_18215,N_17644,N_17844);
xnor U18216 (N_18216,N_17885,N_17713);
xnor U18217 (N_18217,N_17548,N_17641);
nor U18218 (N_18218,N_17842,N_17860);
or U18219 (N_18219,N_17884,N_17873);
or U18220 (N_18220,N_17669,N_17952);
or U18221 (N_18221,N_17820,N_17534);
xnor U18222 (N_18222,N_17796,N_17751);
xor U18223 (N_18223,N_17683,N_17904);
xnor U18224 (N_18224,N_17743,N_17810);
nand U18225 (N_18225,N_17771,N_17652);
nor U18226 (N_18226,N_17932,N_17656);
nand U18227 (N_18227,N_17882,N_17764);
or U18228 (N_18228,N_17716,N_17691);
or U18229 (N_18229,N_17516,N_17502);
nand U18230 (N_18230,N_17557,N_17744);
xor U18231 (N_18231,N_17823,N_17699);
xnor U18232 (N_18232,N_17838,N_17957);
nor U18233 (N_18233,N_17773,N_17676);
xnor U18234 (N_18234,N_17513,N_17889);
nor U18235 (N_18235,N_17994,N_17551);
xnor U18236 (N_18236,N_17960,N_17948);
or U18237 (N_18237,N_17550,N_17558);
xnor U18238 (N_18238,N_17555,N_17584);
nand U18239 (N_18239,N_17537,N_17978);
and U18240 (N_18240,N_17594,N_17897);
nand U18241 (N_18241,N_17850,N_17633);
xnor U18242 (N_18242,N_17799,N_17637);
and U18243 (N_18243,N_17575,N_17712);
nand U18244 (N_18244,N_17753,N_17533);
nor U18245 (N_18245,N_17814,N_17983);
nand U18246 (N_18246,N_17878,N_17845);
xnor U18247 (N_18247,N_17518,N_17784);
xor U18248 (N_18248,N_17679,N_17685);
nand U18249 (N_18249,N_17639,N_17615);
and U18250 (N_18250,N_17992,N_17798);
nand U18251 (N_18251,N_17987,N_17580);
nand U18252 (N_18252,N_17543,N_17590);
xor U18253 (N_18253,N_17970,N_17845);
nor U18254 (N_18254,N_17825,N_17963);
nor U18255 (N_18255,N_17618,N_17632);
nor U18256 (N_18256,N_17759,N_17713);
or U18257 (N_18257,N_17841,N_17822);
and U18258 (N_18258,N_17998,N_17999);
nand U18259 (N_18259,N_17562,N_17880);
and U18260 (N_18260,N_17699,N_17659);
and U18261 (N_18261,N_17623,N_17568);
and U18262 (N_18262,N_17783,N_17865);
or U18263 (N_18263,N_17624,N_17829);
or U18264 (N_18264,N_17845,N_17912);
xnor U18265 (N_18265,N_17503,N_17749);
nand U18266 (N_18266,N_17551,N_17709);
and U18267 (N_18267,N_17785,N_17552);
nor U18268 (N_18268,N_17717,N_17819);
or U18269 (N_18269,N_17636,N_17586);
or U18270 (N_18270,N_17981,N_17886);
nand U18271 (N_18271,N_17507,N_17534);
nand U18272 (N_18272,N_17530,N_17630);
nand U18273 (N_18273,N_17942,N_17618);
and U18274 (N_18274,N_17882,N_17768);
nand U18275 (N_18275,N_17727,N_17933);
nor U18276 (N_18276,N_17830,N_17534);
nor U18277 (N_18277,N_17560,N_17764);
and U18278 (N_18278,N_17578,N_17865);
xor U18279 (N_18279,N_17555,N_17519);
or U18280 (N_18280,N_17738,N_17878);
and U18281 (N_18281,N_17852,N_17739);
nor U18282 (N_18282,N_17579,N_17704);
xor U18283 (N_18283,N_17602,N_17791);
nor U18284 (N_18284,N_17751,N_17560);
and U18285 (N_18285,N_17734,N_17794);
xnor U18286 (N_18286,N_17654,N_17742);
xnor U18287 (N_18287,N_17792,N_17801);
or U18288 (N_18288,N_17725,N_17590);
and U18289 (N_18289,N_17512,N_17789);
and U18290 (N_18290,N_17513,N_17505);
nand U18291 (N_18291,N_17529,N_17699);
and U18292 (N_18292,N_17851,N_17627);
or U18293 (N_18293,N_17801,N_17966);
nand U18294 (N_18294,N_17627,N_17632);
or U18295 (N_18295,N_17922,N_17546);
nand U18296 (N_18296,N_17996,N_17809);
nor U18297 (N_18297,N_17860,N_17895);
or U18298 (N_18298,N_17647,N_17893);
nor U18299 (N_18299,N_17686,N_17511);
nor U18300 (N_18300,N_17846,N_17639);
nand U18301 (N_18301,N_17675,N_17753);
xor U18302 (N_18302,N_17646,N_17589);
nor U18303 (N_18303,N_17630,N_17716);
and U18304 (N_18304,N_17955,N_17908);
and U18305 (N_18305,N_17917,N_17892);
nor U18306 (N_18306,N_17945,N_17697);
nor U18307 (N_18307,N_17986,N_17773);
and U18308 (N_18308,N_17828,N_17571);
or U18309 (N_18309,N_17873,N_17917);
or U18310 (N_18310,N_17914,N_17738);
nor U18311 (N_18311,N_17688,N_17950);
or U18312 (N_18312,N_17841,N_17506);
or U18313 (N_18313,N_17516,N_17912);
or U18314 (N_18314,N_17784,N_17618);
or U18315 (N_18315,N_17540,N_17626);
xnor U18316 (N_18316,N_17884,N_17826);
nor U18317 (N_18317,N_17647,N_17574);
or U18318 (N_18318,N_17695,N_17735);
and U18319 (N_18319,N_17777,N_17858);
nand U18320 (N_18320,N_17758,N_17703);
or U18321 (N_18321,N_17592,N_17926);
xor U18322 (N_18322,N_17602,N_17954);
nand U18323 (N_18323,N_17596,N_17831);
and U18324 (N_18324,N_17766,N_17871);
nand U18325 (N_18325,N_17827,N_17964);
or U18326 (N_18326,N_17717,N_17656);
nor U18327 (N_18327,N_17958,N_17802);
and U18328 (N_18328,N_17607,N_17825);
xor U18329 (N_18329,N_17944,N_17789);
xor U18330 (N_18330,N_17775,N_17743);
nor U18331 (N_18331,N_17760,N_17763);
and U18332 (N_18332,N_17917,N_17935);
nand U18333 (N_18333,N_17831,N_17836);
xnor U18334 (N_18334,N_17666,N_17613);
and U18335 (N_18335,N_17998,N_17793);
nor U18336 (N_18336,N_17501,N_17938);
or U18337 (N_18337,N_17640,N_17768);
nor U18338 (N_18338,N_17552,N_17831);
or U18339 (N_18339,N_17980,N_17967);
xor U18340 (N_18340,N_17881,N_17949);
nand U18341 (N_18341,N_17505,N_17599);
xor U18342 (N_18342,N_17937,N_17563);
or U18343 (N_18343,N_17529,N_17592);
nor U18344 (N_18344,N_17666,N_17929);
nor U18345 (N_18345,N_17519,N_17923);
nor U18346 (N_18346,N_17801,N_17530);
nand U18347 (N_18347,N_17673,N_17899);
and U18348 (N_18348,N_17900,N_17871);
nand U18349 (N_18349,N_17928,N_17644);
xnor U18350 (N_18350,N_17982,N_17967);
xor U18351 (N_18351,N_17895,N_17882);
or U18352 (N_18352,N_17987,N_17815);
nor U18353 (N_18353,N_17628,N_17838);
nand U18354 (N_18354,N_17842,N_17754);
nand U18355 (N_18355,N_17868,N_17774);
xnor U18356 (N_18356,N_17739,N_17835);
nor U18357 (N_18357,N_17810,N_17612);
or U18358 (N_18358,N_17973,N_17709);
nand U18359 (N_18359,N_17945,N_17765);
xnor U18360 (N_18360,N_17569,N_17781);
nor U18361 (N_18361,N_17801,N_17953);
xnor U18362 (N_18362,N_17533,N_17784);
or U18363 (N_18363,N_17980,N_17554);
and U18364 (N_18364,N_17722,N_17742);
xor U18365 (N_18365,N_17996,N_17729);
and U18366 (N_18366,N_17918,N_17905);
nand U18367 (N_18367,N_17615,N_17626);
nor U18368 (N_18368,N_17818,N_17795);
nor U18369 (N_18369,N_17601,N_17549);
nor U18370 (N_18370,N_17567,N_17802);
xor U18371 (N_18371,N_17650,N_17877);
nor U18372 (N_18372,N_17900,N_17760);
and U18373 (N_18373,N_17541,N_17522);
nand U18374 (N_18374,N_17985,N_17796);
and U18375 (N_18375,N_17762,N_17893);
or U18376 (N_18376,N_17743,N_17698);
xor U18377 (N_18377,N_17588,N_17535);
and U18378 (N_18378,N_17784,N_17603);
xor U18379 (N_18379,N_17842,N_17644);
nor U18380 (N_18380,N_17949,N_17998);
nand U18381 (N_18381,N_17901,N_17626);
and U18382 (N_18382,N_17515,N_17743);
and U18383 (N_18383,N_17688,N_17860);
nor U18384 (N_18384,N_17812,N_17612);
nor U18385 (N_18385,N_17750,N_17858);
and U18386 (N_18386,N_17666,N_17622);
nor U18387 (N_18387,N_17903,N_17936);
nand U18388 (N_18388,N_17575,N_17682);
nor U18389 (N_18389,N_17516,N_17603);
nand U18390 (N_18390,N_17769,N_17818);
nor U18391 (N_18391,N_17716,N_17898);
nand U18392 (N_18392,N_17588,N_17751);
nor U18393 (N_18393,N_17512,N_17923);
nand U18394 (N_18394,N_17511,N_17638);
or U18395 (N_18395,N_17866,N_17709);
nor U18396 (N_18396,N_17778,N_17858);
xnor U18397 (N_18397,N_17752,N_17509);
xor U18398 (N_18398,N_17700,N_17675);
nand U18399 (N_18399,N_17879,N_17793);
and U18400 (N_18400,N_17778,N_17542);
nand U18401 (N_18401,N_17936,N_17715);
and U18402 (N_18402,N_17728,N_17901);
nand U18403 (N_18403,N_17552,N_17592);
and U18404 (N_18404,N_17588,N_17571);
nand U18405 (N_18405,N_17999,N_17644);
nor U18406 (N_18406,N_17653,N_17804);
xor U18407 (N_18407,N_17618,N_17762);
and U18408 (N_18408,N_17941,N_17512);
and U18409 (N_18409,N_17500,N_17992);
and U18410 (N_18410,N_17653,N_17954);
xor U18411 (N_18411,N_17585,N_17876);
or U18412 (N_18412,N_17823,N_17946);
nor U18413 (N_18413,N_17698,N_17506);
and U18414 (N_18414,N_17823,N_17884);
and U18415 (N_18415,N_17847,N_17684);
nor U18416 (N_18416,N_17719,N_17715);
xnor U18417 (N_18417,N_17879,N_17736);
or U18418 (N_18418,N_17736,N_17552);
nor U18419 (N_18419,N_17616,N_17702);
nand U18420 (N_18420,N_17898,N_17557);
or U18421 (N_18421,N_17500,N_17599);
and U18422 (N_18422,N_17808,N_17905);
and U18423 (N_18423,N_17715,N_17836);
or U18424 (N_18424,N_17957,N_17913);
nand U18425 (N_18425,N_17832,N_17930);
nand U18426 (N_18426,N_17688,N_17596);
xor U18427 (N_18427,N_17563,N_17670);
nor U18428 (N_18428,N_17603,N_17670);
xnor U18429 (N_18429,N_17555,N_17903);
xor U18430 (N_18430,N_17576,N_17572);
xnor U18431 (N_18431,N_17649,N_17645);
and U18432 (N_18432,N_17970,N_17527);
nand U18433 (N_18433,N_17982,N_17851);
nand U18434 (N_18434,N_17964,N_17925);
xor U18435 (N_18435,N_17693,N_17530);
or U18436 (N_18436,N_17957,N_17963);
or U18437 (N_18437,N_17565,N_17802);
nand U18438 (N_18438,N_17635,N_17772);
nor U18439 (N_18439,N_17548,N_17672);
nand U18440 (N_18440,N_17701,N_17706);
and U18441 (N_18441,N_17982,N_17703);
and U18442 (N_18442,N_17869,N_17579);
xor U18443 (N_18443,N_17690,N_17969);
and U18444 (N_18444,N_17786,N_17920);
or U18445 (N_18445,N_17544,N_17870);
or U18446 (N_18446,N_17815,N_17567);
nor U18447 (N_18447,N_17505,N_17869);
or U18448 (N_18448,N_17972,N_17520);
and U18449 (N_18449,N_17633,N_17687);
nor U18450 (N_18450,N_17938,N_17580);
xnor U18451 (N_18451,N_17537,N_17797);
xor U18452 (N_18452,N_17738,N_17908);
xor U18453 (N_18453,N_17983,N_17637);
nand U18454 (N_18454,N_17964,N_17889);
xnor U18455 (N_18455,N_17970,N_17546);
xnor U18456 (N_18456,N_17653,N_17711);
and U18457 (N_18457,N_17836,N_17706);
xnor U18458 (N_18458,N_17708,N_17926);
nor U18459 (N_18459,N_17949,N_17786);
or U18460 (N_18460,N_17550,N_17511);
nand U18461 (N_18461,N_17772,N_17599);
xnor U18462 (N_18462,N_17712,N_17759);
nor U18463 (N_18463,N_17552,N_17990);
nor U18464 (N_18464,N_17727,N_17741);
or U18465 (N_18465,N_17738,N_17744);
nand U18466 (N_18466,N_17713,N_17526);
or U18467 (N_18467,N_17997,N_17520);
xor U18468 (N_18468,N_17787,N_17541);
or U18469 (N_18469,N_17941,N_17905);
and U18470 (N_18470,N_17805,N_17575);
nor U18471 (N_18471,N_17751,N_17625);
xor U18472 (N_18472,N_17999,N_17560);
or U18473 (N_18473,N_17977,N_17809);
or U18474 (N_18474,N_17933,N_17576);
nand U18475 (N_18475,N_17756,N_17500);
or U18476 (N_18476,N_17589,N_17910);
nand U18477 (N_18477,N_17655,N_17965);
nand U18478 (N_18478,N_17679,N_17853);
or U18479 (N_18479,N_17778,N_17530);
nand U18480 (N_18480,N_17615,N_17876);
or U18481 (N_18481,N_17846,N_17890);
xnor U18482 (N_18482,N_17598,N_17934);
and U18483 (N_18483,N_17980,N_17513);
and U18484 (N_18484,N_17941,N_17835);
nor U18485 (N_18485,N_17724,N_17651);
nor U18486 (N_18486,N_17750,N_17606);
nor U18487 (N_18487,N_17713,N_17529);
nor U18488 (N_18488,N_17614,N_17544);
nand U18489 (N_18489,N_17884,N_17854);
nor U18490 (N_18490,N_17540,N_17650);
nor U18491 (N_18491,N_17598,N_17809);
xnor U18492 (N_18492,N_17608,N_17514);
xnor U18493 (N_18493,N_17765,N_17710);
and U18494 (N_18494,N_17850,N_17687);
nand U18495 (N_18495,N_17908,N_17684);
nand U18496 (N_18496,N_17714,N_17845);
and U18497 (N_18497,N_17932,N_17769);
xor U18498 (N_18498,N_17974,N_17932);
nand U18499 (N_18499,N_17963,N_17749);
or U18500 (N_18500,N_18203,N_18293);
nand U18501 (N_18501,N_18346,N_18042);
nand U18502 (N_18502,N_18123,N_18000);
nor U18503 (N_18503,N_18381,N_18159);
nor U18504 (N_18504,N_18330,N_18396);
and U18505 (N_18505,N_18039,N_18269);
xnor U18506 (N_18506,N_18325,N_18079);
and U18507 (N_18507,N_18316,N_18250);
nand U18508 (N_18508,N_18288,N_18152);
xnor U18509 (N_18509,N_18291,N_18485);
nor U18510 (N_18510,N_18317,N_18248);
and U18511 (N_18511,N_18292,N_18138);
or U18512 (N_18512,N_18400,N_18412);
nor U18513 (N_18513,N_18340,N_18442);
or U18514 (N_18514,N_18484,N_18481);
or U18515 (N_18515,N_18385,N_18022);
xor U18516 (N_18516,N_18093,N_18480);
nor U18517 (N_18517,N_18488,N_18231);
xor U18518 (N_18518,N_18222,N_18227);
or U18519 (N_18519,N_18208,N_18109);
nor U18520 (N_18520,N_18175,N_18472);
and U18521 (N_18521,N_18041,N_18082);
or U18522 (N_18522,N_18392,N_18032);
xnor U18523 (N_18523,N_18394,N_18212);
nand U18524 (N_18524,N_18029,N_18280);
nor U18525 (N_18525,N_18310,N_18060);
nand U18526 (N_18526,N_18077,N_18170);
and U18527 (N_18527,N_18444,N_18278);
nand U18528 (N_18528,N_18424,N_18476);
nand U18529 (N_18529,N_18219,N_18393);
and U18530 (N_18530,N_18179,N_18213);
nand U18531 (N_18531,N_18184,N_18339);
and U18532 (N_18532,N_18144,N_18015);
nor U18533 (N_18533,N_18117,N_18019);
xor U18534 (N_18534,N_18130,N_18341);
nor U18535 (N_18535,N_18220,N_18369);
or U18536 (N_18536,N_18475,N_18191);
xnor U18537 (N_18537,N_18398,N_18092);
or U18538 (N_18538,N_18173,N_18364);
or U18539 (N_18539,N_18172,N_18196);
nand U18540 (N_18540,N_18482,N_18195);
nand U18541 (N_18541,N_18490,N_18096);
and U18542 (N_18542,N_18282,N_18380);
and U18543 (N_18543,N_18433,N_18439);
nand U18544 (N_18544,N_18132,N_18397);
and U18545 (N_18545,N_18352,N_18056);
nor U18546 (N_18546,N_18463,N_18496);
or U18547 (N_18547,N_18379,N_18333);
or U18548 (N_18548,N_18306,N_18491);
and U18549 (N_18549,N_18266,N_18337);
nand U18550 (N_18550,N_18118,N_18073);
nor U18551 (N_18551,N_18155,N_18441);
nand U18552 (N_18552,N_18414,N_18285);
nor U18553 (N_18553,N_18356,N_18299);
nand U18554 (N_18554,N_18202,N_18225);
nand U18555 (N_18555,N_18462,N_18419);
or U18556 (N_18556,N_18193,N_18359);
xor U18557 (N_18557,N_18483,N_18094);
or U18558 (N_18558,N_18067,N_18065);
nor U18559 (N_18559,N_18189,N_18169);
xnor U18560 (N_18560,N_18251,N_18028);
nor U18561 (N_18561,N_18199,N_18088);
xnor U18562 (N_18562,N_18435,N_18160);
xor U18563 (N_18563,N_18360,N_18154);
xor U18564 (N_18564,N_18343,N_18497);
nor U18565 (N_18565,N_18162,N_18194);
xnor U18566 (N_18566,N_18102,N_18091);
or U18567 (N_18567,N_18304,N_18402);
xnor U18568 (N_18568,N_18149,N_18489);
nor U18569 (N_18569,N_18236,N_18426);
nand U18570 (N_18570,N_18284,N_18427);
xor U18571 (N_18571,N_18027,N_18300);
nor U18572 (N_18572,N_18420,N_18072);
nor U18573 (N_18573,N_18009,N_18336);
nand U18574 (N_18574,N_18318,N_18217);
or U18575 (N_18575,N_18097,N_18002);
nand U18576 (N_18576,N_18124,N_18085);
and U18577 (N_18577,N_18302,N_18180);
nand U18578 (N_18578,N_18295,N_18033);
or U18579 (N_18579,N_18450,N_18487);
and U18580 (N_18580,N_18105,N_18255);
nand U18581 (N_18581,N_18366,N_18034);
nand U18582 (N_18582,N_18062,N_18467);
xor U18583 (N_18583,N_18148,N_18498);
nand U18584 (N_18584,N_18466,N_18301);
nand U18585 (N_18585,N_18493,N_18186);
nor U18586 (N_18586,N_18286,N_18342);
nand U18587 (N_18587,N_18246,N_18205);
and U18588 (N_18588,N_18038,N_18308);
nor U18589 (N_18589,N_18030,N_18329);
and U18590 (N_18590,N_18108,N_18014);
nor U18591 (N_18591,N_18171,N_18233);
or U18592 (N_18592,N_18358,N_18110);
and U18593 (N_18593,N_18270,N_18389);
nor U18594 (N_18594,N_18103,N_18201);
nand U18595 (N_18595,N_18150,N_18206);
nand U18596 (N_18596,N_18378,N_18281);
nand U18597 (N_18597,N_18064,N_18406);
or U18598 (N_18598,N_18001,N_18074);
or U18599 (N_18599,N_18120,N_18178);
xor U18600 (N_18600,N_18459,N_18182);
and U18601 (N_18601,N_18020,N_18021);
nand U18602 (N_18602,N_18320,N_18263);
nor U18603 (N_18603,N_18418,N_18101);
nand U18604 (N_18604,N_18107,N_18361);
or U18605 (N_18605,N_18070,N_18478);
nor U18606 (N_18606,N_18239,N_18265);
and U18607 (N_18607,N_18053,N_18164);
nand U18608 (N_18608,N_18453,N_18407);
nand U18609 (N_18609,N_18290,N_18046);
nor U18610 (N_18610,N_18188,N_18365);
nand U18611 (N_18611,N_18113,N_18455);
xor U18612 (N_18612,N_18387,N_18115);
or U18613 (N_18613,N_18452,N_18430);
nor U18614 (N_18614,N_18362,N_18058);
or U18615 (N_18615,N_18357,N_18447);
nand U18616 (N_18616,N_18013,N_18422);
nand U18617 (N_18617,N_18198,N_18168);
nand U18618 (N_18618,N_18440,N_18456);
and U18619 (N_18619,N_18071,N_18176);
nand U18620 (N_18620,N_18134,N_18061);
or U18621 (N_18621,N_18309,N_18068);
and U18622 (N_18622,N_18436,N_18312);
nand U18623 (N_18623,N_18431,N_18147);
and U18624 (N_18624,N_18279,N_18460);
xor U18625 (N_18625,N_18119,N_18010);
nand U18626 (N_18626,N_18273,N_18374);
xnor U18627 (N_18627,N_18238,N_18017);
or U18628 (N_18628,N_18264,N_18298);
nor U18629 (N_18629,N_18363,N_18232);
and U18630 (N_18630,N_18289,N_18224);
nor U18631 (N_18631,N_18388,N_18495);
nor U18632 (N_18632,N_18126,N_18045);
and U18633 (N_18633,N_18187,N_18221);
or U18634 (N_18634,N_18214,N_18040);
nor U18635 (N_18635,N_18458,N_18207);
nand U18636 (N_18636,N_18350,N_18127);
nor U18637 (N_18637,N_18051,N_18276);
xnor U18638 (N_18638,N_18345,N_18254);
nor U18639 (N_18639,N_18125,N_18272);
nand U18640 (N_18640,N_18237,N_18128);
nor U18641 (N_18641,N_18114,N_18314);
nor U18642 (N_18642,N_18408,N_18142);
nor U18643 (N_18643,N_18474,N_18145);
or U18644 (N_18644,N_18401,N_18376);
nor U18645 (N_18645,N_18087,N_18355);
or U18646 (N_18646,N_18253,N_18080);
and U18647 (N_18647,N_18100,N_18157);
and U18648 (N_18648,N_18226,N_18410);
xor U18649 (N_18649,N_18016,N_18216);
or U18650 (N_18650,N_18141,N_18283);
or U18651 (N_18651,N_18025,N_18185);
nand U18652 (N_18652,N_18434,N_18098);
and U18653 (N_18653,N_18090,N_18287);
nand U18654 (N_18654,N_18005,N_18242);
nand U18655 (N_18655,N_18303,N_18031);
and U18656 (N_18656,N_18209,N_18143);
nand U18657 (N_18657,N_18139,N_18305);
nand U18658 (N_18658,N_18324,N_18008);
nor U18659 (N_18659,N_18499,N_18262);
and U18660 (N_18660,N_18129,N_18492);
nor U18661 (N_18661,N_18059,N_18006);
xnor U18662 (N_18662,N_18177,N_18111);
or U18663 (N_18663,N_18390,N_18370);
or U18664 (N_18664,N_18259,N_18223);
or U18665 (N_18665,N_18421,N_18156);
nor U18666 (N_18666,N_18112,N_18383);
nor U18667 (N_18667,N_18234,N_18327);
nor U18668 (N_18668,N_18428,N_18099);
and U18669 (N_18669,N_18146,N_18464);
nor U18670 (N_18670,N_18294,N_18247);
nor U18671 (N_18671,N_18122,N_18245);
nor U18672 (N_18672,N_18136,N_18454);
xnor U18673 (N_18673,N_18399,N_18438);
xnor U18674 (N_18674,N_18429,N_18026);
nor U18675 (N_18675,N_18047,N_18083);
or U18676 (N_18676,N_18432,N_18465);
or U18677 (N_18677,N_18267,N_18161);
nand U18678 (N_18678,N_18004,N_18057);
xor U18679 (N_18679,N_18190,N_18448);
nor U18680 (N_18680,N_18384,N_18081);
xnor U18681 (N_18681,N_18228,N_18425);
nor U18682 (N_18682,N_18382,N_18354);
xnor U18683 (N_18683,N_18271,N_18084);
nand U18684 (N_18684,N_18174,N_18257);
or U18685 (N_18685,N_18323,N_18415);
xnor U18686 (N_18686,N_18375,N_18151);
and U18687 (N_18687,N_18275,N_18069);
and U18688 (N_18688,N_18104,N_18446);
or U18689 (N_18689,N_18048,N_18411);
nand U18690 (N_18690,N_18307,N_18181);
nor U18691 (N_18691,N_18078,N_18066);
xnor U18692 (N_18692,N_18243,N_18404);
nand U18693 (N_18693,N_18121,N_18249);
nand U18694 (N_18694,N_18166,N_18328);
and U18695 (N_18695,N_18391,N_18277);
or U18696 (N_18696,N_18461,N_18252);
nor U18697 (N_18697,N_18204,N_18260);
xor U18698 (N_18698,N_18377,N_18055);
nor U18699 (N_18699,N_18197,N_18200);
nor U18700 (N_18700,N_18445,N_18043);
xnor U18701 (N_18701,N_18274,N_18256);
nand U18702 (N_18702,N_18235,N_18348);
or U18703 (N_18703,N_18437,N_18486);
nor U18704 (N_18704,N_18367,N_18024);
or U18705 (N_18705,N_18395,N_18417);
and U18706 (N_18706,N_18296,N_18211);
or U18707 (N_18707,N_18332,N_18443);
nor U18708 (N_18708,N_18137,N_18268);
and U18709 (N_18709,N_18371,N_18063);
and U18710 (N_18710,N_18322,N_18106);
and U18711 (N_18711,N_18229,N_18409);
nand U18712 (N_18712,N_18405,N_18403);
xor U18713 (N_18713,N_18075,N_18368);
nor U18714 (N_18714,N_18326,N_18479);
nand U18715 (N_18715,N_18449,N_18192);
or U18716 (N_18716,N_18076,N_18473);
xor U18717 (N_18717,N_18469,N_18230);
nand U18718 (N_18718,N_18319,N_18135);
and U18719 (N_18719,N_18315,N_18133);
nand U18720 (N_18720,N_18095,N_18331);
or U18721 (N_18721,N_18037,N_18468);
nand U18722 (N_18722,N_18011,N_18451);
and U18723 (N_18723,N_18086,N_18241);
nand U18724 (N_18724,N_18258,N_18153);
xor U18725 (N_18725,N_18423,N_18494);
and U18726 (N_18726,N_18210,N_18089);
nand U18727 (N_18727,N_18353,N_18334);
xnor U18728 (N_18728,N_18018,N_18052);
xnor U18729 (N_18729,N_18165,N_18050);
nor U18730 (N_18730,N_18471,N_18244);
xnor U18731 (N_18731,N_18140,N_18416);
and U18732 (N_18732,N_18311,N_18373);
or U18733 (N_18733,N_18351,N_18344);
or U18734 (N_18734,N_18321,N_18240);
nor U18735 (N_18735,N_18347,N_18477);
xnor U18736 (N_18736,N_18012,N_18215);
xor U18737 (N_18737,N_18413,N_18054);
xnor U18738 (N_18738,N_18163,N_18297);
and U18739 (N_18739,N_18035,N_18044);
nor U18740 (N_18740,N_18003,N_18313);
nand U18741 (N_18741,N_18049,N_18036);
xnor U18742 (N_18742,N_18335,N_18386);
and U18743 (N_18743,N_18007,N_18183);
and U18744 (N_18744,N_18349,N_18470);
xor U18745 (N_18745,N_18457,N_18023);
xnor U18746 (N_18746,N_18261,N_18338);
nand U18747 (N_18747,N_18218,N_18131);
nor U18748 (N_18748,N_18116,N_18167);
or U18749 (N_18749,N_18372,N_18158);
nand U18750 (N_18750,N_18334,N_18287);
nor U18751 (N_18751,N_18030,N_18125);
nand U18752 (N_18752,N_18384,N_18284);
or U18753 (N_18753,N_18310,N_18334);
nor U18754 (N_18754,N_18131,N_18280);
nor U18755 (N_18755,N_18034,N_18275);
nand U18756 (N_18756,N_18237,N_18477);
or U18757 (N_18757,N_18391,N_18025);
and U18758 (N_18758,N_18121,N_18107);
nor U18759 (N_18759,N_18264,N_18054);
nand U18760 (N_18760,N_18148,N_18497);
xor U18761 (N_18761,N_18411,N_18011);
and U18762 (N_18762,N_18400,N_18358);
xor U18763 (N_18763,N_18494,N_18276);
or U18764 (N_18764,N_18307,N_18140);
xnor U18765 (N_18765,N_18049,N_18168);
or U18766 (N_18766,N_18485,N_18064);
and U18767 (N_18767,N_18426,N_18198);
nor U18768 (N_18768,N_18023,N_18384);
or U18769 (N_18769,N_18098,N_18322);
or U18770 (N_18770,N_18252,N_18023);
xor U18771 (N_18771,N_18172,N_18408);
nor U18772 (N_18772,N_18044,N_18407);
nor U18773 (N_18773,N_18230,N_18074);
nor U18774 (N_18774,N_18095,N_18343);
xor U18775 (N_18775,N_18154,N_18123);
or U18776 (N_18776,N_18132,N_18066);
nor U18777 (N_18777,N_18165,N_18016);
nand U18778 (N_18778,N_18264,N_18021);
nor U18779 (N_18779,N_18385,N_18175);
and U18780 (N_18780,N_18161,N_18186);
or U18781 (N_18781,N_18191,N_18432);
or U18782 (N_18782,N_18453,N_18141);
and U18783 (N_18783,N_18264,N_18491);
and U18784 (N_18784,N_18244,N_18047);
xnor U18785 (N_18785,N_18450,N_18384);
xor U18786 (N_18786,N_18392,N_18093);
xor U18787 (N_18787,N_18029,N_18208);
or U18788 (N_18788,N_18447,N_18378);
nor U18789 (N_18789,N_18165,N_18142);
nor U18790 (N_18790,N_18395,N_18029);
nand U18791 (N_18791,N_18071,N_18416);
or U18792 (N_18792,N_18009,N_18392);
nor U18793 (N_18793,N_18442,N_18322);
xor U18794 (N_18794,N_18404,N_18110);
and U18795 (N_18795,N_18462,N_18069);
or U18796 (N_18796,N_18172,N_18185);
xnor U18797 (N_18797,N_18406,N_18272);
or U18798 (N_18798,N_18131,N_18378);
or U18799 (N_18799,N_18348,N_18046);
xnor U18800 (N_18800,N_18434,N_18092);
or U18801 (N_18801,N_18268,N_18041);
and U18802 (N_18802,N_18150,N_18090);
nor U18803 (N_18803,N_18241,N_18427);
and U18804 (N_18804,N_18342,N_18150);
nand U18805 (N_18805,N_18203,N_18452);
nand U18806 (N_18806,N_18481,N_18299);
xor U18807 (N_18807,N_18313,N_18280);
and U18808 (N_18808,N_18457,N_18434);
or U18809 (N_18809,N_18335,N_18189);
or U18810 (N_18810,N_18192,N_18174);
nor U18811 (N_18811,N_18415,N_18230);
or U18812 (N_18812,N_18347,N_18471);
and U18813 (N_18813,N_18426,N_18154);
xnor U18814 (N_18814,N_18169,N_18454);
or U18815 (N_18815,N_18217,N_18160);
xnor U18816 (N_18816,N_18046,N_18335);
nor U18817 (N_18817,N_18073,N_18371);
and U18818 (N_18818,N_18114,N_18304);
and U18819 (N_18819,N_18082,N_18287);
or U18820 (N_18820,N_18196,N_18324);
or U18821 (N_18821,N_18422,N_18369);
and U18822 (N_18822,N_18430,N_18345);
nand U18823 (N_18823,N_18468,N_18493);
xor U18824 (N_18824,N_18306,N_18348);
xor U18825 (N_18825,N_18133,N_18307);
and U18826 (N_18826,N_18384,N_18427);
xnor U18827 (N_18827,N_18460,N_18065);
and U18828 (N_18828,N_18024,N_18123);
xor U18829 (N_18829,N_18347,N_18089);
xnor U18830 (N_18830,N_18169,N_18363);
nor U18831 (N_18831,N_18085,N_18133);
or U18832 (N_18832,N_18108,N_18200);
nor U18833 (N_18833,N_18439,N_18362);
xor U18834 (N_18834,N_18093,N_18098);
xor U18835 (N_18835,N_18365,N_18189);
and U18836 (N_18836,N_18436,N_18090);
or U18837 (N_18837,N_18223,N_18315);
nand U18838 (N_18838,N_18224,N_18013);
nand U18839 (N_18839,N_18288,N_18257);
nand U18840 (N_18840,N_18036,N_18155);
nor U18841 (N_18841,N_18074,N_18136);
and U18842 (N_18842,N_18032,N_18147);
xnor U18843 (N_18843,N_18291,N_18306);
nor U18844 (N_18844,N_18197,N_18489);
xor U18845 (N_18845,N_18217,N_18149);
and U18846 (N_18846,N_18280,N_18045);
xor U18847 (N_18847,N_18017,N_18204);
xor U18848 (N_18848,N_18451,N_18192);
and U18849 (N_18849,N_18327,N_18232);
nand U18850 (N_18850,N_18414,N_18077);
xor U18851 (N_18851,N_18234,N_18024);
or U18852 (N_18852,N_18271,N_18225);
xor U18853 (N_18853,N_18027,N_18230);
nor U18854 (N_18854,N_18480,N_18149);
and U18855 (N_18855,N_18271,N_18379);
or U18856 (N_18856,N_18033,N_18281);
nor U18857 (N_18857,N_18272,N_18296);
nand U18858 (N_18858,N_18219,N_18489);
and U18859 (N_18859,N_18165,N_18014);
nand U18860 (N_18860,N_18230,N_18499);
xor U18861 (N_18861,N_18423,N_18386);
xor U18862 (N_18862,N_18469,N_18347);
xor U18863 (N_18863,N_18450,N_18470);
and U18864 (N_18864,N_18079,N_18033);
nand U18865 (N_18865,N_18237,N_18103);
nand U18866 (N_18866,N_18138,N_18476);
and U18867 (N_18867,N_18140,N_18057);
or U18868 (N_18868,N_18364,N_18358);
xnor U18869 (N_18869,N_18391,N_18394);
nand U18870 (N_18870,N_18373,N_18029);
or U18871 (N_18871,N_18087,N_18222);
nand U18872 (N_18872,N_18476,N_18245);
xor U18873 (N_18873,N_18328,N_18460);
xnor U18874 (N_18874,N_18139,N_18019);
or U18875 (N_18875,N_18072,N_18241);
nor U18876 (N_18876,N_18044,N_18074);
nor U18877 (N_18877,N_18240,N_18257);
or U18878 (N_18878,N_18148,N_18151);
and U18879 (N_18879,N_18396,N_18233);
or U18880 (N_18880,N_18159,N_18181);
nand U18881 (N_18881,N_18381,N_18141);
nand U18882 (N_18882,N_18048,N_18085);
and U18883 (N_18883,N_18446,N_18058);
or U18884 (N_18884,N_18317,N_18398);
xnor U18885 (N_18885,N_18123,N_18404);
nor U18886 (N_18886,N_18110,N_18478);
and U18887 (N_18887,N_18179,N_18474);
or U18888 (N_18888,N_18011,N_18223);
nor U18889 (N_18889,N_18101,N_18293);
nor U18890 (N_18890,N_18227,N_18018);
nand U18891 (N_18891,N_18177,N_18124);
xnor U18892 (N_18892,N_18172,N_18049);
xor U18893 (N_18893,N_18011,N_18445);
nand U18894 (N_18894,N_18180,N_18084);
nor U18895 (N_18895,N_18356,N_18130);
nand U18896 (N_18896,N_18456,N_18291);
or U18897 (N_18897,N_18353,N_18354);
nand U18898 (N_18898,N_18002,N_18283);
or U18899 (N_18899,N_18334,N_18494);
or U18900 (N_18900,N_18072,N_18463);
or U18901 (N_18901,N_18292,N_18350);
nand U18902 (N_18902,N_18437,N_18326);
nand U18903 (N_18903,N_18332,N_18005);
or U18904 (N_18904,N_18268,N_18465);
or U18905 (N_18905,N_18330,N_18300);
and U18906 (N_18906,N_18093,N_18194);
nand U18907 (N_18907,N_18348,N_18372);
nand U18908 (N_18908,N_18095,N_18315);
nor U18909 (N_18909,N_18216,N_18393);
nand U18910 (N_18910,N_18366,N_18057);
nor U18911 (N_18911,N_18167,N_18293);
nand U18912 (N_18912,N_18457,N_18482);
or U18913 (N_18913,N_18228,N_18033);
and U18914 (N_18914,N_18409,N_18155);
xnor U18915 (N_18915,N_18420,N_18101);
nor U18916 (N_18916,N_18246,N_18338);
and U18917 (N_18917,N_18470,N_18334);
or U18918 (N_18918,N_18199,N_18363);
xnor U18919 (N_18919,N_18284,N_18394);
xor U18920 (N_18920,N_18187,N_18155);
nor U18921 (N_18921,N_18013,N_18360);
and U18922 (N_18922,N_18166,N_18401);
and U18923 (N_18923,N_18199,N_18237);
xnor U18924 (N_18924,N_18421,N_18093);
and U18925 (N_18925,N_18084,N_18164);
nand U18926 (N_18926,N_18410,N_18181);
and U18927 (N_18927,N_18131,N_18335);
nand U18928 (N_18928,N_18163,N_18427);
or U18929 (N_18929,N_18345,N_18049);
or U18930 (N_18930,N_18240,N_18295);
xor U18931 (N_18931,N_18171,N_18372);
or U18932 (N_18932,N_18434,N_18367);
nor U18933 (N_18933,N_18184,N_18418);
nor U18934 (N_18934,N_18175,N_18310);
nor U18935 (N_18935,N_18048,N_18045);
or U18936 (N_18936,N_18359,N_18316);
and U18937 (N_18937,N_18065,N_18263);
xor U18938 (N_18938,N_18229,N_18319);
nor U18939 (N_18939,N_18370,N_18019);
and U18940 (N_18940,N_18284,N_18383);
xnor U18941 (N_18941,N_18138,N_18028);
nor U18942 (N_18942,N_18456,N_18299);
xor U18943 (N_18943,N_18192,N_18407);
and U18944 (N_18944,N_18426,N_18064);
nor U18945 (N_18945,N_18168,N_18316);
and U18946 (N_18946,N_18484,N_18406);
and U18947 (N_18947,N_18345,N_18499);
nand U18948 (N_18948,N_18451,N_18447);
nor U18949 (N_18949,N_18097,N_18199);
and U18950 (N_18950,N_18119,N_18409);
nor U18951 (N_18951,N_18279,N_18168);
or U18952 (N_18952,N_18052,N_18458);
nor U18953 (N_18953,N_18118,N_18361);
or U18954 (N_18954,N_18031,N_18014);
nor U18955 (N_18955,N_18242,N_18493);
nand U18956 (N_18956,N_18129,N_18466);
nor U18957 (N_18957,N_18136,N_18093);
nor U18958 (N_18958,N_18251,N_18279);
nor U18959 (N_18959,N_18457,N_18419);
or U18960 (N_18960,N_18163,N_18251);
nand U18961 (N_18961,N_18110,N_18067);
and U18962 (N_18962,N_18434,N_18233);
and U18963 (N_18963,N_18122,N_18391);
nor U18964 (N_18964,N_18286,N_18133);
or U18965 (N_18965,N_18136,N_18440);
nor U18966 (N_18966,N_18238,N_18485);
or U18967 (N_18967,N_18306,N_18213);
nand U18968 (N_18968,N_18325,N_18036);
or U18969 (N_18969,N_18378,N_18082);
xnor U18970 (N_18970,N_18279,N_18050);
and U18971 (N_18971,N_18291,N_18261);
nand U18972 (N_18972,N_18075,N_18432);
nor U18973 (N_18973,N_18496,N_18016);
xor U18974 (N_18974,N_18357,N_18235);
xor U18975 (N_18975,N_18414,N_18452);
xnor U18976 (N_18976,N_18455,N_18243);
nor U18977 (N_18977,N_18105,N_18224);
and U18978 (N_18978,N_18499,N_18294);
and U18979 (N_18979,N_18169,N_18031);
nand U18980 (N_18980,N_18266,N_18200);
nor U18981 (N_18981,N_18308,N_18263);
nand U18982 (N_18982,N_18140,N_18188);
or U18983 (N_18983,N_18322,N_18423);
nand U18984 (N_18984,N_18034,N_18193);
or U18985 (N_18985,N_18171,N_18157);
nand U18986 (N_18986,N_18210,N_18363);
and U18987 (N_18987,N_18253,N_18284);
nand U18988 (N_18988,N_18126,N_18079);
nand U18989 (N_18989,N_18203,N_18232);
or U18990 (N_18990,N_18044,N_18203);
and U18991 (N_18991,N_18491,N_18131);
and U18992 (N_18992,N_18045,N_18057);
or U18993 (N_18993,N_18434,N_18149);
or U18994 (N_18994,N_18442,N_18160);
nor U18995 (N_18995,N_18294,N_18311);
or U18996 (N_18996,N_18395,N_18447);
nand U18997 (N_18997,N_18137,N_18379);
xnor U18998 (N_18998,N_18428,N_18340);
or U18999 (N_18999,N_18083,N_18068);
xor U19000 (N_19000,N_18510,N_18895);
xor U19001 (N_19001,N_18833,N_18613);
nand U19002 (N_19002,N_18775,N_18847);
or U19003 (N_19003,N_18679,N_18528);
and U19004 (N_19004,N_18907,N_18940);
nor U19005 (N_19005,N_18537,N_18883);
xor U19006 (N_19006,N_18678,N_18608);
nor U19007 (N_19007,N_18952,N_18919);
nand U19008 (N_19008,N_18987,N_18736);
nor U19009 (N_19009,N_18664,N_18655);
and U19010 (N_19010,N_18828,N_18914);
nand U19011 (N_19011,N_18932,N_18688);
nand U19012 (N_19012,N_18646,N_18999);
nand U19013 (N_19013,N_18978,N_18561);
or U19014 (N_19014,N_18665,N_18793);
nor U19015 (N_19015,N_18531,N_18637);
nor U19016 (N_19016,N_18844,N_18909);
xor U19017 (N_19017,N_18929,N_18906);
or U19018 (N_19018,N_18851,N_18603);
and U19019 (N_19019,N_18808,N_18965);
nor U19020 (N_19020,N_18635,N_18506);
nand U19021 (N_19021,N_18894,N_18598);
nand U19022 (N_19022,N_18990,N_18969);
xor U19023 (N_19023,N_18875,N_18609);
xor U19024 (N_19024,N_18873,N_18653);
xnor U19025 (N_19025,N_18810,N_18869);
or U19026 (N_19026,N_18770,N_18681);
and U19027 (N_19027,N_18629,N_18931);
nor U19028 (N_19028,N_18996,N_18755);
and U19029 (N_19029,N_18806,N_18581);
nor U19030 (N_19030,N_18541,N_18955);
xor U19031 (N_19031,N_18960,N_18812);
or U19032 (N_19032,N_18657,N_18804);
nor U19033 (N_19033,N_18795,N_18951);
and U19034 (N_19034,N_18985,N_18625);
or U19035 (N_19035,N_18862,N_18567);
nand U19036 (N_19036,N_18731,N_18831);
nor U19037 (N_19037,N_18902,N_18628);
or U19038 (N_19038,N_18964,N_18887);
xor U19039 (N_19039,N_18607,N_18821);
and U19040 (N_19040,N_18791,N_18939);
nand U19041 (N_19041,N_18675,N_18753);
nor U19042 (N_19042,N_18792,N_18974);
nor U19043 (N_19043,N_18535,N_18935);
nand U19044 (N_19044,N_18687,N_18897);
nor U19045 (N_19045,N_18579,N_18826);
and U19046 (N_19046,N_18942,N_18615);
or U19047 (N_19047,N_18692,N_18995);
nand U19048 (N_19048,N_18778,N_18580);
and U19049 (N_19049,N_18517,N_18602);
nand U19050 (N_19050,N_18839,N_18604);
or U19051 (N_19051,N_18976,N_18515);
or U19052 (N_19052,N_18893,N_18570);
xnor U19053 (N_19053,N_18714,N_18924);
nand U19054 (N_19054,N_18724,N_18658);
xor U19055 (N_19055,N_18986,N_18583);
nor U19056 (N_19056,N_18536,N_18533);
or U19057 (N_19057,N_18549,N_18972);
and U19058 (N_19058,N_18956,N_18761);
and U19059 (N_19059,N_18502,N_18915);
or U19060 (N_19060,N_18560,N_18758);
or U19061 (N_19061,N_18944,N_18538);
nor U19062 (N_19062,N_18728,N_18740);
nand U19063 (N_19063,N_18959,N_18565);
and U19064 (N_19064,N_18641,N_18689);
and U19065 (N_19065,N_18747,N_18624);
xnor U19066 (N_19066,N_18866,N_18648);
or U19067 (N_19067,N_18882,N_18846);
nand U19068 (N_19068,N_18558,N_18966);
or U19069 (N_19069,N_18691,N_18546);
nor U19070 (N_19070,N_18763,N_18864);
nand U19071 (N_19071,N_18874,N_18977);
xnor U19072 (N_19072,N_18988,N_18733);
nand U19073 (N_19073,N_18814,N_18879);
and U19074 (N_19074,N_18671,N_18920);
xor U19075 (N_19075,N_18837,N_18654);
nor U19076 (N_19076,N_18863,N_18899);
nor U19077 (N_19077,N_18950,N_18835);
xor U19078 (N_19078,N_18695,N_18601);
nor U19079 (N_19079,N_18680,N_18889);
nor U19080 (N_19080,N_18975,N_18922);
xnor U19081 (N_19081,N_18813,N_18872);
and U19082 (N_19082,N_18627,N_18534);
nand U19083 (N_19083,N_18910,N_18656);
nand U19084 (N_19084,N_18962,N_18521);
and U19085 (N_19085,N_18871,N_18584);
or U19086 (N_19086,N_18519,N_18830);
nand U19087 (N_19087,N_18711,N_18709);
or U19088 (N_19088,N_18784,N_18704);
xnor U19089 (N_19089,N_18732,N_18717);
nand U19090 (N_19090,N_18762,N_18652);
or U19091 (N_19091,N_18600,N_18721);
xnor U19092 (N_19092,N_18632,N_18997);
and U19093 (N_19093,N_18578,N_18557);
nand U19094 (N_19094,N_18746,N_18504);
or U19095 (N_19095,N_18823,N_18781);
or U19096 (N_19096,N_18530,N_18788);
nor U19097 (N_19097,N_18945,N_18794);
nor U19098 (N_19098,N_18766,N_18551);
nor U19099 (N_19099,N_18880,N_18735);
and U19100 (N_19100,N_18553,N_18722);
nand U19101 (N_19101,N_18824,N_18550);
nor U19102 (N_19102,N_18660,N_18759);
or U19103 (N_19103,N_18968,N_18649);
or U19104 (N_19104,N_18957,N_18529);
xnor U19105 (N_19105,N_18981,N_18523);
nand U19106 (N_19106,N_18760,N_18597);
or U19107 (N_19107,N_18797,N_18890);
nand U19108 (N_19108,N_18838,N_18850);
or U19109 (N_19109,N_18564,N_18522);
or U19110 (N_19110,N_18858,N_18514);
or U19111 (N_19111,N_18619,N_18905);
xor U19112 (N_19112,N_18562,N_18822);
nand U19113 (N_19113,N_18937,N_18511);
nor U19114 (N_19114,N_18507,N_18668);
nor U19115 (N_19115,N_18694,N_18983);
nand U19116 (N_19116,N_18661,N_18768);
nand U19117 (N_19117,N_18789,N_18903);
xor U19118 (N_19118,N_18832,N_18650);
xnor U19119 (N_19119,N_18991,N_18727);
or U19120 (N_19120,N_18685,N_18622);
nor U19121 (N_19121,N_18738,N_18848);
nand U19122 (N_19122,N_18908,N_18803);
xnor U19123 (N_19123,N_18585,N_18706);
nor U19124 (N_19124,N_18720,N_18936);
nor U19125 (N_19125,N_18749,N_18734);
nor U19126 (N_19126,N_18904,N_18786);
nor U19127 (N_19127,N_18643,N_18702);
nand U19128 (N_19128,N_18593,N_18690);
or U19129 (N_19129,N_18911,N_18647);
and U19130 (N_19130,N_18672,N_18563);
and U19131 (N_19131,N_18539,N_18925);
nor U19132 (N_19132,N_18693,N_18750);
nand U19133 (N_19133,N_18820,N_18540);
and U19134 (N_19134,N_18765,N_18855);
nor U19135 (N_19135,N_18913,N_18626);
nor U19136 (N_19136,N_18928,N_18742);
and U19137 (N_19137,N_18898,N_18730);
xor U19138 (N_19138,N_18699,N_18620);
xnor U19139 (N_19139,N_18973,N_18774);
or U19140 (N_19140,N_18712,N_18860);
and U19141 (N_19141,N_18994,N_18670);
nand U19142 (N_19142,N_18663,N_18642);
nor U19143 (N_19143,N_18548,N_18623);
and U19144 (N_19144,N_18769,N_18667);
xor U19145 (N_19145,N_18982,N_18923);
nand U19146 (N_19146,N_18917,N_18638);
nor U19147 (N_19147,N_18644,N_18729);
or U19148 (N_19148,N_18841,N_18543);
and U19149 (N_19149,N_18927,N_18958);
nand U19150 (N_19150,N_18980,N_18586);
nor U19151 (N_19151,N_18568,N_18989);
nor U19152 (N_19152,N_18612,N_18885);
and U19153 (N_19153,N_18787,N_18816);
nand U19154 (N_19154,N_18518,N_18503);
xnor U19155 (N_19155,N_18777,N_18916);
or U19156 (N_19156,N_18859,N_18509);
or U19157 (N_19157,N_18544,N_18798);
nor U19158 (N_19158,N_18817,N_18707);
xor U19159 (N_19159,N_18870,N_18590);
xnor U19160 (N_19160,N_18713,N_18520);
nor U19161 (N_19161,N_18500,N_18809);
xor U19162 (N_19162,N_18595,N_18877);
nand U19163 (N_19163,N_18834,N_18737);
and U19164 (N_19164,N_18524,N_18633);
nor U19165 (N_19165,N_18884,N_18516);
nand U19166 (N_19166,N_18552,N_18805);
nand U19167 (N_19167,N_18556,N_18881);
xnor U19168 (N_19168,N_18849,N_18751);
or U19169 (N_19169,N_18948,N_18811);
xor U19170 (N_19170,N_18545,N_18616);
nor U19171 (N_19171,N_18697,N_18576);
xor U19172 (N_19172,N_18926,N_18611);
nand U19173 (N_19173,N_18606,N_18780);
nand U19174 (N_19174,N_18527,N_18949);
and U19175 (N_19175,N_18577,N_18569);
nor U19176 (N_19176,N_18963,N_18745);
or U19177 (N_19177,N_18621,N_18998);
or U19178 (N_19178,N_18748,N_18796);
and U19179 (N_19179,N_18825,N_18992);
xnor U19180 (N_19180,N_18630,N_18840);
nor U19181 (N_19181,N_18930,N_18512);
nand U19182 (N_19182,N_18505,N_18744);
or U19183 (N_19183,N_18571,N_18573);
or U19184 (N_19184,N_18631,N_18900);
nand U19185 (N_19185,N_18961,N_18934);
or U19186 (N_19186,N_18659,N_18921);
xnor U19187 (N_19187,N_18971,N_18861);
or U19188 (N_19188,N_18979,N_18617);
nand U19189 (N_19189,N_18715,N_18852);
or U19190 (N_19190,N_18842,N_18891);
nor U19191 (N_19191,N_18754,N_18708);
nand U19192 (N_19192,N_18912,N_18856);
xnor U19193 (N_19193,N_18526,N_18896);
and U19194 (N_19194,N_18943,N_18764);
or U19195 (N_19195,N_18686,N_18634);
or U19196 (N_19196,N_18718,N_18799);
nand U19197 (N_19197,N_18547,N_18572);
and U19198 (N_19198,N_18741,N_18676);
xor U19199 (N_19199,N_18843,N_18867);
and U19200 (N_19200,N_18888,N_18554);
or U19201 (N_19201,N_18865,N_18710);
nand U19202 (N_19202,N_18639,N_18614);
and U19203 (N_19203,N_18501,N_18984);
and U19204 (N_19204,N_18779,N_18705);
or U19205 (N_19205,N_18698,N_18723);
xnor U19206 (N_19206,N_18640,N_18941);
or U19207 (N_19207,N_18947,N_18782);
nand U19208 (N_19208,N_18574,N_18773);
xnor U19209 (N_19209,N_18599,N_18589);
or U19210 (N_19210,N_18725,N_18807);
xor U19211 (N_19211,N_18684,N_18771);
nand U19212 (N_19212,N_18818,N_18610);
xnor U19213 (N_19213,N_18756,N_18636);
and U19214 (N_19214,N_18800,N_18582);
nand U19215 (N_19215,N_18701,N_18892);
nand U19216 (N_19216,N_18669,N_18790);
xnor U19217 (N_19217,N_18967,N_18783);
or U19218 (N_19218,N_18683,N_18513);
nand U19219 (N_19219,N_18605,N_18566);
nor U19220 (N_19220,N_18845,N_18696);
and U19221 (N_19221,N_18525,N_18802);
nand U19222 (N_19222,N_18651,N_18752);
xor U19223 (N_19223,N_18954,N_18993);
xor U19224 (N_19224,N_18836,N_18739);
xnor U19225 (N_19225,N_18716,N_18886);
xnor U19226 (N_19226,N_18829,N_18508);
nor U19227 (N_19227,N_18677,N_18853);
and U19228 (N_19228,N_18776,N_18618);
nor U19229 (N_19229,N_18946,N_18662);
xnor U19230 (N_19230,N_18592,N_18726);
and U19231 (N_19231,N_18719,N_18596);
or U19232 (N_19232,N_18757,N_18819);
nor U19233 (N_19233,N_18588,N_18555);
xnor U19234 (N_19234,N_18970,N_18587);
xor U19235 (N_19235,N_18857,N_18674);
nor U19236 (N_19236,N_18785,N_18878);
and U19237 (N_19237,N_18594,N_18938);
xor U19238 (N_19238,N_18767,N_18645);
nor U19239 (N_19239,N_18901,N_18575);
nand U19240 (N_19240,N_18700,N_18542);
nand U19241 (N_19241,N_18743,N_18703);
nor U19242 (N_19242,N_18933,N_18559);
and U19243 (N_19243,N_18591,N_18854);
nor U19244 (N_19244,N_18673,N_18827);
or U19245 (N_19245,N_18953,N_18876);
or U19246 (N_19246,N_18815,N_18918);
or U19247 (N_19247,N_18532,N_18772);
or U19248 (N_19248,N_18682,N_18666);
and U19249 (N_19249,N_18868,N_18801);
nand U19250 (N_19250,N_18901,N_18622);
or U19251 (N_19251,N_18585,N_18519);
nor U19252 (N_19252,N_18648,N_18726);
nand U19253 (N_19253,N_18942,N_18920);
or U19254 (N_19254,N_18509,N_18530);
nand U19255 (N_19255,N_18921,N_18972);
nand U19256 (N_19256,N_18519,N_18558);
nand U19257 (N_19257,N_18888,N_18611);
nand U19258 (N_19258,N_18546,N_18896);
and U19259 (N_19259,N_18657,N_18953);
and U19260 (N_19260,N_18770,N_18898);
xor U19261 (N_19261,N_18637,N_18932);
xnor U19262 (N_19262,N_18854,N_18622);
nor U19263 (N_19263,N_18689,N_18527);
or U19264 (N_19264,N_18837,N_18645);
xor U19265 (N_19265,N_18779,N_18871);
nor U19266 (N_19266,N_18584,N_18605);
nor U19267 (N_19267,N_18745,N_18887);
or U19268 (N_19268,N_18949,N_18899);
nand U19269 (N_19269,N_18918,N_18966);
nand U19270 (N_19270,N_18834,N_18846);
nand U19271 (N_19271,N_18815,N_18791);
or U19272 (N_19272,N_18760,N_18862);
xnor U19273 (N_19273,N_18737,N_18718);
and U19274 (N_19274,N_18518,N_18898);
or U19275 (N_19275,N_18504,N_18981);
and U19276 (N_19276,N_18525,N_18909);
nor U19277 (N_19277,N_18749,N_18910);
nand U19278 (N_19278,N_18744,N_18991);
and U19279 (N_19279,N_18528,N_18784);
or U19280 (N_19280,N_18982,N_18897);
nand U19281 (N_19281,N_18553,N_18943);
nor U19282 (N_19282,N_18942,N_18862);
nor U19283 (N_19283,N_18618,N_18888);
and U19284 (N_19284,N_18591,N_18566);
nand U19285 (N_19285,N_18941,N_18598);
xnor U19286 (N_19286,N_18898,N_18775);
or U19287 (N_19287,N_18812,N_18780);
nand U19288 (N_19288,N_18816,N_18583);
or U19289 (N_19289,N_18961,N_18553);
nor U19290 (N_19290,N_18879,N_18801);
nand U19291 (N_19291,N_18782,N_18612);
nor U19292 (N_19292,N_18861,N_18902);
or U19293 (N_19293,N_18623,N_18593);
nand U19294 (N_19294,N_18816,N_18784);
nand U19295 (N_19295,N_18833,N_18891);
xor U19296 (N_19296,N_18924,N_18692);
nand U19297 (N_19297,N_18849,N_18847);
nand U19298 (N_19298,N_18871,N_18736);
xnor U19299 (N_19299,N_18646,N_18617);
and U19300 (N_19300,N_18983,N_18641);
nand U19301 (N_19301,N_18685,N_18853);
xor U19302 (N_19302,N_18978,N_18846);
and U19303 (N_19303,N_18824,N_18982);
or U19304 (N_19304,N_18564,N_18530);
and U19305 (N_19305,N_18744,N_18868);
nor U19306 (N_19306,N_18670,N_18725);
nor U19307 (N_19307,N_18607,N_18624);
nor U19308 (N_19308,N_18687,N_18941);
or U19309 (N_19309,N_18636,N_18716);
nand U19310 (N_19310,N_18545,N_18506);
nand U19311 (N_19311,N_18927,N_18696);
xor U19312 (N_19312,N_18532,N_18718);
nand U19313 (N_19313,N_18846,N_18604);
or U19314 (N_19314,N_18531,N_18723);
nor U19315 (N_19315,N_18652,N_18630);
nand U19316 (N_19316,N_18961,N_18906);
nor U19317 (N_19317,N_18611,N_18560);
xor U19318 (N_19318,N_18672,N_18561);
or U19319 (N_19319,N_18859,N_18966);
nor U19320 (N_19320,N_18875,N_18753);
xor U19321 (N_19321,N_18601,N_18919);
xnor U19322 (N_19322,N_18947,N_18800);
and U19323 (N_19323,N_18765,N_18851);
or U19324 (N_19324,N_18757,N_18845);
nand U19325 (N_19325,N_18901,N_18674);
nor U19326 (N_19326,N_18587,N_18809);
nand U19327 (N_19327,N_18788,N_18584);
nor U19328 (N_19328,N_18659,N_18656);
or U19329 (N_19329,N_18585,N_18878);
or U19330 (N_19330,N_18510,N_18574);
nor U19331 (N_19331,N_18666,N_18798);
xor U19332 (N_19332,N_18862,N_18737);
nor U19333 (N_19333,N_18737,N_18799);
and U19334 (N_19334,N_18757,N_18927);
and U19335 (N_19335,N_18683,N_18964);
nor U19336 (N_19336,N_18971,N_18588);
or U19337 (N_19337,N_18726,N_18533);
nor U19338 (N_19338,N_18767,N_18591);
nand U19339 (N_19339,N_18747,N_18857);
or U19340 (N_19340,N_18894,N_18501);
nor U19341 (N_19341,N_18578,N_18959);
and U19342 (N_19342,N_18617,N_18764);
or U19343 (N_19343,N_18982,N_18861);
nor U19344 (N_19344,N_18532,N_18928);
nand U19345 (N_19345,N_18894,N_18726);
or U19346 (N_19346,N_18889,N_18639);
xnor U19347 (N_19347,N_18890,N_18533);
or U19348 (N_19348,N_18801,N_18839);
and U19349 (N_19349,N_18932,N_18603);
and U19350 (N_19350,N_18694,N_18717);
or U19351 (N_19351,N_18678,N_18663);
nor U19352 (N_19352,N_18542,N_18525);
nor U19353 (N_19353,N_18665,N_18834);
and U19354 (N_19354,N_18527,N_18922);
or U19355 (N_19355,N_18549,N_18848);
nand U19356 (N_19356,N_18709,N_18525);
xor U19357 (N_19357,N_18547,N_18823);
xor U19358 (N_19358,N_18730,N_18722);
xor U19359 (N_19359,N_18929,N_18720);
and U19360 (N_19360,N_18535,N_18833);
nand U19361 (N_19361,N_18718,N_18650);
and U19362 (N_19362,N_18995,N_18601);
nor U19363 (N_19363,N_18899,N_18580);
or U19364 (N_19364,N_18738,N_18975);
and U19365 (N_19365,N_18967,N_18574);
nand U19366 (N_19366,N_18735,N_18703);
or U19367 (N_19367,N_18668,N_18513);
or U19368 (N_19368,N_18619,N_18665);
xnor U19369 (N_19369,N_18566,N_18872);
or U19370 (N_19370,N_18965,N_18756);
and U19371 (N_19371,N_18768,N_18796);
or U19372 (N_19372,N_18574,N_18699);
nor U19373 (N_19373,N_18759,N_18588);
and U19374 (N_19374,N_18624,N_18510);
or U19375 (N_19375,N_18709,N_18516);
xnor U19376 (N_19376,N_18539,N_18883);
and U19377 (N_19377,N_18774,N_18668);
xor U19378 (N_19378,N_18855,N_18933);
nor U19379 (N_19379,N_18903,N_18966);
or U19380 (N_19380,N_18680,N_18672);
nor U19381 (N_19381,N_18715,N_18632);
nor U19382 (N_19382,N_18680,N_18838);
nand U19383 (N_19383,N_18834,N_18645);
nor U19384 (N_19384,N_18670,N_18667);
nand U19385 (N_19385,N_18588,N_18842);
and U19386 (N_19386,N_18677,N_18603);
and U19387 (N_19387,N_18622,N_18972);
or U19388 (N_19388,N_18712,N_18954);
nand U19389 (N_19389,N_18878,N_18870);
nor U19390 (N_19390,N_18587,N_18737);
nor U19391 (N_19391,N_18595,N_18840);
xor U19392 (N_19392,N_18662,N_18900);
xor U19393 (N_19393,N_18889,N_18992);
nor U19394 (N_19394,N_18597,N_18581);
nor U19395 (N_19395,N_18861,N_18690);
or U19396 (N_19396,N_18675,N_18655);
nor U19397 (N_19397,N_18585,N_18543);
xnor U19398 (N_19398,N_18606,N_18953);
xnor U19399 (N_19399,N_18570,N_18980);
and U19400 (N_19400,N_18807,N_18895);
and U19401 (N_19401,N_18790,N_18789);
and U19402 (N_19402,N_18778,N_18523);
and U19403 (N_19403,N_18891,N_18661);
xor U19404 (N_19404,N_18981,N_18566);
xnor U19405 (N_19405,N_18716,N_18877);
xor U19406 (N_19406,N_18724,N_18911);
or U19407 (N_19407,N_18677,N_18631);
nor U19408 (N_19408,N_18572,N_18635);
nor U19409 (N_19409,N_18623,N_18531);
and U19410 (N_19410,N_18681,N_18778);
and U19411 (N_19411,N_18618,N_18829);
nand U19412 (N_19412,N_18924,N_18941);
nand U19413 (N_19413,N_18930,N_18793);
nor U19414 (N_19414,N_18795,N_18630);
and U19415 (N_19415,N_18827,N_18983);
or U19416 (N_19416,N_18876,N_18649);
or U19417 (N_19417,N_18561,N_18767);
xnor U19418 (N_19418,N_18662,N_18760);
nor U19419 (N_19419,N_18667,N_18998);
nor U19420 (N_19420,N_18659,N_18651);
nand U19421 (N_19421,N_18772,N_18913);
or U19422 (N_19422,N_18919,N_18618);
nand U19423 (N_19423,N_18777,N_18998);
nor U19424 (N_19424,N_18870,N_18545);
or U19425 (N_19425,N_18921,N_18984);
and U19426 (N_19426,N_18892,N_18810);
and U19427 (N_19427,N_18832,N_18737);
and U19428 (N_19428,N_18612,N_18680);
xnor U19429 (N_19429,N_18876,N_18686);
or U19430 (N_19430,N_18832,N_18594);
or U19431 (N_19431,N_18633,N_18891);
nand U19432 (N_19432,N_18547,N_18659);
or U19433 (N_19433,N_18627,N_18617);
and U19434 (N_19434,N_18714,N_18581);
xor U19435 (N_19435,N_18683,N_18644);
nor U19436 (N_19436,N_18928,N_18901);
and U19437 (N_19437,N_18576,N_18895);
and U19438 (N_19438,N_18554,N_18738);
xnor U19439 (N_19439,N_18726,N_18852);
nand U19440 (N_19440,N_18810,N_18978);
or U19441 (N_19441,N_18985,N_18755);
xor U19442 (N_19442,N_18872,N_18863);
nand U19443 (N_19443,N_18868,N_18649);
xnor U19444 (N_19444,N_18905,N_18669);
or U19445 (N_19445,N_18760,N_18855);
and U19446 (N_19446,N_18856,N_18939);
nor U19447 (N_19447,N_18863,N_18956);
or U19448 (N_19448,N_18897,N_18616);
xor U19449 (N_19449,N_18744,N_18778);
xor U19450 (N_19450,N_18923,N_18795);
and U19451 (N_19451,N_18924,N_18878);
xor U19452 (N_19452,N_18779,N_18602);
nor U19453 (N_19453,N_18898,N_18960);
xnor U19454 (N_19454,N_18611,N_18980);
and U19455 (N_19455,N_18861,N_18547);
and U19456 (N_19456,N_18884,N_18986);
and U19457 (N_19457,N_18885,N_18807);
xor U19458 (N_19458,N_18934,N_18775);
and U19459 (N_19459,N_18594,N_18990);
nand U19460 (N_19460,N_18782,N_18961);
or U19461 (N_19461,N_18514,N_18510);
nand U19462 (N_19462,N_18596,N_18936);
or U19463 (N_19463,N_18784,N_18735);
nand U19464 (N_19464,N_18838,N_18968);
or U19465 (N_19465,N_18731,N_18737);
and U19466 (N_19466,N_18601,N_18769);
and U19467 (N_19467,N_18891,N_18989);
xnor U19468 (N_19468,N_18989,N_18634);
or U19469 (N_19469,N_18646,N_18671);
nand U19470 (N_19470,N_18710,N_18994);
nand U19471 (N_19471,N_18566,N_18935);
xor U19472 (N_19472,N_18690,N_18603);
xor U19473 (N_19473,N_18720,N_18647);
xnor U19474 (N_19474,N_18972,N_18730);
nand U19475 (N_19475,N_18550,N_18512);
and U19476 (N_19476,N_18812,N_18667);
nor U19477 (N_19477,N_18735,N_18628);
nand U19478 (N_19478,N_18816,N_18872);
and U19479 (N_19479,N_18572,N_18902);
nand U19480 (N_19480,N_18528,N_18688);
and U19481 (N_19481,N_18839,N_18688);
and U19482 (N_19482,N_18957,N_18726);
xnor U19483 (N_19483,N_18516,N_18616);
or U19484 (N_19484,N_18714,N_18684);
nor U19485 (N_19485,N_18791,N_18596);
nor U19486 (N_19486,N_18563,N_18878);
nand U19487 (N_19487,N_18774,N_18529);
and U19488 (N_19488,N_18913,N_18939);
xnor U19489 (N_19489,N_18696,N_18943);
xor U19490 (N_19490,N_18591,N_18820);
xnor U19491 (N_19491,N_18528,N_18750);
and U19492 (N_19492,N_18677,N_18872);
xnor U19493 (N_19493,N_18981,N_18743);
nor U19494 (N_19494,N_18995,N_18788);
or U19495 (N_19495,N_18974,N_18518);
and U19496 (N_19496,N_18501,N_18932);
or U19497 (N_19497,N_18602,N_18793);
or U19498 (N_19498,N_18997,N_18948);
or U19499 (N_19499,N_18522,N_18565);
and U19500 (N_19500,N_19192,N_19333);
and U19501 (N_19501,N_19083,N_19411);
and U19502 (N_19502,N_19232,N_19498);
and U19503 (N_19503,N_19127,N_19357);
nor U19504 (N_19504,N_19334,N_19254);
nand U19505 (N_19505,N_19032,N_19121);
nor U19506 (N_19506,N_19466,N_19362);
or U19507 (N_19507,N_19123,N_19265);
nor U19508 (N_19508,N_19188,N_19463);
nor U19509 (N_19509,N_19157,N_19026);
nor U19510 (N_19510,N_19247,N_19181);
and U19511 (N_19511,N_19170,N_19143);
and U19512 (N_19512,N_19483,N_19383);
and U19513 (N_19513,N_19251,N_19271);
or U19514 (N_19514,N_19344,N_19320);
nor U19515 (N_19515,N_19057,N_19093);
and U19516 (N_19516,N_19231,N_19211);
xor U19517 (N_19517,N_19115,N_19212);
or U19518 (N_19518,N_19112,N_19124);
or U19519 (N_19519,N_19243,N_19087);
nor U19520 (N_19520,N_19052,N_19216);
nor U19521 (N_19521,N_19240,N_19282);
xnor U19522 (N_19522,N_19384,N_19287);
xor U19523 (N_19523,N_19108,N_19142);
and U19524 (N_19524,N_19060,N_19015);
xor U19525 (N_19525,N_19474,N_19202);
nand U19526 (N_19526,N_19033,N_19224);
nand U19527 (N_19527,N_19402,N_19494);
and U19528 (N_19528,N_19013,N_19377);
nand U19529 (N_19529,N_19488,N_19173);
nor U19530 (N_19530,N_19058,N_19332);
or U19531 (N_19531,N_19397,N_19199);
nand U19532 (N_19532,N_19046,N_19230);
nor U19533 (N_19533,N_19117,N_19272);
nand U19534 (N_19534,N_19329,N_19130);
or U19535 (N_19535,N_19414,N_19423);
and U19536 (N_19536,N_19473,N_19063);
nor U19537 (N_19537,N_19183,N_19338);
and U19538 (N_19538,N_19492,N_19210);
and U19539 (N_19539,N_19168,N_19040);
and U19540 (N_19540,N_19159,N_19128);
or U19541 (N_19541,N_19234,N_19480);
xor U19542 (N_19542,N_19074,N_19141);
and U19543 (N_19543,N_19438,N_19138);
or U19544 (N_19544,N_19252,N_19053);
or U19545 (N_19545,N_19499,N_19311);
nor U19546 (N_19546,N_19069,N_19394);
and U19547 (N_19547,N_19286,N_19289);
and U19548 (N_19548,N_19491,N_19253);
nand U19549 (N_19549,N_19431,N_19244);
nor U19550 (N_19550,N_19261,N_19072);
and U19551 (N_19551,N_19184,N_19007);
or U19552 (N_19552,N_19082,N_19324);
nand U19553 (N_19553,N_19160,N_19449);
nor U19554 (N_19554,N_19070,N_19442);
nand U19555 (N_19555,N_19154,N_19398);
nand U19556 (N_19556,N_19386,N_19430);
and U19557 (N_19557,N_19493,N_19229);
nand U19558 (N_19558,N_19061,N_19169);
xor U19559 (N_19559,N_19393,N_19054);
nand U19560 (N_19560,N_19443,N_19204);
and U19561 (N_19561,N_19217,N_19413);
nor U19562 (N_19562,N_19385,N_19328);
nor U19563 (N_19563,N_19429,N_19167);
and U19564 (N_19564,N_19018,N_19441);
nand U19565 (N_19565,N_19428,N_19484);
and U19566 (N_19566,N_19045,N_19487);
xnor U19567 (N_19567,N_19369,N_19301);
nand U19568 (N_19568,N_19291,N_19309);
or U19569 (N_19569,N_19303,N_19129);
nand U19570 (N_19570,N_19350,N_19312);
and U19571 (N_19571,N_19379,N_19178);
nand U19572 (N_19572,N_19360,N_19479);
nand U19573 (N_19573,N_19283,N_19064);
nand U19574 (N_19574,N_19023,N_19470);
nand U19575 (N_19575,N_19034,N_19279);
nand U19576 (N_19576,N_19006,N_19408);
or U19577 (N_19577,N_19485,N_19118);
nand U19578 (N_19578,N_19177,N_19073);
nor U19579 (N_19579,N_19455,N_19161);
nor U19580 (N_19580,N_19445,N_19010);
or U19581 (N_19581,N_19246,N_19315);
or U19582 (N_19582,N_19353,N_19077);
xnor U19583 (N_19583,N_19342,N_19260);
nand U19584 (N_19584,N_19144,N_19381);
and U19585 (N_19585,N_19102,N_19292);
nor U19586 (N_19586,N_19266,N_19120);
xor U19587 (N_19587,N_19456,N_19076);
and U19588 (N_19588,N_19462,N_19049);
xor U19589 (N_19589,N_19314,N_19364);
xnor U19590 (N_19590,N_19255,N_19444);
and U19591 (N_19591,N_19335,N_19495);
xor U19592 (N_19592,N_19215,N_19062);
and U19593 (N_19593,N_19136,N_19290);
nor U19594 (N_19594,N_19203,N_19318);
and U19595 (N_19595,N_19080,N_19294);
nand U19596 (N_19596,N_19317,N_19158);
nor U19597 (N_19597,N_19425,N_19476);
or U19598 (N_19598,N_19196,N_19280);
xor U19599 (N_19599,N_19078,N_19024);
xnor U19600 (N_19600,N_19276,N_19106);
xnor U19601 (N_19601,N_19351,N_19306);
xor U19602 (N_19602,N_19222,N_19081);
xor U19603 (N_19603,N_19002,N_19099);
nor U19604 (N_19604,N_19179,N_19304);
and U19605 (N_19605,N_19417,N_19037);
nand U19606 (N_19606,N_19004,N_19162);
nand U19607 (N_19607,N_19238,N_19194);
or U19608 (N_19608,N_19305,N_19302);
or U19609 (N_19609,N_19446,N_19050);
nor U19610 (N_19610,N_19091,N_19307);
nand U19611 (N_19611,N_19259,N_19469);
or U19612 (N_19612,N_19156,N_19009);
xnor U19613 (N_19613,N_19405,N_19263);
xnor U19614 (N_19614,N_19088,N_19206);
nand U19615 (N_19615,N_19436,N_19126);
xnor U19616 (N_19616,N_19191,N_19207);
nor U19617 (N_19617,N_19270,N_19137);
nand U19618 (N_19618,N_19086,N_19225);
or U19619 (N_19619,N_19134,N_19012);
xor U19620 (N_19620,N_19109,N_19047);
and U19621 (N_19621,N_19092,N_19005);
xnor U19622 (N_19622,N_19075,N_19481);
xor U19623 (N_19623,N_19331,N_19223);
or U19624 (N_19624,N_19450,N_19003);
and U19625 (N_19625,N_19415,N_19275);
nor U19626 (N_19626,N_19299,N_19400);
nand U19627 (N_19627,N_19226,N_19163);
nand U19628 (N_19628,N_19281,N_19375);
and U19629 (N_19629,N_19457,N_19453);
or U19630 (N_19630,N_19490,N_19395);
nand U19631 (N_19631,N_19391,N_19042);
nor U19632 (N_19632,N_19349,N_19296);
and U19633 (N_19633,N_19201,N_19475);
nor U19634 (N_19634,N_19104,N_19298);
or U19635 (N_19635,N_19418,N_19187);
or U19636 (N_19636,N_19147,N_19008);
nor U19637 (N_19637,N_19327,N_19084);
nand U19638 (N_19638,N_19267,N_19094);
and U19639 (N_19639,N_19348,N_19451);
xnor U19640 (N_19640,N_19020,N_19482);
and U19641 (N_19641,N_19343,N_19175);
nor U19642 (N_19642,N_19472,N_19354);
and U19643 (N_19643,N_19101,N_19110);
or U19644 (N_19644,N_19363,N_19021);
nor U19645 (N_19645,N_19111,N_19239);
xnor U19646 (N_19646,N_19326,N_19310);
nand U19647 (N_19647,N_19366,N_19464);
or U19648 (N_19648,N_19030,N_19345);
and U19649 (N_19649,N_19218,N_19460);
xor U19650 (N_19650,N_19347,N_19434);
or U19651 (N_19651,N_19432,N_19209);
xnor U19652 (N_19652,N_19416,N_19300);
and U19653 (N_19653,N_19262,N_19389);
nand U19654 (N_19654,N_19257,N_19146);
xor U19655 (N_19655,N_19219,N_19268);
and U19656 (N_19656,N_19245,N_19036);
nor U19657 (N_19657,N_19330,N_19103);
and U19658 (N_19658,N_19471,N_19017);
nor U19659 (N_19659,N_19352,N_19424);
or U19660 (N_19660,N_19153,N_19228);
or U19661 (N_19661,N_19241,N_19486);
xor U19662 (N_19662,N_19155,N_19149);
and U19663 (N_19663,N_19139,N_19233);
or U19664 (N_19664,N_19025,N_19195);
xnor U19665 (N_19665,N_19105,N_19370);
nor U19666 (N_19666,N_19237,N_19358);
xor U19667 (N_19667,N_19097,N_19264);
xor U19668 (N_19668,N_19337,N_19410);
or U19669 (N_19669,N_19447,N_19068);
or U19670 (N_19670,N_19185,N_19277);
xor U19671 (N_19671,N_19467,N_19421);
and U19672 (N_19672,N_19131,N_19113);
nor U19673 (N_19673,N_19433,N_19227);
nand U19674 (N_19674,N_19284,N_19107);
or U19675 (N_19675,N_19190,N_19039);
xor U19676 (N_19676,N_19197,N_19412);
and U19677 (N_19677,N_19182,N_19171);
nand U19678 (N_19678,N_19396,N_19001);
nand U19679 (N_19679,N_19346,N_19140);
or U19680 (N_19680,N_19341,N_19308);
and U19681 (N_19681,N_19269,N_19373);
xor U19682 (N_19682,N_19193,N_19458);
nand U19683 (N_19683,N_19114,N_19014);
or U19684 (N_19684,N_19387,N_19249);
and U19685 (N_19685,N_19392,N_19096);
nand U19686 (N_19686,N_19371,N_19221);
and U19687 (N_19687,N_19340,N_19066);
nor U19688 (N_19688,N_19055,N_19372);
or U19689 (N_19689,N_19019,N_19031);
nand U19690 (N_19690,N_19205,N_19213);
nor U19691 (N_19691,N_19166,N_19100);
xor U19692 (N_19692,N_19079,N_19321);
nand U19693 (N_19693,N_19465,N_19355);
nand U19694 (N_19694,N_19016,N_19059);
and U19695 (N_19695,N_19095,N_19085);
xor U19696 (N_19696,N_19089,N_19145);
nor U19697 (N_19697,N_19043,N_19090);
nand U19698 (N_19698,N_19011,N_19151);
and U19699 (N_19699,N_19388,N_19407);
xnor U19700 (N_19700,N_19048,N_19478);
xnor U19701 (N_19701,N_19250,N_19258);
or U19702 (N_19702,N_19319,N_19133);
xor U19703 (N_19703,N_19098,N_19489);
nor U19704 (N_19704,N_19165,N_19119);
nand U19705 (N_19705,N_19273,N_19420);
nor U19706 (N_19706,N_19236,N_19390);
and U19707 (N_19707,N_19051,N_19477);
or U19708 (N_19708,N_19367,N_19041);
and U19709 (N_19709,N_19454,N_19409);
nor U19710 (N_19710,N_19378,N_19176);
xor U19711 (N_19711,N_19022,N_19404);
xor U19712 (N_19712,N_19406,N_19316);
nor U19713 (N_19713,N_19422,N_19497);
xnor U19714 (N_19714,N_19440,N_19116);
or U19715 (N_19715,N_19132,N_19180);
nand U19716 (N_19716,N_19365,N_19468);
or U19717 (N_19717,N_19380,N_19071);
nand U19718 (N_19718,N_19189,N_19427);
and U19719 (N_19719,N_19452,N_19285);
nor U19720 (N_19720,N_19459,N_19248);
xor U19721 (N_19721,N_19496,N_19419);
and U19722 (N_19722,N_19065,N_19186);
nand U19723 (N_19723,N_19382,N_19323);
nor U19724 (N_19724,N_19374,N_19000);
nor U19725 (N_19725,N_19399,N_19359);
or U19726 (N_19726,N_19437,N_19368);
xor U19727 (N_19727,N_19235,N_19403);
xor U19728 (N_19728,N_19208,N_19293);
nor U19729 (N_19729,N_19122,N_19164);
or U19730 (N_19730,N_19056,N_19401);
and U19731 (N_19731,N_19339,N_19035);
or U19732 (N_19732,N_19148,N_19028);
or U19733 (N_19733,N_19435,N_19198);
and U19734 (N_19734,N_19152,N_19461);
nand U19735 (N_19735,N_19376,N_19336);
nor U19736 (N_19736,N_19278,N_19448);
or U19737 (N_19737,N_19322,N_19044);
nand U19738 (N_19738,N_19135,N_19426);
and U19739 (N_19739,N_19150,N_19439);
and U19740 (N_19740,N_19288,N_19313);
or U19741 (N_19741,N_19242,N_19295);
or U19742 (N_19742,N_19214,N_19297);
nor U19743 (N_19743,N_19038,N_19067);
nor U19744 (N_19744,N_19125,N_19256);
nand U19745 (N_19745,N_19274,N_19027);
or U19746 (N_19746,N_19174,N_19325);
nor U19747 (N_19747,N_19200,N_19172);
xor U19748 (N_19748,N_19220,N_19029);
or U19749 (N_19749,N_19356,N_19361);
and U19750 (N_19750,N_19209,N_19420);
and U19751 (N_19751,N_19274,N_19410);
and U19752 (N_19752,N_19062,N_19400);
nand U19753 (N_19753,N_19314,N_19127);
nor U19754 (N_19754,N_19240,N_19166);
and U19755 (N_19755,N_19462,N_19498);
xnor U19756 (N_19756,N_19021,N_19040);
or U19757 (N_19757,N_19144,N_19256);
xor U19758 (N_19758,N_19359,N_19051);
nand U19759 (N_19759,N_19254,N_19461);
nand U19760 (N_19760,N_19198,N_19196);
xor U19761 (N_19761,N_19399,N_19225);
nor U19762 (N_19762,N_19171,N_19081);
or U19763 (N_19763,N_19112,N_19472);
and U19764 (N_19764,N_19256,N_19232);
or U19765 (N_19765,N_19444,N_19106);
or U19766 (N_19766,N_19497,N_19382);
xnor U19767 (N_19767,N_19353,N_19059);
xor U19768 (N_19768,N_19378,N_19311);
or U19769 (N_19769,N_19417,N_19022);
nor U19770 (N_19770,N_19390,N_19048);
nor U19771 (N_19771,N_19110,N_19164);
or U19772 (N_19772,N_19164,N_19270);
and U19773 (N_19773,N_19349,N_19145);
nor U19774 (N_19774,N_19380,N_19115);
nand U19775 (N_19775,N_19321,N_19370);
or U19776 (N_19776,N_19109,N_19175);
nand U19777 (N_19777,N_19081,N_19354);
nand U19778 (N_19778,N_19381,N_19361);
and U19779 (N_19779,N_19135,N_19315);
and U19780 (N_19780,N_19442,N_19198);
nor U19781 (N_19781,N_19288,N_19330);
nor U19782 (N_19782,N_19048,N_19258);
and U19783 (N_19783,N_19034,N_19392);
xor U19784 (N_19784,N_19199,N_19165);
and U19785 (N_19785,N_19039,N_19256);
or U19786 (N_19786,N_19114,N_19022);
and U19787 (N_19787,N_19361,N_19236);
or U19788 (N_19788,N_19347,N_19245);
and U19789 (N_19789,N_19428,N_19268);
nand U19790 (N_19790,N_19142,N_19464);
or U19791 (N_19791,N_19346,N_19481);
or U19792 (N_19792,N_19285,N_19344);
nand U19793 (N_19793,N_19273,N_19264);
or U19794 (N_19794,N_19132,N_19497);
nor U19795 (N_19795,N_19320,N_19448);
or U19796 (N_19796,N_19490,N_19445);
xnor U19797 (N_19797,N_19498,N_19460);
and U19798 (N_19798,N_19210,N_19243);
or U19799 (N_19799,N_19393,N_19204);
nand U19800 (N_19800,N_19278,N_19416);
xnor U19801 (N_19801,N_19070,N_19254);
nor U19802 (N_19802,N_19421,N_19437);
and U19803 (N_19803,N_19293,N_19015);
nor U19804 (N_19804,N_19085,N_19199);
xor U19805 (N_19805,N_19296,N_19008);
xnor U19806 (N_19806,N_19163,N_19359);
xor U19807 (N_19807,N_19206,N_19123);
nand U19808 (N_19808,N_19142,N_19038);
or U19809 (N_19809,N_19079,N_19309);
or U19810 (N_19810,N_19025,N_19405);
nand U19811 (N_19811,N_19207,N_19222);
and U19812 (N_19812,N_19195,N_19188);
nand U19813 (N_19813,N_19382,N_19292);
or U19814 (N_19814,N_19011,N_19175);
or U19815 (N_19815,N_19225,N_19137);
nor U19816 (N_19816,N_19347,N_19066);
nand U19817 (N_19817,N_19334,N_19055);
xor U19818 (N_19818,N_19218,N_19164);
or U19819 (N_19819,N_19296,N_19403);
or U19820 (N_19820,N_19198,N_19026);
nand U19821 (N_19821,N_19007,N_19423);
and U19822 (N_19822,N_19468,N_19329);
or U19823 (N_19823,N_19338,N_19172);
nor U19824 (N_19824,N_19465,N_19346);
or U19825 (N_19825,N_19116,N_19093);
and U19826 (N_19826,N_19405,N_19485);
and U19827 (N_19827,N_19195,N_19331);
or U19828 (N_19828,N_19140,N_19116);
and U19829 (N_19829,N_19181,N_19445);
or U19830 (N_19830,N_19202,N_19382);
nor U19831 (N_19831,N_19362,N_19206);
or U19832 (N_19832,N_19032,N_19301);
nand U19833 (N_19833,N_19020,N_19231);
and U19834 (N_19834,N_19258,N_19444);
and U19835 (N_19835,N_19393,N_19110);
nor U19836 (N_19836,N_19044,N_19388);
or U19837 (N_19837,N_19366,N_19468);
nor U19838 (N_19838,N_19470,N_19010);
and U19839 (N_19839,N_19022,N_19107);
nand U19840 (N_19840,N_19086,N_19213);
and U19841 (N_19841,N_19022,N_19225);
xnor U19842 (N_19842,N_19155,N_19467);
nand U19843 (N_19843,N_19312,N_19364);
and U19844 (N_19844,N_19418,N_19448);
nand U19845 (N_19845,N_19272,N_19195);
nand U19846 (N_19846,N_19163,N_19446);
and U19847 (N_19847,N_19471,N_19346);
nand U19848 (N_19848,N_19383,N_19239);
nor U19849 (N_19849,N_19092,N_19196);
and U19850 (N_19850,N_19468,N_19075);
nand U19851 (N_19851,N_19044,N_19380);
nor U19852 (N_19852,N_19089,N_19294);
nor U19853 (N_19853,N_19483,N_19413);
xor U19854 (N_19854,N_19487,N_19411);
or U19855 (N_19855,N_19151,N_19432);
or U19856 (N_19856,N_19093,N_19040);
nand U19857 (N_19857,N_19043,N_19164);
nand U19858 (N_19858,N_19432,N_19025);
and U19859 (N_19859,N_19185,N_19384);
nor U19860 (N_19860,N_19382,N_19096);
nand U19861 (N_19861,N_19429,N_19466);
nor U19862 (N_19862,N_19330,N_19006);
nor U19863 (N_19863,N_19253,N_19252);
and U19864 (N_19864,N_19431,N_19013);
xnor U19865 (N_19865,N_19033,N_19171);
nand U19866 (N_19866,N_19399,N_19189);
or U19867 (N_19867,N_19110,N_19122);
nor U19868 (N_19868,N_19000,N_19459);
or U19869 (N_19869,N_19406,N_19416);
nand U19870 (N_19870,N_19166,N_19127);
nor U19871 (N_19871,N_19331,N_19102);
or U19872 (N_19872,N_19189,N_19005);
or U19873 (N_19873,N_19490,N_19411);
nand U19874 (N_19874,N_19008,N_19424);
nand U19875 (N_19875,N_19451,N_19059);
nor U19876 (N_19876,N_19318,N_19019);
or U19877 (N_19877,N_19085,N_19220);
or U19878 (N_19878,N_19081,N_19243);
xor U19879 (N_19879,N_19005,N_19186);
nand U19880 (N_19880,N_19330,N_19425);
or U19881 (N_19881,N_19087,N_19000);
xnor U19882 (N_19882,N_19089,N_19352);
xnor U19883 (N_19883,N_19105,N_19380);
or U19884 (N_19884,N_19414,N_19020);
and U19885 (N_19885,N_19451,N_19052);
xor U19886 (N_19886,N_19144,N_19061);
or U19887 (N_19887,N_19470,N_19209);
nor U19888 (N_19888,N_19289,N_19254);
xnor U19889 (N_19889,N_19033,N_19143);
or U19890 (N_19890,N_19250,N_19376);
xnor U19891 (N_19891,N_19226,N_19171);
nor U19892 (N_19892,N_19016,N_19153);
and U19893 (N_19893,N_19017,N_19472);
or U19894 (N_19894,N_19442,N_19157);
nand U19895 (N_19895,N_19486,N_19394);
or U19896 (N_19896,N_19268,N_19091);
nor U19897 (N_19897,N_19453,N_19099);
or U19898 (N_19898,N_19262,N_19325);
nand U19899 (N_19899,N_19446,N_19362);
nor U19900 (N_19900,N_19107,N_19187);
xnor U19901 (N_19901,N_19493,N_19245);
and U19902 (N_19902,N_19391,N_19141);
nand U19903 (N_19903,N_19284,N_19367);
nand U19904 (N_19904,N_19124,N_19258);
nor U19905 (N_19905,N_19040,N_19470);
or U19906 (N_19906,N_19377,N_19208);
and U19907 (N_19907,N_19004,N_19272);
and U19908 (N_19908,N_19183,N_19408);
nand U19909 (N_19909,N_19309,N_19294);
or U19910 (N_19910,N_19413,N_19259);
nand U19911 (N_19911,N_19220,N_19403);
nand U19912 (N_19912,N_19143,N_19181);
nand U19913 (N_19913,N_19048,N_19458);
nor U19914 (N_19914,N_19219,N_19222);
nand U19915 (N_19915,N_19196,N_19261);
nor U19916 (N_19916,N_19424,N_19247);
and U19917 (N_19917,N_19437,N_19431);
nand U19918 (N_19918,N_19261,N_19055);
and U19919 (N_19919,N_19006,N_19299);
or U19920 (N_19920,N_19201,N_19164);
and U19921 (N_19921,N_19496,N_19230);
and U19922 (N_19922,N_19362,N_19449);
nor U19923 (N_19923,N_19396,N_19321);
or U19924 (N_19924,N_19292,N_19097);
nor U19925 (N_19925,N_19497,N_19351);
and U19926 (N_19926,N_19407,N_19415);
or U19927 (N_19927,N_19432,N_19184);
and U19928 (N_19928,N_19336,N_19152);
or U19929 (N_19929,N_19068,N_19420);
nor U19930 (N_19930,N_19048,N_19435);
xor U19931 (N_19931,N_19045,N_19223);
or U19932 (N_19932,N_19174,N_19278);
xnor U19933 (N_19933,N_19073,N_19314);
xor U19934 (N_19934,N_19111,N_19310);
xnor U19935 (N_19935,N_19010,N_19179);
nor U19936 (N_19936,N_19058,N_19428);
xor U19937 (N_19937,N_19074,N_19471);
or U19938 (N_19938,N_19020,N_19460);
nor U19939 (N_19939,N_19467,N_19299);
and U19940 (N_19940,N_19405,N_19251);
nand U19941 (N_19941,N_19211,N_19101);
or U19942 (N_19942,N_19307,N_19421);
or U19943 (N_19943,N_19377,N_19272);
or U19944 (N_19944,N_19013,N_19272);
and U19945 (N_19945,N_19357,N_19418);
and U19946 (N_19946,N_19042,N_19420);
or U19947 (N_19947,N_19228,N_19444);
nand U19948 (N_19948,N_19169,N_19065);
or U19949 (N_19949,N_19075,N_19255);
nor U19950 (N_19950,N_19268,N_19311);
xor U19951 (N_19951,N_19314,N_19206);
or U19952 (N_19952,N_19442,N_19096);
nor U19953 (N_19953,N_19339,N_19499);
or U19954 (N_19954,N_19394,N_19215);
and U19955 (N_19955,N_19339,N_19204);
or U19956 (N_19956,N_19242,N_19169);
or U19957 (N_19957,N_19360,N_19072);
xnor U19958 (N_19958,N_19166,N_19248);
or U19959 (N_19959,N_19193,N_19147);
xor U19960 (N_19960,N_19307,N_19435);
or U19961 (N_19961,N_19050,N_19221);
nand U19962 (N_19962,N_19082,N_19204);
xor U19963 (N_19963,N_19130,N_19364);
and U19964 (N_19964,N_19461,N_19398);
or U19965 (N_19965,N_19355,N_19304);
nand U19966 (N_19966,N_19109,N_19307);
nor U19967 (N_19967,N_19146,N_19249);
nand U19968 (N_19968,N_19145,N_19293);
nand U19969 (N_19969,N_19238,N_19065);
xor U19970 (N_19970,N_19295,N_19025);
nand U19971 (N_19971,N_19095,N_19327);
and U19972 (N_19972,N_19053,N_19398);
and U19973 (N_19973,N_19248,N_19289);
xnor U19974 (N_19974,N_19264,N_19231);
nand U19975 (N_19975,N_19386,N_19060);
and U19976 (N_19976,N_19323,N_19056);
and U19977 (N_19977,N_19394,N_19488);
or U19978 (N_19978,N_19367,N_19438);
or U19979 (N_19979,N_19399,N_19472);
nor U19980 (N_19980,N_19342,N_19129);
xnor U19981 (N_19981,N_19289,N_19468);
xnor U19982 (N_19982,N_19347,N_19069);
or U19983 (N_19983,N_19383,N_19074);
xor U19984 (N_19984,N_19224,N_19470);
or U19985 (N_19985,N_19274,N_19480);
and U19986 (N_19986,N_19094,N_19374);
nand U19987 (N_19987,N_19198,N_19159);
and U19988 (N_19988,N_19378,N_19049);
and U19989 (N_19989,N_19118,N_19035);
nor U19990 (N_19990,N_19028,N_19335);
or U19991 (N_19991,N_19394,N_19137);
or U19992 (N_19992,N_19239,N_19234);
nor U19993 (N_19993,N_19439,N_19302);
or U19994 (N_19994,N_19370,N_19483);
and U19995 (N_19995,N_19278,N_19352);
nand U19996 (N_19996,N_19200,N_19328);
or U19997 (N_19997,N_19051,N_19080);
nand U19998 (N_19998,N_19286,N_19278);
nor U19999 (N_19999,N_19110,N_19208);
xnor UO_0 (O_0,N_19669,N_19931);
xor UO_1 (O_1,N_19622,N_19711);
nor UO_2 (O_2,N_19876,N_19507);
and UO_3 (O_3,N_19524,N_19728);
nand UO_4 (O_4,N_19924,N_19839);
or UO_5 (O_5,N_19937,N_19883);
xor UO_6 (O_6,N_19988,N_19590);
or UO_7 (O_7,N_19872,N_19692);
nor UO_8 (O_8,N_19897,N_19849);
or UO_9 (O_9,N_19996,N_19782);
xnor UO_10 (O_10,N_19701,N_19861);
xnor UO_11 (O_11,N_19962,N_19573);
or UO_12 (O_12,N_19626,N_19617);
and UO_13 (O_13,N_19793,N_19623);
xor UO_14 (O_14,N_19655,N_19762);
nand UO_15 (O_15,N_19614,N_19824);
nand UO_16 (O_16,N_19856,N_19620);
and UO_17 (O_17,N_19994,N_19847);
nand UO_18 (O_18,N_19564,N_19645);
nor UO_19 (O_19,N_19726,N_19791);
and UO_20 (O_20,N_19775,N_19990);
nand UO_21 (O_21,N_19680,N_19739);
nand UO_22 (O_22,N_19902,N_19664);
nor UO_23 (O_23,N_19577,N_19826);
nand UO_24 (O_24,N_19621,N_19950);
or UO_25 (O_25,N_19991,N_19871);
xnor UO_26 (O_26,N_19596,N_19732);
and UO_27 (O_27,N_19607,N_19853);
xor UO_28 (O_28,N_19539,N_19820);
or UO_29 (O_29,N_19636,N_19979);
and UO_30 (O_30,N_19719,N_19867);
nor UO_31 (O_31,N_19699,N_19986);
or UO_32 (O_32,N_19689,N_19909);
and UO_33 (O_33,N_19709,N_19629);
nor UO_34 (O_34,N_19541,N_19803);
nand UO_35 (O_35,N_19521,N_19500);
nor UO_36 (O_36,N_19570,N_19850);
nor UO_37 (O_37,N_19748,N_19965);
and UO_38 (O_38,N_19956,N_19764);
xnor UO_39 (O_39,N_19684,N_19603);
nor UO_40 (O_40,N_19651,N_19890);
xnor UO_41 (O_41,N_19633,N_19835);
and UO_42 (O_42,N_19566,N_19503);
and UO_43 (O_43,N_19634,N_19823);
nand UO_44 (O_44,N_19722,N_19955);
nand UO_45 (O_45,N_19836,N_19501);
and UO_46 (O_46,N_19892,N_19553);
or UO_47 (O_47,N_19683,N_19885);
xnor UO_48 (O_48,N_19925,N_19713);
nand UO_49 (O_49,N_19825,N_19505);
or UO_50 (O_50,N_19877,N_19630);
or UO_51 (O_51,N_19884,N_19671);
xor UO_52 (O_52,N_19949,N_19720);
and UO_53 (O_53,N_19589,N_19679);
nand UO_54 (O_54,N_19543,N_19637);
or UO_55 (O_55,N_19646,N_19592);
and UO_56 (O_56,N_19518,N_19881);
nand UO_57 (O_57,N_19754,N_19802);
and UO_58 (O_58,N_19661,N_19591);
xnor UO_59 (O_59,N_19814,N_19790);
nand UO_60 (O_60,N_19960,N_19536);
nor UO_61 (O_61,N_19674,N_19611);
or UO_62 (O_62,N_19852,N_19992);
and UO_63 (O_63,N_19968,N_19773);
nand UO_64 (O_64,N_19615,N_19801);
xnor UO_65 (O_65,N_19690,N_19708);
and UO_66 (O_66,N_19586,N_19723);
xnor UO_67 (O_67,N_19567,N_19675);
nand UO_68 (O_68,N_19588,N_19602);
nand UO_69 (O_69,N_19941,N_19612);
nand UO_70 (O_70,N_19783,N_19687);
nor UO_71 (O_71,N_19800,N_19542);
nand UO_72 (O_72,N_19917,N_19788);
and UO_73 (O_73,N_19627,N_19812);
and UO_74 (O_74,N_19742,N_19842);
or UO_75 (O_75,N_19923,N_19863);
nor UO_76 (O_76,N_19747,N_19868);
or UO_77 (O_77,N_19795,N_19625);
xnor UO_78 (O_78,N_19963,N_19854);
xor UO_79 (O_79,N_19668,N_19736);
nor UO_80 (O_80,N_19753,N_19695);
or UO_81 (O_81,N_19571,N_19656);
nand UO_82 (O_82,N_19860,N_19821);
nand UO_83 (O_83,N_19817,N_19658);
and UO_84 (O_84,N_19947,N_19880);
nor UO_85 (O_85,N_19616,N_19506);
nand UO_86 (O_86,N_19523,N_19927);
nand UO_87 (O_87,N_19584,N_19580);
xnor UO_88 (O_88,N_19828,N_19562);
nor UO_89 (O_89,N_19517,N_19557);
nor UO_90 (O_90,N_19918,N_19551);
nand UO_91 (O_91,N_19698,N_19933);
and UO_92 (O_92,N_19516,N_19705);
and UO_93 (O_93,N_19756,N_19948);
or UO_94 (O_94,N_19830,N_19741);
and UO_95 (O_95,N_19799,N_19903);
or UO_96 (O_96,N_19905,N_19600);
nor UO_97 (O_97,N_19743,N_19544);
nand UO_98 (O_98,N_19792,N_19766);
or UO_99 (O_99,N_19889,N_19982);
nand UO_100 (O_100,N_19976,N_19534);
or UO_101 (O_101,N_19575,N_19993);
and UO_102 (O_102,N_19735,N_19650);
nand UO_103 (O_103,N_19777,N_19998);
nand UO_104 (O_104,N_19789,N_19707);
xor UO_105 (O_105,N_19938,N_19961);
or UO_106 (O_106,N_19816,N_19632);
xor UO_107 (O_107,N_19599,N_19737);
nor UO_108 (O_108,N_19749,N_19638);
and UO_109 (O_109,N_19601,N_19914);
nor UO_110 (O_110,N_19797,N_19858);
or UO_111 (O_111,N_19921,N_19727);
nor UO_112 (O_112,N_19900,N_19840);
or UO_113 (O_113,N_19529,N_19606);
xor UO_114 (O_114,N_19581,N_19663);
nand UO_115 (O_115,N_19971,N_19647);
nor UO_116 (O_116,N_19966,N_19526);
or UO_117 (O_117,N_19718,N_19780);
or UO_118 (O_118,N_19696,N_19970);
xor UO_119 (O_119,N_19916,N_19846);
xor UO_120 (O_120,N_19869,N_19662);
nand UO_121 (O_121,N_19893,N_19710);
or UO_122 (O_122,N_19672,N_19745);
or UO_123 (O_123,N_19535,N_19659);
nand UO_124 (O_124,N_19832,N_19904);
nor UO_125 (O_125,N_19755,N_19700);
xnor UO_126 (O_126,N_19843,N_19932);
xnor UO_127 (O_127,N_19779,N_19653);
or UO_128 (O_128,N_19528,N_19583);
nor UO_129 (O_129,N_19978,N_19827);
and UO_130 (O_130,N_19758,N_19731);
xnor UO_131 (O_131,N_19578,N_19702);
nand UO_132 (O_132,N_19538,N_19572);
xor UO_133 (O_133,N_19746,N_19922);
nor UO_134 (O_134,N_19547,N_19935);
and UO_135 (O_135,N_19787,N_19857);
nand UO_136 (O_136,N_19587,N_19502);
nor UO_137 (O_137,N_19894,N_19714);
nand UO_138 (O_138,N_19886,N_19525);
xor UO_139 (O_139,N_19665,N_19763);
or UO_140 (O_140,N_19769,N_19810);
and UO_141 (O_141,N_19974,N_19652);
nor UO_142 (O_142,N_19644,N_19997);
xor UO_143 (O_143,N_19911,N_19555);
nor UO_144 (O_144,N_19530,N_19765);
or UO_145 (O_145,N_19818,N_19729);
nand UO_146 (O_146,N_19673,N_19648);
xnor UO_147 (O_147,N_19660,N_19907);
xor UO_148 (O_148,N_19569,N_19838);
nor UO_149 (O_149,N_19759,N_19510);
nor UO_150 (O_150,N_19608,N_19981);
nand UO_151 (O_151,N_19896,N_19781);
nor UO_152 (O_152,N_19806,N_19550);
xnor UO_153 (O_153,N_19964,N_19940);
nor UO_154 (O_154,N_19953,N_19957);
nand UO_155 (O_155,N_19770,N_19666);
or UO_156 (O_156,N_19560,N_19667);
nor UO_157 (O_157,N_19715,N_19865);
and UO_158 (O_158,N_19678,N_19576);
and UO_159 (O_159,N_19942,N_19724);
or UO_160 (O_160,N_19685,N_19734);
xnor UO_161 (O_161,N_19631,N_19855);
or UO_162 (O_162,N_19604,N_19595);
and UO_163 (O_163,N_19784,N_19563);
or UO_164 (O_164,N_19899,N_19951);
nand UO_165 (O_165,N_19831,N_19598);
and UO_166 (O_166,N_19624,N_19859);
or UO_167 (O_167,N_19813,N_19643);
xor UO_168 (O_168,N_19805,N_19509);
xnor UO_169 (O_169,N_19677,N_19767);
nor UO_170 (O_170,N_19654,N_19717);
and UO_171 (O_171,N_19670,N_19874);
nand UO_172 (O_172,N_19833,N_19969);
xor UO_173 (O_173,N_19511,N_19915);
and UO_174 (O_174,N_19681,N_19841);
and UO_175 (O_175,N_19987,N_19697);
and UO_176 (O_176,N_19768,N_19559);
nor UO_177 (O_177,N_19794,N_19891);
or UO_178 (O_178,N_19778,N_19504);
nand UO_179 (O_179,N_19887,N_19989);
and UO_180 (O_180,N_19808,N_19983);
xor UO_181 (O_181,N_19558,N_19597);
or UO_182 (O_182,N_19657,N_19811);
nor UO_183 (O_183,N_19878,N_19546);
xnor UO_184 (O_184,N_19848,N_19751);
nor UO_185 (O_185,N_19774,N_19930);
xor UO_186 (O_186,N_19527,N_19515);
nand UO_187 (O_187,N_19552,N_19958);
nand UO_188 (O_188,N_19613,N_19815);
or UO_189 (O_189,N_19760,N_19798);
nor UO_190 (O_190,N_19866,N_19879);
or UO_191 (O_191,N_19906,N_19785);
and UO_192 (O_192,N_19642,N_19875);
and UO_193 (O_193,N_19786,N_19628);
and UO_194 (O_194,N_19761,N_19531);
xnor UO_195 (O_195,N_19776,N_19733);
or UO_196 (O_196,N_19508,N_19851);
xnor UO_197 (O_197,N_19640,N_19554);
or UO_198 (O_198,N_19944,N_19999);
nor UO_199 (O_199,N_19834,N_19936);
and UO_200 (O_200,N_19959,N_19712);
nand UO_201 (O_201,N_19972,N_19888);
or UO_202 (O_202,N_19882,N_19556);
or UO_203 (O_203,N_19946,N_19740);
nand UO_204 (O_204,N_19837,N_19561);
and UO_205 (O_205,N_19537,N_19919);
or UO_206 (O_206,N_19738,N_19618);
nor UO_207 (O_207,N_19934,N_19594);
or UO_208 (O_208,N_19549,N_19574);
nand UO_209 (O_209,N_19895,N_19829);
xor UO_210 (O_210,N_19864,N_19752);
or UO_211 (O_211,N_19721,N_19635);
or UO_212 (O_212,N_19582,N_19926);
nor UO_213 (O_213,N_19920,N_19977);
and UO_214 (O_214,N_19519,N_19822);
nand UO_215 (O_215,N_19706,N_19725);
nor UO_216 (O_216,N_19844,N_19682);
xor UO_217 (O_217,N_19513,N_19639);
or UO_218 (O_218,N_19676,N_19512);
nor UO_219 (O_219,N_19796,N_19744);
or UO_220 (O_220,N_19862,N_19532);
or UO_221 (O_221,N_19688,N_19730);
and UO_222 (O_222,N_19514,N_19954);
and UO_223 (O_223,N_19975,N_19804);
nand UO_224 (O_224,N_19704,N_19703);
or UO_225 (O_225,N_19540,N_19649);
xnor UO_226 (O_226,N_19819,N_19910);
and UO_227 (O_227,N_19929,N_19912);
nand UO_228 (O_228,N_19610,N_19522);
nand UO_229 (O_229,N_19980,N_19995);
and UO_230 (O_230,N_19908,N_19716);
and UO_231 (O_231,N_19807,N_19809);
nor UO_232 (O_232,N_19913,N_19693);
and UO_233 (O_233,N_19694,N_19641);
or UO_234 (O_234,N_19973,N_19928);
or UO_235 (O_235,N_19605,N_19548);
and UO_236 (O_236,N_19772,N_19943);
xor UO_237 (O_237,N_19609,N_19691);
and UO_238 (O_238,N_19901,N_19585);
xnor UO_239 (O_239,N_19568,N_19750);
nand UO_240 (O_240,N_19593,N_19967);
and UO_241 (O_241,N_19873,N_19945);
and UO_242 (O_242,N_19984,N_19771);
nor UO_243 (O_243,N_19845,N_19898);
nor UO_244 (O_244,N_19985,N_19757);
xor UO_245 (O_245,N_19870,N_19545);
xor UO_246 (O_246,N_19619,N_19533);
nor UO_247 (O_247,N_19686,N_19565);
nand UO_248 (O_248,N_19952,N_19520);
nor UO_249 (O_249,N_19939,N_19579);
nand UO_250 (O_250,N_19661,N_19685);
and UO_251 (O_251,N_19850,N_19953);
nor UO_252 (O_252,N_19572,N_19727);
nor UO_253 (O_253,N_19505,N_19943);
nand UO_254 (O_254,N_19952,N_19760);
and UO_255 (O_255,N_19921,N_19809);
and UO_256 (O_256,N_19519,N_19790);
xnor UO_257 (O_257,N_19981,N_19914);
and UO_258 (O_258,N_19931,N_19984);
xnor UO_259 (O_259,N_19631,N_19600);
or UO_260 (O_260,N_19560,N_19803);
nor UO_261 (O_261,N_19609,N_19587);
xnor UO_262 (O_262,N_19892,N_19519);
nand UO_263 (O_263,N_19620,N_19876);
nand UO_264 (O_264,N_19630,N_19512);
or UO_265 (O_265,N_19541,N_19704);
or UO_266 (O_266,N_19598,N_19908);
nor UO_267 (O_267,N_19854,N_19862);
nand UO_268 (O_268,N_19615,N_19689);
nand UO_269 (O_269,N_19586,N_19775);
nor UO_270 (O_270,N_19589,N_19929);
nor UO_271 (O_271,N_19787,N_19719);
and UO_272 (O_272,N_19792,N_19500);
nand UO_273 (O_273,N_19860,N_19739);
or UO_274 (O_274,N_19966,N_19584);
nor UO_275 (O_275,N_19910,N_19814);
xor UO_276 (O_276,N_19650,N_19585);
nand UO_277 (O_277,N_19880,N_19996);
xor UO_278 (O_278,N_19808,N_19556);
nand UO_279 (O_279,N_19901,N_19709);
nor UO_280 (O_280,N_19662,N_19506);
or UO_281 (O_281,N_19588,N_19697);
nand UO_282 (O_282,N_19865,N_19749);
and UO_283 (O_283,N_19569,N_19576);
xor UO_284 (O_284,N_19797,N_19740);
nor UO_285 (O_285,N_19958,N_19878);
and UO_286 (O_286,N_19660,N_19590);
and UO_287 (O_287,N_19842,N_19961);
nand UO_288 (O_288,N_19511,N_19903);
or UO_289 (O_289,N_19595,N_19866);
nor UO_290 (O_290,N_19917,N_19927);
nand UO_291 (O_291,N_19805,N_19680);
xor UO_292 (O_292,N_19997,N_19717);
nand UO_293 (O_293,N_19696,N_19644);
and UO_294 (O_294,N_19530,N_19904);
or UO_295 (O_295,N_19627,N_19981);
or UO_296 (O_296,N_19505,N_19889);
nor UO_297 (O_297,N_19960,N_19998);
and UO_298 (O_298,N_19562,N_19982);
and UO_299 (O_299,N_19664,N_19642);
nand UO_300 (O_300,N_19761,N_19646);
xnor UO_301 (O_301,N_19807,N_19530);
xnor UO_302 (O_302,N_19938,N_19945);
nor UO_303 (O_303,N_19821,N_19996);
nand UO_304 (O_304,N_19563,N_19606);
and UO_305 (O_305,N_19773,N_19618);
or UO_306 (O_306,N_19966,N_19802);
or UO_307 (O_307,N_19754,N_19668);
nor UO_308 (O_308,N_19970,N_19856);
nor UO_309 (O_309,N_19639,N_19959);
xnor UO_310 (O_310,N_19788,N_19695);
nor UO_311 (O_311,N_19869,N_19643);
or UO_312 (O_312,N_19777,N_19930);
nand UO_313 (O_313,N_19618,N_19908);
or UO_314 (O_314,N_19770,N_19728);
or UO_315 (O_315,N_19883,N_19701);
xnor UO_316 (O_316,N_19985,N_19949);
and UO_317 (O_317,N_19877,N_19890);
xor UO_318 (O_318,N_19555,N_19755);
and UO_319 (O_319,N_19627,N_19718);
xnor UO_320 (O_320,N_19803,N_19716);
xor UO_321 (O_321,N_19511,N_19907);
and UO_322 (O_322,N_19578,N_19567);
xnor UO_323 (O_323,N_19821,N_19727);
nand UO_324 (O_324,N_19672,N_19949);
and UO_325 (O_325,N_19729,N_19881);
xnor UO_326 (O_326,N_19953,N_19807);
or UO_327 (O_327,N_19952,N_19649);
and UO_328 (O_328,N_19510,N_19508);
nand UO_329 (O_329,N_19677,N_19826);
xnor UO_330 (O_330,N_19854,N_19765);
xor UO_331 (O_331,N_19525,N_19536);
nand UO_332 (O_332,N_19752,N_19901);
nand UO_333 (O_333,N_19822,N_19700);
nand UO_334 (O_334,N_19696,N_19774);
and UO_335 (O_335,N_19643,N_19908);
xnor UO_336 (O_336,N_19669,N_19995);
or UO_337 (O_337,N_19804,N_19779);
or UO_338 (O_338,N_19680,N_19917);
and UO_339 (O_339,N_19629,N_19523);
xor UO_340 (O_340,N_19901,N_19620);
nand UO_341 (O_341,N_19693,N_19518);
nor UO_342 (O_342,N_19657,N_19880);
and UO_343 (O_343,N_19821,N_19920);
and UO_344 (O_344,N_19954,N_19562);
and UO_345 (O_345,N_19948,N_19729);
nand UO_346 (O_346,N_19817,N_19575);
xnor UO_347 (O_347,N_19749,N_19693);
nor UO_348 (O_348,N_19933,N_19952);
nor UO_349 (O_349,N_19878,N_19777);
and UO_350 (O_350,N_19710,N_19805);
or UO_351 (O_351,N_19708,N_19631);
xor UO_352 (O_352,N_19914,N_19755);
nand UO_353 (O_353,N_19712,N_19722);
and UO_354 (O_354,N_19711,N_19887);
nor UO_355 (O_355,N_19590,N_19573);
xor UO_356 (O_356,N_19553,N_19861);
xor UO_357 (O_357,N_19732,N_19804);
nor UO_358 (O_358,N_19690,N_19838);
nand UO_359 (O_359,N_19757,N_19815);
nor UO_360 (O_360,N_19904,N_19623);
and UO_361 (O_361,N_19850,N_19848);
or UO_362 (O_362,N_19666,N_19835);
nand UO_363 (O_363,N_19742,N_19559);
or UO_364 (O_364,N_19777,N_19879);
or UO_365 (O_365,N_19600,N_19636);
or UO_366 (O_366,N_19831,N_19917);
or UO_367 (O_367,N_19763,N_19547);
xnor UO_368 (O_368,N_19643,N_19520);
nand UO_369 (O_369,N_19999,N_19998);
or UO_370 (O_370,N_19584,N_19776);
and UO_371 (O_371,N_19672,N_19941);
nor UO_372 (O_372,N_19842,N_19597);
xor UO_373 (O_373,N_19922,N_19992);
nor UO_374 (O_374,N_19902,N_19515);
xnor UO_375 (O_375,N_19919,N_19981);
nand UO_376 (O_376,N_19766,N_19917);
or UO_377 (O_377,N_19620,N_19969);
nor UO_378 (O_378,N_19548,N_19932);
and UO_379 (O_379,N_19710,N_19771);
xor UO_380 (O_380,N_19534,N_19575);
or UO_381 (O_381,N_19755,N_19539);
nand UO_382 (O_382,N_19896,N_19613);
nor UO_383 (O_383,N_19647,N_19692);
nor UO_384 (O_384,N_19732,N_19650);
or UO_385 (O_385,N_19514,N_19899);
nand UO_386 (O_386,N_19930,N_19510);
nor UO_387 (O_387,N_19642,N_19707);
nor UO_388 (O_388,N_19714,N_19977);
nor UO_389 (O_389,N_19828,N_19676);
xnor UO_390 (O_390,N_19734,N_19736);
or UO_391 (O_391,N_19719,N_19722);
or UO_392 (O_392,N_19562,N_19991);
or UO_393 (O_393,N_19529,N_19755);
nor UO_394 (O_394,N_19924,N_19866);
xor UO_395 (O_395,N_19651,N_19542);
xor UO_396 (O_396,N_19872,N_19658);
xor UO_397 (O_397,N_19557,N_19573);
nor UO_398 (O_398,N_19848,N_19754);
nor UO_399 (O_399,N_19931,N_19784);
nor UO_400 (O_400,N_19740,N_19529);
nor UO_401 (O_401,N_19655,N_19888);
and UO_402 (O_402,N_19559,N_19642);
or UO_403 (O_403,N_19680,N_19542);
nor UO_404 (O_404,N_19862,N_19989);
nand UO_405 (O_405,N_19503,N_19608);
or UO_406 (O_406,N_19995,N_19649);
and UO_407 (O_407,N_19828,N_19618);
nor UO_408 (O_408,N_19721,N_19943);
and UO_409 (O_409,N_19946,N_19695);
or UO_410 (O_410,N_19697,N_19919);
or UO_411 (O_411,N_19906,N_19724);
nand UO_412 (O_412,N_19749,N_19533);
nor UO_413 (O_413,N_19544,N_19796);
and UO_414 (O_414,N_19816,N_19542);
nand UO_415 (O_415,N_19640,N_19696);
or UO_416 (O_416,N_19885,N_19875);
nand UO_417 (O_417,N_19750,N_19527);
nand UO_418 (O_418,N_19644,N_19699);
nor UO_419 (O_419,N_19856,N_19780);
nand UO_420 (O_420,N_19957,N_19608);
or UO_421 (O_421,N_19611,N_19691);
nor UO_422 (O_422,N_19795,N_19504);
and UO_423 (O_423,N_19670,N_19762);
nor UO_424 (O_424,N_19574,N_19729);
or UO_425 (O_425,N_19559,N_19517);
nor UO_426 (O_426,N_19524,N_19787);
xnor UO_427 (O_427,N_19700,N_19760);
nor UO_428 (O_428,N_19898,N_19719);
nor UO_429 (O_429,N_19637,N_19626);
or UO_430 (O_430,N_19955,N_19905);
nor UO_431 (O_431,N_19797,N_19893);
nor UO_432 (O_432,N_19929,N_19590);
nand UO_433 (O_433,N_19697,N_19944);
or UO_434 (O_434,N_19723,N_19502);
or UO_435 (O_435,N_19564,N_19966);
nor UO_436 (O_436,N_19999,N_19908);
and UO_437 (O_437,N_19746,N_19916);
or UO_438 (O_438,N_19682,N_19821);
nand UO_439 (O_439,N_19844,N_19567);
nand UO_440 (O_440,N_19747,N_19653);
xnor UO_441 (O_441,N_19704,N_19523);
nor UO_442 (O_442,N_19986,N_19779);
nor UO_443 (O_443,N_19663,N_19818);
and UO_444 (O_444,N_19844,N_19803);
nand UO_445 (O_445,N_19797,N_19957);
xor UO_446 (O_446,N_19672,N_19784);
or UO_447 (O_447,N_19954,N_19528);
and UO_448 (O_448,N_19820,N_19764);
nand UO_449 (O_449,N_19992,N_19856);
and UO_450 (O_450,N_19737,N_19543);
nor UO_451 (O_451,N_19897,N_19674);
or UO_452 (O_452,N_19929,N_19562);
and UO_453 (O_453,N_19954,N_19745);
and UO_454 (O_454,N_19599,N_19979);
nor UO_455 (O_455,N_19848,N_19963);
nor UO_456 (O_456,N_19788,N_19771);
and UO_457 (O_457,N_19519,N_19835);
nor UO_458 (O_458,N_19612,N_19898);
or UO_459 (O_459,N_19509,N_19784);
xor UO_460 (O_460,N_19520,N_19788);
xor UO_461 (O_461,N_19663,N_19743);
or UO_462 (O_462,N_19761,N_19767);
nand UO_463 (O_463,N_19895,N_19574);
or UO_464 (O_464,N_19895,N_19722);
and UO_465 (O_465,N_19765,N_19950);
xor UO_466 (O_466,N_19550,N_19961);
nor UO_467 (O_467,N_19906,N_19702);
or UO_468 (O_468,N_19686,N_19760);
or UO_469 (O_469,N_19843,N_19845);
nand UO_470 (O_470,N_19506,N_19923);
nor UO_471 (O_471,N_19734,N_19501);
xnor UO_472 (O_472,N_19985,N_19951);
nand UO_473 (O_473,N_19612,N_19685);
or UO_474 (O_474,N_19947,N_19969);
or UO_475 (O_475,N_19997,N_19836);
nor UO_476 (O_476,N_19670,N_19714);
and UO_477 (O_477,N_19734,N_19716);
nor UO_478 (O_478,N_19621,N_19522);
nand UO_479 (O_479,N_19532,N_19748);
xnor UO_480 (O_480,N_19711,N_19835);
nor UO_481 (O_481,N_19935,N_19613);
and UO_482 (O_482,N_19746,N_19627);
or UO_483 (O_483,N_19696,N_19595);
xor UO_484 (O_484,N_19510,N_19910);
and UO_485 (O_485,N_19707,N_19967);
nand UO_486 (O_486,N_19932,N_19532);
nand UO_487 (O_487,N_19507,N_19969);
or UO_488 (O_488,N_19776,N_19813);
xor UO_489 (O_489,N_19958,N_19866);
nor UO_490 (O_490,N_19982,N_19672);
and UO_491 (O_491,N_19532,N_19872);
xor UO_492 (O_492,N_19556,N_19609);
nor UO_493 (O_493,N_19622,N_19952);
xnor UO_494 (O_494,N_19995,N_19799);
xor UO_495 (O_495,N_19826,N_19601);
nor UO_496 (O_496,N_19835,N_19720);
nand UO_497 (O_497,N_19929,N_19577);
nand UO_498 (O_498,N_19714,N_19824);
xor UO_499 (O_499,N_19886,N_19640);
nand UO_500 (O_500,N_19571,N_19812);
xor UO_501 (O_501,N_19946,N_19729);
nor UO_502 (O_502,N_19870,N_19705);
and UO_503 (O_503,N_19967,N_19876);
nor UO_504 (O_504,N_19843,N_19614);
nor UO_505 (O_505,N_19793,N_19527);
and UO_506 (O_506,N_19595,N_19892);
and UO_507 (O_507,N_19829,N_19537);
or UO_508 (O_508,N_19946,N_19909);
nor UO_509 (O_509,N_19716,N_19976);
nor UO_510 (O_510,N_19566,N_19786);
nor UO_511 (O_511,N_19872,N_19924);
xor UO_512 (O_512,N_19584,N_19939);
xnor UO_513 (O_513,N_19797,N_19801);
and UO_514 (O_514,N_19514,N_19936);
xor UO_515 (O_515,N_19952,N_19601);
or UO_516 (O_516,N_19656,N_19867);
nor UO_517 (O_517,N_19936,N_19809);
nor UO_518 (O_518,N_19634,N_19837);
nor UO_519 (O_519,N_19617,N_19713);
and UO_520 (O_520,N_19934,N_19665);
nor UO_521 (O_521,N_19928,N_19594);
or UO_522 (O_522,N_19659,N_19731);
xnor UO_523 (O_523,N_19593,N_19975);
nor UO_524 (O_524,N_19788,N_19764);
or UO_525 (O_525,N_19547,N_19984);
nor UO_526 (O_526,N_19611,N_19870);
xor UO_527 (O_527,N_19795,N_19884);
nor UO_528 (O_528,N_19950,N_19662);
nor UO_529 (O_529,N_19623,N_19509);
and UO_530 (O_530,N_19982,N_19941);
nand UO_531 (O_531,N_19647,N_19703);
nand UO_532 (O_532,N_19986,N_19615);
or UO_533 (O_533,N_19866,N_19881);
nand UO_534 (O_534,N_19583,N_19960);
xnor UO_535 (O_535,N_19695,N_19771);
nor UO_536 (O_536,N_19547,N_19526);
nor UO_537 (O_537,N_19826,N_19673);
and UO_538 (O_538,N_19626,N_19894);
nand UO_539 (O_539,N_19531,N_19724);
xnor UO_540 (O_540,N_19764,N_19564);
or UO_541 (O_541,N_19603,N_19524);
and UO_542 (O_542,N_19574,N_19857);
or UO_543 (O_543,N_19745,N_19569);
nor UO_544 (O_544,N_19721,N_19898);
and UO_545 (O_545,N_19587,N_19917);
nand UO_546 (O_546,N_19682,N_19764);
nand UO_547 (O_547,N_19896,N_19709);
xor UO_548 (O_548,N_19828,N_19843);
and UO_549 (O_549,N_19702,N_19604);
xnor UO_550 (O_550,N_19672,N_19963);
nand UO_551 (O_551,N_19574,N_19870);
nand UO_552 (O_552,N_19968,N_19820);
xnor UO_553 (O_553,N_19820,N_19646);
xnor UO_554 (O_554,N_19844,N_19845);
or UO_555 (O_555,N_19750,N_19871);
xnor UO_556 (O_556,N_19662,N_19907);
nor UO_557 (O_557,N_19674,N_19966);
nor UO_558 (O_558,N_19728,N_19584);
nand UO_559 (O_559,N_19680,N_19584);
nor UO_560 (O_560,N_19711,N_19982);
nor UO_561 (O_561,N_19514,N_19631);
nor UO_562 (O_562,N_19641,N_19982);
and UO_563 (O_563,N_19720,N_19787);
nor UO_564 (O_564,N_19965,N_19523);
xor UO_565 (O_565,N_19808,N_19745);
xnor UO_566 (O_566,N_19901,N_19757);
xnor UO_567 (O_567,N_19920,N_19997);
and UO_568 (O_568,N_19897,N_19728);
xnor UO_569 (O_569,N_19592,N_19927);
nand UO_570 (O_570,N_19843,N_19547);
nor UO_571 (O_571,N_19737,N_19644);
nand UO_572 (O_572,N_19553,N_19922);
nor UO_573 (O_573,N_19719,N_19501);
or UO_574 (O_574,N_19766,N_19935);
xnor UO_575 (O_575,N_19687,N_19840);
xor UO_576 (O_576,N_19697,N_19632);
or UO_577 (O_577,N_19888,N_19837);
and UO_578 (O_578,N_19570,N_19987);
nor UO_579 (O_579,N_19814,N_19544);
and UO_580 (O_580,N_19656,N_19617);
xnor UO_581 (O_581,N_19899,N_19609);
nand UO_582 (O_582,N_19857,N_19527);
xor UO_583 (O_583,N_19944,N_19604);
nor UO_584 (O_584,N_19965,N_19605);
xor UO_585 (O_585,N_19589,N_19548);
nor UO_586 (O_586,N_19861,N_19570);
and UO_587 (O_587,N_19705,N_19933);
and UO_588 (O_588,N_19550,N_19653);
nand UO_589 (O_589,N_19802,N_19995);
or UO_590 (O_590,N_19809,N_19796);
or UO_591 (O_591,N_19520,N_19821);
xor UO_592 (O_592,N_19514,N_19798);
nor UO_593 (O_593,N_19671,N_19822);
and UO_594 (O_594,N_19567,N_19965);
xor UO_595 (O_595,N_19830,N_19807);
nand UO_596 (O_596,N_19948,N_19941);
nor UO_597 (O_597,N_19895,N_19508);
xnor UO_598 (O_598,N_19579,N_19974);
nand UO_599 (O_599,N_19516,N_19680);
and UO_600 (O_600,N_19630,N_19594);
and UO_601 (O_601,N_19571,N_19980);
nor UO_602 (O_602,N_19611,N_19578);
and UO_603 (O_603,N_19608,N_19690);
and UO_604 (O_604,N_19550,N_19883);
and UO_605 (O_605,N_19963,N_19505);
nor UO_606 (O_606,N_19590,N_19685);
and UO_607 (O_607,N_19748,N_19525);
xnor UO_608 (O_608,N_19585,N_19624);
nor UO_609 (O_609,N_19774,N_19569);
or UO_610 (O_610,N_19979,N_19691);
nand UO_611 (O_611,N_19906,N_19510);
nand UO_612 (O_612,N_19986,N_19571);
nor UO_613 (O_613,N_19532,N_19826);
nand UO_614 (O_614,N_19885,N_19798);
xor UO_615 (O_615,N_19966,N_19984);
nor UO_616 (O_616,N_19977,N_19606);
nand UO_617 (O_617,N_19721,N_19792);
and UO_618 (O_618,N_19945,N_19842);
or UO_619 (O_619,N_19733,N_19871);
nand UO_620 (O_620,N_19893,N_19642);
or UO_621 (O_621,N_19658,N_19735);
or UO_622 (O_622,N_19511,N_19965);
and UO_623 (O_623,N_19914,N_19882);
nand UO_624 (O_624,N_19549,N_19960);
or UO_625 (O_625,N_19926,N_19765);
or UO_626 (O_626,N_19949,N_19786);
xnor UO_627 (O_627,N_19574,N_19530);
nand UO_628 (O_628,N_19828,N_19912);
nand UO_629 (O_629,N_19939,N_19630);
nor UO_630 (O_630,N_19855,N_19615);
or UO_631 (O_631,N_19643,N_19983);
or UO_632 (O_632,N_19633,N_19979);
xor UO_633 (O_633,N_19528,N_19587);
nand UO_634 (O_634,N_19526,N_19525);
and UO_635 (O_635,N_19575,N_19830);
xnor UO_636 (O_636,N_19563,N_19673);
nor UO_637 (O_637,N_19510,N_19899);
or UO_638 (O_638,N_19910,N_19827);
nand UO_639 (O_639,N_19564,N_19900);
or UO_640 (O_640,N_19869,N_19529);
nand UO_641 (O_641,N_19670,N_19598);
and UO_642 (O_642,N_19987,N_19958);
and UO_643 (O_643,N_19654,N_19743);
or UO_644 (O_644,N_19875,N_19641);
xor UO_645 (O_645,N_19746,N_19598);
and UO_646 (O_646,N_19993,N_19956);
nor UO_647 (O_647,N_19614,N_19766);
or UO_648 (O_648,N_19647,N_19584);
nand UO_649 (O_649,N_19987,N_19935);
nor UO_650 (O_650,N_19870,N_19504);
and UO_651 (O_651,N_19894,N_19928);
or UO_652 (O_652,N_19617,N_19812);
nor UO_653 (O_653,N_19780,N_19683);
nor UO_654 (O_654,N_19838,N_19853);
and UO_655 (O_655,N_19534,N_19821);
nand UO_656 (O_656,N_19992,N_19594);
nand UO_657 (O_657,N_19507,N_19553);
nor UO_658 (O_658,N_19546,N_19725);
or UO_659 (O_659,N_19836,N_19820);
and UO_660 (O_660,N_19512,N_19716);
nor UO_661 (O_661,N_19675,N_19502);
nand UO_662 (O_662,N_19815,N_19680);
nand UO_663 (O_663,N_19889,N_19938);
nand UO_664 (O_664,N_19692,N_19547);
and UO_665 (O_665,N_19656,N_19992);
or UO_666 (O_666,N_19613,N_19839);
and UO_667 (O_667,N_19876,N_19542);
or UO_668 (O_668,N_19648,N_19714);
nor UO_669 (O_669,N_19873,N_19547);
nand UO_670 (O_670,N_19836,N_19996);
xor UO_671 (O_671,N_19721,N_19665);
nand UO_672 (O_672,N_19750,N_19649);
and UO_673 (O_673,N_19982,N_19535);
and UO_674 (O_674,N_19843,N_19673);
nor UO_675 (O_675,N_19846,N_19546);
and UO_676 (O_676,N_19836,N_19764);
and UO_677 (O_677,N_19575,N_19949);
or UO_678 (O_678,N_19734,N_19965);
or UO_679 (O_679,N_19968,N_19897);
xnor UO_680 (O_680,N_19784,N_19621);
xor UO_681 (O_681,N_19513,N_19935);
or UO_682 (O_682,N_19814,N_19798);
nor UO_683 (O_683,N_19900,N_19978);
nor UO_684 (O_684,N_19740,N_19775);
and UO_685 (O_685,N_19836,N_19974);
and UO_686 (O_686,N_19526,N_19538);
xnor UO_687 (O_687,N_19643,N_19513);
or UO_688 (O_688,N_19623,N_19891);
xor UO_689 (O_689,N_19575,N_19645);
and UO_690 (O_690,N_19939,N_19603);
and UO_691 (O_691,N_19871,N_19710);
or UO_692 (O_692,N_19712,N_19676);
nor UO_693 (O_693,N_19550,N_19608);
nor UO_694 (O_694,N_19918,N_19895);
nand UO_695 (O_695,N_19709,N_19747);
nand UO_696 (O_696,N_19882,N_19943);
or UO_697 (O_697,N_19916,N_19791);
or UO_698 (O_698,N_19534,N_19636);
and UO_699 (O_699,N_19799,N_19645);
and UO_700 (O_700,N_19657,N_19763);
or UO_701 (O_701,N_19797,N_19573);
and UO_702 (O_702,N_19652,N_19955);
and UO_703 (O_703,N_19806,N_19612);
nor UO_704 (O_704,N_19918,N_19519);
and UO_705 (O_705,N_19770,N_19988);
and UO_706 (O_706,N_19631,N_19836);
and UO_707 (O_707,N_19691,N_19684);
and UO_708 (O_708,N_19593,N_19506);
nand UO_709 (O_709,N_19985,N_19990);
nand UO_710 (O_710,N_19820,N_19521);
nor UO_711 (O_711,N_19924,N_19601);
nor UO_712 (O_712,N_19587,N_19963);
and UO_713 (O_713,N_19728,N_19864);
and UO_714 (O_714,N_19669,N_19956);
or UO_715 (O_715,N_19588,N_19773);
nor UO_716 (O_716,N_19675,N_19727);
nand UO_717 (O_717,N_19774,N_19851);
and UO_718 (O_718,N_19790,N_19808);
nor UO_719 (O_719,N_19574,N_19715);
xnor UO_720 (O_720,N_19764,N_19983);
nand UO_721 (O_721,N_19843,N_19504);
nand UO_722 (O_722,N_19632,N_19811);
nand UO_723 (O_723,N_19702,N_19932);
nand UO_724 (O_724,N_19971,N_19929);
nor UO_725 (O_725,N_19862,N_19642);
xor UO_726 (O_726,N_19811,N_19543);
and UO_727 (O_727,N_19639,N_19813);
xnor UO_728 (O_728,N_19887,N_19625);
or UO_729 (O_729,N_19805,N_19588);
xor UO_730 (O_730,N_19581,N_19582);
nand UO_731 (O_731,N_19953,N_19673);
nor UO_732 (O_732,N_19886,N_19709);
nand UO_733 (O_733,N_19574,N_19920);
or UO_734 (O_734,N_19569,N_19894);
and UO_735 (O_735,N_19991,N_19781);
or UO_736 (O_736,N_19919,N_19836);
nor UO_737 (O_737,N_19722,N_19780);
nand UO_738 (O_738,N_19598,N_19750);
or UO_739 (O_739,N_19947,N_19711);
and UO_740 (O_740,N_19866,N_19986);
xnor UO_741 (O_741,N_19521,N_19705);
nor UO_742 (O_742,N_19958,N_19689);
xnor UO_743 (O_743,N_19853,N_19868);
and UO_744 (O_744,N_19856,N_19761);
and UO_745 (O_745,N_19822,N_19535);
nand UO_746 (O_746,N_19763,N_19895);
or UO_747 (O_747,N_19607,N_19715);
and UO_748 (O_748,N_19900,N_19705);
xnor UO_749 (O_749,N_19624,N_19790);
nand UO_750 (O_750,N_19507,N_19574);
xnor UO_751 (O_751,N_19633,N_19919);
nor UO_752 (O_752,N_19886,N_19923);
nand UO_753 (O_753,N_19710,N_19786);
xor UO_754 (O_754,N_19799,N_19874);
nand UO_755 (O_755,N_19604,N_19845);
nor UO_756 (O_756,N_19504,N_19708);
nor UO_757 (O_757,N_19632,N_19589);
nor UO_758 (O_758,N_19624,N_19687);
nor UO_759 (O_759,N_19678,N_19890);
and UO_760 (O_760,N_19767,N_19603);
and UO_761 (O_761,N_19514,N_19616);
or UO_762 (O_762,N_19701,N_19702);
and UO_763 (O_763,N_19909,N_19826);
nand UO_764 (O_764,N_19598,N_19936);
or UO_765 (O_765,N_19975,N_19649);
and UO_766 (O_766,N_19691,N_19956);
nand UO_767 (O_767,N_19911,N_19761);
xor UO_768 (O_768,N_19720,N_19986);
xor UO_769 (O_769,N_19790,N_19911);
or UO_770 (O_770,N_19835,N_19535);
nor UO_771 (O_771,N_19924,N_19834);
or UO_772 (O_772,N_19869,N_19782);
and UO_773 (O_773,N_19576,N_19725);
and UO_774 (O_774,N_19618,N_19910);
nor UO_775 (O_775,N_19804,N_19714);
nand UO_776 (O_776,N_19622,N_19908);
xnor UO_777 (O_777,N_19836,N_19970);
nor UO_778 (O_778,N_19648,N_19601);
and UO_779 (O_779,N_19856,N_19518);
or UO_780 (O_780,N_19960,N_19573);
xor UO_781 (O_781,N_19642,N_19775);
and UO_782 (O_782,N_19834,N_19591);
or UO_783 (O_783,N_19577,N_19540);
xor UO_784 (O_784,N_19623,N_19749);
and UO_785 (O_785,N_19507,N_19572);
xnor UO_786 (O_786,N_19617,N_19673);
nor UO_787 (O_787,N_19565,N_19880);
and UO_788 (O_788,N_19822,N_19921);
nor UO_789 (O_789,N_19761,N_19837);
nor UO_790 (O_790,N_19663,N_19610);
nor UO_791 (O_791,N_19972,N_19890);
xor UO_792 (O_792,N_19637,N_19995);
nor UO_793 (O_793,N_19834,N_19598);
nand UO_794 (O_794,N_19713,N_19627);
and UO_795 (O_795,N_19575,N_19718);
and UO_796 (O_796,N_19905,N_19759);
and UO_797 (O_797,N_19718,N_19733);
or UO_798 (O_798,N_19641,N_19770);
and UO_799 (O_799,N_19558,N_19512);
and UO_800 (O_800,N_19659,N_19792);
or UO_801 (O_801,N_19938,N_19627);
xor UO_802 (O_802,N_19953,N_19504);
and UO_803 (O_803,N_19617,N_19540);
xnor UO_804 (O_804,N_19539,N_19878);
nand UO_805 (O_805,N_19825,N_19668);
or UO_806 (O_806,N_19808,N_19585);
xnor UO_807 (O_807,N_19819,N_19766);
nand UO_808 (O_808,N_19942,N_19888);
or UO_809 (O_809,N_19995,N_19927);
nand UO_810 (O_810,N_19535,N_19721);
and UO_811 (O_811,N_19816,N_19847);
or UO_812 (O_812,N_19599,N_19960);
nand UO_813 (O_813,N_19587,N_19983);
or UO_814 (O_814,N_19702,N_19704);
nand UO_815 (O_815,N_19642,N_19686);
nand UO_816 (O_816,N_19533,N_19963);
and UO_817 (O_817,N_19639,N_19923);
and UO_818 (O_818,N_19560,N_19697);
and UO_819 (O_819,N_19895,N_19540);
or UO_820 (O_820,N_19863,N_19948);
nor UO_821 (O_821,N_19769,N_19680);
xor UO_822 (O_822,N_19610,N_19509);
and UO_823 (O_823,N_19556,N_19966);
nand UO_824 (O_824,N_19737,N_19746);
and UO_825 (O_825,N_19901,N_19944);
or UO_826 (O_826,N_19654,N_19815);
nor UO_827 (O_827,N_19607,N_19943);
nand UO_828 (O_828,N_19589,N_19935);
xnor UO_829 (O_829,N_19622,N_19819);
and UO_830 (O_830,N_19961,N_19625);
nand UO_831 (O_831,N_19543,N_19542);
and UO_832 (O_832,N_19628,N_19565);
nor UO_833 (O_833,N_19543,N_19501);
and UO_834 (O_834,N_19771,N_19936);
or UO_835 (O_835,N_19598,N_19817);
xnor UO_836 (O_836,N_19911,N_19539);
or UO_837 (O_837,N_19615,N_19883);
and UO_838 (O_838,N_19970,N_19971);
xnor UO_839 (O_839,N_19850,N_19885);
and UO_840 (O_840,N_19971,N_19945);
xor UO_841 (O_841,N_19866,N_19853);
nand UO_842 (O_842,N_19764,N_19511);
nor UO_843 (O_843,N_19868,N_19511);
and UO_844 (O_844,N_19821,N_19970);
or UO_845 (O_845,N_19643,N_19673);
nand UO_846 (O_846,N_19766,N_19946);
nand UO_847 (O_847,N_19944,N_19555);
nor UO_848 (O_848,N_19913,N_19794);
nor UO_849 (O_849,N_19951,N_19924);
nor UO_850 (O_850,N_19792,N_19884);
or UO_851 (O_851,N_19997,N_19645);
nor UO_852 (O_852,N_19793,N_19956);
nor UO_853 (O_853,N_19595,N_19876);
xor UO_854 (O_854,N_19533,N_19518);
xor UO_855 (O_855,N_19973,N_19929);
nor UO_856 (O_856,N_19922,N_19584);
and UO_857 (O_857,N_19949,N_19702);
nor UO_858 (O_858,N_19982,N_19762);
nor UO_859 (O_859,N_19868,N_19899);
xor UO_860 (O_860,N_19879,N_19508);
and UO_861 (O_861,N_19866,N_19787);
nor UO_862 (O_862,N_19695,N_19694);
nor UO_863 (O_863,N_19815,N_19500);
nand UO_864 (O_864,N_19769,N_19798);
or UO_865 (O_865,N_19665,N_19509);
or UO_866 (O_866,N_19513,N_19696);
xnor UO_867 (O_867,N_19918,N_19968);
and UO_868 (O_868,N_19654,N_19733);
or UO_869 (O_869,N_19768,N_19915);
nand UO_870 (O_870,N_19611,N_19793);
nor UO_871 (O_871,N_19679,N_19766);
and UO_872 (O_872,N_19980,N_19947);
nor UO_873 (O_873,N_19938,N_19724);
or UO_874 (O_874,N_19595,N_19586);
nor UO_875 (O_875,N_19701,N_19704);
nand UO_876 (O_876,N_19819,N_19873);
nand UO_877 (O_877,N_19719,N_19841);
or UO_878 (O_878,N_19880,N_19525);
or UO_879 (O_879,N_19836,N_19693);
or UO_880 (O_880,N_19791,N_19689);
nor UO_881 (O_881,N_19890,N_19748);
or UO_882 (O_882,N_19788,N_19769);
nand UO_883 (O_883,N_19532,N_19676);
or UO_884 (O_884,N_19520,N_19765);
nand UO_885 (O_885,N_19703,N_19543);
nand UO_886 (O_886,N_19889,N_19552);
or UO_887 (O_887,N_19641,N_19721);
and UO_888 (O_888,N_19663,N_19733);
nor UO_889 (O_889,N_19624,N_19582);
nor UO_890 (O_890,N_19872,N_19887);
nor UO_891 (O_891,N_19622,N_19703);
nor UO_892 (O_892,N_19615,N_19840);
and UO_893 (O_893,N_19889,N_19604);
xor UO_894 (O_894,N_19590,N_19530);
or UO_895 (O_895,N_19918,N_19719);
nand UO_896 (O_896,N_19942,N_19860);
xor UO_897 (O_897,N_19810,N_19630);
and UO_898 (O_898,N_19838,N_19959);
and UO_899 (O_899,N_19740,N_19748);
or UO_900 (O_900,N_19581,N_19980);
and UO_901 (O_901,N_19888,N_19879);
nand UO_902 (O_902,N_19882,N_19653);
or UO_903 (O_903,N_19544,N_19516);
nor UO_904 (O_904,N_19789,N_19961);
and UO_905 (O_905,N_19550,N_19860);
nor UO_906 (O_906,N_19592,N_19725);
xnor UO_907 (O_907,N_19815,N_19808);
or UO_908 (O_908,N_19816,N_19856);
nor UO_909 (O_909,N_19539,N_19658);
and UO_910 (O_910,N_19510,N_19850);
and UO_911 (O_911,N_19792,N_19804);
nor UO_912 (O_912,N_19840,N_19543);
or UO_913 (O_913,N_19541,N_19827);
nand UO_914 (O_914,N_19721,N_19863);
nor UO_915 (O_915,N_19626,N_19904);
and UO_916 (O_916,N_19799,N_19953);
or UO_917 (O_917,N_19685,N_19836);
and UO_918 (O_918,N_19566,N_19903);
xor UO_919 (O_919,N_19858,N_19571);
nor UO_920 (O_920,N_19956,N_19531);
and UO_921 (O_921,N_19771,N_19527);
nand UO_922 (O_922,N_19672,N_19923);
and UO_923 (O_923,N_19504,N_19625);
nand UO_924 (O_924,N_19754,N_19899);
or UO_925 (O_925,N_19792,N_19621);
or UO_926 (O_926,N_19556,N_19785);
nand UO_927 (O_927,N_19864,N_19682);
nor UO_928 (O_928,N_19545,N_19724);
or UO_929 (O_929,N_19805,N_19989);
or UO_930 (O_930,N_19632,N_19825);
or UO_931 (O_931,N_19569,N_19508);
nand UO_932 (O_932,N_19644,N_19852);
or UO_933 (O_933,N_19813,N_19500);
and UO_934 (O_934,N_19969,N_19723);
or UO_935 (O_935,N_19550,N_19834);
nand UO_936 (O_936,N_19783,N_19930);
nor UO_937 (O_937,N_19830,N_19685);
nand UO_938 (O_938,N_19865,N_19881);
xor UO_939 (O_939,N_19787,N_19722);
xor UO_940 (O_940,N_19724,N_19579);
nor UO_941 (O_941,N_19903,N_19699);
xor UO_942 (O_942,N_19759,N_19626);
and UO_943 (O_943,N_19885,N_19688);
nand UO_944 (O_944,N_19541,N_19900);
or UO_945 (O_945,N_19843,N_19970);
or UO_946 (O_946,N_19508,N_19869);
or UO_947 (O_947,N_19563,N_19839);
or UO_948 (O_948,N_19693,N_19666);
nor UO_949 (O_949,N_19701,N_19582);
nor UO_950 (O_950,N_19528,N_19526);
nand UO_951 (O_951,N_19850,N_19525);
or UO_952 (O_952,N_19688,N_19526);
nand UO_953 (O_953,N_19917,N_19795);
xor UO_954 (O_954,N_19545,N_19761);
xor UO_955 (O_955,N_19749,N_19511);
nor UO_956 (O_956,N_19579,N_19922);
and UO_957 (O_957,N_19689,N_19596);
and UO_958 (O_958,N_19509,N_19778);
xor UO_959 (O_959,N_19575,N_19910);
xnor UO_960 (O_960,N_19960,N_19713);
or UO_961 (O_961,N_19525,N_19944);
or UO_962 (O_962,N_19718,N_19965);
and UO_963 (O_963,N_19852,N_19702);
or UO_964 (O_964,N_19697,N_19799);
nand UO_965 (O_965,N_19681,N_19609);
xor UO_966 (O_966,N_19796,N_19536);
nor UO_967 (O_967,N_19891,N_19552);
and UO_968 (O_968,N_19624,N_19715);
xnor UO_969 (O_969,N_19621,N_19862);
nor UO_970 (O_970,N_19996,N_19534);
or UO_971 (O_971,N_19823,N_19977);
xor UO_972 (O_972,N_19688,N_19886);
xor UO_973 (O_973,N_19687,N_19915);
nand UO_974 (O_974,N_19979,N_19529);
nand UO_975 (O_975,N_19825,N_19893);
and UO_976 (O_976,N_19599,N_19916);
or UO_977 (O_977,N_19973,N_19555);
nor UO_978 (O_978,N_19891,N_19798);
or UO_979 (O_979,N_19677,N_19957);
nand UO_980 (O_980,N_19886,N_19612);
xnor UO_981 (O_981,N_19686,N_19667);
xor UO_982 (O_982,N_19597,N_19779);
or UO_983 (O_983,N_19687,N_19625);
xnor UO_984 (O_984,N_19929,N_19576);
and UO_985 (O_985,N_19513,N_19899);
and UO_986 (O_986,N_19864,N_19567);
nor UO_987 (O_987,N_19551,N_19795);
nand UO_988 (O_988,N_19713,N_19593);
or UO_989 (O_989,N_19776,N_19822);
nor UO_990 (O_990,N_19714,N_19598);
or UO_991 (O_991,N_19637,N_19956);
or UO_992 (O_992,N_19821,N_19744);
nand UO_993 (O_993,N_19765,N_19969);
and UO_994 (O_994,N_19747,N_19702);
or UO_995 (O_995,N_19642,N_19939);
nor UO_996 (O_996,N_19622,N_19593);
xnor UO_997 (O_997,N_19820,N_19805);
and UO_998 (O_998,N_19901,N_19815);
xnor UO_999 (O_999,N_19887,N_19868);
or UO_1000 (O_1000,N_19549,N_19709);
nand UO_1001 (O_1001,N_19548,N_19684);
or UO_1002 (O_1002,N_19608,N_19560);
xor UO_1003 (O_1003,N_19533,N_19704);
nor UO_1004 (O_1004,N_19835,N_19860);
xor UO_1005 (O_1005,N_19980,N_19715);
and UO_1006 (O_1006,N_19906,N_19649);
and UO_1007 (O_1007,N_19794,N_19935);
nor UO_1008 (O_1008,N_19559,N_19745);
xor UO_1009 (O_1009,N_19743,N_19842);
nand UO_1010 (O_1010,N_19757,N_19740);
and UO_1011 (O_1011,N_19866,N_19817);
nand UO_1012 (O_1012,N_19741,N_19843);
and UO_1013 (O_1013,N_19727,N_19689);
xnor UO_1014 (O_1014,N_19502,N_19949);
nand UO_1015 (O_1015,N_19828,N_19621);
or UO_1016 (O_1016,N_19530,N_19816);
xor UO_1017 (O_1017,N_19758,N_19739);
nand UO_1018 (O_1018,N_19780,N_19574);
xnor UO_1019 (O_1019,N_19949,N_19953);
nor UO_1020 (O_1020,N_19658,N_19786);
and UO_1021 (O_1021,N_19551,N_19765);
or UO_1022 (O_1022,N_19981,N_19951);
or UO_1023 (O_1023,N_19659,N_19876);
or UO_1024 (O_1024,N_19903,N_19668);
and UO_1025 (O_1025,N_19527,N_19848);
or UO_1026 (O_1026,N_19861,N_19640);
nor UO_1027 (O_1027,N_19766,N_19970);
nand UO_1028 (O_1028,N_19749,N_19692);
xor UO_1029 (O_1029,N_19892,N_19629);
nand UO_1030 (O_1030,N_19562,N_19780);
nand UO_1031 (O_1031,N_19926,N_19798);
and UO_1032 (O_1032,N_19872,N_19753);
nand UO_1033 (O_1033,N_19993,N_19921);
or UO_1034 (O_1034,N_19725,N_19777);
and UO_1035 (O_1035,N_19665,N_19992);
nand UO_1036 (O_1036,N_19719,N_19636);
nand UO_1037 (O_1037,N_19568,N_19664);
xor UO_1038 (O_1038,N_19878,N_19914);
or UO_1039 (O_1039,N_19940,N_19674);
xnor UO_1040 (O_1040,N_19678,N_19844);
or UO_1041 (O_1041,N_19641,N_19511);
nand UO_1042 (O_1042,N_19849,N_19508);
xnor UO_1043 (O_1043,N_19599,N_19827);
xor UO_1044 (O_1044,N_19503,N_19515);
and UO_1045 (O_1045,N_19696,N_19966);
or UO_1046 (O_1046,N_19994,N_19904);
nor UO_1047 (O_1047,N_19699,N_19776);
nor UO_1048 (O_1048,N_19949,N_19844);
and UO_1049 (O_1049,N_19687,N_19850);
and UO_1050 (O_1050,N_19832,N_19973);
nor UO_1051 (O_1051,N_19965,N_19674);
nand UO_1052 (O_1052,N_19705,N_19552);
or UO_1053 (O_1053,N_19792,N_19620);
nor UO_1054 (O_1054,N_19689,N_19735);
xor UO_1055 (O_1055,N_19778,N_19711);
xor UO_1056 (O_1056,N_19680,N_19727);
nand UO_1057 (O_1057,N_19561,N_19833);
xor UO_1058 (O_1058,N_19623,N_19867);
nand UO_1059 (O_1059,N_19780,N_19675);
xor UO_1060 (O_1060,N_19678,N_19959);
nand UO_1061 (O_1061,N_19774,N_19784);
or UO_1062 (O_1062,N_19502,N_19990);
nor UO_1063 (O_1063,N_19622,N_19802);
or UO_1064 (O_1064,N_19936,N_19562);
nand UO_1065 (O_1065,N_19612,N_19759);
or UO_1066 (O_1066,N_19972,N_19968);
nor UO_1067 (O_1067,N_19931,N_19838);
nand UO_1068 (O_1068,N_19581,N_19677);
and UO_1069 (O_1069,N_19506,N_19510);
nand UO_1070 (O_1070,N_19806,N_19784);
and UO_1071 (O_1071,N_19687,N_19931);
nor UO_1072 (O_1072,N_19510,N_19707);
and UO_1073 (O_1073,N_19904,N_19512);
xor UO_1074 (O_1074,N_19748,N_19968);
xor UO_1075 (O_1075,N_19956,N_19976);
nor UO_1076 (O_1076,N_19560,N_19616);
nand UO_1077 (O_1077,N_19547,N_19808);
or UO_1078 (O_1078,N_19710,N_19801);
xnor UO_1079 (O_1079,N_19998,N_19698);
xor UO_1080 (O_1080,N_19859,N_19584);
nand UO_1081 (O_1081,N_19902,N_19669);
xor UO_1082 (O_1082,N_19748,N_19619);
nor UO_1083 (O_1083,N_19848,N_19954);
and UO_1084 (O_1084,N_19937,N_19745);
or UO_1085 (O_1085,N_19593,N_19584);
nor UO_1086 (O_1086,N_19725,N_19820);
nor UO_1087 (O_1087,N_19781,N_19888);
and UO_1088 (O_1088,N_19710,N_19980);
and UO_1089 (O_1089,N_19750,N_19960);
and UO_1090 (O_1090,N_19846,N_19578);
nor UO_1091 (O_1091,N_19537,N_19875);
xnor UO_1092 (O_1092,N_19595,N_19954);
nor UO_1093 (O_1093,N_19578,N_19571);
nand UO_1094 (O_1094,N_19689,N_19533);
nand UO_1095 (O_1095,N_19615,N_19519);
and UO_1096 (O_1096,N_19937,N_19713);
nor UO_1097 (O_1097,N_19593,N_19529);
and UO_1098 (O_1098,N_19841,N_19751);
or UO_1099 (O_1099,N_19504,N_19709);
nand UO_1100 (O_1100,N_19571,N_19917);
nand UO_1101 (O_1101,N_19584,N_19651);
nand UO_1102 (O_1102,N_19507,N_19920);
xnor UO_1103 (O_1103,N_19512,N_19730);
nor UO_1104 (O_1104,N_19867,N_19750);
and UO_1105 (O_1105,N_19840,N_19517);
and UO_1106 (O_1106,N_19552,N_19946);
nor UO_1107 (O_1107,N_19801,N_19544);
nor UO_1108 (O_1108,N_19885,N_19871);
xnor UO_1109 (O_1109,N_19610,N_19665);
nand UO_1110 (O_1110,N_19606,N_19549);
or UO_1111 (O_1111,N_19757,N_19588);
nand UO_1112 (O_1112,N_19878,N_19900);
nand UO_1113 (O_1113,N_19858,N_19743);
or UO_1114 (O_1114,N_19586,N_19578);
xnor UO_1115 (O_1115,N_19579,N_19701);
nand UO_1116 (O_1116,N_19937,N_19910);
and UO_1117 (O_1117,N_19993,N_19660);
xor UO_1118 (O_1118,N_19538,N_19836);
nor UO_1119 (O_1119,N_19871,N_19746);
and UO_1120 (O_1120,N_19938,N_19858);
nor UO_1121 (O_1121,N_19987,N_19604);
nor UO_1122 (O_1122,N_19523,N_19738);
or UO_1123 (O_1123,N_19877,N_19973);
nor UO_1124 (O_1124,N_19544,N_19925);
xor UO_1125 (O_1125,N_19943,N_19908);
xnor UO_1126 (O_1126,N_19526,N_19555);
nand UO_1127 (O_1127,N_19515,N_19973);
nand UO_1128 (O_1128,N_19633,N_19903);
nor UO_1129 (O_1129,N_19755,N_19927);
or UO_1130 (O_1130,N_19947,N_19583);
nor UO_1131 (O_1131,N_19930,N_19772);
xnor UO_1132 (O_1132,N_19959,N_19645);
xnor UO_1133 (O_1133,N_19649,N_19584);
nand UO_1134 (O_1134,N_19743,N_19977);
nor UO_1135 (O_1135,N_19921,N_19867);
or UO_1136 (O_1136,N_19798,N_19810);
xnor UO_1137 (O_1137,N_19671,N_19808);
nor UO_1138 (O_1138,N_19624,N_19631);
or UO_1139 (O_1139,N_19516,N_19525);
and UO_1140 (O_1140,N_19575,N_19912);
nand UO_1141 (O_1141,N_19676,N_19571);
nand UO_1142 (O_1142,N_19832,N_19782);
or UO_1143 (O_1143,N_19839,N_19641);
or UO_1144 (O_1144,N_19547,N_19558);
or UO_1145 (O_1145,N_19878,N_19807);
and UO_1146 (O_1146,N_19627,N_19602);
xnor UO_1147 (O_1147,N_19842,N_19512);
or UO_1148 (O_1148,N_19605,N_19822);
or UO_1149 (O_1149,N_19552,N_19999);
nor UO_1150 (O_1150,N_19960,N_19600);
nor UO_1151 (O_1151,N_19984,N_19623);
or UO_1152 (O_1152,N_19952,N_19818);
xor UO_1153 (O_1153,N_19904,N_19606);
or UO_1154 (O_1154,N_19867,N_19543);
nor UO_1155 (O_1155,N_19849,N_19507);
or UO_1156 (O_1156,N_19803,N_19652);
nand UO_1157 (O_1157,N_19548,N_19623);
xor UO_1158 (O_1158,N_19713,N_19981);
or UO_1159 (O_1159,N_19957,N_19609);
or UO_1160 (O_1160,N_19774,N_19543);
nand UO_1161 (O_1161,N_19944,N_19562);
nand UO_1162 (O_1162,N_19673,N_19909);
nor UO_1163 (O_1163,N_19522,N_19981);
nand UO_1164 (O_1164,N_19872,N_19842);
xnor UO_1165 (O_1165,N_19991,N_19705);
and UO_1166 (O_1166,N_19966,N_19504);
xnor UO_1167 (O_1167,N_19861,N_19738);
nand UO_1168 (O_1168,N_19624,N_19534);
nand UO_1169 (O_1169,N_19542,N_19624);
or UO_1170 (O_1170,N_19509,N_19804);
xor UO_1171 (O_1171,N_19823,N_19882);
nor UO_1172 (O_1172,N_19538,N_19779);
nand UO_1173 (O_1173,N_19514,N_19938);
or UO_1174 (O_1174,N_19973,N_19504);
nand UO_1175 (O_1175,N_19667,N_19834);
and UO_1176 (O_1176,N_19502,N_19821);
or UO_1177 (O_1177,N_19902,N_19516);
or UO_1178 (O_1178,N_19554,N_19690);
or UO_1179 (O_1179,N_19565,N_19511);
nand UO_1180 (O_1180,N_19621,N_19559);
and UO_1181 (O_1181,N_19723,N_19530);
nand UO_1182 (O_1182,N_19989,N_19865);
xor UO_1183 (O_1183,N_19593,N_19735);
and UO_1184 (O_1184,N_19543,N_19786);
nor UO_1185 (O_1185,N_19541,N_19843);
xnor UO_1186 (O_1186,N_19501,N_19735);
or UO_1187 (O_1187,N_19613,N_19923);
nor UO_1188 (O_1188,N_19930,N_19842);
and UO_1189 (O_1189,N_19892,N_19722);
nor UO_1190 (O_1190,N_19694,N_19967);
xor UO_1191 (O_1191,N_19890,N_19744);
xor UO_1192 (O_1192,N_19676,N_19680);
nand UO_1193 (O_1193,N_19564,N_19515);
or UO_1194 (O_1194,N_19579,N_19946);
nor UO_1195 (O_1195,N_19570,N_19645);
and UO_1196 (O_1196,N_19936,N_19783);
nand UO_1197 (O_1197,N_19536,N_19514);
nor UO_1198 (O_1198,N_19736,N_19672);
xor UO_1199 (O_1199,N_19966,N_19607);
nand UO_1200 (O_1200,N_19562,N_19974);
and UO_1201 (O_1201,N_19761,N_19714);
nor UO_1202 (O_1202,N_19534,N_19855);
nor UO_1203 (O_1203,N_19737,N_19595);
and UO_1204 (O_1204,N_19891,N_19652);
nor UO_1205 (O_1205,N_19855,N_19938);
nor UO_1206 (O_1206,N_19746,N_19773);
nand UO_1207 (O_1207,N_19769,N_19920);
and UO_1208 (O_1208,N_19793,N_19635);
nor UO_1209 (O_1209,N_19752,N_19917);
or UO_1210 (O_1210,N_19885,N_19629);
and UO_1211 (O_1211,N_19908,N_19793);
xnor UO_1212 (O_1212,N_19921,N_19585);
and UO_1213 (O_1213,N_19885,N_19724);
nor UO_1214 (O_1214,N_19722,N_19893);
nor UO_1215 (O_1215,N_19760,N_19642);
and UO_1216 (O_1216,N_19622,N_19807);
nor UO_1217 (O_1217,N_19695,N_19608);
or UO_1218 (O_1218,N_19822,N_19951);
nor UO_1219 (O_1219,N_19555,N_19793);
or UO_1220 (O_1220,N_19849,N_19935);
nor UO_1221 (O_1221,N_19557,N_19781);
xnor UO_1222 (O_1222,N_19698,N_19768);
nand UO_1223 (O_1223,N_19949,N_19779);
nand UO_1224 (O_1224,N_19657,N_19922);
or UO_1225 (O_1225,N_19871,N_19557);
and UO_1226 (O_1226,N_19978,N_19544);
and UO_1227 (O_1227,N_19672,N_19688);
or UO_1228 (O_1228,N_19897,N_19604);
or UO_1229 (O_1229,N_19867,N_19833);
nor UO_1230 (O_1230,N_19639,N_19799);
xnor UO_1231 (O_1231,N_19961,N_19627);
and UO_1232 (O_1232,N_19841,N_19601);
or UO_1233 (O_1233,N_19538,N_19856);
nand UO_1234 (O_1234,N_19634,N_19697);
and UO_1235 (O_1235,N_19584,N_19644);
nor UO_1236 (O_1236,N_19738,N_19583);
nor UO_1237 (O_1237,N_19819,N_19617);
xor UO_1238 (O_1238,N_19692,N_19984);
nand UO_1239 (O_1239,N_19930,N_19682);
or UO_1240 (O_1240,N_19987,N_19524);
nor UO_1241 (O_1241,N_19793,N_19612);
and UO_1242 (O_1242,N_19784,N_19988);
nand UO_1243 (O_1243,N_19773,N_19514);
or UO_1244 (O_1244,N_19554,N_19541);
nand UO_1245 (O_1245,N_19888,N_19614);
nor UO_1246 (O_1246,N_19576,N_19907);
or UO_1247 (O_1247,N_19586,N_19605);
nor UO_1248 (O_1248,N_19671,N_19971);
nand UO_1249 (O_1249,N_19686,N_19656);
nor UO_1250 (O_1250,N_19673,N_19755);
nor UO_1251 (O_1251,N_19678,N_19617);
and UO_1252 (O_1252,N_19623,N_19516);
or UO_1253 (O_1253,N_19623,N_19565);
nor UO_1254 (O_1254,N_19971,N_19511);
nand UO_1255 (O_1255,N_19695,N_19540);
xor UO_1256 (O_1256,N_19518,N_19759);
nor UO_1257 (O_1257,N_19964,N_19780);
nor UO_1258 (O_1258,N_19646,N_19931);
or UO_1259 (O_1259,N_19936,N_19983);
xor UO_1260 (O_1260,N_19840,N_19719);
and UO_1261 (O_1261,N_19687,N_19588);
nand UO_1262 (O_1262,N_19692,N_19953);
nand UO_1263 (O_1263,N_19994,N_19920);
nand UO_1264 (O_1264,N_19971,N_19576);
nor UO_1265 (O_1265,N_19749,N_19889);
nor UO_1266 (O_1266,N_19977,N_19877);
or UO_1267 (O_1267,N_19507,N_19836);
nor UO_1268 (O_1268,N_19542,N_19608);
nand UO_1269 (O_1269,N_19586,N_19695);
nor UO_1270 (O_1270,N_19865,N_19755);
nor UO_1271 (O_1271,N_19950,N_19571);
nor UO_1272 (O_1272,N_19813,N_19778);
nand UO_1273 (O_1273,N_19802,N_19698);
and UO_1274 (O_1274,N_19926,N_19810);
nand UO_1275 (O_1275,N_19586,N_19915);
and UO_1276 (O_1276,N_19926,N_19873);
xor UO_1277 (O_1277,N_19987,N_19843);
and UO_1278 (O_1278,N_19678,N_19612);
and UO_1279 (O_1279,N_19794,N_19850);
and UO_1280 (O_1280,N_19727,N_19779);
nor UO_1281 (O_1281,N_19889,N_19947);
nor UO_1282 (O_1282,N_19706,N_19781);
and UO_1283 (O_1283,N_19737,N_19757);
nor UO_1284 (O_1284,N_19644,N_19542);
nand UO_1285 (O_1285,N_19747,N_19835);
or UO_1286 (O_1286,N_19573,N_19636);
nand UO_1287 (O_1287,N_19945,N_19899);
and UO_1288 (O_1288,N_19744,N_19853);
nand UO_1289 (O_1289,N_19863,N_19890);
xor UO_1290 (O_1290,N_19902,N_19620);
nor UO_1291 (O_1291,N_19714,N_19984);
nor UO_1292 (O_1292,N_19939,N_19891);
nand UO_1293 (O_1293,N_19568,N_19674);
or UO_1294 (O_1294,N_19635,N_19942);
nor UO_1295 (O_1295,N_19509,N_19847);
xor UO_1296 (O_1296,N_19857,N_19862);
nand UO_1297 (O_1297,N_19559,N_19698);
and UO_1298 (O_1298,N_19582,N_19647);
nor UO_1299 (O_1299,N_19694,N_19903);
or UO_1300 (O_1300,N_19978,N_19562);
xnor UO_1301 (O_1301,N_19884,N_19863);
nand UO_1302 (O_1302,N_19740,N_19943);
nand UO_1303 (O_1303,N_19943,N_19715);
nand UO_1304 (O_1304,N_19644,N_19949);
nor UO_1305 (O_1305,N_19959,N_19891);
or UO_1306 (O_1306,N_19653,N_19706);
xnor UO_1307 (O_1307,N_19942,N_19966);
or UO_1308 (O_1308,N_19870,N_19917);
or UO_1309 (O_1309,N_19706,N_19931);
and UO_1310 (O_1310,N_19803,N_19710);
and UO_1311 (O_1311,N_19754,N_19687);
nor UO_1312 (O_1312,N_19508,N_19782);
nor UO_1313 (O_1313,N_19894,N_19672);
nand UO_1314 (O_1314,N_19756,N_19546);
or UO_1315 (O_1315,N_19649,N_19665);
nor UO_1316 (O_1316,N_19532,N_19803);
nor UO_1317 (O_1317,N_19989,N_19795);
nor UO_1318 (O_1318,N_19807,N_19933);
and UO_1319 (O_1319,N_19720,N_19640);
and UO_1320 (O_1320,N_19704,N_19584);
nand UO_1321 (O_1321,N_19976,N_19917);
or UO_1322 (O_1322,N_19829,N_19898);
and UO_1323 (O_1323,N_19821,N_19701);
nor UO_1324 (O_1324,N_19958,N_19941);
or UO_1325 (O_1325,N_19893,N_19791);
and UO_1326 (O_1326,N_19968,N_19794);
or UO_1327 (O_1327,N_19622,N_19912);
nor UO_1328 (O_1328,N_19870,N_19685);
or UO_1329 (O_1329,N_19880,N_19511);
and UO_1330 (O_1330,N_19630,N_19963);
nand UO_1331 (O_1331,N_19712,N_19502);
nor UO_1332 (O_1332,N_19942,N_19640);
and UO_1333 (O_1333,N_19569,N_19778);
nor UO_1334 (O_1334,N_19928,N_19519);
and UO_1335 (O_1335,N_19735,N_19661);
nand UO_1336 (O_1336,N_19960,N_19911);
xnor UO_1337 (O_1337,N_19763,N_19528);
nor UO_1338 (O_1338,N_19586,N_19975);
nand UO_1339 (O_1339,N_19704,N_19988);
nor UO_1340 (O_1340,N_19912,N_19818);
nand UO_1341 (O_1341,N_19928,N_19949);
or UO_1342 (O_1342,N_19691,N_19520);
and UO_1343 (O_1343,N_19729,N_19860);
or UO_1344 (O_1344,N_19821,N_19992);
or UO_1345 (O_1345,N_19827,N_19816);
xnor UO_1346 (O_1346,N_19701,N_19520);
nor UO_1347 (O_1347,N_19547,N_19898);
and UO_1348 (O_1348,N_19997,N_19759);
nand UO_1349 (O_1349,N_19812,N_19572);
xnor UO_1350 (O_1350,N_19768,N_19549);
nand UO_1351 (O_1351,N_19656,N_19897);
nor UO_1352 (O_1352,N_19706,N_19520);
nand UO_1353 (O_1353,N_19784,N_19657);
nand UO_1354 (O_1354,N_19822,N_19769);
and UO_1355 (O_1355,N_19876,N_19888);
nand UO_1356 (O_1356,N_19779,N_19729);
nor UO_1357 (O_1357,N_19712,N_19922);
and UO_1358 (O_1358,N_19613,N_19776);
nor UO_1359 (O_1359,N_19673,N_19853);
or UO_1360 (O_1360,N_19952,N_19583);
nand UO_1361 (O_1361,N_19620,N_19714);
nand UO_1362 (O_1362,N_19636,N_19939);
or UO_1363 (O_1363,N_19747,N_19810);
and UO_1364 (O_1364,N_19506,N_19577);
nor UO_1365 (O_1365,N_19993,N_19877);
xor UO_1366 (O_1366,N_19502,N_19661);
nand UO_1367 (O_1367,N_19722,N_19897);
and UO_1368 (O_1368,N_19600,N_19673);
nand UO_1369 (O_1369,N_19805,N_19744);
nor UO_1370 (O_1370,N_19500,N_19698);
and UO_1371 (O_1371,N_19598,N_19901);
nor UO_1372 (O_1372,N_19946,N_19775);
nor UO_1373 (O_1373,N_19893,N_19941);
nand UO_1374 (O_1374,N_19893,N_19943);
nor UO_1375 (O_1375,N_19824,N_19563);
xnor UO_1376 (O_1376,N_19852,N_19669);
nand UO_1377 (O_1377,N_19973,N_19643);
or UO_1378 (O_1378,N_19795,N_19736);
nor UO_1379 (O_1379,N_19908,N_19713);
and UO_1380 (O_1380,N_19773,N_19676);
nor UO_1381 (O_1381,N_19721,N_19973);
nand UO_1382 (O_1382,N_19818,N_19832);
xor UO_1383 (O_1383,N_19956,N_19518);
nor UO_1384 (O_1384,N_19599,N_19939);
and UO_1385 (O_1385,N_19761,N_19535);
nand UO_1386 (O_1386,N_19568,N_19545);
or UO_1387 (O_1387,N_19557,N_19542);
nor UO_1388 (O_1388,N_19926,N_19794);
nor UO_1389 (O_1389,N_19919,N_19680);
or UO_1390 (O_1390,N_19687,N_19945);
or UO_1391 (O_1391,N_19788,N_19875);
xnor UO_1392 (O_1392,N_19937,N_19842);
and UO_1393 (O_1393,N_19974,N_19526);
nor UO_1394 (O_1394,N_19909,N_19666);
xor UO_1395 (O_1395,N_19900,N_19502);
and UO_1396 (O_1396,N_19528,N_19898);
xor UO_1397 (O_1397,N_19896,N_19807);
or UO_1398 (O_1398,N_19691,N_19834);
xnor UO_1399 (O_1399,N_19545,N_19882);
nand UO_1400 (O_1400,N_19670,N_19795);
xor UO_1401 (O_1401,N_19697,N_19555);
and UO_1402 (O_1402,N_19858,N_19512);
or UO_1403 (O_1403,N_19693,N_19790);
nor UO_1404 (O_1404,N_19737,N_19698);
nand UO_1405 (O_1405,N_19570,N_19984);
nor UO_1406 (O_1406,N_19726,N_19786);
nor UO_1407 (O_1407,N_19757,N_19785);
or UO_1408 (O_1408,N_19905,N_19664);
nand UO_1409 (O_1409,N_19514,N_19955);
nor UO_1410 (O_1410,N_19606,N_19653);
and UO_1411 (O_1411,N_19536,N_19547);
or UO_1412 (O_1412,N_19649,N_19981);
nor UO_1413 (O_1413,N_19644,N_19731);
nor UO_1414 (O_1414,N_19697,N_19843);
xor UO_1415 (O_1415,N_19683,N_19938);
or UO_1416 (O_1416,N_19504,N_19684);
nor UO_1417 (O_1417,N_19753,N_19809);
xnor UO_1418 (O_1418,N_19622,N_19987);
and UO_1419 (O_1419,N_19952,N_19896);
xnor UO_1420 (O_1420,N_19930,N_19762);
nand UO_1421 (O_1421,N_19527,N_19652);
xor UO_1422 (O_1422,N_19574,N_19865);
nand UO_1423 (O_1423,N_19726,N_19709);
nor UO_1424 (O_1424,N_19640,N_19772);
nor UO_1425 (O_1425,N_19819,N_19706);
nor UO_1426 (O_1426,N_19688,N_19650);
nor UO_1427 (O_1427,N_19688,N_19746);
nor UO_1428 (O_1428,N_19618,N_19768);
or UO_1429 (O_1429,N_19876,N_19616);
nor UO_1430 (O_1430,N_19776,N_19570);
nor UO_1431 (O_1431,N_19663,N_19869);
nor UO_1432 (O_1432,N_19759,N_19532);
nand UO_1433 (O_1433,N_19707,N_19767);
nand UO_1434 (O_1434,N_19626,N_19635);
nor UO_1435 (O_1435,N_19741,N_19699);
or UO_1436 (O_1436,N_19777,N_19766);
or UO_1437 (O_1437,N_19667,N_19893);
nor UO_1438 (O_1438,N_19708,N_19791);
nor UO_1439 (O_1439,N_19951,N_19651);
or UO_1440 (O_1440,N_19592,N_19843);
nand UO_1441 (O_1441,N_19839,N_19948);
and UO_1442 (O_1442,N_19949,N_19888);
xor UO_1443 (O_1443,N_19765,N_19502);
or UO_1444 (O_1444,N_19820,N_19802);
or UO_1445 (O_1445,N_19921,N_19505);
xnor UO_1446 (O_1446,N_19762,N_19926);
xor UO_1447 (O_1447,N_19588,N_19538);
or UO_1448 (O_1448,N_19862,N_19577);
nor UO_1449 (O_1449,N_19538,N_19721);
nor UO_1450 (O_1450,N_19796,N_19810);
or UO_1451 (O_1451,N_19609,N_19794);
nor UO_1452 (O_1452,N_19750,N_19536);
xor UO_1453 (O_1453,N_19504,N_19727);
or UO_1454 (O_1454,N_19987,N_19674);
nand UO_1455 (O_1455,N_19930,N_19896);
and UO_1456 (O_1456,N_19691,N_19833);
nand UO_1457 (O_1457,N_19736,N_19628);
nor UO_1458 (O_1458,N_19657,N_19872);
nand UO_1459 (O_1459,N_19610,N_19933);
and UO_1460 (O_1460,N_19602,N_19942);
xor UO_1461 (O_1461,N_19946,N_19623);
or UO_1462 (O_1462,N_19889,N_19856);
nor UO_1463 (O_1463,N_19657,N_19917);
xnor UO_1464 (O_1464,N_19959,N_19524);
or UO_1465 (O_1465,N_19981,N_19651);
xnor UO_1466 (O_1466,N_19558,N_19796);
and UO_1467 (O_1467,N_19797,N_19668);
and UO_1468 (O_1468,N_19984,N_19849);
nand UO_1469 (O_1469,N_19711,N_19686);
nor UO_1470 (O_1470,N_19602,N_19540);
nand UO_1471 (O_1471,N_19760,N_19860);
nand UO_1472 (O_1472,N_19887,N_19514);
xnor UO_1473 (O_1473,N_19805,N_19833);
xor UO_1474 (O_1474,N_19637,N_19846);
xnor UO_1475 (O_1475,N_19733,N_19525);
or UO_1476 (O_1476,N_19525,N_19847);
xnor UO_1477 (O_1477,N_19956,N_19844);
nand UO_1478 (O_1478,N_19715,N_19985);
or UO_1479 (O_1479,N_19715,N_19691);
nor UO_1480 (O_1480,N_19591,N_19924);
xnor UO_1481 (O_1481,N_19941,N_19559);
or UO_1482 (O_1482,N_19500,N_19942);
xnor UO_1483 (O_1483,N_19643,N_19770);
or UO_1484 (O_1484,N_19752,N_19951);
or UO_1485 (O_1485,N_19602,N_19573);
or UO_1486 (O_1486,N_19633,N_19820);
nand UO_1487 (O_1487,N_19753,N_19564);
xor UO_1488 (O_1488,N_19801,N_19795);
or UO_1489 (O_1489,N_19896,N_19843);
nand UO_1490 (O_1490,N_19586,N_19881);
or UO_1491 (O_1491,N_19982,N_19876);
xor UO_1492 (O_1492,N_19649,N_19809);
nor UO_1493 (O_1493,N_19542,N_19732);
and UO_1494 (O_1494,N_19674,N_19653);
and UO_1495 (O_1495,N_19934,N_19519);
and UO_1496 (O_1496,N_19600,N_19518);
or UO_1497 (O_1497,N_19650,N_19929);
nand UO_1498 (O_1498,N_19784,N_19731);
and UO_1499 (O_1499,N_19805,N_19547);
nor UO_1500 (O_1500,N_19908,N_19910);
nor UO_1501 (O_1501,N_19880,N_19787);
nand UO_1502 (O_1502,N_19716,N_19556);
and UO_1503 (O_1503,N_19630,N_19540);
nand UO_1504 (O_1504,N_19824,N_19631);
nor UO_1505 (O_1505,N_19895,N_19710);
or UO_1506 (O_1506,N_19531,N_19744);
or UO_1507 (O_1507,N_19928,N_19883);
or UO_1508 (O_1508,N_19924,N_19940);
nand UO_1509 (O_1509,N_19882,N_19890);
xnor UO_1510 (O_1510,N_19749,N_19550);
and UO_1511 (O_1511,N_19703,N_19672);
nand UO_1512 (O_1512,N_19830,N_19950);
or UO_1513 (O_1513,N_19631,N_19589);
xnor UO_1514 (O_1514,N_19731,N_19955);
nand UO_1515 (O_1515,N_19951,N_19890);
nand UO_1516 (O_1516,N_19591,N_19562);
and UO_1517 (O_1517,N_19518,N_19990);
xor UO_1518 (O_1518,N_19522,N_19705);
or UO_1519 (O_1519,N_19591,N_19559);
nor UO_1520 (O_1520,N_19878,N_19960);
or UO_1521 (O_1521,N_19750,N_19805);
or UO_1522 (O_1522,N_19847,N_19826);
nor UO_1523 (O_1523,N_19524,N_19775);
xor UO_1524 (O_1524,N_19997,N_19928);
nand UO_1525 (O_1525,N_19620,N_19913);
nand UO_1526 (O_1526,N_19555,N_19921);
and UO_1527 (O_1527,N_19522,N_19710);
and UO_1528 (O_1528,N_19929,N_19826);
nor UO_1529 (O_1529,N_19964,N_19846);
xnor UO_1530 (O_1530,N_19875,N_19993);
nand UO_1531 (O_1531,N_19547,N_19937);
xnor UO_1532 (O_1532,N_19537,N_19930);
xnor UO_1533 (O_1533,N_19884,N_19738);
or UO_1534 (O_1534,N_19647,N_19558);
nor UO_1535 (O_1535,N_19912,N_19935);
and UO_1536 (O_1536,N_19802,N_19562);
and UO_1537 (O_1537,N_19538,N_19980);
or UO_1538 (O_1538,N_19788,N_19792);
and UO_1539 (O_1539,N_19941,N_19579);
nor UO_1540 (O_1540,N_19676,N_19579);
or UO_1541 (O_1541,N_19693,N_19976);
or UO_1542 (O_1542,N_19913,N_19627);
or UO_1543 (O_1543,N_19617,N_19831);
nor UO_1544 (O_1544,N_19657,N_19954);
nor UO_1545 (O_1545,N_19708,N_19636);
nor UO_1546 (O_1546,N_19991,N_19619);
and UO_1547 (O_1547,N_19611,N_19899);
xor UO_1548 (O_1548,N_19668,N_19960);
or UO_1549 (O_1549,N_19905,N_19705);
nand UO_1550 (O_1550,N_19941,N_19696);
or UO_1551 (O_1551,N_19773,N_19538);
nor UO_1552 (O_1552,N_19693,N_19822);
nor UO_1553 (O_1553,N_19765,N_19880);
or UO_1554 (O_1554,N_19761,N_19992);
nand UO_1555 (O_1555,N_19994,N_19785);
nand UO_1556 (O_1556,N_19768,N_19602);
or UO_1557 (O_1557,N_19719,N_19524);
xnor UO_1558 (O_1558,N_19933,N_19546);
and UO_1559 (O_1559,N_19765,N_19861);
nor UO_1560 (O_1560,N_19672,N_19515);
xor UO_1561 (O_1561,N_19738,N_19999);
xor UO_1562 (O_1562,N_19663,N_19910);
nand UO_1563 (O_1563,N_19500,N_19888);
xnor UO_1564 (O_1564,N_19757,N_19775);
nor UO_1565 (O_1565,N_19706,N_19686);
or UO_1566 (O_1566,N_19650,N_19839);
or UO_1567 (O_1567,N_19760,N_19959);
nor UO_1568 (O_1568,N_19614,N_19946);
xnor UO_1569 (O_1569,N_19900,N_19735);
xnor UO_1570 (O_1570,N_19904,N_19943);
xnor UO_1571 (O_1571,N_19668,N_19664);
and UO_1572 (O_1572,N_19664,N_19543);
nand UO_1573 (O_1573,N_19980,N_19572);
or UO_1574 (O_1574,N_19845,N_19908);
and UO_1575 (O_1575,N_19587,N_19666);
nand UO_1576 (O_1576,N_19726,N_19956);
xnor UO_1577 (O_1577,N_19939,N_19525);
and UO_1578 (O_1578,N_19863,N_19817);
or UO_1579 (O_1579,N_19779,N_19766);
nand UO_1580 (O_1580,N_19582,N_19504);
and UO_1581 (O_1581,N_19517,N_19914);
xor UO_1582 (O_1582,N_19836,N_19773);
xor UO_1583 (O_1583,N_19659,N_19516);
nand UO_1584 (O_1584,N_19775,N_19967);
xnor UO_1585 (O_1585,N_19545,N_19713);
xor UO_1586 (O_1586,N_19632,N_19940);
xnor UO_1587 (O_1587,N_19950,N_19700);
nand UO_1588 (O_1588,N_19600,N_19686);
or UO_1589 (O_1589,N_19797,N_19735);
nand UO_1590 (O_1590,N_19634,N_19992);
or UO_1591 (O_1591,N_19824,N_19909);
xnor UO_1592 (O_1592,N_19949,N_19822);
or UO_1593 (O_1593,N_19686,N_19580);
or UO_1594 (O_1594,N_19670,N_19674);
and UO_1595 (O_1595,N_19775,N_19706);
nand UO_1596 (O_1596,N_19939,N_19571);
nand UO_1597 (O_1597,N_19552,N_19588);
nand UO_1598 (O_1598,N_19595,N_19607);
and UO_1599 (O_1599,N_19506,N_19758);
and UO_1600 (O_1600,N_19999,N_19913);
nor UO_1601 (O_1601,N_19667,N_19734);
nand UO_1602 (O_1602,N_19638,N_19700);
and UO_1603 (O_1603,N_19816,N_19686);
xnor UO_1604 (O_1604,N_19987,N_19768);
and UO_1605 (O_1605,N_19714,N_19731);
and UO_1606 (O_1606,N_19537,N_19932);
and UO_1607 (O_1607,N_19623,N_19733);
nand UO_1608 (O_1608,N_19803,N_19931);
nor UO_1609 (O_1609,N_19893,N_19548);
or UO_1610 (O_1610,N_19519,N_19951);
or UO_1611 (O_1611,N_19732,N_19597);
and UO_1612 (O_1612,N_19907,N_19966);
or UO_1613 (O_1613,N_19705,N_19635);
and UO_1614 (O_1614,N_19541,N_19981);
nand UO_1615 (O_1615,N_19760,N_19572);
and UO_1616 (O_1616,N_19793,N_19632);
xor UO_1617 (O_1617,N_19920,N_19790);
and UO_1618 (O_1618,N_19515,N_19743);
and UO_1619 (O_1619,N_19676,N_19872);
or UO_1620 (O_1620,N_19962,N_19562);
xor UO_1621 (O_1621,N_19845,N_19967);
and UO_1622 (O_1622,N_19594,N_19937);
nor UO_1623 (O_1623,N_19740,N_19636);
nor UO_1624 (O_1624,N_19959,N_19852);
or UO_1625 (O_1625,N_19644,N_19736);
and UO_1626 (O_1626,N_19911,N_19869);
or UO_1627 (O_1627,N_19924,N_19993);
or UO_1628 (O_1628,N_19675,N_19665);
or UO_1629 (O_1629,N_19830,N_19874);
xnor UO_1630 (O_1630,N_19725,N_19564);
and UO_1631 (O_1631,N_19938,N_19621);
xor UO_1632 (O_1632,N_19687,N_19577);
nor UO_1633 (O_1633,N_19893,N_19579);
or UO_1634 (O_1634,N_19696,N_19534);
nand UO_1635 (O_1635,N_19524,N_19793);
and UO_1636 (O_1636,N_19639,N_19675);
xnor UO_1637 (O_1637,N_19582,N_19807);
or UO_1638 (O_1638,N_19866,N_19758);
nor UO_1639 (O_1639,N_19715,N_19587);
and UO_1640 (O_1640,N_19502,N_19516);
xor UO_1641 (O_1641,N_19925,N_19707);
nor UO_1642 (O_1642,N_19703,N_19801);
xnor UO_1643 (O_1643,N_19890,N_19812);
or UO_1644 (O_1644,N_19803,N_19525);
nor UO_1645 (O_1645,N_19629,N_19836);
and UO_1646 (O_1646,N_19936,N_19806);
nor UO_1647 (O_1647,N_19645,N_19998);
xnor UO_1648 (O_1648,N_19935,N_19566);
and UO_1649 (O_1649,N_19800,N_19932);
or UO_1650 (O_1650,N_19756,N_19914);
xor UO_1651 (O_1651,N_19850,N_19612);
nor UO_1652 (O_1652,N_19746,N_19752);
nand UO_1653 (O_1653,N_19619,N_19850);
nand UO_1654 (O_1654,N_19755,N_19864);
xor UO_1655 (O_1655,N_19937,N_19620);
and UO_1656 (O_1656,N_19500,N_19569);
nand UO_1657 (O_1657,N_19817,N_19891);
xor UO_1658 (O_1658,N_19948,N_19696);
xnor UO_1659 (O_1659,N_19683,N_19831);
nand UO_1660 (O_1660,N_19612,N_19719);
or UO_1661 (O_1661,N_19907,N_19602);
or UO_1662 (O_1662,N_19616,N_19908);
xnor UO_1663 (O_1663,N_19613,N_19581);
and UO_1664 (O_1664,N_19543,N_19624);
xor UO_1665 (O_1665,N_19949,N_19747);
nor UO_1666 (O_1666,N_19626,N_19652);
xnor UO_1667 (O_1667,N_19880,N_19520);
xor UO_1668 (O_1668,N_19552,N_19626);
xor UO_1669 (O_1669,N_19630,N_19883);
or UO_1670 (O_1670,N_19994,N_19658);
nand UO_1671 (O_1671,N_19575,N_19799);
xnor UO_1672 (O_1672,N_19607,N_19603);
nor UO_1673 (O_1673,N_19791,N_19819);
or UO_1674 (O_1674,N_19943,N_19594);
nor UO_1675 (O_1675,N_19857,N_19571);
and UO_1676 (O_1676,N_19507,N_19520);
xnor UO_1677 (O_1677,N_19675,N_19794);
nand UO_1678 (O_1678,N_19578,N_19958);
and UO_1679 (O_1679,N_19879,N_19909);
nor UO_1680 (O_1680,N_19958,N_19691);
or UO_1681 (O_1681,N_19884,N_19523);
nor UO_1682 (O_1682,N_19956,N_19707);
or UO_1683 (O_1683,N_19680,N_19724);
or UO_1684 (O_1684,N_19600,N_19741);
and UO_1685 (O_1685,N_19940,N_19994);
xor UO_1686 (O_1686,N_19846,N_19832);
and UO_1687 (O_1687,N_19596,N_19550);
or UO_1688 (O_1688,N_19759,N_19709);
and UO_1689 (O_1689,N_19566,N_19844);
and UO_1690 (O_1690,N_19520,N_19590);
nand UO_1691 (O_1691,N_19936,N_19769);
xor UO_1692 (O_1692,N_19835,N_19920);
or UO_1693 (O_1693,N_19810,N_19749);
nor UO_1694 (O_1694,N_19980,N_19731);
nand UO_1695 (O_1695,N_19668,N_19888);
or UO_1696 (O_1696,N_19605,N_19635);
xnor UO_1697 (O_1697,N_19819,N_19936);
nor UO_1698 (O_1698,N_19871,N_19613);
xnor UO_1699 (O_1699,N_19725,N_19569);
or UO_1700 (O_1700,N_19779,N_19970);
nor UO_1701 (O_1701,N_19907,N_19640);
nand UO_1702 (O_1702,N_19643,N_19631);
and UO_1703 (O_1703,N_19515,N_19965);
or UO_1704 (O_1704,N_19935,N_19964);
xnor UO_1705 (O_1705,N_19536,N_19822);
nor UO_1706 (O_1706,N_19962,N_19942);
xnor UO_1707 (O_1707,N_19685,N_19771);
nor UO_1708 (O_1708,N_19877,N_19736);
and UO_1709 (O_1709,N_19905,N_19830);
or UO_1710 (O_1710,N_19865,N_19947);
or UO_1711 (O_1711,N_19866,N_19936);
xnor UO_1712 (O_1712,N_19913,N_19863);
xor UO_1713 (O_1713,N_19638,N_19985);
and UO_1714 (O_1714,N_19820,N_19888);
or UO_1715 (O_1715,N_19531,N_19955);
nand UO_1716 (O_1716,N_19610,N_19530);
or UO_1717 (O_1717,N_19755,N_19765);
xor UO_1718 (O_1718,N_19953,N_19812);
xor UO_1719 (O_1719,N_19979,N_19931);
nand UO_1720 (O_1720,N_19688,N_19838);
nand UO_1721 (O_1721,N_19906,N_19813);
or UO_1722 (O_1722,N_19909,N_19610);
nand UO_1723 (O_1723,N_19993,N_19823);
nor UO_1724 (O_1724,N_19807,N_19838);
xnor UO_1725 (O_1725,N_19558,N_19641);
nand UO_1726 (O_1726,N_19758,N_19635);
nor UO_1727 (O_1727,N_19574,N_19587);
nand UO_1728 (O_1728,N_19568,N_19811);
or UO_1729 (O_1729,N_19740,N_19542);
and UO_1730 (O_1730,N_19519,N_19718);
nor UO_1731 (O_1731,N_19762,N_19792);
xnor UO_1732 (O_1732,N_19674,N_19529);
nor UO_1733 (O_1733,N_19609,N_19521);
and UO_1734 (O_1734,N_19750,N_19566);
or UO_1735 (O_1735,N_19981,N_19695);
and UO_1736 (O_1736,N_19853,N_19501);
or UO_1737 (O_1737,N_19852,N_19936);
nand UO_1738 (O_1738,N_19640,N_19650);
nor UO_1739 (O_1739,N_19917,N_19674);
or UO_1740 (O_1740,N_19779,N_19642);
nand UO_1741 (O_1741,N_19943,N_19785);
and UO_1742 (O_1742,N_19903,N_19963);
or UO_1743 (O_1743,N_19747,N_19699);
nand UO_1744 (O_1744,N_19891,N_19543);
and UO_1745 (O_1745,N_19607,N_19507);
nand UO_1746 (O_1746,N_19896,N_19543);
nand UO_1747 (O_1747,N_19594,N_19988);
or UO_1748 (O_1748,N_19640,N_19875);
or UO_1749 (O_1749,N_19645,N_19540);
nor UO_1750 (O_1750,N_19887,N_19985);
nand UO_1751 (O_1751,N_19807,N_19923);
and UO_1752 (O_1752,N_19711,N_19500);
nor UO_1753 (O_1753,N_19877,N_19758);
or UO_1754 (O_1754,N_19562,N_19844);
and UO_1755 (O_1755,N_19738,N_19957);
and UO_1756 (O_1756,N_19769,N_19557);
nand UO_1757 (O_1757,N_19796,N_19548);
nand UO_1758 (O_1758,N_19822,N_19517);
nor UO_1759 (O_1759,N_19550,N_19949);
nor UO_1760 (O_1760,N_19618,N_19779);
and UO_1761 (O_1761,N_19615,N_19676);
and UO_1762 (O_1762,N_19662,N_19976);
and UO_1763 (O_1763,N_19753,N_19605);
and UO_1764 (O_1764,N_19680,N_19706);
nor UO_1765 (O_1765,N_19876,N_19743);
nand UO_1766 (O_1766,N_19612,N_19624);
nor UO_1767 (O_1767,N_19652,N_19691);
and UO_1768 (O_1768,N_19512,N_19766);
xnor UO_1769 (O_1769,N_19853,N_19803);
xor UO_1770 (O_1770,N_19546,N_19950);
nand UO_1771 (O_1771,N_19766,N_19587);
xnor UO_1772 (O_1772,N_19750,N_19776);
or UO_1773 (O_1773,N_19546,N_19567);
nor UO_1774 (O_1774,N_19658,N_19501);
nor UO_1775 (O_1775,N_19697,N_19573);
or UO_1776 (O_1776,N_19572,N_19778);
and UO_1777 (O_1777,N_19671,N_19934);
nand UO_1778 (O_1778,N_19910,N_19643);
nand UO_1779 (O_1779,N_19842,N_19596);
xor UO_1780 (O_1780,N_19875,N_19541);
xor UO_1781 (O_1781,N_19905,N_19740);
nor UO_1782 (O_1782,N_19779,N_19719);
xor UO_1783 (O_1783,N_19500,N_19573);
xor UO_1784 (O_1784,N_19619,N_19710);
or UO_1785 (O_1785,N_19565,N_19838);
or UO_1786 (O_1786,N_19794,N_19808);
nor UO_1787 (O_1787,N_19767,N_19709);
or UO_1788 (O_1788,N_19968,N_19906);
nor UO_1789 (O_1789,N_19775,N_19624);
nand UO_1790 (O_1790,N_19922,N_19733);
xor UO_1791 (O_1791,N_19732,N_19790);
and UO_1792 (O_1792,N_19897,N_19889);
or UO_1793 (O_1793,N_19876,N_19742);
or UO_1794 (O_1794,N_19519,N_19626);
nor UO_1795 (O_1795,N_19916,N_19881);
or UO_1796 (O_1796,N_19911,N_19642);
or UO_1797 (O_1797,N_19649,N_19609);
and UO_1798 (O_1798,N_19505,N_19502);
xor UO_1799 (O_1799,N_19676,N_19816);
nand UO_1800 (O_1800,N_19877,N_19652);
xnor UO_1801 (O_1801,N_19768,N_19565);
nand UO_1802 (O_1802,N_19719,N_19509);
nor UO_1803 (O_1803,N_19716,N_19703);
nor UO_1804 (O_1804,N_19838,N_19519);
nor UO_1805 (O_1805,N_19789,N_19980);
or UO_1806 (O_1806,N_19627,N_19518);
and UO_1807 (O_1807,N_19756,N_19866);
and UO_1808 (O_1808,N_19933,N_19741);
xnor UO_1809 (O_1809,N_19663,N_19578);
xnor UO_1810 (O_1810,N_19638,N_19920);
nor UO_1811 (O_1811,N_19619,N_19799);
nand UO_1812 (O_1812,N_19863,N_19520);
and UO_1813 (O_1813,N_19700,N_19730);
xnor UO_1814 (O_1814,N_19923,N_19705);
nand UO_1815 (O_1815,N_19668,N_19859);
nor UO_1816 (O_1816,N_19714,N_19847);
or UO_1817 (O_1817,N_19753,N_19621);
nand UO_1818 (O_1818,N_19709,N_19850);
or UO_1819 (O_1819,N_19984,N_19654);
or UO_1820 (O_1820,N_19678,N_19619);
xnor UO_1821 (O_1821,N_19629,N_19583);
nand UO_1822 (O_1822,N_19538,N_19754);
and UO_1823 (O_1823,N_19932,N_19940);
and UO_1824 (O_1824,N_19855,N_19985);
and UO_1825 (O_1825,N_19571,N_19855);
and UO_1826 (O_1826,N_19652,N_19654);
xnor UO_1827 (O_1827,N_19998,N_19679);
xnor UO_1828 (O_1828,N_19648,N_19610);
nand UO_1829 (O_1829,N_19640,N_19784);
and UO_1830 (O_1830,N_19791,N_19534);
and UO_1831 (O_1831,N_19990,N_19620);
xor UO_1832 (O_1832,N_19695,N_19958);
nand UO_1833 (O_1833,N_19861,N_19642);
and UO_1834 (O_1834,N_19804,N_19997);
and UO_1835 (O_1835,N_19814,N_19951);
and UO_1836 (O_1836,N_19670,N_19998);
xor UO_1837 (O_1837,N_19706,N_19526);
nor UO_1838 (O_1838,N_19730,N_19974);
nor UO_1839 (O_1839,N_19757,N_19780);
or UO_1840 (O_1840,N_19813,N_19685);
nor UO_1841 (O_1841,N_19795,N_19518);
xnor UO_1842 (O_1842,N_19625,N_19617);
or UO_1843 (O_1843,N_19933,N_19980);
and UO_1844 (O_1844,N_19740,N_19690);
nand UO_1845 (O_1845,N_19946,N_19869);
nor UO_1846 (O_1846,N_19525,N_19796);
and UO_1847 (O_1847,N_19723,N_19505);
or UO_1848 (O_1848,N_19641,N_19637);
nand UO_1849 (O_1849,N_19577,N_19706);
and UO_1850 (O_1850,N_19794,N_19767);
nor UO_1851 (O_1851,N_19576,N_19959);
or UO_1852 (O_1852,N_19638,N_19534);
and UO_1853 (O_1853,N_19650,N_19693);
and UO_1854 (O_1854,N_19859,N_19789);
and UO_1855 (O_1855,N_19660,N_19874);
xor UO_1856 (O_1856,N_19603,N_19786);
or UO_1857 (O_1857,N_19738,N_19793);
xor UO_1858 (O_1858,N_19998,N_19693);
xor UO_1859 (O_1859,N_19889,N_19751);
or UO_1860 (O_1860,N_19579,N_19822);
or UO_1861 (O_1861,N_19986,N_19911);
or UO_1862 (O_1862,N_19713,N_19715);
and UO_1863 (O_1863,N_19611,N_19552);
xnor UO_1864 (O_1864,N_19512,N_19704);
xor UO_1865 (O_1865,N_19669,N_19633);
nand UO_1866 (O_1866,N_19798,N_19666);
nor UO_1867 (O_1867,N_19778,N_19684);
nand UO_1868 (O_1868,N_19982,N_19893);
and UO_1869 (O_1869,N_19692,N_19612);
nor UO_1870 (O_1870,N_19585,N_19753);
nor UO_1871 (O_1871,N_19673,N_19671);
or UO_1872 (O_1872,N_19638,N_19518);
or UO_1873 (O_1873,N_19910,N_19641);
nor UO_1874 (O_1874,N_19513,N_19511);
nand UO_1875 (O_1875,N_19862,N_19841);
or UO_1876 (O_1876,N_19667,N_19984);
nand UO_1877 (O_1877,N_19536,N_19924);
and UO_1878 (O_1878,N_19969,N_19786);
and UO_1879 (O_1879,N_19593,N_19687);
nor UO_1880 (O_1880,N_19653,N_19875);
xor UO_1881 (O_1881,N_19580,N_19613);
or UO_1882 (O_1882,N_19662,N_19834);
and UO_1883 (O_1883,N_19784,N_19837);
nor UO_1884 (O_1884,N_19951,N_19959);
xnor UO_1885 (O_1885,N_19732,N_19997);
or UO_1886 (O_1886,N_19727,N_19987);
nor UO_1887 (O_1887,N_19894,N_19833);
or UO_1888 (O_1888,N_19599,N_19771);
nor UO_1889 (O_1889,N_19791,N_19624);
xor UO_1890 (O_1890,N_19966,N_19633);
xnor UO_1891 (O_1891,N_19570,N_19827);
xor UO_1892 (O_1892,N_19987,N_19745);
nor UO_1893 (O_1893,N_19709,N_19843);
xnor UO_1894 (O_1894,N_19947,N_19975);
xnor UO_1895 (O_1895,N_19723,N_19754);
and UO_1896 (O_1896,N_19926,N_19604);
and UO_1897 (O_1897,N_19711,N_19605);
nor UO_1898 (O_1898,N_19684,N_19853);
nand UO_1899 (O_1899,N_19525,N_19829);
or UO_1900 (O_1900,N_19769,N_19690);
nand UO_1901 (O_1901,N_19736,N_19618);
xnor UO_1902 (O_1902,N_19541,N_19672);
nand UO_1903 (O_1903,N_19632,N_19835);
and UO_1904 (O_1904,N_19911,N_19518);
nor UO_1905 (O_1905,N_19783,N_19513);
xor UO_1906 (O_1906,N_19813,N_19669);
nor UO_1907 (O_1907,N_19784,N_19547);
or UO_1908 (O_1908,N_19974,N_19969);
xnor UO_1909 (O_1909,N_19642,N_19997);
nand UO_1910 (O_1910,N_19868,N_19722);
nor UO_1911 (O_1911,N_19584,N_19980);
nor UO_1912 (O_1912,N_19626,N_19644);
xnor UO_1913 (O_1913,N_19501,N_19676);
or UO_1914 (O_1914,N_19583,N_19730);
xnor UO_1915 (O_1915,N_19640,N_19635);
nand UO_1916 (O_1916,N_19653,N_19899);
nor UO_1917 (O_1917,N_19690,N_19813);
nand UO_1918 (O_1918,N_19976,N_19688);
nand UO_1919 (O_1919,N_19640,N_19614);
nand UO_1920 (O_1920,N_19842,N_19992);
nor UO_1921 (O_1921,N_19933,N_19701);
nand UO_1922 (O_1922,N_19628,N_19530);
nand UO_1923 (O_1923,N_19990,N_19983);
or UO_1924 (O_1924,N_19573,N_19999);
xor UO_1925 (O_1925,N_19564,N_19757);
nand UO_1926 (O_1926,N_19799,N_19857);
and UO_1927 (O_1927,N_19926,N_19831);
nor UO_1928 (O_1928,N_19750,N_19994);
nor UO_1929 (O_1929,N_19754,N_19873);
or UO_1930 (O_1930,N_19671,N_19897);
xor UO_1931 (O_1931,N_19928,N_19965);
xnor UO_1932 (O_1932,N_19560,N_19614);
and UO_1933 (O_1933,N_19820,N_19528);
nand UO_1934 (O_1934,N_19915,N_19872);
xor UO_1935 (O_1935,N_19550,N_19579);
or UO_1936 (O_1936,N_19847,N_19643);
or UO_1937 (O_1937,N_19873,N_19794);
nand UO_1938 (O_1938,N_19663,N_19642);
or UO_1939 (O_1939,N_19730,N_19729);
nor UO_1940 (O_1940,N_19946,N_19612);
xnor UO_1941 (O_1941,N_19573,N_19907);
or UO_1942 (O_1942,N_19988,N_19924);
nor UO_1943 (O_1943,N_19750,N_19828);
xnor UO_1944 (O_1944,N_19886,N_19782);
and UO_1945 (O_1945,N_19639,N_19579);
or UO_1946 (O_1946,N_19958,N_19543);
nand UO_1947 (O_1947,N_19622,N_19764);
nor UO_1948 (O_1948,N_19604,N_19862);
or UO_1949 (O_1949,N_19779,N_19579);
or UO_1950 (O_1950,N_19743,N_19828);
and UO_1951 (O_1951,N_19609,N_19916);
xor UO_1952 (O_1952,N_19962,N_19751);
nand UO_1953 (O_1953,N_19705,N_19619);
or UO_1954 (O_1954,N_19711,N_19866);
nand UO_1955 (O_1955,N_19728,N_19973);
nand UO_1956 (O_1956,N_19834,N_19713);
and UO_1957 (O_1957,N_19707,N_19579);
and UO_1958 (O_1958,N_19832,N_19829);
and UO_1959 (O_1959,N_19597,N_19935);
nand UO_1960 (O_1960,N_19582,N_19859);
nor UO_1961 (O_1961,N_19917,N_19679);
xnor UO_1962 (O_1962,N_19853,N_19948);
nor UO_1963 (O_1963,N_19939,N_19625);
and UO_1964 (O_1964,N_19840,N_19505);
or UO_1965 (O_1965,N_19582,N_19755);
xor UO_1966 (O_1966,N_19745,N_19687);
and UO_1967 (O_1967,N_19663,N_19894);
xnor UO_1968 (O_1968,N_19926,N_19782);
nor UO_1969 (O_1969,N_19711,N_19768);
nor UO_1970 (O_1970,N_19982,N_19946);
nor UO_1971 (O_1971,N_19645,N_19850);
and UO_1972 (O_1972,N_19535,N_19973);
nor UO_1973 (O_1973,N_19821,N_19588);
and UO_1974 (O_1974,N_19826,N_19911);
xor UO_1975 (O_1975,N_19577,N_19544);
nand UO_1976 (O_1976,N_19696,N_19580);
and UO_1977 (O_1977,N_19939,N_19684);
and UO_1978 (O_1978,N_19918,N_19832);
xnor UO_1979 (O_1979,N_19671,N_19504);
nor UO_1980 (O_1980,N_19573,N_19794);
or UO_1981 (O_1981,N_19544,N_19535);
and UO_1982 (O_1982,N_19920,N_19537);
or UO_1983 (O_1983,N_19997,N_19522);
and UO_1984 (O_1984,N_19828,N_19891);
xor UO_1985 (O_1985,N_19774,N_19650);
nand UO_1986 (O_1986,N_19607,N_19880);
or UO_1987 (O_1987,N_19566,N_19530);
or UO_1988 (O_1988,N_19575,N_19630);
nand UO_1989 (O_1989,N_19561,N_19796);
or UO_1990 (O_1990,N_19969,N_19823);
nand UO_1991 (O_1991,N_19826,N_19845);
nand UO_1992 (O_1992,N_19582,N_19529);
nor UO_1993 (O_1993,N_19608,N_19605);
nand UO_1994 (O_1994,N_19945,N_19598);
nand UO_1995 (O_1995,N_19940,N_19740);
xor UO_1996 (O_1996,N_19716,N_19655);
nand UO_1997 (O_1997,N_19839,N_19826);
nand UO_1998 (O_1998,N_19817,N_19777);
xnor UO_1999 (O_1999,N_19760,N_19926);
xnor UO_2000 (O_2000,N_19824,N_19888);
or UO_2001 (O_2001,N_19651,N_19952);
nor UO_2002 (O_2002,N_19709,N_19831);
nand UO_2003 (O_2003,N_19737,N_19710);
and UO_2004 (O_2004,N_19629,N_19876);
nor UO_2005 (O_2005,N_19625,N_19785);
and UO_2006 (O_2006,N_19743,N_19624);
or UO_2007 (O_2007,N_19969,N_19843);
nand UO_2008 (O_2008,N_19938,N_19508);
and UO_2009 (O_2009,N_19978,N_19982);
and UO_2010 (O_2010,N_19692,N_19602);
nor UO_2011 (O_2011,N_19703,N_19744);
and UO_2012 (O_2012,N_19615,N_19660);
nor UO_2013 (O_2013,N_19591,N_19600);
xnor UO_2014 (O_2014,N_19681,N_19578);
nand UO_2015 (O_2015,N_19908,N_19984);
and UO_2016 (O_2016,N_19500,N_19966);
nand UO_2017 (O_2017,N_19725,N_19910);
or UO_2018 (O_2018,N_19839,N_19611);
nor UO_2019 (O_2019,N_19870,N_19771);
or UO_2020 (O_2020,N_19508,N_19636);
or UO_2021 (O_2021,N_19524,N_19914);
nand UO_2022 (O_2022,N_19818,N_19715);
nor UO_2023 (O_2023,N_19835,N_19830);
and UO_2024 (O_2024,N_19946,N_19932);
and UO_2025 (O_2025,N_19581,N_19916);
or UO_2026 (O_2026,N_19538,N_19865);
nor UO_2027 (O_2027,N_19760,N_19852);
nor UO_2028 (O_2028,N_19974,N_19949);
nor UO_2029 (O_2029,N_19947,N_19626);
or UO_2030 (O_2030,N_19935,N_19600);
nand UO_2031 (O_2031,N_19791,N_19927);
and UO_2032 (O_2032,N_19807,N_19628);
and UO_2033 (O_2033,N_19850,N_19950);
and UO_2034 (O_2034,N_19717,N_19977);
or UO_2035 (O_2035,N_19929,N_19939);
nor UO_2036 (O_2036,N_19909,N_19904);
or UO_2037 (O_2037,N_19859,N_19529);
xnor UO_2038 (O_2038,N_19988,N_19661);
nor UO_2039 (O_2039,N_19844,N_19838);
nor UO_2040 (O_2040,N_19537,N_19757);
nor UO_2041 (O_2041,N_19805,N_19564);
and UO_2042 (O_2042,N_19793,N_19596);
nor UO_2043 (O_2043,N_19929,N_19648);
and UO_2044 (O_2044,N_19673,N_19989);
or UO_2045 (O_2045,N_19521,N_19633);
nor UO_2046 (O_2046,N_19761,N_19516);
and UO_2047 (O_2047,N_19605,N_19767);
and UO_2048 (O_2048,N_19564,N_19683);
nand UO_2049 (O_2049,N_19598,N_19781);
nand UO_2050 (O_2050,N_19508,N_19687);
nor UO_2051 (O_2051,N_19870,N_19752);
and UO_2052 (O_2052,N_19724,N_19604);
xnor UO_2053 (O_2053,N_19763,N_19546);
nand UO_2054 (O_2054,N_19783,N_19639);
nor UO_2055 (O_2055,N_19959,N_19984);
nand UO_2056 (O_2056,N_19649,N_19982);
or UO_2057 (O_2057,N_19689,N_19782);
nor UO_2058 (O_2058,N_19842,N_19717);
and UO_2059 (O_2059,N_19545,N_19907);
xor UO_2060 (O_2060,N_19687,N_19661);
xor UO_2061 (O_2061,N_19944,N_19900);
nand UO_2062 (O_2062,N_19707,N_19660);
nand UO_2063 (O_2063,N_19729,N_19559);
nor UO_2064 (O_2064,N_19740,N_19858);
nor UO_2065 (O_2065,N_19618,N_19596);
xnor UO_2066 (O_2066,N_19542,N_19547);
or UO_2067 (O_2067,N_19576,N_19989);
nand UO_2068 (O_2068,N_19814,N_19719);
xnor UO_2069 (O_2069,N_19881,N_19939);
and UO_2070 (O_2070,N_19695,N_19646);
and UO_2071 (O_2071,N_19952,N_19713);
and UO_2072 (O_2072,N_19657,N_19530);
and UO_2073 (O_2073,N_19678,N_19638);
xor UO_2074 (O_2074,N_19980,N_19998);
and UO_2075 (O_2075,N_19959,N_19915);
and UO_2076 (O_2076,N_19780,N_19865);
and UO_2077 (O_2077,N_19756,N_19951);
or UO_2078 (O_2078,N_19886,N_19733);
nor UO_2079 (O_2079,N_19676,N_19965);
nor UO_2080 (O_2080,N_19596,N_19688);
nand UO_2081 (O_2081,N_19870,N_19839);
nor UO_2082 (O_2082,N_19943,N_19999);
or UO_2083 (O_2083,N_19658,N_19760);
nor UO_2084 (O_2084,N_19960,N_19928);
nor UO_2085 (O_2085,N_19844,N_19708);
xnor UO_2086 (O_2086,N_19859,N_19870);
xor UO_2087 (O_2087,N_19713,N_19853);
xnor UO_2088 (O_2088,N_19941,N_19955);
nand UO_2089 (O_2089,N_19515,N_19720);
nor UO_2090 (O_2090,N_19520,N_19565);
and UO_2091 (O_2091,N_19670,N_19790);
xor UO_2092 (O_2092,N_19817,N_19688);
xnor UO_2093 (O_2093,N_19524,N_19707);
nor UO_2094 (O_2094,N_19745,N_19831);
or UO_2095 (O_2095,N_19657,N_19519);
or UO_2096 (O_2096,N_19718,N_19557);
and UO_2097 (O_2097,N_19960,N_19829);
nor UO_2098 (O_2098,N_19779,N_19990);
nand UO_2099 (O_2099,N_19779,N_19685);
nand UO_2100 (O_2100,N_19994,N_19722);
and UO_2101 (O_2101,N_19749,N_19794);
xnor UO_2102 (O_2102,N_19763,N_19676);
nand UO_2103 (O_2103,N_19908,N_19642);
xnor UO_2104 (O_2104,N_19568,N_19854);
or UO_2105 (O_2105,N_19985,N_19577);
nand UO_2106 (O_2106,N_19857,N_19860);
nor UO_2107 (O_2107,N_19574,N_19571);
nor UO_2108 (O_2108,N_19873,N_19884);
or UO_2109 (O_2109,N_19775,N_19774);
nand UO_2110 (O_2110,N_19548,N_19569);
and UO_2111 (O_2111,N_19812,N_19940);
nand UO_2112 (O_2112,N_19634,N_19748);
and UO_2113 (O_2113,N_19939,N_19951);
and UO_2114 (O_2114,N_19794,N_19632);
xnor UO_2115 (O_2115,N_19926,N_19829);
and UO_2116 (O_2116,N_19521,N_19825);
nor UO_2117 (O_2117,N_19891,N_19627);
and UO_2118 (O_2118,N_19601,N_19906);
or UO_2119 (O_2119,N_19749,N_19714);
nor UO_2120 (O_2120,N_19516,N_19997);
nor UO_2121 (O_2121,N_19818,N_19616);
nor UO_2122 (O_2122,N_19792,N_19704);
xor UO_2123 (O_2123,N_19810,N_19603);
or UO_2124 (O_2124,N_19680,N_19857);
or UO_2125 (O_2125,N_19515,N_19859);
nand UO_2126 (O_2126,N_19659,N_19946);
nor UO_2127 (O_2127,N_19519,N_19602);
nand UO_2128 (O_2128,N_19842,N_19566);
nand UO_2129 (O_2129,N_19746,N_19708);
and UO_2130 (O_2130,N_19972,N_19897);
or UO_2131 (O_2131,N_19835,N_19635);
nor UO_2132 (O_2132,N_19864,N_19560);
nand UO_2133 (O_2133,N_19565,N_19834);
nand UO_2134 (O_2134,N_19522,N_19903);
nand UO_2135 (O_2135,N_19680,N_19610);
and UO_2136 (O_2136,N_19901,N_19963);
nor UO_2137 (O_2137,N_19660,N_19555);
or UO_2138 (O_2138,N_19550,N_19632);
nor UO_2139 (O_2139,N_19531,N_19813);
nor UO_2140 (O_2140,N_19626,N_19787);
and UO_2141 (O_2141,N_19692,N_19858);
and UO_2142 (O_2142,N_19633,N_19829);
xor UO_2143 (O_2143,N_19642,N_19817);
xor UO_2144 (O_2144,N_19746,N_19625);
nand UO_2145 (O_2145,N_19903,N_19772);
nor UO_2146 (O_2146,N_19637,N_19749);
nor UO_2147 (O_2147,N_19760,N_19573);
and UO_2148 (O_2148,N_19509,N_19672);
nor UO_2149 (O_2149,N_19551,N_19806);
and UO_2150 (O_2150,N_19647,N_19669);
nand UO_2151 (O_2151,N_19986,N_19799);
xor UO_2152 (O_2152,N_19826,N_19533);
or UO_2153 (O_2153,N_19841,N_19698);
and UO_2154 (O_2154,N_19810,N_19918);
nor UO_2155 (O_2155,N_19848,N_19586);
nor UO_2156 (O_2156,N_19666,N_19627);
nand UO_2157 (O_2157,N_19619,N_19600);
and UO_2158 (O_2158,N_19833,N_19798);
or UO_2159 (O_2159,N_19903,N_19848);
xor UO_2160 (O_2160,N_19873,N_19842);
xor UO_2161 (O_2161,N_19512,N_19543);
nand UO_2162 (O_2162,N_19769,N_19563);
xor UO_2163 (O_2163,N_19783,N_19942);
xnor UO_2164 (O_2164,N_19908,N_19929);
or UO_2165 (O_2165,N_19524,N_19588);
and UO_2166 (O_2166,N_19740,N_19778);
nor UO_2167 (O_2167,N_19954,N_19806);
nor UO_2168 (O_2168,N_19559,N_19749);
nor UO_2169 (O_2169,N_19500,N_19677);
nand UO_2170 (O_2170,N_19760,N_19887);
and UO_2171 (O_2171,N_19723,N_19651);
or UO_2172 (O_2172,N_19772,N_19669);
and UO_2173 (O_2173,N_19565,N_19818);
or UO_2174 (O_2174,N_19834,N_19897);
xnor UO_2175 (O_2175,N_19846,N_19901);
xor UO_2176 (O_2176,N_19688,N_19511);
nand UO_2177 (O_2177,N_19889,N_19586);
xor UO_2178 (O_2178,N_19670,N_19531);
nand UO_2179 (O_2179,N_19928,N_19747);
or UO_2180 (O_2180,N_19749,N_19884);
or UO_2181 (O_2181,N_19602,N_19567);
or UO_2182 (O_2182,N_19829,N_19556);
and UO_2183 (O_2183,N_19801,N_19912);
and UO_2184 (O_2184,N_19846,N_19987);
and UO_2185 (O_2185,N_19610,N_19686);
xnor UO_2186 (O_2186,N_19789,N_19590);
nand UO_2187 (O_2187,N_19685,N_19547);
or UO_2188 (O_2188,N_19951,N_19685);
and UO_2189 (O_2189,N_19729,N_19719);
nand UO_2190 (O_2190,N_19677,N_19952);
nor UO_2191 (O_2191,N_19995,N_19930);
nor UO_2192 (O_2192,N_19712,N_19664);
nor UO_2193 (O_2193,N_19981,N_19852);
and UO_2194 (O_2194,N_19608,N_19791);
and UO_2195 (O_2195,N_19785,N_19800);
nand UO_2196 (O_2196,N_19893,N_19751);
xnor UO_2197 (O_2197,N_19608,N_19874);
and UO_2198 (O_2198,N_19709,N_19844);
nor UO_2199 (O_2199,N_19903,N_19706);
or UO_2200 (O_2200,N_19984,N_19626);
nor UO_2201 (O_2201,N_19512,N_19639);
and UO_2202 (O_2202,N_19961,N_19628);
xnor UO_2203 (O_2203,N_19830,N_19509);
or UO_2204 (O_2204,N_19530,N_19685);
nor UO_2205 (O_2205,N_19682,N_19511);
and UO_2206 (O_2206,N_19578,N_19575);
and UO_2207 (O_2207,N_19594,N_19775);
or UO_2208 (O_2208,N_19947,N_19912);
or UO_2209 (O_2209,N_19802,N_19677);
nand UO_2210 (O_2210,N_19784,N_19986);
xnor UO_2211 (O_2211,N_19805,N_19565);
xor UO_2212 (O_2212,N_19743,N_19809);
nor UO_2213 (O_2213,N_19681,N_19860);
nand UO_2214 (O_2214,N_19899,N_19953);
and UO_2215 (O_2215,N_19984,N_19880);
nor UO_2216 (O_2216,N_19918,N_19596);
or UO_2217 (O_2217,N_19709,N_19579);
nand UO_2218 (O_2218,N_19936,N_19787);
and UO_2219 (O_2219,N_19846,N_19886);
or UO_2220 (O_2220,N_19862,N_19919);
and UO_2221 (O_2221,N_19700,N_19621);
or UO_2222 (O_2222,N_19518,N_19585);
or UO_2223 (O_2223,N_19529,N_19780);
and UO_2224 (O_2224,N_19902,N_19780);
xor UO_2225 (O_2225,N_19903,N_19656);
xnor UO_2226 (O_2226,N_19999,N_19864);
xor UO_2227 (O_2227,N_19852,N_19544);
nand UO_2228 (O_2228,N_19532,N_19724);
or UO_2229 (O_2229,N_19871,N_19940);
and UO_2230 (O_2230,N_19945,N_19689);
or UO_2231 (O_2231,N_19817,N_19630);
xor UO_2232 (O_2232,N_19845,N_19793);
nor UO_2233 (O_2233,N_19544,N_19923);
or UO_2234 (O_2234,N_19646,N_19898);
or UO_2235 (O_2235,N_19983,N_19685);
nor UO_2236 (O_2236,N_19510,N_19830);
nor UO_2237 (O_2237,N_19815,N_19842);
xnor UO_2238 (O_2238,N_19788,N_19794);
or UO_2239 (O_2239,N_19898,N_19661);
and UO_2240 (O_2240,N_19658,N_19679);
nor UO_2241 (O_2241,N_19679,N_19863);
xor UO_2242 (O_2242,N_19634,N_19603);
nor UO_2243 (O_2243,N_19684,N_19809);
and UO_2244 (O_2244,N_19513,N_19803);
nand UO_2245 (O_2245,N_19682,N_19628);
and UO_2246 (O_2246,N_19964,N_19970);
and UO_2247 (O_2247,N_19669,N_19706);
nand UO_2248 (O_2248,N_19647,N_19622);
nor UO_2249 (O_2249,N_19502,N_19897);
nor UO_2250 (O_2250,N_19943,N_19633);
or UO_2251 (O_2251,N_19697,N_19682);
nor UO_2252 (O_2252,N_19530,N_19880);
nand UO_2253 (O_2253,N_19821,N_19977);
or UO_2254 (O_2254,N_19691,N_19661);
and UO_2255 (O_2255,N_19758,N_19887);
or UO_2256 (O_2256,N_19814,N_19872);
xnor UO_2257 (O_2257,N_19923,N_19664);
nor UO_2258 (O_2258,N_19958,N_19540);
xor UO_2259 (O_2259,N_19877,N_19842);
or UO_2260 (O_2260,N_19504,N_19731);
or UO_2261 (O_2261,N_19891,N_19886);
nor UO_2262 (O_2262,N_19823,N_19503);
xor UO_2263 (O_2263,N_19516,N_19518);
or UO_2264 (O_2264,N_19527,N_19835);
nand UO_2265 (O_2265,N_19593,N_19635);
nand UO_2266 (O_2266,N_19840,N_19590);
nor UO_2267 (O_2267,N_19538,N_19675);
and UO_2268 (O_2268,N_19925,N_19785);
nor UO_2269 (O_2269,N_19749,N_19939);
and UO_2270 (O_2270,N_19848,N_19863);
xnor UO_2271 (O_2271,N_19683,N_19738);
and UO_2272 (O_2272,N_19982,N_19784);
nand UO_2273 (O_2273,N_19821,N_19839);
nand UO_2274 (O_2274,N_19784,N_19840);
xor UO_2275 (O_2275,N_19865,N_19948);
nor UO_2276 (O_2276,N_19812,N_19648);
nor UO_2277 (O_2277,N_19941,N_19524);
and UO_2278 (O_2278,N_19783,N_19701);
and UO_2279 (O_2279,N_19885,N_19926);
and UO_2280 (O_2280,N_19870,N_19786);
and UO_2281 (O_2281,N_19909,N_19741);
and UO_2282 (O_2282,N_19671,N_19566);
xnor UO_2283 (O_2283,N_19972,N_19529);
nor UO_2284 (O_2284,N_19513,N_19637);
or UO_2285 (O_2285,N_19967,N_19915);
nand UO_2286 (O_2286,N_19526,N_19782);
nor UO_2287 (O_2287,N_19511,N_19894);
and UO_2288 (O_2288,N_19943,N_19936);
or UO_2289 (O_2289,N_19636,N_19566);
and UO_2290 (O_2290,N_19558,N_19749);
or UO_2291 (O_2291,N_19754,N_19890);
nor UO_2292 (O_2292,N_19960,N_19991);
nand UO_2293 (O_2293,N_19727,N_19594);
nand UO_2294 (O_2294,N_19907,N_19972);
nand UO_2295 (O_2295,N_19755,N_19629);
or UO_2296 (O_2296,N_19894,N_19880);
nor UO_2297 (O_2297,N_19501,N_19592);
and UO_2298 (O_2298,N_19875,N_19553);
or UO_2299 (O_2299,N_19531,N_19632);
and UO_2300 (O_2300,N_19868,N_19657);
nand UO_2301 (O_2301,N_19592,N_19836);
nand UO_2302 (O_2302,N_19792,N_19972);
xnor UO_2303 (O_2303,N_19726,N_19913);
or UO_2304 (O_2304,N_19511,N_19872);
nand UO_2305 (O_2305,N_19841,N_19996);
nor UO_2306 (O_2306,N_19948,N_19829);
nor UO_2307 (O_2307,N_19747,N_19778);
nand UO_2308 (O_2308,N_19726,N_19932);
and UO_2309 (O_2309,N_19647,N_19696);
nand UO_2310 (O_2310,N_19763,N_19641);
nor UO_2311 (O_2311,N_19680,N_19583);
and UO_2312 (O_2312,N_19610,N_19751);
nor UO_2313 (O_2313,N_19700,N_19506);
xnor UO_2314 (O_2314,N_19595,N_19772);
nand UO_2315 (O_2315,N_19869,N_19985);
or UO_2316 (O_2316,N_19558,N_19636);
or UO_2317 (O_2317,N_19923,N_19703);
xnor UO_2318 (O_2318,N_19952,N_19909);
xor UO_2319 (O_2319,N_19675,N_19998);
nor UO_2320 (O_2320,N_19927,N_19502);
nand UO_2321 (O_2321,N_19949,N_19986);
nor UO_2322 (O_2322,N_19938,N_19545);
xnor UO_2323 (O_2323,N_19500,N_19709);
or UO_2324 (O_2324,N_19639,N_19645);
nor UO_2325 (O_2325,N_19862,N_19730);
xor UO_2326 (O_2326,N_19799,N_19831);
nor UO_2327 (O_2327,N_19939,N_19835);
or UO_2328 (O_2328,N_19845,N_19821);
nor UO_2329 (O_2329,N_19856,N_19942);
or UO_2330 (O_2330,N_19662,N_19792);
or UO_2331 (O_2331,N_19605,N_19948);
and UO_2332 (O_2332,N_19616,N_19600);
nor UO_2333 (O_2333,N_19631,N_19915);
xnor UO_2334 (O_2334,N_19841,N_19709);
xnor UO_2335 (O_2335,N_19649,N_19683);
nor UO_2336 (O_2336,N_19733,N_19562);
xor UO_2337 (O_2337,N_19932,N_19614);
xor UO_2338 (O_2338,N_19630,N_19803);
or UO_2339 (O_2339,N_19798,N_19864);
xor UO_2340 (O_2340,N_19848,N_19950);
xnor UO_2341 (O_2341,N_19827,N_19825);
and UO_2342 (O_2342,N_19770,N_19781);
or UO_2343 (O_2343,N_19852,N_19887);
xnor UO_2344 (O_2344,N_19706,N_19829);
nand UO_2345 (O_2345,N_19888,N_19919);
nand UO_2346 (O_2346,N_19909,N_19987);
or UO_2347 (O_2347,N_19757,N_19820);
nor UO_2348 (O_2348,N_19993,N_19777);
or UO_2349 (O_2349,N_19541,N_19651);
xor UO_2350 (O_2350,N_19952,N_19537);
or UO_2351 (O_2351,N_19647,N_19770);
nor UO_2352 (O_2352,N_19913,N_19554);
or UO_2353 (O_2353,N_19548,N_19584);
or UO_2354 (O_2354,N_19758,N_19812);
xnor UO_2355 (O_2355,N_19811,N_19596);
xnor UO_2356 (O_2356,N_19931,N_19771);
nor UO_2357 (O_2357,N_19621,N_19715);
nor UO_2358 (O_2358,N_19914,N_19929);
or UO_2359 (O_2359,N_19823,N_19629);
nand UO_2360 (O_2360,N_19769,N_19795);
nand UO_2361 (O_2361,N_19765,N_19929);
xor UO_2362 (O_2362,N_19728,N_19631);
nor UO_2363 (O_2363,N_19698,N_19911);
or UO_2364 (O_2364,N_19967,N_19999);
xor UO_2365 (O_2365,N_19924,N_19618);
nor UO_2366 (O_2366,N_19859,N_19738);
nor UO_2367 (O_2367,N_19905,N_19693);
nand UO_2368 (O_2368,N_19708,N_19814);
or UO_2369 (O_2369,N_19839,N_19636);
nand UO_2370 (O_2370,N_19743,N_19952);
xor UO_2371 (O_2371,N_19900,N_19813);
xor UO_2372 (O_2372,N_19877,N_19975);
nor UO_2373 (O_2373,N_19920,N_19970);
nand UO_2374 (O_2374,N_19663,N_19890);
xor UO_2375 (O_2375,N_19859,N_19711);
nor UO_2376 (O_2376,N_19871,N_19661);
nand UO_2377 (O_2377,N_19890,N_19980);
and UO_2378 (O_2378,N_19541,N_19626);
or UO_2379 (O_2379,N_19876,N_19644);
xor UO_2380 (O_2380,N_19551,N_19728);
xnor UO_2381 (O_2381,N_19872,N_19844);
or UO_2382 (O_2382,N_19983,N_19915);
nand UO_2383 (O_2383,N_19966,N_19647);
nand UO_2384 (O_2384,N_19550,N_19644);
or UO_2385 (O_2385,N_19569,N_19542);
and UO_2386 (O_2386,N_19802,N_19932);
nand UO_2387 (O_2387,N_19700,N_19975);
xnor UO_2388 (O_2388,N_19726,N_19724);
and UO_2389 (O_2389,N_19728,N_19579);
or UO_2390 (O_2390,N_19760,N_19905);
nor UO_2391 (O_2391,N_19683,N_19640);
xnor UO_2392 (O_2392,N_19967,N_19633);
nor UO_2393 (O_2393,N_19573,N_19745);
nand UO_2394 (O_2394,N_19548,N_19786);
xor UO_2395 (O_2395,N_19831,N_19995);
xnor UO_2396 (O_2396,N_19758,N_19507);
or UO_2397 (O_2397,N_19813,N_19510);
nand UO_2398 (O_2398,N_19601,N_19842);
nand UO_2399 (O_2399,N_19593,N_19514);
nor UO_2400 (O_2400,N_19670,N_19882);
nor UO_2401 (O_2401,N_19707,N_19508);
nand UO_2402 (O_2402,N_19525,N_19793);
nor UO_2403 (O_2403,N_19717,N_19754);
xnor UO_2404 (O_2404,N_19754,N_19948);
nor UO_2405 (O_2405,N_19668,N_19751);
nand UO_2406 (O_2406,N_19603,N_19670);
nand UO_2407 (O_2407,N_19946,N_19808);
nand UO_2408 (O_2408,N_19994,N_19936);
nand UO_2409 (O_2409,N_19678,N_19541);
and UO_2410 (O_2410,N_19582,N_19592);
nand UO_2411 (O_2411,N_19678,N_19879);
xor UO_2412 (O_2412,N_19621,N_19878);
nand UO_2413 (O_2413,N_19839,N_19575);
nor UO_2414 (O_2414,N_19918,N_19908);
xnor UO_2415 (O_2415,N_19571,N_19864);
xor UO_2416 (O_2416,N_19959,N_19659);
nand UO_2417 (O_2417,N_19627,N_19956);
or UO_2418 (O_2418,N_19650,N_19827);
and UO_2419 (O_2419,N_19920,N_19513);
and UO_2420 (O_2420,N_19743,N_19914);
and UO_2421 (O_2421,N_19850,N_19995);
and UO_2422 (O_2422,N_19565,N_19645);
xnor UO_2423 (O_2423,N_19849,N_19763);
xor UO_2424 (O_2424,N_19906,N_19771);
xor UO_2425 (O_2425,N_19611,N_19988);
and UO_2426 (O_2426,N_19886,N_19888);
nor UO_2427 (O_2427,N_19539,N_19874);
nor UO_2428 (O_2428,N_19561,N_19570);
xor UO_2429 (O_2429,N_19554,N_19691);
or UO_2430 (O_2430,N_19721,N_19581);
and UO_2431 (O_2431,N_19753,N_19869);
nand UO_2432 (O_2432,N_19625,N_19779);
or UO_2433 (O_2433,N_19774,N_19568);
nor UO_2434 (O_2434,N_19508,N_19583);
and UO_2435 (O_2435,N_19585,N_19578);
xnor UO_2436 (O_2436,N_19870,N_19947);
and UO_2437 (O_2437,N_19785,N_19798);
or UO_2438 (O_2438,N_19782,N_19962);
xnor UO_2439 (O_2439,N_19582,N_19650);
xor UO_2440 (O_2440,N_19693,N_19672);
nor UO_2441 (O_2441,N_19761,N_19678);
xnor UO_2442 (O_2442,N_19619,N_19534);
xnor UO_2443 (O_2443,N_19984,N_19929);
or UO_2444 (O_2444,N_19575,N_19657);
or UO_2445 (O_2445,N_19797,N_19984);
and UO_2446 (O_2446,N_19815,N_19797);
nor UO_2447 (O_2447,N_19978,N_19710);
nor UO_2448 (O_2448,N_19676,N_19568);
xnor UO_2449 (O_2449,N_19974,N_19747);
and UO_2450 (O_2450,N_19688,N_19840);
nor UO_2451 (O_2451,N_19821,N_19917);
nand UO_2452 (O_2452,N_19954,N_19674);
and UO_2453 (O_2453,N_19565,N_19561);
xnor UO_2454 (O_2454,N_19649,N_19679);
or UO_2455 (O_2455,N_19534,N_19665);
and UO_2456 (O_2456,N_19592,N_19754);
xor UO_2457 (O_2457,N_19522,N_19985);
nor UO_2458 (O_2458,N_19665,N_19955);
nor UO_2459 (O_2459,N_19534,N_19905);
or UO_2460 (O_2460,N_19633,N_19897);
xor UO_2461 (O_2461,N_19513,N_19656);
nor UO_2462 (O_2462,N_19969,N_19863);
xor UO_2463 (O_2463,N_19747,N_19758);
nand UO_2464 (O_2464,N_19773,N_19702);
or UO_2465 (O_2465,N_19574,N_19921);
and UO_2466 (O_2466,N_19934,N_19654);
nor UO_2467 (O_2467,N_19905,N_19667);
or UO_2468 (O_2468,N_19629,N_19661);
or UO_2469 (O_2469,N_19832,N_19717);
nor UO_2470 (O_2470,N_19940,N_19754);
nand UO_2471 (O_2471,N_19978,N_19787);
and UO_2472 (O_2472,N_19854,N_19825);
nor UO_2473 (O_2473,N_19945,N_19946);
and UO_2474 (O_2474,N_19871,N_19952);
nor UO_2475 (O_2475,N_19739,N_19791);
nor UO_2476 (O_2476,N_19947,N_19990);
nor UO_2477 (O_2477,N_19688,N_19815);
xor UO_2478 (O_2478,N_19653,N_19982);
nor UO_2479 (O_2479,N_19791,N_19772);
xor UO_2480 (O_2480,N_19832,N_19542);
nand UO_2481 (O_2481,N_19574,N_19815);
and UO_2482 (O_2482,N_19996,N_19997);
nor UO_2483 (O_2483,N_19840,N_19853);
or UO_2484 (O_2484,N_19606,N_19698);
and UO_2485 (O_2485,N_19605,N_19536);
nand UO_2486 (O_2486,N_19719,N_19899);
or UO_2487 (O_2487,N_19757,N_19860);
nor UO_2488 (O_2488,N_19610,N_19727);
nand UO_2489 (O_2489,N_19843,N_19588);
nor UO_2490 (O_2490,N_19637,N_19950);
nor UO_2491 (O_2491,N_19895,N_19695);
nor UO_2492 (O_2492,N_19786,N_19966);
nand UO_2493 (O_2493,N_19804,N_19757);
and UO_2494 (O_2494,N_19785,N_19980);
or UO_2495 (O_2495,N_19732,N_19788);
xnor UO_2496 (O_2496,N_19508,N_19550);
or UO_2497 (O_2497,N_19779,N_19603);
xnor UO_2498 (O_2498,N_19634,N_19831);
nor UO_2499 (O_2499,N_19923,N_19637);
endmodule