module basic_3000_30000_3500_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_259,In_1477);
nand U1 (N_1,In_2305,In_1647);
nand U2 (N_2,In_2278,In_484);
nand U3 (N_3,In_965,In_446);
nand U4 (N_4,In_186,In_1870);
nand U5 (N_5,In_2119,In_2042);
nand U6 (N_6,In_2641,In_788);
nor U7 (N_7,In_312,In_885);
and U8 (N_8,In_2389,In_2002);
nand U9 (N_9,In_1707,In_1979);
and U10 (N_10,In_599,In_2744);
nor U11 (N_11,In_1257,In_757);
nor U12 (N_12,In_225,In_117);
or U13 (N_13,In_1432,In_2829);
nor U14 (N_14,In_1172,In_1997);
or U15 (N_15,In_1832,In_2909);
and U16 (N_16,In_2104,In_985);
nor U17 (N_17,In_1671,In_1759);
or U18 (N_18,In_2133,In_2337);
nor U19 (N_19,In_986,In_724);
or U20 (N_20,In_2738,In_2822);
xor U21 (N_21,In_2523,In_1680);
and U22 (N_22,In_1496,In_2825);
and U23 (N_23,In_1561,In_419);
and U24 (N_24,In_461,In_503);
nor U25 (N_25,In_1460,In_465);
or U26 (N_26,In_379,In_64);
and U27 (N_27,In_2379,In_1925);
xor U28 (N_28,In_410,In_118);
and U29 (N_29,In_262,In_2984);
xor U30 (N_30,In_2053,In_2481);
and U31 (N_31,In_899,In_295);
xnor U32 (N_32,In_2244,In_1139);
or U33 (N_33,In_1327,In_148);
xnor U34 (N_34,In_1623,In_2114);
or U35 (N_35,In_1977,In_2680);
xor U36 (N_36,In_2480,In_391);
nand U37 (N_37,In_1350,In_2232);
or U38 (N_38,In_1904,In_632);
or U39 (N_39,In_2025,In_1417);
nor U40 (N_40,In_2227,In_839);
nor U41 (N_41,In_2638,In_10);
xnor U42 (N_42,In_2218,In_2646);
nor U43 (N_43,In_252,In_611);
or U44 (N_44,In_523,In_1193);
xor U45 (N_45,In_2761,In_293);
or U46 (N_46,In_1634,In_1800);
and U47 (N_47,In_881,In_218);
and U48 (N_48,In_1975,In_91);
nor U49 (N_49,In_2125,In_713);
nor U50 (N_50,In_2078,In_2037);
and U51 (N_51,In_1377,In_2540);
xor U52 (N_52,In_417,In_918);
nand U53 (N_53,In_324,In_404);
or U54 (N_54,In_1912,In_113);
nand U55 (N_55,In_2221,In_2383);
xnor U56 (N_56,In_1365,In_1873);
xor U57 (N_57,In_2277,In_2211);
nand U58 (N_58,In_332,In_1787);
nor U59 (N_59,In_289,In_313);
and U60 (N_60,In_668,In_192);
nand U61 (N_61,In_427,In_1211);
nand U62 (N_62,In_745,In_2422);
nor U63 (N_63,In_1546,In_984);
nor U64 (N_64,In_385,In_1494);
nand U65 (N_65,In_1041,In_1272);
nor U66 (N_66,In_2720,In_2351);
nor U67 (N_67,In_1027,In_2685);
nand U68 (N_68,In_1326,In_2110);
and U69 (N_69,In_2183,In_1716);
and U70 (N_70,In_999,In_2722);
or U71 (N_71,In_2173,In_1370);
xor U72 (N_72,In_2459,In_2556);
xnor U73 (N_73,In_1059,In_209);
and U74 (N_74,In_2513,In_1499);
nand U75 (N_75,In_1543,In_2484);
nor U76 (N_76,In_778,In_1711);
and U77 (N_77,In_2349,In_2327);
nor U78 (N_78,In_1118,In_1701);
nand U79 (N_79,In_700,In_2387);
nor U80 (N_80,In_600,In_2805);
nand U81 (N_81,In_2189,In_1210);
or U82 (N_82,In_445,In_927);
nor U83 (N_83,In_1345,In_257);
nand U84 (N_84,In_2315,In_2317);
or U85 (N_85,In_1306,In_1132);
nor U86 (N_86,In_854,In_2694);
and U87 (N_87,In_2979,In_342);
nor U88 (N_88,In_1259,In_1497);
and U89 (N_89,In_2156,In_1905);
or U90 (N_90,In_634,In_304);
nand U91 (N_91,In_1444,In_2295);
nor U92 (N_92,In_1094,In_2592);
nor U93 (N_93,In_1849,In_2157);
xnor U94 (N_94,In_1673,In_892);
nand U95 (N_95,In_1104,In_2191);
and U96 (N_96,In_860,In_1751);
xnor U97 (N_97,In_1303,In_2094);
or U98 (N_98,In_2443,In_143);
and U99 (N_99,In_2085,In_516);
nand U100 (N_100,In_637,In_684);
nand U101 (N_101,In_916,In_462);
nor U102 (N_102,In_2151,In_644);
and U103 (N_103,In_2759,In_1750);
nor U104 (N_104,In_801,In_2879);
nor U105 (N_105,In_1710,In_2099);
nand U106 (N_106,In_1167,In_493);
nor U107 (N_107,In_1770,In_1681);
and U108 (N_108,In_2742,In_1741);
nand U109 (N_109,In_451,In_478);
nor U110 (N_110,In_229,In_105);
or U111 (N_111,In_2981,In_1605);
nor U112 (N_112,In_2370,In_1422);
nand U113 (N_113,In_942,In_1334);
nand U114 (N_114,In_331,In_1322);
xor U115 (N_115,In_1974,In_2139);
and U116 (N_116,In_2036,In_2033);
nand U117 (N_117,In_469,In_2455);
nand U118 (N_118,In_2795,In_907);
nand U119 (N_119,In_169,In_1944);
or U120 (N_120,In_2771,In_578);
nand U121 (N_121,In_2171,In_1552);
or U122 (N_122,In_426,In_551);
and U123 (N_123,In_1380,In_2920);
nand U124 (N_124,In_335,In_1168);
or U125 (N_125,In_2165,In_2194);
and U126 (N_126,In_2617,In_1713);
nand U127 (N_127,In_787,In_572);
nor U128 (N_128,In_1248,In_2535);
and U129 (N_129,In_1699,In_1379);
and U130 (N_130,In_1233,In_1451);
nand U131 (N_131,In_2529,In_1544);
or U132 (N_132,In_2441,In_2915);
nor U133 (N_133,In_760,In_1061);
xor U134 (N_134,In_2753,In_1789);
or U135 (N_135,In_2869,In_1060);
and U136 (N_136,In_337,In_240);
nor U137 (N_137,In_1079,In_2276);
nand U138 (N_138,In_1698,In_26);
xnor U139 (N_139,In_152,In_318);
or U140 (N_140,In_1956,In_2862);
and U141 (N_141,In_255,In_766);
nand U142 (N_142,In_2854,In_977);
nor U143 (N_143,In_2539,In_934);
nor U144 (N_144,In_2326,In_1984);
nand U145 (N_145,In_587,In_2615);
or U146 (N_146,In_153,In_1833);
or U147 (N_147,In_2973,In_1113);
nand U148 (N_148,In_167,In_2774);
xnor U149 (N_149,In_1164,In_1186);
nand U150 (N_150,In_455,In_2187);
and U151 (N_151,In_13,In_2384);
xor U152 (N_152,In_2666,In_2091);
xnor U153 (N_153,In_1766,In_1029);
nand U154 (N_154,In_279,In_1892);
nor U155 (N_155,In_73,In_974);
or U156 (N_156,In_2161,In_548);
nand U157 (N_157,In_1403,In_2813);
or U158 (N_158,In_2634,In_2279);
xnor U159 (N_159,In_1578,In_1449);
xor U160 (N_160,In_998,In_2385);
and U161 (N_161,In_1057,In_2982);
and U162 (N_162,In_938,In_2560);
or U163 (N_163,In_301,In_349);
nor U164 (N_164,In_2288,In_1495);
and U165 (N_165,In_489,In_1369);
nand U166 (N_166,In_889,In_2275);
nand U167 (N_167,In_730,In_2164);
or U168 (N_168,In_690,In_2782);
xor U169 (N_169,In_2308,In_502);
or U170 (N_170,In_1919,In_57);
xnor U171 (N_171,In_359,In_1091);
and U172 (N_172,In_1674,In_1313);
nor U173 (N_173,In_884,In_651);
or U174 (N_174,In_1913,In_2180);
nor U175 (N_175,In_912,In_2581);
nor U176 (N_176,In_2645,In_464);
xor U177 (N_177,In_1626,In_61);
nand U178 (N_178,In_2236,In_1388);
and U179 (N_179,In_563,In_2153);
nor U180 (N_180,In_996,In_1706);
and U181 (N_181,In_2328,In_1646);
or U182 (N_182,In_278,In_165);
and U183 (N_183,In_2301,In_32);
and U184 (N_184,In_1315,In_2258);
nor U185 (N_185,In_490,In_1243);
and U186 (N_186,In_1428,In_1344);
xor U187 (N_187,In_1721,In_1074);
xor U188 (N_188,In_1840,In_2494);
nor U189 (N_189,In_1607,In_2663);
and U190 (N_190,In_2054,In_807);
xnor U191 (N_191,In_2280,In_1328);
nor U192 (N_192,In_640,In_1360);
xnor U193 (N_193,In_505,In_2587);
and U194 (N_194,In_183,In_360);
and U195 (N_195,In_1105,In_580);
or U196 (N_196,In_1858,In_2642);
nor U197 (N_197,In_2439,In_2371);
nor U198 (N_198,In_1252,In_1547);
and U199 (N_199,In_2150,In_876);
nand U200 (N_200,In_647,In_2927);
nand U201 (N_201,In_2514,In_1875);
nor U202 (N_202,In_1719,In_1159);
nor U203 (N_203,In_532,In_1114);
xnor U204 (N_204,In_1485,In_2606);
xor U205 (N_205,In_865,In_2237);
nand U206 (N_206,In_1932,In_188);
nand U207 (N_207,In_2014,In_1943);
and U208 (N_208,In_957,In_2291);
or U209 (N_209,In_836,In_1385);
and U210 (N_210,In_1448,In_137);
nand U211 (N_211,In_2791,In_592);
nor U212 (N_212,In_2034,In_2743);
nand U213 (N_213,In_1968,In_1670);
or U214 (N_214,In_1465,In_1346);
xnor U215 (N_215,In_2250,In_2269);
and U216 (N_216,In_444,In_995);
xor U217 (N_217,In_2947,In_191);
and U218 (N_218,In_2671,In_2294);
xnor U219 (N_219,In_717,In_1280);
or U220 (N_220,In_1479,In_2541);
or U221 (N_221,In_2576,In_1430);
xor U222 (N_222,In_1249,In_2418);
nor U223 (N_223,In_2223,In_2284);
nand U224 (N_224,In_1250,In_1372);
nand U225 (N_225,In_115,In_702);
and U226 (N_226,In_768,In_1207);
or U227 (N_227,In_1008,In_2167);
xnor U228 (N_228,In_2787,In_1416);
and U229 (N_229,In_935,In_649);
nor U230 (N_230,In_852,In_298);
xor U231 (N_231,In_425,In_394);
nor U232 (N_232,In_721,In_2597);
and U233 (N_233,In_796,In_16);
or U234 (N_234,In_657,In_900);
nor U235 (N_235,In_2620,In_2550);
xor U236 (N_236,In_1046,In_1583);
and U237 (N_237,In_2528,In_1765);
nand U238 (N_238,In_878,In_2292);
or U239 (N_239,In_2346,In_2045);
nand U240 (N_240,In_1933,In_2404);
and U241 (N_241,In_2548,In_1763);
and U242 (N_242,In_628,In_575);
or U243 (N_243,In_1400,In_1361);
or U244 (N_244,In_2135,In_120);
nand U245 (N_245,In_1898,In_2354);
nand U246 (N_246,In_406,In_2719);
nor U247 (N_247,In_937,In_1879);
or U248 (N_248,In_557,In_1198);
and U249 (N_249,In_1539,In_1160);
xor U250 (N_250,In_2444,In_1631);
nand U251 (N_251,In_973,In_2971);
nor U252 (N_252,In_753,In_1266);
or U253 (N_253,In_1540,In_2883);
and U254 (N_254,In_1237,In_1777);
nor U255 (N_255,In_2565,In_2381);
xor U256 (N_256,In_1938,In_232);
nor U257 (N_257,In_1799,In_726);
and U258 (N_258,In_930,In_2695);
nand U259 (N_259,In_762,In_2059);
or U260 (N_260,In_1505,In_2056);
or U261 (N_261,In_2533,In_2919);
nand U262 (N_262,In_1817,In_824);
and U263 (N_263,In_577,In_1704);
or U264 (N_264,In_2248,In_1426);
nand U265 (N_265,In_686,In_509);
xnor U266 (N_266,In_2922,In_1503);
nor U267 (N_267,In_2797,In_761);
or U268 (N_268,In_864,In_564);
xnor U269 (N_269,In_1402,In_441);
xnor U270 (N_270,In_2380,In_988);
nor U271 (N_271,In_1573,In_1827);
xor U272 (N_272,In_2736,In_2249);
nor U273 (N_273,In_1953,In_1086);
nand U274 (N_274,In_2071,In_364);
nor U275 (N_275,In_47,In_1881);
or U276 (N_276,In_140,In_68);
nor U277 (N_277,In_888,In_2409);
and U278 (N_278,In_1924,In_2811);
nor U279 (N_279,In_519,In_2457);
xnor U280 (N_280,In_1125,In_1021);
nor U281 (N_281,In_499,In_841);
or U282 (N_282,In_334,In_1915);
xnor U283 (N_283,In_1204,In_24);
nand U284 (N_284,In_645,In_1131);
or U285 (N_285,In_2911,In_693);
nand U286 (N_286,In_2307,In_1696);
and U287 (N_287,In_2509,In_87);
xnor U288 (N_288,In_1731,In_2281);
xnor U289 (N_289,In_650,In_2618);
xor U290 (N_290,In_1183,In_2259);
nand U291 (N_291,In_1043,In_800);
or U292 (N_292,In_483,In_228);
nor U293 (N_293,In_1216,In_413);
or U294 (N_294,In_1464,In_1876);
xnor U295 (N_295,In_2599,In_2878);
nor U296 (N_296,In_1419,In_323);
nand U297 (N_297,In_2487,In_831);
and U298 (N_298,In_2423,In_1174);
or U299 (N_299,In_420,In_939);
xor U300 (N_300,In_2679,In_689);
or U301 (N_301,In_1302,In_748);
nand U302 (N_302,In_2109,In_859);
nand U303 (N_303,In_565,In_254);
and U304 (N_304,In_2076,In_2001);
and U305 (N_305,In_1439,In_1140);
or U306 (N_306,In_740,In_2375);
and U307 (N_307,In_504,In_1175);
nor U308 (N_308,In_387,In_194);
xnor U309 (N_309,In_843,In_2230);
or U310 (N_310,In_466,In_193);
and U311 (N_311,In_2020,In_615);
nand U312 (N_312,In_211,In_2543);
and U313 (N_313,In_2362,In_2704);
or U314 (N_314,In_2092,In_861);
and U315 (N_315,In_2516,In_6);
and U316 (N_316,In_928,In_2029);
xor U317 (N_317,In_1054,In_2894);
and U318 (N_318,In_936,In_952);
xnor U319 (N_319,In_2298,In_1900);
or U320 (N_320,In_11,In_1025);
or U321 (N_321,In_2152,In_877);
nor U322 (N_322,In_513,In_1851);
nor U323 (N_323,In_749,In_2584);
nand U324 (N_324,In_1893,In_2160);
xor U325 (N_325,In_1232,In_400);
or U326 (N_326,In_1507,In_1577);
and U327 (N_327,In_2425,In_236);
or U328 (N_328,In_2814,In_2340);
nor U329 (N_329,In_1429,In_1611);
nand U330 (N_330,In_1047,In_1729);
nand U331 (N_331,In_1685,In_173);
nand U332 (N_332,In_879,In_1032);
nor U333 (N_333,In_2500,In_2413);
or U334 (N_334,In_1,In_2473);
nor U335 (N_335,In_1071,In_2974);
nor U336 (N_336,In_785,In_386);
and U337 (N_337,In_8,In_1040);
nor U338 (N_338,In_1981,In_1812);
or U339 (N_339,In_555,In_2926);
and U340 (N_340,In_1628,In_1392);
or U341 (N_341,In_1512,In_2339);
or U342 (N_342,In_1959,In_904);
nand U343 (N_343,In_1620,In_1070);
or U344 (N_344,In_1614,In_821);
nor U345 (N_345,In_2579,In_1220);
and U346 (N_346,In_277,In_1431);
and U347 (N_347,In_1003,In_438);
xnor U348 (N_348,In_2283,In_2953);
nand U349 (N_349,In_1147,In_573);
xor U350 (N_350,In_1106,In_2011);
nor U351 (N_351,In_1309,In_2692);
or U352 (N_352,In_951,In_2834);
or U353 (N_353,In_2239,In_2873);
xor U354 (N_354,In_1045,In_2806);
nand U355 (N_355,In_1459,In_2257);
or U356 (N_356,In_2828,In_975);
or U357 (N_357,In_1148,In_1409);
xor U358 (N_358,In_1846,In_2235);
xnor U359 (N_359,In_529,In_742);
nor U360 (N_360,In_2469,In_1241);
nand U361 (N_361,In_1276,In_827);
xor U362 (N_362,In_2670,In_1324);
and U363 (N_363,In_1121,In_1571);
xnor U364 (N_364,In_2386,In_1410);
nor U365 (N_365,In_2388,In_2746);
xor U366 (N_366,In_2703,In_773);
nand U367 (N_367,In_1686,In_45);
nand U368 (N_368,In_468,In_189);
nand U369 (N_369,In_2923,In_2408);
and U370 (N_370,In_127,In_834);
and U371 (N_371,In_74,In_2286);
xor U372 (N_372,In_2038,In_1589);
nand U373 (N_373,In_82,In_1053);
and U374 (N_374,In_2976,In_160);
nor U375 (N_375,In_2735,In_823);
xnor U376 (N_376,In_798,In_956);
and U377 (N_377,In_1834,In_409);
and U378 (N_378,In_913,In_1299);
nor U379 (N_379,In_2016,In_1602);
xor U380 (N_380,In_245,In_1095);
xor U381 (N_381,In_2776,In_2426);
and U382 (N_382,In_2136,In_2783);
nand U383 (N_383,In_2318,In_2185);
nor U384 (N_384,In_1387,In_1829);
nand U385 (N_385,In_1935,In_813);
or U386 (N_386,In_1194,In_149);
xor U387 (N_387,In_620,In_1942);
and U388 (N_388,In_2306,In_2192);
nor U389 (N_389,In_52,In_2453);
and U390 (N_390,In_2740,In_1854);
nand U391 (N_391,In_2009,In_808);
nand U392 (N_392,In_1407,In_56);
xnor U393 (N_393,In_2954,In_1384);
nand U394 (N_394,In_948,In_867);
xnor U395 (N_395,In_2763,In_339);
nand U396 (N_396,In_97,In_2905);
nor U397 (N_397,In_804,In_2940);
and U398 (N_398,In_352,In_1764);
or U399 (N_399,In_2366,In_1285);
and U400 (N_400,In_1773,In_1373);
nand U401 (N_401,In_1691,In_1518);
xnor U402 (N_402,In_2637,In_2570);
nor U403 (N_403,In_2843,In_828);
or U404 (N_404,In_402,In_2062);
nor U405 (N_405,In_7,In_2519);
nor U406 (N_406,In_2598,In_1378);
or U407 (N_407,In_2534,In_1600);
and U408 (N_408,In_1287,In_2470);
nor U409 (N_409,In_1488,In_688);
nand U410 (N_410,In_1238,In_1447);
nor U411 (N_411,In_388,In_2737);
xnor U412 (N_412,In_2367,In_1155);
or U413 (N_413,In_2005,In_2522);
nor U414 (N_414,In_695,In_1511);
and U415 (N_415,In_1790,In_1170);
or U416 (N_416,In_2665,In_1267);
nor U417 (N_417,In_1754,In_537);
or U418 (N_418,In_849,In_2324);
nor U419 (N_419,In_1049,In_2983);
nand U420 (N_420,In_2093,In_1917);
xnor U421 (N_421,In_207,In_2510);
nand U422 (N_422,In_698,In_273);
xor U423 (N_423,In_1726,In_161);
or U424 (N_424,In_2147,In_491);
or U425 (N_425,In_763,In_1591);
nor U426 (N_426,In_1971,In_2415);
xor U427 (N_427,In_1093,In_424);
nor U428 (N_428,In_38,In_2043);
and U429 (N_429,In_2137,In_1668);
or U430 (N_430,In_2547,In_1217);
and U431 (N_431,In_1484,In_518);
nor U432 (N_432,In_2867,In_177);
and U433 (N_433,In_2962,In_1970);
nand U434 (N_434,In_2952,In_622);
nor U435 (N_435,In_2325,In_447);
nand U436 (N_436,In_126,In_1990);
nor U437 (N_437,In_2553,In_754);
xnor U438 (N_438,In_2901,In_283);
and U439 (N_439,In_909,In_723);
nand U440 (N_440,In_826,In_381);
nand U441 (N_441,In_1087,In_1277);
nand U442 (N_442,In_85,In_1270);
nand U443 (N_443,In_2348,In_674);
and U444 (N_444,In_1796,In_1742);
nand U445 (N_445,In_2488,In_1821);
nor U446 (N_446,In_579,In_2495);
nor U447 (N_447,In_2378,In_1520);
and U448 (N_448,In_134,In_80);
and U449 (N_449,In_1895,In_2098);
nand U450 (N_450,In_1076,In_2332);
nor U451 (N_451,In_405,In_131);
nand U452 (N_452,In_2461,In_560);
and U453 (N_453,In_2272,In_2177);
xnor U454 (N_454,In_1633,In_1531);
and U455 (N_455,In_1482,In_508);
xnor U456 (N_456,In_752,In_2698);
nand U457 (N_457,In_1251,In_990);
nor U458 (N_458,In_1794,In_736);
xnor U459 (N_459,In_543,In_554);
and U460 (N_460,In_317,In_1149);
nor U461 (N_461,In_60,In_1228);
xnor U462 (N_462,In_2158,In_1031);
or U463 (N_463,In_1650,In_2312);
or U464 (N_464,In_1782,In_1335);
nor U465 (N_465,In_212,In_2992);
nor U466 (N_466,In_2718,In_423);
nor U467 (N_467,In_1594,In_2585);
or U468 (N_468,In_515,In_1097);
nor U469 (N_469,In_2985,In_2405);
nor U470 (N_470,In_2891,In_2299);
or U471 (N_471,In_78,In_1213);
nand U472 (N_472,In_2662,In_65);
or U473 (N_473,In_2830,In_2086);
or U474 (N_474,In_2347,In_1154);
or U475 (N_475,In_2730,In_1985);
xnor U476 (N_476,In_588,In_1080);
nand U477 (N_477,In_2639,In_1024);
xor U478 (N_478,In_2655,In_1354);
and U479 (N_479,In_1470,In_1848);
xnor U480 (N_480,In_2356,In_2731);
or U481 (N_481,In_1100,In_2079);
xor U482 (N_482,In_1877,In_660);
nor U483 (N_483,In_1037,In_418);
nand U484 (N_484,In_2364,In_1949);
nand U485 (N_485,In_1208,In_811);
or U486 (N_486,In_964,In_2588);
or U487 (N_487,In_1934,In_1993);
xor U488 (N_488,In_1158,In_1362);
xnor U489 (N_489,In_408,In_114);
nand U490 (N_490,In_830,In_2892);
and U491 (N_491,In_157,In_1058);
nand U492 (N_492,In_1414,In_2577);
nand U493 (N_493,In_2857,In_2452);
and U494 (N_494,In_1929,In_2392);
or U495 (N_495,In_1513,In_2474);
nor U496 (N_496,In_138,In_1928);
and U497 (N_497,In_2603,In_1036);
and U498 (N_498,In_2688,In_2228);
nor U499 (N_499,In_1206,In_1542);
nor U500 (N_500,In_2246,In_1261);
or U501 (N_501,In_2849,In_1013);
nand U502 (N_502,In_1918,In_1077);
xnor U503 (N_503,In_583,In_2101);
xnor U504 (N_504,In_2499,In_549);
and U505 (N_505,In_210,In_2395);
xor U506 (N_506,In_1535,In_363);
nand U507 (N_507,In_2414,In_2496);
nand U508 (N_508,In_1242,In_1618);
and U509 (N_509,In_1475,In_2106);
nand U510 (N_510,In_1500,In_917);
and U511 (N_511,In_2842,In_397);
nand U512 (N_512,In_822,In_1941);
nor U513 (N_513,In_1826,In_2214);
and U514 (N_514,In_21,In_710);
or U515 (N_515,In_1240,In_2437);
or U516 (N_516,In_103,In_1418);
nor U517 (N_517,In_915,In_1708);
or U518 (N_518,In_49,In_1382);
xor U519 (N_519,In_119,In_372);
nor U520 (N_520,In_914,In_1824);
and U521 (N_521,In_2105,In_2026);
xor U522 (N_522,In_781,In_15);
or U523 (N_523,In_1964,In_42);
nand U524 (N_524,In_1016,In_163);
xnor U525 (N_525,In_1639,In_661);
or U526 (N_526,In_539,In_471);
nor U527 (N_527,In_214,In_2711);
or U528 (N_528,In_1693,In_1493);
nand U529 (N_529,In_2069,In_1785);
xor U530 (N_530,In_2734,In_1438);
nor U531 (N_531,In_2626,In_2066);
nor U532 (N_532,In_2296,In_527);
nand U533 (N_533,In_2376,In_2166);
nand U534 (N_534,In_2779,In_992);
nor U535 (N_535,In_2572,In_66);
or U536 (N_536,In_2573,In_1569);
and U537 (N_537,In_180,In_472);
or U538 (N_538,In_2142,In_500);
and U539 (N_539,In_2451,In_1136);
or U540 (N_540,In_1218,In_1397);
and U541 (N_541,In_924,In_2921);
and U542 (N_542,In_2571,In_1958);
nand U543 (N_543,In_2096,In_1596);
and U544 (N_544,In_2460,In_817);
and U545 (N_545,In_1492,In_1014);
xor U546 (N_546,In_393,In_223);
nand U547 (N_547,In_594,In_978);
xnor U548 (N_548,In_213,In_2868);
or U549 (N_549,In_2225,In_528);
or U550 (N_550,In_979,In_2506);
xnor U551 (N_551,In_863,In_2758);
xnor U552 (N_552,In_1712,In_2254);
or U553 (N_553,In_1481,In_1615);
or U554 (N_554,In_102,In_751);
or U555 (N_555,In_2916,In_1572);
nand U556 (N_556,In_1376,In_1509);
xor U557 (N_557,In_806,In_2068);
or U558 (N_558,In_2546,In_158);
and U559 (N_559,In_411,In_2908);
and U560 (N_560,In_416,In_737);
and U561 (N_561,In_2789,In_1978);
nand U562 (N_562,In_1343,In_2827);
nand U563 (N_563,In_1660,In_586);
nand U564 (N_564,In_1203,In_1568);
nor U565 (N_565,In_1735,In_641);
nand U566 (N_566,In_2697,In_1294);
or U567 (N_567,In_421,In_2118);
xnor U568 (N_568,In_2112,In_2330);
nand U569 (N_569,In_1371,In_2126);
xor U570 (N_570,In_1404,In_1176);
or U571 (N_571,In_1359,In_1722);
and U572 (N_572,In_2937,In_1102);
or U573 (N_573,In_1896,In_2723);
nand U574 (N_574,In_480,In_1275);
xor U575 (N_575,In_2213,In_2240);
nand U576 (N_576,In_2100,In_2417);
xor U577 (N_577,In_244,In_1560);
nand U578 (N_578,In_125,In_562);
or U579 (N_579,In_1316,In_890);
xnor U580 (N_580,In_1133,In_2262);
and U581 (N_581,In_1521,In_1115);
nand U582 (N_582,In_853,In_1101);
and U583 (N_583,In_1588,In_275);
nand U584 (N_584,In_415,In_692);
xor U585 (N_585,In_2807,In_270);
nand U586 (N_586,In_1586,In_2181);
nand U587 (N_587,In_282,In_609);
xnor U588 (N_588,In_2216,In_1188);
or U589 (N_589,In_705,In_2130);
or U590 (N_590,In_2661,In_187);
nor U591 (N_591,In_707,In_1916);
and U592 (N_592,In_1635,In_2933);
nor U593 (N_593,In_1453,In_2052);
or U594 (N_594,In_683,In_1026);
and U595 (N_595,In_2640,In_2304);
or U596 (N_596,In_171,In_154);
nand U597 (N_597,In_1471,In_1524);
nor U598 (N_598,In_1069,In_2683);
nor U599 (N_599,In_1966,In_1996);
nor U600 (N_600,In_1000,In_2566);
and U601 (N_601,In_199,In_607);
xnor U602 (N_602,In_475,In_2700);
nor U603 (N_603,In_1830,In_2712);
or U604 (N_604,In_2654,In_873);
or U605 (N_605,In_746,In_2872);
nor U606 (N_606,In_2319,In_1649);
nor U607 (N_607,In_2752,In_1127);
or U608 (N_608,In_1995,In_486);
and U609 (N_609,In_1271,In_2810);
xnor U610 (N_610,In_1697,In_307);
nor U611 (N_611,In_2604,In_448);
and U612 (N_612,In_2690,In_1555);
or U613 (N_613,In_1055,In_2608);
nor U614 (N_614,In_67,In_2321);
nor U615 (N_615,In_124,In_2950);
or U616 (N_616,In_1857,In_901);
nand U617 (N_617,In_994,In_2204);
or U618 (N_618,In_389,In_2087);
nand U619 (N_619,In_734,In_969);
xnor U620 (N_620,In_1957,In_604);
nor U621 (N_621,In_2607,In_963);
nand U622 (N_622,In_2880,In_959);
and U623 (N_623,In_2401,In_2003);
xnor U624 (N_624,In_911,In_2890);
or U625 (N_625,In_2335,In_2682);
or U626 (N_626,In_708,In_2959);
nand U627 (N_627,In_1469,In_1677);
nor U628 (N_628,In_308,In_2051);
or U629 (N_629,In_2845,In_1084);
xnor U630 (N_630,In_666,In_2412);
and U631 (N_631,In_2559,In_369);
or U632 (N_632,In_2442,In_1538);
nor U633 (N_633,In_2792,In_1580);
or U634 (N_634,In_1926,In_1135);
and U635 (N_635,In_1641,In_1202);
nor U636 (N_636,In_2140,In_2251);
and U637 (N_637,In_883,In_2208);
nor U638 (N_638,In_2707,In_1063);
xor U639 (N_639,In_2353,In_1843);
and U640 (N_640,In_2567,In_699);
nand U641 (N_641,In_835,In_2398);
nand U642 (N_642,In_2310,In_814);
nand U643 (N_643,In_224,In_2070);
or U644 (N_644,In_1235,In_2400);
or U645 (N_645,In_732,In_1321);
nor U646 (N_646,In_1011,In_1065);
nand U647 (N_647,In_2021,In_2800);
nor U648 (N_648,In_812,In_1342);
nor U649 (N_649,In_568,In_1556);
nand U650 (N_650,In_2032,In_1563);
or U651 (N_651,In_1643,In_2762);
or U652 (N_652,In_84,In_2635);
or U653 (N_653,In_584,In_2861);
nand U654 (N_654,In_2526,In_846);
and U655 (N_655,In_374,In_1911);
nand U656 (N_656,In_128,In_2515);
and U657 (N_657,In_894,In_2613);
xor U658 (N_658,In_2929,In_1050);
or U659 (N_659,In_1301,In_2936);
nor U660 (N_660,In_772,In_1749);
and U661 (N_661,In_989,In_2206);
xor U662 (N_662,In_1487,In_2231);
and U663 (N_663,In_531,In_1412);
or U664 (N_664,In_2438,In_933);
or U665 (N_665,In_2562,In_886);
or U666 (N_666,In_251,In_1654);
and U667 (N_667,In_1336,In_1473);
nand U668 (N_668,In_2313,In_1557);
nand U669 (N_669,In_1579,In_847);
nor U670 (N_670,In_242,In_655);
xor U671 (N_671,In_2636,In_932);
xnor U672 (N_672,In_1278,In_2479);
nand U673 (N_673,In_1405,In_243);
and U674 (N_674,In_1068,In_2058);
xnor U675 (N_675,In_59,In_2082);
nor U676 (N_676,In_625,In_2817);
xnor U677 (N_677,In_2583,In_2888);
nor U678 (N_678,In_1466,In_1806);
nor U679 (N_679,In_2102,In_2586);
and U680 (N_680,In_287,In_2050);
nor U681 (N_681,In_1421,In_2289);
nand U682 (N_682,In_442,In_1141);
or U683 (N_683,In_1659,In_1111);
nor U684 (N_684,In_178,In_2912);
nand U685 (N_685,In_81,In_2061);
xnor U686 (N_686,In_145,In_1679);
nor U687 (N_687,In_1886,In_98);
xnor U688 (N_688,In_2017,In_235);
nand U689 (N_689,In_1119,In_1440);
xor U690 (N_690,In_2593,In_810);
or U691 (N_691,In_570,In_582);
nand U692 (N_692,In_1089,In_1955);
xor U693 (N_693,In_305,In_832);
nand U694 (N_694,In_2876,In_2574);
nor U695 (N_695,In_2411,In_2575);
and U696 (N_696,In_1260,In_1525);
nand U697 (N_697,In_1502,In_727);
xor U698 (N_698,In_2266,In_2175);
xnor U699 (N_699,In_921,In_598);
and U700 (N_700,In_1399,In_1746);
nor U701 (N_701,In_2823,In_1355);
nor U702 (N_702,In_106,In_844);
or U703 (N_703,In_2788,In_1107);
xor U704 (N_704,In_2846,In_2747);
xnor U705 (N_705,In_2837,In_1720);
nand U706 (N_706,In_910,In_237);
nor U707 (N_707,In_2989,In_2172);
nor U708 (N_708,In_2420,In_501);
or U709 (N_709,In_875,In_1180);
and U710 (N_710,In_2490,In_770);
nor U711 (N_711,In_146,In_792);
and U712 (N_712,In_2938,In_276);
nor U713 (N_713,In_1802,In_2421);
nor U714 (N_714,In_2468,In_1640);
nor U715 (N_715,In_524,In_2975);
nand U716 (N_716,In_2373,In_1813);
or U717 (N_717,In_1437,In_2935);
or U718 (N_718,In_2115,In_2958);
and U719 (N_719,In_327,In_2893);
and U720 (N_720,In_2755,In_1744);
and U721 (N_721,In_2633,In_76);
xor U722 (N_722,In_263,In_1728);
and U723 (N_723,In_2949,In_943);
or U724 (N_724,In_2203,In_2178);
nor U725 (N_725,In_2416,In_432);
xor U726 (N_726,In_566,In_453);
nor U727 (N_727,In_2174,In_2551);
xnor U728 (N_728,In_1161,In_159);
nor U729 (N_729,In_1018,In_286);
nor U730 (N_730,In_997,In_487);
and U731 (N_731,In_1672,In_2088);
or U732 (N_732,In_2906,In_222);
xnor U733 (N_733,In_967,In_1368);
xor U734 (N_734,In_1733,In_1205);
xnor U735 (N_735,In_1536,In_1601);
xnor U736 (N_736,In_1855,In_2396);
xnor U737 (N_737,In_2724,In_1288);
xor U738 (N_738,In_664,In_46);
and U739 (N_739,In_23,In_2693);
xnor U740 (N_740,In_1856,In_1020);
nand U741 (N_741,In_2875,In_371);
and U742 (N_742,In_2803,In_1700);
or U743 (N_743,In_802,In_2903);
or U744 (N_744,In_9,In_2138);
and U745 (N_745,In_1396,In_1795);
nor U746 (N_746,In_1075,In_1364);
nand U747 (N_747,In_1117,In_1394);
nand U748 (N_748,In_488,In_496);
and U749 (N_749,In_340,In_1338);
and U750 (N_750,In_819,In_51);
nor U751 (N_751,In_2904,In_285);
xnor U752 (N_752,In_2991,In_48);
nor U753 (N_753,In_220,In_593);
nand U754 (N_754,In_1375,In_1022);
and U755 (N_755,In_2524,In_164);
xnor U756 (N_756,In_1406,In_1666);
xor U757 (N_757,In_320,In_1311);
and U758 (N_758,In_2095,In_440);
nor U759 (N_759,In_201,In_2812);
xor U760 (N_760,In_2899,In_1667);
xor U761 (N_761,In_1861,In_422);
and U762 (N_762,In_1226,In_1163);
nor U763 (N_763,In_2199,In_544);
nand U764 (N_764,In_2344,In_2311);
xor U765 (N_765,In_711,In_434);
and U766 (N_766,In_35,In_40);
nor U767 (N_767,In_3,In_2856);
nand U768 (N_768,In_1028,In_1907);
or U769 (N_769,In_1347,In_2219);
or U770 (N_770,In_2019,In_981);
nand U771 (N_771,In_1887,In_1566);
or U772 (N_772,In_2928,In_771);
and U773 (N_773,In_41,In_1033);
and U774 (N_774,In_1715,In_896);
nor U775 (N_775,In_791,In_1305);
or U776 (N_776,In_510,In_373);
xor U777 (N_777,In_2748,In_1644);
or U778 (N_778,In_2394,In_1108);
nor U779 (N_779,In_2841,In_1550);
nor U780 (N_780,In_2018,In_2467);
nand U781 (N_781,In_1190,In_1819);
nand U782 (N_782,In_1433,In_506);
nand U783 (N_783,In_109,In_93);
and U784 (N_784,In_1352,In_2063);
nor U785 (N_785,In_325,In_2083);
and U786 (N_786,In_2508,In_2123);
and U787 (N_787,In_2433,In_1947);
xnor U788 (N_788,In_215,In_1743);
xnor U789 (N_789,In_2309,In_2859);
nor U790 (N_790,In_2732,In_665);
nor U791 (N_791,In_71,In_477);
or U792 (N_792,In_29,In_1860);
and U793 (N_793,In_1663,In_1807);
nand U794 (N_794,In_482,In_2667);
nor U795 (N_795,In_2941,In_735);
or U796 (N_796,In_1081,In_1835);
and U797 (N_797,In_1797,In_147);
and U798 (N_798,In_2833,In_629);
and U799 (N_799,In_365,In_1329);
nand U800 (N_800,In_2333,In_2220);
and U801 (N_801,In_1863,In_99);
nand U802 (N_802,In_355,In_694);
or U803 (N_803,In_681,In_971);
xnor U804 (N_804,In_1012,In_2839);
xor U805 (N_805,In_2860,In_1395);
and U806 (N_806,In_1587,In_2134);
xnor U807 (N_807,In_1529,In_2132);
nand U808 (N_808,In_2024,In_249);
or U809 (N_809,In_1462,In_2648);
nor U810 (N_810,In_2882,In_1688);
nor U811 (N_811,In_2041,In_292);
or U812 (N_812,In_1209,In_458);
nand U813 (N_813,In_2794,In_362);
nand U814 (N_814,In_2943,In_361);
nand U815 (N_815,In_1675,In_1909);
or U816 (N_816,In_1793,In_1212);
nand U817 (N_817,In_1816,In_1885);
or U818 (N_818,In_1386,In_1778);
and U819 (N_819,In_19,In_2832);
nor U820 (N_820,In_1630,In_310);
nand U821 (N_821,In_1468,In_682);
nor U822 (N_822,In_980,In_1989);
and U823 (N_823,In_1142,In_1178);
xor U824 (N_824,In_2659,In_1262);
nand U825 (N_825,In_2374,In_1078);
nor U826 (N_826,In_1828,In_2502);
xor U827 (N_827,In_2558,In_1908);
or U828 (N_828,In_676,In_112);
xor U829 (N_829,In_1230,In_1922);
nand U830 (N_830,In_1541,In_642);
nand U831 (N_831,In_1774,In_2557);
nand U832 (N_832,In_643,In_1954);
and U833 (N_833,In_618,In_1201);
nor U834 (N_834,In_53,In_750);
or U835 (N_835,In_176,In_718);
or U836 (N_836,In_2767,In_1357);
or U837 (N_837,In_1268,In_987);
nor U838 (N_838,In_2532,In_2610);
and U839 (N_839,In_241,In_2612);
or U840 (N_840,In_403,In_2628);
and U841 (N_841,In_2031,In_2363);
xnor U842 (N_842,In_1224,In_116);
or U843 (N_843,In_522,In_2580);
and U844 (N_844,In_820,In_780);
and U845 (N_845,In_454,In_922);
xor U846 (N_846,In_536,In_635);
or U847 (N_847,In_958,In_2360);
xnor U848 (N_848,In_2342,In_1349);
nor U849 (N_849,In_1651,In_1510);
nand U850 (N_850,In_1332,In_2007);
and U851 (N_851,In_925,In_1581);
nor U852 (N_852,In_1831,In_414);
nand U853 (N_853,In_1562,In_196);
nor U854 (N_854,In_1776,In_816);
nor U855 (N_855,In_2836,In_2672);
nor U856 (N_856,In_2699,In_142);
xnor U857 (N_857,In_264,In_1798);
nand U858 (N_858,In_1300,In_837);
nand U859 (N_859,In_633,In_691);
or U860 (N_860,In_1002,In_1156);
nand U861 (N_861,In_2255,In_1991);
nand U862 (N_862,In_1980,In_306);
xnor U863 (N_863,In_2410,In_328);
or U864 (N_864,In_2631,In_2497);
and U865 (N_865,In_670,In_517);
or U866 (N_866,In_1312,In_654);
or U867 (N_867,In_1737,In_1897);
nor U868 (N_868,In_268,In_976);
xor U869 (N_869,In_297,In_1424);
and U870 (N_870,In_1665,In_2852);
nand U871 (N_871,In_2334,In_36);
or U872 (N_872,In_2701,In_893);
nor U873 (N_873,In_2544,In_2902);
nand U874 (N_874,In_2676,In_1637);
nor U875 (N_875,In_1593,In_1374);
and U876 (N_876,In_1129,In_382);
nor U877 (N_877,In_2650,In_2170);
nand U878 (N_878,In_1109,In_2749);
or U879 (N_879,In_2564,In_1199);
and U880 (N_880,In_733,In_696);
or U881 (N_881,In_1823,In_2039);
or U882 (N_882,In_1039,In_2047);
xnor U883 (N_883,In_1914,In_2715);
xor U884 (N_884,In_27,In_433);
or U885 (N_885,In_443,In_1221);
nor U886 (N_886,In_1609,In_284);
xor U887 (N_887,In_908,In_1690);
nand U888 (N_888,In_1804,In_302);
nand U889 (N_889,In_195,In_2530);
xor U890 (N_890,In_2361,In_2709);
nor U891 (N_891,In_1757,In_1227);
or U892 (N_892,In_687,In_2103);
or U893 (N_893,In_1222,In_858);
and U894 (N_894,In_95,In_1169);
xnor U895 (N_895,In_923,In_2207);
nor U896 (N_896,In_613,In_1005);
nand U897 (N_897,In_1786,In_2475);
xor U898 (N_898,In_2369,In_1717);
nand U899 (N_899,In_1514,In_2129);
nand U900 (N_900,In_2957,In_630);
or U901 (N_901,In_1627,In_1874);
or U902 (N_902,In_2622,In_2716);
nand U903 (N_903,In_1072,In_2790);
or U904 (N_904,In_1151,In_2939);
nand U905 (N_905,In_55,In_1705);
xnor U906 (N_906,In_1454,In_2706);
and U907 (N_907,In_2820,In_34);
or U908 (N_908,In_2089,In_77);
xnor U909 (N_909,In_571,In_12);
nand U910 (N_910,In_764,In_166);
and U911 (N_911,In_208,In_100);
xor U912 (N_912,In_2871,In_2464);
nor U913 (N_913,In_1181,In_1508);
or U914 (N_914,In_1490,In_1653);
nand U915 (N_915,In_2431,In_2511);
nand U916 (N_916,In_136,In_2297);
nor U917 (N_917,In_2270,In_759);
nor U918 (N_918,In_1727,In_833);
nand U919 (N_919,In_874,In_460);
and U920 (N_920,In_1692,In_1565);
nor U921 (N_921,In_2993,In_2644);
or U922 (N_922,In_2478,In_1189);
xnor U923 (N_923,In_1413,In_931);
nand U924 (N_924,In_1341,In_1567);
nand U925 (N_925,In_2256,In_715);
and U926 (N_926,In_107,In_398);
nor U927 (N_927,In_1732,In_1951);
xnor U928 (N_928,In_2247,In_2517);
xnor U929 (N_929,In_2930,In_970);
and U930 (N_930,In_961,In_2472);
or U931 (N_931,In_1987,In_43);
and U932 (N_932,In_669,In_1110);
nand U933 (N_933,In_2424,In_39);
nand U934 (N_934,In_75,In_567);
nand U935 (N_935,In_150,In_1682);
xnor U936 (N_936,In_1165,In_2729);
nor U937 (N_937,In_982,In_174);
or U938 (N_938,In_2146,In_1767);
nor U939 (N_939,In_2594,In_680);
or U940 (N_940,In_1195,In_2447);
and U941 (N_941,In_1062,In_1425);
xnor U942 (N_942,In_1636,In_2717);
or U943 (N_943,In_2602,In_774);
xor U944 (N_944,In_712,In_428);
and U945 (N_945,In_2995,In_829);
and U946 (N_946,In_1570,In_1678);
or U947 (N_947,In_2960,In_2267);
and U948 (N_948,In_1755,In_767);
and U949 (N_949,In_1884,In_2012);
or U950 (N_950,In_1761,In_2065);
nand U951 (N_951,In_1963,In_2741);
nor U952 (N_952,In_2121,In_1491);
and U953 (N_953,In_795,In_765);
and U954 (N_954,In_2946,In_882);
nor U955 (N_955,In_673,In_185);
nand U956 (N_956,In_1246,In_1652);
and U957 (N_957,In_2162,In_1962);
xnor U958 (N_958,In_2826,In_2990);
or U959 (N_959,In_2601,In_2554);
nand U960 (N_960,In_818,In_2435);
xor U961 (N_961,In_2972,In_887);
and U962 (N_962,In_706,In_1839);
and U963 (N_963,In_2691,In_1269);
nor U964 (N_964,In_2463,In_2786);
and U965 (N_965,In_1498,In_1655);
or U966 (N_966,In_2197,In_474);
nor U967 (N_967,In_1598,In_2141);
xor U968 (N_968,In_350,In_722);
nor U969 (N_969,In_857,In_784);
and U970 (N_970,In_30,In_1187);
nor U971 (N_971,In_1657,In_1617);
or U972 (N_972,In_1792,In_1007);
nor U973 (N_973,In_1948,In_2205);
and U974 (N_974,In_139,In_1501);
xnor U975 (N_975,In_2955,In_2799);
or U976 (N_976,In_815,In_253);
xor U977 (N_977,In_2864,In_2996);
nor U978 (N_978,In_610,In_2393);
xnor U979 (N_979,In_1092,In_716);
nor U980 (N_980,In_2855,In_983);
nand U981 (N_981,In_1780,In_2874);
nand U982 (N_982,In_396,In_1103);
nor U983 (N_983,In_652,In_351);
nor U984 (N_984,In_2229,In_2647);
nand U985 (N_985,In_1869,In_2483);
nand U986 (N_986,In_1825,In_2840);
nand U987 (N_987,In_891,In_1621);
nand U988 (N_988,In_1282,In_535);
xnor U989 (N_989,In_966,In_1263);
or U990 (N_990,In_90,In_1184);
xnor U991 (N_991,In_1606,In_1295);
nand U992 (N_992,In_2004,In_58);
nor U993 (N_993,In_463,In_2084);
nor U994 (N_994,In_946,In_2127);
nand U995 (N_995,In_597,In_953);
nand U996 (N_996,In_345,In_2320);
xnor U997 (N_997,In_558,In_2831);
and U998 (N_998,In_2,In_2844);
or U999 (N_999,In_1290,In_1890);
nand U1000 (N_1000,In_1023,In_258);
nor U1001 (N_1001,In_2209,In_2804);
nand U1002 (N_1002,In_230,In_541);
xor U1003 (N_1003,In_2450,In_206);
nor U1004 (N_1004,In_1116,In_86);
nor U1005 (N_1005,In_1576,In_659);
nand U1006 (N_1006,In_2200,In_569);
nand U1007 (N_1007,In_2627,In_1803);
nor U1008 (N_1008,In_2777,In_1356);
or U1009 (N_1009,In_2080,In_1822);
and U1010 (N_1010,In_18,In_2624);
nand U1011 (N_1011,In_288,In_1865);
or U1012 (N_1012,In_906,In_356);
nor U1013 (N_1013,In_376,In_294);
nor U1014 (N_1014,In_2397,In_1937);
nor U1015 (N_1015,In_954,In_1458);
xnor U1016 (N_1016,In_333,In_1730);
nor U1017 (N_1017,In_1196,In_135);
nand U1018 (N_1018,In_1946,In_179);
or U1019 (N_1019,In_2668,In_22);
or U1020 (N_1020,In_1134,In_2186);
nor U1021 (N_1021,In_354,In_1923);
or U1022 (N_1022,In_175,In_2678);
nand U1023 (N_1023,In_658,In_368);
nor U1024 (N_1024,In_1320,In_2365);
or U1025 (N_1025,In_412,In_2674);
nor U1026 (N_1026,In_133,In_2714);
and U1027 (N_1027,In_481,In_2090);
xnor U1028 (N_1028,In_1197,In_1351);
xnor U1029 (N_1029,In_1748,In_2035);
or U1030 (N_1030,In_521,In_221);
nor U1031 (N_1031,In_542,In_2000);
nor U1032 (N_1032,In_1866,In_1850);
nor U1033 (N_1033,In_2537,In_1483);
nand U1034 (N_1034,In_540,In_697);
or U1035 (N_1035,In_1530,In_2030);
and U1036 (N_1036,In_1853,In_430);
and U1037 (N_1037,In_202,In_2924);
xor U1038 (N_1038,In_2801,In_1714);
or U1039 (N_1039,In_2163,In_182);
nor U1040 (N_1040,In_1445,In_639);
nand U1041 (N_1041,In_1709,In_231);
xnor U1042 (N_1042,In_1658,In_2427);
nand U1043 (N_1043,In_2656,In_37);
or U1044 (N_1044,In_1138,In_2925);
and U1045 (N_1045,In_2149,In_2851);
nor U1046 (N_1046,In_1515,In_2781);
nand U1047 (N_1047,In_601,In_132);
xnor U1048 (N_1048,In_25,In_2798);
nand U1049 (N_1049,In_871,In_743);
xnor U1050 (N_1050,In_631,In_111);
xor U1051 (N_1051,In_547,In_2590);
or U1052 (N_1052,In_2057,In_2866);
xnor U1053 (N_1053,In_1998,In_2595);
and U1054 (N_1054,In_1899,In_1599);
xor U1055 (N_1055,In_2198,In_2917);
or U1056 (N_1056,In_2436,In_1972);
or U1057 (N_1057,In_2113,In_1389);
or U1058 (N_1058,In_390,In_1401);
or U1059 (N_1059,In_2848,In_2252);
nor U1060 (N_1060,In_450,In_2895);
and U1061 (N_1061,In_296,In_2122);
and U1062 (N_1062,In_789,In_2600);
nor U1063 (N_1063,In_2210,In_367);
or U1064 (N_1064,In_614,In_2815);
nand U1065 (N_1065,In_1339,In_239);
xor U1066 (N_1066,In_1391,In_991);
or U1067 (N_1067,In_2780,In_2233);
and U1068 (N_1068,In_2476,In_2944);
or U1069 (N_1069,In_2702,In_1809);
xnor U1070 (N_1070,In_2784,In_1532);
nor U1071 (N_1071,In_1738,In_1936);
nor U1072 (N_1072,In_520,In_2073);
nand U1073 (N_1073,In_1096,In_1130);
xor U1074 (N_1074,In_2064,In_2358);
nand U1075 (N_1075,In_156,In_870);
nor U1076 (N_1076,In_2705,In_2006);
or U1077 (N_1077,In_2458,In_512);
nor U1078 (N_1078,In_2552,In_2316);
nand U1079 (N_1079,In_1906,In_407);
or U1080 (N_1080,In_1340,In_1772);
nor U1081 (N_1081,In_1185,In_1323);
and U1082 (N_1082,In_671,In_940);
nand U1083 (N_1083,In_2967,In_776);
and U1084 (N_1084,In_1927,In_494);
and U1085 (N_1085,In_1842,In_2406);
or U1086 (N_1086,In_1867,In_1891);
xor U1087 (N_1087,In_344,In_663);
or U1088 (N_1088,In_2368,In_129);
and U1089 (N_1089,In_2884,In_2445);
and U1090 (N_1090,In_2159,In_2055);
nor U1091 (N_1091,In_1783,In_383);
nand U1092 (N_1092,In_2226,In_1358);
or U1093 (N_1093,In_1085,In_31);
or U1094 (N_1094,In_2195,In_2858);
nand U1095 (N_1095,In_2687,In_1258);
xor U1096 (N_1096,In_2751,In_2621);
or U1097 (N_1097,In_452,In_1592);
nand U1098 (N_1098,In_1740,In_662);
xor U1099 (N_1099,In_217,In_2684);
nor U1100 (N_1100,In_851,In_1363);
nor U1101 (N_1101,In_1779,In_1656);
nand U1102 (N_1102,In_2201,In_2816);
or U1103 (N_1103,In_260,In_1318);
nand U1104 (N_1104,In_2144,In_1610);
nand U1105 (N_1105,In_2945,In_2793);
nand U1106 (N_1106,In_2462,In_2120);
nand U1107 (N_1107,In_1223,In_2824);
and U1108 (N_1108,In_1952,In_731);
and U1109 (N_1109,In_1004,In_2507);
xor U1110 (N_1110,In_719,In_130);
and U1111 (N_1111,In_2486,In_1517);
xor U1112 (N_1112,In_1010,In_850);
and U1113 (N_1113,In_897,In_2986);
or U1114 (N_1114,In_648,In_1903);
and U1115 (N_1115,In_1811,In_1982);
and U1116 (N_1116,In_2503,In_370);
and U1117 (N_1117,In_2504,In_2193);
or U1118 (N_1118,In_1847,In_2341);
nor U1119 (N_1119,In_1420,In_319);
and U1120 (N_1120,In_271,In_2287);
and U1121 (N_1121,In_2726,In_955);
and U1122 (N_1122,In_2377,In_2619);
and U1123 (N_1123,In_2887,In_246);
nor U1124 (N_1124,In_1120,In_265);
and U1125 (N_1125,In_2910,In_155);
xor U1126 (N_1126,In_703,In_905);
or U1127 (N_1127,In_5,In_121);
and U1128 (N_1128,In_2563,In_2074);
xnor U1129 (N_1129,In_2261,In_1034);
nand U1130 (N_1130,In_2531,In_1398);
nand U1131 (N_1131,In_1752,In_1177);
and U1132 (N_1132,In_2253,In_556);
xnor U1133 (N_1133,In_1836,In_793);
and U1134 (N_1134,In_1791,In_2658);
or U1135 (N_1135,In_1808,In_1009);
nand U1136 (N_1136,In_1463,In_2768);
nand U1137 (N_1137,In_1253,In_326);
nor U1138 (N_1138,In_1128,In_1367);
nor U1139 (N_1139,In_2616,In_2015);
or U1140 (N_1140,In_1872,In_2942);
or U1141 (N_1141,In_2302,In_2263);
and U1142 (N_1142,In_2075,In_1945);
nor U1143 (N_1143,In_2721,In_842);
nor U1144 (N_1144,In_2434,In_2215);
or U1145 (N_1145,In_2931,In_623);
and U1146 (N_1146,In_1381,In_2111);
nor U1147 (N_1147,In_358,In_1331);
nand U1148 (N_1148,In_2419,In_1265);
and U1149 (N_1149,In_2900,In_1664);
and U1150 (N_1150,In_550,In_110);
nor U1151 (N_1151,In_1612,In_1126);
or U1152 (N_1152,In_595,In_2964);
nand U1153 (N_1153,In_2760,In_2998);
nand U1154 (N_1154,In_790,In_291);
and U1155 (N_1155,In_1489,In_1684);
nand U1156 (N_1156,In_2591,In_856);
or U1157 (N_1157,In_2399,In_250);
or U1158 (N_1158,In_848,In_2168);
xor U1159 (N_1159,In_1124,In_1478);
and U1160 (N_1160,In_2343,In_638);
or U1161 (N_1161,In_720,In_2493);
nand U1162 (N_1162,In_2745,In_2673);
nand U1163 (N_1163,In_1038,In_399);
and U1164 (N_1164,In_1474,In_1516);
and U1165 (N_1165,In_1247,In_2331);
nand U1166 (N_1166,In_920,In_2629);
nand U1167 (N_1167,In_1064,In_2853);
nand U1168 (N_1168,In_1756,In_1083);
nand U1169 (N_1169,In_2664,In_17);
and U1170 (N_1170,In_2501,In_2322);
nand U1171 (N_1171,In_1452,In_2907);
or U1172 (N_1172,In_782,In_2934);
xor U1173 (N_1173,In_2605,In_2630);
nand U1174 (N_1174,In_2838,In_1969);
xnor U1175 (N_1175,In_1545,In_1153);
or U1176 (N_1176,In_1642,In_1528);
xnor U1177 (N_1177,In_92,In_709);
or U1178 (N_1178,In_2403,In_1582);
and U1179 (N_1179,In_1553,In_1781);
and U1180 (N_1180,In_395,In_2865);
and U1181 (N_1181,In_1775,In_20);
nand U1182 (N_1182,In_162,In_2885);
and U1183 (N_1183,In_1537,In_1976);
nor U1184 (N_1184,In_2429,In_576);
or U1185 (N_1185,In_533,In_738);
and U1186 (N_1186,In_2124,In_2809);
or U1187 (N_1187,In_2632,In_1676);
xor U1188 (N_1188,In_2350,In_2273);
and U1189 (N_1189,In_758,In_704);
or U1190 (N_1190,In_1986,In_2796);
and U1191 (N_1191,In_585,In_574);
nand U1192 (N_1192,In_1805,In_2881);
nand U1193 (N_1193,In_949,In_1522);
nand U1194 (N_1194,In_2897,In_678);
or U1195 (N_1195,In_605,In_2107);
or U1196 (N_1196,In_1455,In_1456);
xnor U1197 (N_1197,In_1901,In_1880);
or U1198 (N_1198,In_2449,In_794);
xnor U1199 (N_1199,In_2067,In_2739);
nand U1200 (N_1200,In_744,In_261);
nand U1201 (N_1201,In_2757,In_596);
or U1202 (N_1202,In_756,In_1304);
xnor U1203 (N_1203,In_203,In_769);
nor U1204 (N_1204,In_1052,In_626);
and U1205 (N_1205,In_2918,In_962);
nand U1206 (N_1206,In_1292,In_2963);
nand U1207 (N_1207,In_485,In_872);
or U1208 (N_1208,In_993,In_2217);
nand U1209 (N_1209,In_1122,In_2492);
nor U1210 (N_1210,In_170,In_300);
or U1211 (N_1211,In_2969,In_1308);
xnor U1212 (N_1212,In_2446,In_1801);
and U1213 (N_1213,In_1734,In_2027);
xor U1214 (N_1214,In_1661,In_2440);
nand U1215 (N_1215,In_2521,In_2681);
nand U1216 (N_1216,In_589,In_1931);
xnor U1217 (N_1217,In_1669,In_2402);
or U1218 (N_1218,In_1298,In_2686);
nand U1219 (N_1219,In_2355,In_1725);
and U1220 (N_1220,In_314,In_1042);
or U1221 (N_1221,In_280,In_862);
and U1222 (N_1222,In_1526,In_2241);
xor U1223 (N_1223,In_2196,In_1254);
and U1224 (N_1224,In_1724,In_1067);
xnor U1225 (N_1225,In_216,In_184);
xnor U1226 (N_1226,In_54,In_1245);
nand U1227 (N_1227,In_435,In_2527);
xor U1228 (N_1228,In_1098,In_1137);
nand U1229 (N_1229,In_2224,In_1622);
nor U1230 (N_1230,In_1472,In_2710);
nand U1231 (N_1231,In_316,In_1859);
nor U1232 (N_1232,In_2913,In_366);
xor U1233 (N_1233,In_1608,In_1784);
nor U1234 (N_1234,In_559,In_1868);
xnor U1235 (N_1235,In_2970,In_2116);
nor U1236 (N_1236,In_1939,In_1291);
nand U1237 (N_1237,In_1435,In_840);
xor U1238 (N_1238,In_63,In_1930);
nand U1239 (N_1239,In_88,In_1307);
nor U1240 (N_1240,In_1619,In_321);
or U1241 (N_1241,In_2491,In_1051);
nor U1242 (N_1242,In_2202,In_701);
and U1243 (N_1243,In_1574,In_2265);
nand U1244 (N_1244,In_1604,In_2212);
or U1245 (N_1245,In_272,In_1019);
xnor U1246 (N_1246,In_197,In_1297);
nand U1247 (N_1247,In_755,In_2728);
nor U1248 (N_1248,In_1992,In_1736);
nor U1249 (N_1249,In_2525,In_2769);
nand U1250 (N_1250,In_2657,In_1035);
xor U1251 (N_1251,In_2948,In_1317);
and U1252 (N_1252,In_1888,In_612);
and U1253 (N_1253,In_281,In_2407);
xnor U1254 (N_1254,In_28,In_2896);
or U1255 (N_1255,In_2482,In_2708);
xor U1256 (N_1256,In_1112,In_2456);
xnor U1257 (N_1257,In_2542,In_401);
and U1258 (N_1258,In_2245,In_1145);
xor U1259 (N_1259,In_1325,In_1638);
nor U1260 (N_1260,In_1841,In_2303);
and U1261 (N_1261,In_1314,In_880);
and U1262 (N_1262,In_2466,In_2010);
or U1263 (N_1263,In_473,In_2271);
nand U1264 (N_1264,In_1467,In_903);
nand U1265 (N_1265,In_303,In_234);
nand U1266 (N_1266,In_2785,In_1143);
and U1267 (N_1267,In_1852,In_2023);
and U1268 (N_1268,In_439,In_1215);
or U1269 (N_1269,In_677,In_1585);
xor U1270 (N_1270,In_636,In_2870);
and U1271 (N_1271,In_431,In_2060);
nand U1272 (N_1272,In_653,In_2643);
xnor U1273 (N_1273,In_1788,In_2978);
and U1274 (N_1274,In_2008,In_2260);
and U1275 (N_1275,In_1166,In_2727);
or U1276 (N_1276,In_248,In_1838);
and U1277 (N_1277,In_322,In_2625);
xnor U1278 (N_1278,In_1200,In_1006);
nor U1279 (N_1279,In_2072,In_2040);
and U1280 (N_1280,In_624,In_89);
xnor U1281 (N_1281,In_101,In_2117);
xnor U1282 (N_1282,In_1179,In_902);
and U1283 (N_1283,In_429,In_2609);
xor U1284 (N_1284,In_2555,In_1330);
nand U1285 (N_1285,In_1920,In_2489);
and U1286 (N_1286,In_1519,In_1192);
nand U1287 (N_1287,In_511,In_1088);
and U1288 (N_1288,In_2802,In_2818);
nand U1289 (N_1289,In_219,In_1965);
nand U1290 (N_1290,In_2432,In_1436);
xnor U1291 (N_1291,In_1162,In_545);
nor U1292 (N_1292,In_2336,In_1648);
or U1293 (N_1293,In_1239,In_141);
nand U1294 (N_1294,In_603,In_1739);
nor U1295 (N_1295,In_1066,In_1689);
nand U1296 (N_1296,In_1319,In_1815);
or U1297 (N_1297,In_714,In_855);
and U1298 (N_1298,In_1480,In_2268);
or U1299 (N_1299,In_728,In_602);
nand U1300 (N_1300,In_2754,In_204);
or U1301 (N_1301,In_1695,In_2518);
nor U1302 (N_1302,In_534,In_1862);
and U1303 (N_1303,In_1293,In_656);
and U1304 (N_1304,In_2545,In_33);
or U1305 (N_1305,In_2184,In_941);
xor U1306 (N_1306,In_1082,In_470);
xor U1307 (N_1307,In_2182,In_2293);
nand U1308 (N_1308,In_1283,In_1015);
or U1309 (N_1309,In_1973,In_1476);
and U1310 (N_1310,In_2465,In_2611);
or U1311 (N_1311,In_1348,In_1256);
or U1312 (N_1312,In_1173,In_1383);
and U1313 (N_1313,In_456,In_2932);
xnor U1314 (N_1314,In_1506,In_1533);
xor U1315 (N_1315,In_2819,In_1048);
nand U1316 (N_1316,In_2077,In_1960);
and U1317 (N_1317,In_256,In_1753);
or U1318 (N_1318,In_94,In_2154);
nor U1319 (N_1319,In_2725,In_2536);
nor U1320 (N_1320,In_1001,In_144);
nor U1321 (N_1321,In_729,In_2454);
or U1322 (N_1322,In_1144,In_1244);
xor U1323 (N_1323,In_2448,In_1284);
xnor U1324 (N_1324,In_1279,In_2190);
and U1325 (N_1325,In_1616,In_667);
and U1326 (N_1326,In_805,In_2677);
nor U1327 (N_1327,In_1191,In_2961);
or U1328 (N_1328,In_2145,In_299);
nor U1329 (N_1329,In_2713,In_198);
nand U1330 (N_1330,In_553,In_1597);
nor U1331 (N_1331,In_1910,In_2048);
nor U1332 (N_1332,In_1814,In_2651);
xnor U1333 (N_1333,In_2898,In_621);
or U1334 (N_1334,In_1845,In_1434);
nand U1335 (N_1335,In_507,In_1575);
xnor U1336 (N_1336,In_200,In_1182);
nand U1337 (N_1337,In_2108,In_1559);
and U1338 (N_1338,In_1044,In_2773);
nor U1339 (N_1339,In_2391,In_1551);
and U1340 (N_1340,In_2561,In_2323);
xnor U1341 (N_1341,In_672,In_346);
xor U1342 (N_1342,In_2956,In_495);
nor U1343 (N_1343,In_2568,In_50);
or U1344 (N_1344,In_2382,In_2485);
nor U1345 (N_1345,In_797,In_2889);
xnor U1346 (N_1346,In_1820,In_1625);
nor U1347 (N_1347,In_329,In_449);
xnor U1348 (N_1348,In_1281,In_467);
xnor U1349 (N_1349,In_1446,In_1527);
xor U1350 (N_1350,In_378,In_581);
nor U1351 (N_1351,In_122,In_2359);
nor U1352 (N_1352,In_1225,In_2243);
and U1353 (N_1353,In_2994,In_1289);
or U1354 (N_1354,In_1150,In_205);
nor U1355 (N_1355,In_895,In_1255);
nand U1356 (N_1356,In_2022,In_1411);
nand U1357 (N_1357,In_538,In_1296);
and U1358 (N_1358,In_96,In_2951);
and U1359 (N_1359,In_348,In_1662);
nand U1360 (N_1360,In_2169,In_384);
nor U1361 (N_1361,In_2997,In_2234);
nand U1362 (N_1362,In_2675,In_2242);
nor U1363 (N_1363,In_1264,In_1234);
xor U1364 (N_1364,In_330,In_898);
and U1365 (N_1365,In_1558,In_2733);
or U1366 (N_1366,In_266,In_561);
nor U1367 (N_1367,In_2128,In_1229);
nand U1368 (N_1368,In_2966,In_1461);
xor U1369 (N_1369,In_1902,In_2987);
nand U1370 (N_1370,In_2614,In_70);
or U1371 (N_1371,In_1353,In_123);
and U1372 (N_1372,In_2863,In_72);
or U1373 (N_1373,In_1595,In_79);
xnor U1374 (N_1374,In_380,In_968);
nor U1375 (N_1375,In_1603,In_479);
nor U1376 (N_1376,In_1450,In_1940);
xnor U1377 (N_1377,In_1273,In_2049);
nor U1378 (N_1378,In_290,In_2300);
nand U1379 (N_1379,In_947,In_238);
or U1380 (N_1380,In_2770,In_2914);
xor U1381 (N_1381,In_1864,In_457);
or U1382 (N_1382,In_247,In_311);
or U1383 (N_1383,In_608,In_1871);
nand U1384 (N_1384,In_1441,In_226);
and U1385 (N_1385,In_2046,In_2314);
or U1386 (N_1386,In_2044,In_436);
or U1387 (N_1387,In_2097,In_2352);
nor U1388 (N_1388,In_2778,In_1810);
nor U1389 (N_1389,In_2148,In_944);
or U1390 (N_1390,In_1687,In_739);
nand U1391 (N_1391,In_498,In_526);
and U1392 (N_1392,In_2689,In_779);
and U1393 (N_1393,In_2977,In_1703);
nand U1394 (N_1394,In_2750,In_1486);
nor U1395 (N_1395,In_514,In_1415);
nor U1396 (N_1396,In_546,In_1745);
or U1397 (N_1397,In_0,In_838);
xor U1398 (N_1398,In_476,In_315);
or U1399 (N_1399,In_343,In_679);
and U1400 (N_1400,In_1723,In_1549);
xnor U1401 (N_1401,In_1883,In_357);
xor U1402 (N_1402,In_2669,In_1961);
nand U1403 (N_1403,In_619,In_777);
or U1404 (N_1404,In_2582,In_2596);
xor U1405 (N_1405,In_1427,In_2264);
or U1406 (N_1406,In_2660,In_2143);
or U1407 (N_1407,In_1921,In_2238);
and U1408 (N_1408,In_1994,In_2653);
xor U1409 (N_1409,In_2549,In_2430);
xnor U1410 (N_1410,In_267,In_2569);
or U1411 (N_1411,In_1457,In_606);
and U1412 (N_1412,In_336,In_799);
nor U1413 (N_1413,In_1629,In_616);
and U1414 (N_1414,In_1564,In_1632);
or U1415 (N_1415,In_2155,In_2968);
and U1416 (N_1416,In_646,In_1762);
and U1417 (N_1417,In_950,In_2505);
nor U1418 (N_1418,In_353,In_2179);
xnor U1419 (N_1419,In_1747,In_1878);
nor U1420 (N_1420,In_783,In_2498);
or U1421 (N_1421,In_2980,In_2850);
xnor U1422 (N_1422,In_1333,In_190);
nand U1423 (N_1423,In_1073,In_1882);
nor U1424 (N_1424,In_2765,In_1548);
or U1425 (N_1425,In_926,In_2808);
xnor U1426 (N_1426,In_309,In_1988);
nand U1427 (N_1427,In_825,In_2965);
xor U1428 (N_1428,In_1090,In_945);
nand U1429 (N_1429,In_1171,In_1423);
or U1430 (N_1430,In_552,In_1768);
xnor U1431 (N_1431,In_181,In_2188);
and U1432 (N_1432,In_2471,In_1769);
or U1433 (N_1433,In_104,In_1231);
and U1434 (N_1434,In_2696,In_2372);
or U1435 (N_1435,In_591,In_2652);
and U1436 (N_1436,In_83,In_1214);
nor U1437 (N_1437,In_2764,In_69);
and U1438 (N_1438,In_1157,In_2329);
nor U1439 (N_1439,In_1771,In_2338);
or U1440 (N_1440,In_1718,In_269);
and U1441 (N_1441,In_1056,In_437);
or U1442 (N_1442,In_392,In_2623);
or U1443 (N_1443,In_375,In_2766);
nor U1444 (N_1444,In_62,In_1554);
nand U1445 (N_1445,In_747,In_1702);
and U1446 (N_1446,In_2835,In_2756);
and U1447 (N_1447,In_1624,In_2649);
nand U1448 (N_1448,In_775,In_1393);
nand U1449 (N_1449,In_459,In_2428);
or U1450 (N_1450,In_2988,In_1274);
or U1451 (N_1451,In_685,In_2589);
xnor U1452 (N_1452,In_1017,In_525);
nand U1453 (N_1453,In_2847,In_960);
nand U1454 (N_1454,In_2081,In_338);
or U1455 (N_1455,In_2274,In_2886);
nand U1456 (N_1456,In_1999,In_2357);
nor U1457 (N_1457,In_2285,In_1894);
and U1458 (N_1458,In_972,In_2290);
xor U1459 (N_1459,In_2222,In_2477);
nor U1460 (N_1460,In_725,In_2538);
nor U1461 (N_1461,In_2821,In_786);
nand U1462 (N_1462,In_1694,In_1219);
xor U1463 (N_1463,In_919,In_675);
nand U1464 (N_1464,In_2775,In_868);
or U1465 (N_1465,In_929,In_1683);
nand U1466 (N_1466,In_845,In_1950);
or U1467 (N_1467,In_590,In_1099);
nand U1468 (N_1468,In_1146,In_1844);
or U1469 (N_1469,In_44,In_1523);
or U1470 (N_1470,In_227,In_347);
and U1471 (N_1471,In_741,In_1837);
nand U1472 (N_1472,In_274,In_377);
nand U1473 (N_1473,In_4,In_1584);
xor U1474 (N_1474,In_2028,In_1408);
nand U1475 (N_1475,In_2345,In_1152);
or U1476 (N_1476,In_1123,In_809);
or U1477 (N_1477,In_1645,In_866);
or U1478 (N_1478,In_1236,In_2999);
or U1479 (N_1479,In_869,In_2176);
nor U1480 (N_1480,In_1967,In_341);
xor U1481 (N_1481,In_1390,In_14);
or U1482 (N_1482,In_1818,In_617);
and U1483 (N_1483,In_2520,In_627);
and U1484 (N_1484,In_1286,In_151);
or U1485 (N_1485,In_2131,In_1310);
nand U1486 (N_1486,In_803,In_1760);
and U1487 (N_1487,In_1443,In_492);
nand U1488 (N_1488,In_2013,In_168);
xor U1489 (N_1489,In_1030,In_2390);
nor U1490 (N_1490,In_1613,In_1366);
or U1491 (N_1491,In_233,In_1504);
nand U1492 (N_1492,In_1442,In_530);
nand U1493 (N_1493,In_1337,In_1534);
nor U1494 (N_1494,In_1983,In_2512);
nor U1495 (N_1495,In_2877,In_1889);
or U1496 (N_1496,In_497,In_2772);
and U1497 (N_1497,In_172,In_2282);
nand U1498 (N_1498,In_1590,In_2578);
nor U1499 (N_1499,In_1758,In_108);
and U1500 (N_1500,In_2178,In_2596);
nor U1501 (N_1501,In_2435,In_1332);
and U1502 (N_1502,In_1740,In_333);
xnor U1503 (N_1503,In_1087,In_603);
and U1504 (N_1504,In_2299,In_1922);
xnor U1505 (N_1505,In_1166,In_1409);
xnor U1506 (N_1506,In_2724,In_2482);
and U1507 (N_1507,In_286,In_1386);
xor U1508 (N_1508,In_2376,In_1280);
nor U1509 (N_1509,In_716,In_230);
or U1510 (N_1510,In_673,In_168);
and U1511 (N_1511,In_1815,In_798);
or U1512 (N_1512,In_207,In_1348);
and U1513 (N_1513,In_1346,In_2946);
xnor U1514 (N_1514,In_9,In_2790);
nor U1515 (N_1515,In_745,In_2273);
and U1516 (N_1516,In_2758,In_1133);
xnor U1517 (N_1517,In_1156,In_2290);
nor U1518 (N_1518,In_1088,In_1894);
xnor U1519 (N_1519,In_1567,In_649);
nor U1520 (N_1520,In_514,In_1262);
and U1521 (N_1521,In_840,In_1457);
nand U1522 (N_1522,In_2646,In_320);
and U1523 (N_1523,In_2010,In_1116);
nor U1524 (N_1524,In_981,In_2391);
nor U1525 (N_1525,In_2490,In_1140);
nor U1526 (N_1526,In_1749,In_1043);
nor U1527 (N_1527,In_1330,In_1333);
xor U1528 (N_1528,In_645,In_673);
xnor U1529 (N_1529,In_1120,In_1654);
and U1530 (N_1530,In_2135,In_2520);
or U1531 (N_1531,In_2560,In_2959);
xor U1532 (N_1532,In_2181,In_2066);
or U1533 (N_1533,In_2953,In_2763);
xor U1534 (N_1534,In_1919,In_2245);
nor U1535 (N_1535,In_918,In_468);
and U1536 (N_1536,In_2974,In_158);
xnor U1537 (N_1537,In_1728,In_1406);
and U1538 (N_1538,In_2016,In_976);
xnor U1539 (N_1539,In_747,In_1342);
nor U1540 (N_1540,In_1516,In_919);
nand U1541 (N_1541,In_2939,In_701);
and U1542 (N_1542,In_1674,In_794);
nand U1543 (N_1543,In_2627,In_2971);
or U1544 (N_1544,In_1185,In_2621);
nor U1545 (N_1545,In_1522,In_591);
nand U1546 (N_1546,In_242,In_1655);
or U1547 (N_1547,In_586,In_2368);
or U1548 (N_1548,In_1495,In_2233);
nand U1549 (N_1549,In_2571,In_726);
or U1550 (N_1550,In_2077,In_738);
and U1551 (N_1551,In_556,In_1031);
or U1552 (N_1552,In_2863,In_1646);
nor U1553 (N_1553,In_417,In_874);
or U1554 (N_1554,In_531,In_474);
nor U1555 (N_1555,In_2662,In_484);
nand U1556 (N_1556,In_2703,In_172);
and U1557 (N_1557,In_779,In_2302);
and U1558 (N_1558,In_2650,In_1167);
or U1559 (N_1559,In_2726,In_1777);
and U1560 (N_1560,In_2458,In_613);
nand U1561 (N_1561,In_1439,In_2041);
nor U1562 (N_1562,In_1668,In_422);
or U1563 (N_1563,In_2049,In_2982);
and U1564 (N_1564,In_626,In_170);
nand U1565 (N_1565,In_794,In_1997);
nor U1566 (N_1566,In_434,In_1231);
and U1567 (N_1567,In_2410,In_767);
nor U1568 (N_1568,In_143,In_2649);
nor U1569 (N_1569,In_362,In_425);
nor U1570 (N_1570,In_139,In_2271);
or U1571 (N_1571,In_2987,In_2349);
xor U1572 (N_1572,In_2100,In_1344);
nor U1573 (N_1573,In_1162,In_1152);
xor U1574 (N_1574,In_2984,In_963);
and U1575 (N_1575,In_1848,In_2973);
nand U1576 (N_1576,In_119,In_1874);
and U1577 (N_1577,In_2559,In_896);
and U1578 (N_1578,In_1092,In_1709);
xor U1579 (N_1579,In_498,In_888);
nor U1580 (N_1580,In_1460,In_298);
nor U1581 (N_1581,In_134,In_444);
nor U1582 (N_1582,In_1057,In_541);
nor U1583 (N_1583,In_419,In_1218);
nor U1584 (N_1584,In_2631,In_1752);
and U1585 (N_1585,In_944,In_1401);
or U1586 (N_1586,In_881,In_467);
nand U1587 (N_1587,In_1600,In_272);
nor U1588 (N_1588,In_1925,In_1816);
or U1589 (N_1589,In_414,In_291);
or U1590 (N_1590,In_1569,In_2794);
or U1591 (N_1591,In_1770,In_2411);
or U1592 (N_1592,In_447,In_1620);
xor U1593 (N_1593,In_686,In_2599);
xnor U1594 (N_1594,In_2122,In_2064);
nor U1595 (N_1595,In_643,In_1311);
nand U1596 (N_1596,In_2748,In_149);
xor U1597 (N_1597,In_2366,In_311);
or U1598 (N_1598,In_2946,In_2928);
nand U1599 (N_1599,In_1693,In_2036);
or U1600 (N_1600,In_712,In_2979);
or U1601 (N_1601,In_133,In_2365);
xnor U1602 (N_1602,In_2135,In_2094);
xnor U1603 (N_1603,In_1641,In_1932);
and U1604 (N_1604,In_2407,In_1130);
xor U1605 (N_1605,In_1439,In_1776);
and U1606 (N_1606,In_915,In_2411);
xor U1607 (N_1607,In_2576,In_779);
nand U1608 (N_1608,In_2473,In_2710);
nand U1609 (N_1609,In_2885,In_2386);
nand U1610 (N_1610,In_1010,In_2644);
nor U1611 (N_1611,In_314,In_1410);
xnor U1612 (N_1612,In_2616,In_2031);
xnor U1613 (N_1613,In_1129,In_718);
nand U1614 (N_1614,In_1598,In_1160);
nand U1615 (N_1615,In_2812,In_212);
xnor U1616 (N_1616,In_162,In_815);
xnor U1617 (N_1617,In_191,In_290);
nor U1618 (N_1618,In_1633,In_2958);
and U1619 (N_1619,In_2036,In_356);
nor U1620 (N_1620,In_1761,In_2738);
nand U1621 (N_1621,In_2364,In_1412);
nand U1622 (N_1622,In_2719,In_804);
and U1623 (N_1623,In_1300,In_1343);
xnor U1624 (N_1624,In_2157,In_685);
xor U1625 (N_1625,In_2696,In_801);
xor U1626 (N_1626,In_337,In_2381);
and U1627 (N_1627,In_521,In_2849);
nand U1628 (N_1628,In_692,In_1030);
nor U1629 (N_1629,In_1835,In_2925);
nand U1630 (N_1630,In_2519,In_198);
nor U1631 (N_1631,In_1592,In_271);
xnor U1632 (N_1632,In_2469,In_1353);
xor U1633 (N_1633,In_2046,In_1401);
nand U1634 (N_1634,In_1750,In_825);
nand U1635 (N_1635,In_2869,In_1598);
and U1636 (N_1636,In_1686,In_2878);
nand U1637 (N_1637,In_184,In_2743);
nand U1638 (N_1638,In_921,In_1547);
or U1639 (N_1639,In_52,In_509);
or U1640 (N_1640,In_2858,In_2772);
nor U1641 (N_1641,In_2467,In_483);
nand U1642 (N_1642,In_2326,In_1671);
xnor U1643 (N_1643,In_930,In_746);
or U1644 (N_1644,In_1220,In_2721);
xor U1645 (N_1645,In_882,In_2158);
or U1646 (N_1646,In_1800,In_1000);
xnor U1647 (N_1647,In_2043,In_2647);
xnor U1648 (N_1648,In_2555,In_758);
and U1649 (N_1649,In_2680,In_2758);
xnor U1650 (N_1650,In_452,In_2583);
or U1651 (N_1651,In_2440,In_165);
or U1652 (N_1652,In_344,In_88);
or U1653 (N_1653,In_1319,In_384);
and U1654 (N_1654,In_1152,In_2139);
nor U1655 (N_1655,In_2195,In_1768);
or U1656 (N_1656,In_805,In_1574);
nor U1657 (N_1657,In_813,In_963);
nand U1658 (N_1658,In_2230,In_2590);
and U1659 (N_1659,In_1650,In_59);
and U1660 (N_1660,In_665,In_921);
or U1661 (N_1661,In_2646,In_262);
nor U1662 (N_1662,In_590,In_563);
and U1663 (N_1663,In_1242,In_424);
nand U1664 (N_1664,In_429,In_2732);
xnor U1665 (N_1665,In_692,In_1391);
and U1666 (N_1666,In_301,In_54);
nand U1667 (N_1667,In_1314,In_327);
xnor U1668 (N_1668,In_2885,In_2248);
nand U1669 (N_1669,In_1038,In_2644);
nor U1670 (N_1670,In_1677,In_2274);
xnor U1671 (N_1671,In_436,In_2107);
nand U1672 (N_1672,In_1154,In_1573);
or U1673 (N_1673,In_396,In_2987);
nand U1674 (N_1674,In_2815,In_311);
and U1675 (N_1675,In_2922,In_2857);
nor U1676 (N_1676,In_1883,In_1813);
or U1677 (N_1677,In_1453,In_1104);
nor U1678 (N_1678,In_1829,In_1904);
nand U1679 (N_1679,In_561,In_2054);
xnor U1680 (N_1680,In_2872,In_158);
or U1681 (N_1681,In_1000,In_1311);
or U1682 (N_1682,In_2836,In_2304);
or U1683 (N_1683,In_2817,In_713);
or U1684 (N_1684,In_232,In_2989);
nor U1685 (N_1685,In_688,In_2278);
or U1686 (N_1686,In_635,In_2883);
and U1687 (N_1687,In_2255,In_2560);
or U1688 (N_1688,In_1095,In_176);
or U1689 (N_1689,In_1628,In_606);
xor U1690 (N_1690,In_2541,In_2067);
nand U1691 (N_1691,In_519,In_1437);
nand U1692 (N_1692,In_998,In_305);
xnor U1693 (N_1693,In_875,In_2151);
nand U1694 (N_1694,In_1529,In_498);
nor U1695 (N_1695,In_228,In_1104);
or U1696 (N_1696,In_1989,In_1741);
nand U1697 (N_1697,In_1661,In_53);
and U1698 (N_1698,In_2608,In_620);
and U1699 (N_1699,In_2973,In_2763);
and U1700 (N_1700,In_28,In_2694);
and U1701 (N_1701,In_1901,In_2089);
or U1702 (N_1702,In_2940,In_822);
and U1703 (N_1703,In_1118,In_2855);
nand U1704 (N_1704,In_2083,In_261);
xor U1705 (N_1705,In_1192,In_558);
nor U1706 (N_1706,In_1026,In_1109);
nand U1707 (N_1707,In_21,In_540);
nor U1708 (N_1708,In_1185,In_2000);
and U1709 (N_1709,In_239,In_357);
xor U1710 (N_1710,In_2840,In_1805);
nor U1711 (N_1711,In_1362,In_166);
xnor U1712 (N_1712,In_79,In_162);
or U1713 (N_1713,In_1798,In_439);
nor U1714 (N_1714,In_1614,In_1671);
nor U1715 (N_1715,In_1319,In_137);
and U1716 (N_1716,In_1319,In_2783);
nor U1717 (N_1717,In_7,In_2938);
and U1718 (N_1718,In_2319,In_2663);
xor U1719 (N_1719,In_85,In_614);
nor U1720 (N_1720,In_1934,In_1056);
nor U1721 (N_1721,In_1450,In_2882);
and U1722 (N_1722,In_2613,In_1617);
or U1723 (N_1723,In_241,In_2386);
xnor U1724 (N_1724,In_885,In_2207);
xnor U1725 (N_1725,In_691,In_192);
nand U1726 (N_1726,In_1506,In_2794);
xor U1727 (N_1727,In_2123,In_100);
nor U1728 (N_1728,In_1831,In_2537);
nor U1729 (N_1729,In_1726,In_815);
and U1730 (N_1730,In_1978,In_204);
or U1731 (N_1731,In_1187,In_277);
nand U1732 (N_1732,In_1489,In_687);
nor U1733 (N_1733,In_364,In_2643);
and U1734 (N_1734,In_1450,In_1331);
xor U1735 (N_1735,In_1354,In_2046);
nand U1736 (N_1736,In_302,In_179);
nand U1737 (N_1737,In_1001,In_1105);
or U1738 (N_1738,In_2602,In_2436);
and U1739 (N_1739,In_37,In_446);
and U1740 (N_1740,In_1423,In_563);
nor U1741 (N_1741,In_2345,In_1947);
and U1742 (N_1742,In_1283,In_928);
or U1743 (N_1743,In_2076,In_2971);
nor U1744 (N_1744,In_138,In_1253);
nand U1745 (N_1745,In_2264,In_170);
or U1746 (N_1746,In_2194,In_883);
and U1747 (N_1747,In_1804,In_1358);
nor U1748 (N_1748,In_361,In_1611);
nor U1749 (N_1749,In_699,In_1676);
or U1750 (N_1750,In_2250,In_2346);
xnor U1751 (N_1751,In_459,In_1622);
xor U1752 (N_1752,In_2501,In_1776);
nand U1753 (N_1753,In_1867,In_607);
or U1754 (N_1754,In_202,In_419);
nor U1755 (N_1755,In_933,In_495);
xnor U1756 (N_1756,In_358,In_371);
and U1757 (N_1757,In_2465,In_2582);
nand U1758 (N_1758,In_2973,In_1410);
nand U1759 (N_1759,In_1334,In_2251);
xnor U1760 (N_1760,In_1862,In_2834);
nor U1761 (N_1761,In_659,In_2489);
nor U1762 (N_1762,In_1304,In_375);
xnor U1763 (N_1763,In_205,In_2251);
xnor U1764 (N_1764,In_285,In_2143);
or U1765 (N_1765,In_1574,In_2740);
nor U1766 (N_1766,In_731,In_90);
xor U1767 (N_1767,In_895,In_2426);
nor U1768 (N_1768,In_2445,In_1813);
nand U1769 (N_1769,In_1220,In_2766);
or U1770 (N_1770,In_851,In_1502);
and U1771 (N_1771,In_1682,In_1317);
nand U1772 (N_1772,In_2589,In_681);
and U1773 (N_1773,In_2873,In_2544);
nor U1774 (N_1774,In_1116,In_1387);
nand U1775 (N_1775,In_1551,In_1048);
nor U1776 (N_1776,In_1568,In_2022);
xor U1777 (N_1777,In_2508,In_2240);
xnor U1778 (N_1778,In_2990,In_1065);
xor U1779 (N_1779,In_1532,In_477);
and U1780 (N_1780,In_232,In_70);
nor U1781 (N_1781,In_2487,In_2872);
or U1782 (N_1782,In_404,In_1313);
and U1783 (N_1783,In_341,In_1625);
or U1784 (N_1784,In_856,In_2731);
nand U1785 (N_1785,In_1942,In_1458);
nand U1786 (N_1786,In_318,In_545);
or U1787 (N_1787,In_1610,In_1146);
or U1788 (N_1788,In_1013,In_1024);
and U1789 (N_1789,In_387,In_2551);
nand U1790 (N_1790,In_586,In_1337);
or U1791 (N_1791,In_1626,In_1163);
nand U1792 (N_1792,In_2136,In_198);
or U1793 (N_1793,In_603,In_2420);
nor U1794 (N_1794,In_2891,In_545);
or U1795 (N_1795,In_2180,In_2691);
nor U1796 (N_1796,In_2672,In_268);
nand U1797 (N_1797,In_1534,In_1817);
or U1798 (N_1798,In_1299,In_1577);
nor U1799 (N_1799,In_1061,In_2492);
and U1800 (N_1800,In_165,In_2296);
or U1801 (N_1801,In_470,In_1763);
xnor U1802 (N_1802,In_1201,In_2183);
and U1803 (N_1803,In_1638,In_2613);
xor U1804 (N_1804,In_2021,In_535);
xnor U1805 (N_1805,In_1971,In_676);
xnor U1806 (N_1806,In_2646,In_1207);
or U1807 (N_1807,In_1721,In_1245);
nand U1808 (N_1808,In_1053,In_2042);
and U1809 (N_1809,In_28,In_764);
xor U1810 (N_1810,In_580,In_1963);
or U1811 (N_1811,In_2121,In_2932);
or U1812 (N_1812,In_2405,In_1370);
and U1813 (N_1813,In_1709,In_1304);
and U1814 (N_1814,In_2087,In_1064);
nand U1815 (N_1815,In_1566,In_1366);
nor U1816 (N_1816,In_523,In_2427);
or U1817 (N_1817,In_1216,In_914);
nand U1818 (N_1818,In_2681,In_2137);
nand U1819 (N_1819,In_2922,In_2144);
nand U1820 (N_1820,In_2260,In_2769);
nor U1821 (N_1821,In_1866,In_2767);
nor U1822 (N_1822,In_2871,In_2602);
or U1823 (N_1823,In_2093,In_606);
nor U1824 (N_1824,In_1986,In_1784);
xor U1825 (N_1825,In_2340,In_809);
xnor U1826 (N_1826,In_149,In_2386);
and U1827 (N_1827,In_739,In_2706);
or U1828 (N_1828,In_1293,In_1475);
nand U1829 (N_1829,In_833,In_2744);
xnor U1830 (N_1830,In_999,In_2298);
nor U1831 (N_1831,In_1495,In_452);
nor U1832 (N_1832,In_335,In_928);
nor U1833 (N_1833,In_2492,In_2121);
xnor U1834 (N_1834,In_914,In_1871);
and U1835 (N_1835,In_889,In_343);
xnor U1836 (N_1836,In_2439,In_2259);
xor U1837 (N_1837,In_2690,In_754);
or U1838 (N_1838,In_1764,In_2151);
and U1839 (N_1839,In_778,In_587);
nor U1840 (N_1840,In_137,In_899);
nand U1841 (N_1841,In_2174,In_1673);
nor U1842 (N_1842,In_671,In_146);
nand U1843 (N_1843,In_2791,In_2129);
nand U1844 (N_1844,In_426,In_2258);
nor U1845 (N_1845,In_1020,In_1237);
xnor U1846 (N_1846,In_1689,In_2346);
or U1847 (N_1847,In_264,In_2003);
nand U1848 (N_1848,In_2419,In_1378);
and U1849 (N_1849,In_1119,In_725);
nand U1850 (N_1850,In_467,In_2965);
xnor U1851 (N_1851,In_2884,In_1728);
nand U1852 (N_1852,In_2019,In_1282);
or U1853 (N_1853,In_958,In_2573);
and U1854 (N_1854,In_2851,In_1299);
nand U1855 (N_1855,In_2498,In_1098);
nand U1856 (N_1856,In_509,In_1573);
nand U1857 (N_1857,In_269,In_1188);
xor U1858 (N_1858,In_1420,In_1659);
nand U1859 (N_1859,In_1367,In_427);
or U1860 (N_1860,In_922,In_862);
and U1861 (N_1861,In_1777,In_2009);
and U1862 (N_1862,In_262,In_668);
xnor U1863 (N_1863,In_2960,In_2138);
or U1864 (N_1864,In_2062,In_2872);
and U1865 (N_1865,In_600,In_418);
xor U1866 (N_1866,In_1359,In_1799);
nand U1867 (N_1867,In_2364,In_2979);
and U1868 (N_1868,In_1318,In_1680);
xor U1869 (N_1869,In_810,In_793);
and U1870 (N_1870,In_946,In_1801);
nor U1871 (N_1871,In_1112,In_1047);
and U1872 (N_1872,In_942,In_677);
nand U1873 (N_1873,In_2159,In_2931);
and U1874 (N_1874,In_2328,In_673);
nor U1875 (N_1875,In_1762,In_626);
nand U1876 (N_1876,In_286,In_1658);
and U1877 (N_1877,In_1101,In_2190);
xnor U1878 (N_1878,In_1770,In_1583);
nor U1879 (N_1879,In_141,In_1439);
and U1880 (N_1880,In_1141,In_1698);
or U1881 (N_1881,In_2619,In_958);
nand U1882 (N_1882,In_436,In_1212);
and U1883 (N_1883,In_2395,In_323);
and U1884 (N_1884,In_32,In_1861);
nand U1885 (N_1885,In_1037,In_1176);
nor U1886 (N_1886,In_346,In_1638);
xor U1887 (N_1887,In_2633,In_165);
xor U1888 (N_1888,In_11,In_1324);
and U1889 (N_1889,In_220,In_2934);
nor U1890 (N_1890,In_2856,In_2925);
nand U1891 (N_1891,In_1934,In_2910);
and U1892 (N_1892,In_734,In_977);
nand U1893 (N_1893,In_1627,In_435);
nor U1894 (N_1894,In_2092,In_436);
nand U1895 (N_1895,In_420,In_2965);
xor U1896 (N_1896,In_2803,In_771);
or U1897 (N_1897,In_2114,In_2865);
nor U1898 (N_1898,In_9,In_1800);
xor U1899 (N_1899,In_2931,In_1177);
xor U1900 (N_1900,In_977,In_546);
or U1901 (N_1901,In_1376,In_1144);
nand U1902 (N_1902,In_2797,In_2955);
and U1903 (N_1903,In_1257,In_2703);
and U1904 (N_1904,In_1913,In_1014);
and U1905 (N_1905,In_996,In_30);
and U1906 (N_1906,In_1602,In_1202);
nor U1907 (N_1907,In_832,In_276);
nand U1908 (N_1908,In_2860,In_2421);
or U1909 (N_1909,In_1698,In_2434);
and U1910 (N_1910,In_1864,In_2277);
nor U1911 (N_1911,In_1855,In_692);
xor U1912 (N_1912,In_1393,In_1852);
xnor U1913 (N_1913,In_1741,In_2237);
xor U1914 (N_1914,In_1909,In_2467);
nor U1915 (N_1915,In_576,In_497);
or U1916 (N_1916,In_1611,In_2758);
or U1917 (N_1917,In_2876,In_2274);
nand U1918 (N_1918,In_1829,In_738);
nand U1919 (N_1919,In_962,In_2732);
or U1920 (N_1920,In_2274,In_2639);
xnor U1921 (N_1921,In_2052,In_1550);
xor U1922 (N_1922,In_2262,In_139);
or U1923 (N_1923,In_481,In_416);
nor U1924 (N_1924,In_1507,In_1553);
nor U1925 (N_1925,In_62,In_384);
xor U1926 (N_1926,In_1121,In_430);
and U1927 (N_1927,In_845,In_937);
or U1928 (N_1928,In_955,In_1795);
nor U1929 (N_1929,In_1347,In_2571);
nand U1930 (N_1930,In_2715,In_406);
xor U1931 (N_1931,In_1715,In_156);
nand U1932 (N_1932,In_1556,In_969);
xnor U1933 (N_1933,In_305,In_2443);
nand U1934 (N_1934,In_2075,In_501);
nand U1935 (N_1935,In_1920,In_2085);
or U1936 (N_1936,In_1053,In_1552);
xor U1937 (N_1937,In_2485,In_2642);
xor U1938 (N_1938,In_1941,In_1557);
or U1939 (N_1939,In_2205,In_473);
and U1940 (N_1940,In_2783,In_679);
xor U1941 (N_1941,In_1536,In_1452);
xor U1942 (N_1942,In_1955,In_2489);
nor U1943 (N_1943,In_2077,In_2180);
nand U1944 (N_1944,In_868,In_1770);
or U1945 (N_1945,In_544,In_2124);
nand U1946 (N_1946,In_1367,In_312);
or U1947 (N_1947,In_1151,In_580);
nor U1948 (N_1948,In_1912,In_2511);
nand U1949 (N_1949,In_377,In_947);
nor U1950 (N_1950,In_1588,In_1867);
and U1951 (N_1951,In_2931,In_1243);
xnor U1952 (N_1952,In_528,In_2892);
nor U1953 (N_1953,In_2422,In_2972);
nand U1954 (N_1954,In_277,In_729);
nor U1955 (N_1955,In_2753,In_2551);
nand U1956 (N_1956,In_1453,In_977);
and U1957 (N_1957,In_2899,In_144);
and U1958 (N_1958,In_532,In_1172);
nor U1959 (N_1959,In_2866,In_1519);
and U1960 (N_1960,In_2220,In_2983);
nand U1961 (N_1961,In_62,In_611);
or U1962 (N_1962,In_2009,In_76);
nor U1963 (N_1963,In_1391,In_2691);
and U1964 (N_1964,In_652,In_31);
nand U1965 (N_1965,In_1150,In_113);
nand U1966 (N_1966,In_58,In_84);
nor U1967 (N_1967,In_1686,In_2343);
nand U1968 (N_1968,In_346,In_2812);
xor U1969 (N_1969,In_166,In_1100);
xnor U1970 (N_1970,In_1280,In_237);
and U1971 (N_1971,In_2147,In_2389);
nor U1972 (N_1972,In_1798,In_585);
nand U1973 (N_1973,In_2508,In_2433);
nor U1974 (N_1974,In_2665,In_1095);
nor U1975 (N_1975,In_1476,In_1831);
xor U1976 (N_1976,In_106,In_2638);
nor U1977 (N_1977,In_2105,In_2179);
and U1978 (N_1978,In_1677,In_1483);
and U1979 (N_1979,In_2752,In_2377);
xor U1980 (N_1980,In_2363,In_2449);
xor U1981 (N_1981,In_298,In_2242);
and U1982 (N_1982,In_1137,In_1184);
or U1983 (N_1983,In_928,In_872);
and U1984 (N_1984,In_1426,In_1395);
xor U1985 (N_1985,In_1915,In_1695);
xnor U1986 (N_1986,In_2967,In_1175);
xor U1987 (N_1987,In_167,In_1752);
nor U1988 (N_1988,In_2592,In_665);
xnor U1989 (N_1989,In_2287,In_2785);
nand U1990 (N_1990,In_2040,In_1744);
or U1991 (N_1991,In_1888,In_2714);
xor U1992 (N_1992,In_501,In_2132);
nor U1993 (N_1993,In_2937,In_2340);
nand U1994 (N_1994,In_126,In_1487);
xnor U1995 (N_1995,In_2389,In_2675);
or U1996 (N_1996,In_2562,In_2494);
xnor U1997 (N_1997,In_411,In_1673);
xor U1998 (N_1998,In_2765,In_1947);
or U1999 (N_1999,In_712,In_739);
and U2000 (N_2000,In_328,In_817);
nand U2001 (N_2001,In_807,In_458);
nand U2002 (N_2002,In_2963,In_2886);
nor U2003 (N_2003,In_2564,In_1193);
and U2004 (N_2004,In_1440,In_2851);
xnor U2005 (N_2005,In_940,In_1315);
or U2006 (N_2006,In_802,In_2974);
and U2007 (N_2007,In_2700,In_29);
nand U2008 (N_2008,In_2567,In_2419);
nor U2009 (N_2009,In_1472,In_1113);
xor U2010 (N_2010,In_1101,In_59);
or U2011 (N_2011,In_242,In_2573);
xor U2012 (N_2012,In_1937,In_1247);
nor U2013 (N_2013,In_2662,In_2170);
or U2014 (N_2014,In_994,In_2184);
nand U2015 (N_2015,In_61,In_2770);
nand U2016 (N_2016,In_2640,In_271);
and U2017 (N_2017,In_773,In_1447);
nor U2018 (N_2018,In_651,In_1126);
or U2019 (N_2019,In_195,In_821);
or U2020 (N_2020,In_226,In_211);
nor U2021 (N_2021,In_64,In_2767);
nor U2022 (N_2022,In_1358,In_641);
xor U2023 (N_2023,In_627,In_282);
or U2024 (N_2024,In_2453,In_1353);
xnor U2025 (N_2025,In_1161,In_675);
xor U2026 (N_2026,In_2004,In_2413);
nor U2027 (N_2027,In_921,In_1974);
nand U2028 (N_2028,In_107,In_1101);
nor U2029 (N_2029,In_2766,In_228);
or U2030 (N_2030,In_2116,In_873);
or U2031 (N_2031,In_2300,In_1764);
nor U2032 (N_2032,In_1858,In_259);
xnor U2033 (N_2033,In_1153,In_582);
and U2034 (N_2034,In_1377,In_1077);
nor U2035 (N_2035,In_1039,In_1341);
nor U2036 (N_2036,In_1074,In_845);
nand U2037 (N_2037,In_2282,In_1419);
or U2038 (N_2038,In_1156,In_2717);
or U2039 (N_2039,In_1169,In_568);
xnor U2040 (N_2040,In_2906,In_731);
and U2041 (N_2041,In_2115,In_1955);
nand U2042 (N_2042,In_1183,In_1103);
and U2043 (N_2043,In_2848,In_1475);
nor U2044 (N_2044,In_1916,In_2658);
xnor U2045 (N_2045,In_2426,In_2621);
xnor U2046 (N_2046,In_1046,In_1332);
and U2047 (N_2047,In_1433,In_1564);
nand U2048 (N_2048,In_445,In_418);
xor U2049 (N_2049,In_2306,In_164);
and U2050 (N_2050,In_2130,In_2374);
xnor U2051 (N_2051,In_1637,In_672);
or U2052 (N_2052,In_1166,In_2032);
nor U2053 (N_2053,In_907,In_1730);
or U2054 (N_2054,In_2624,In_2732);
xor U2055 (N_2055,In_1768,In_2115);
or U2056 (N_2056,In_1244,In_847);
nor U2057 (N_2057,In_1367,In_1484);
or U2058 (N_2058,In_686,In_1384);
and U2059 (N_2059,In_2535,In_1904);
xor U2060 (N_2060,In_2876,In_843);
xor U2061 (N_2061,In_901,In_914);
and U2062 (N_2062,In_194,In_2932);
nor U2063 (N_2063,In_2929,In_618);
nor U2064 (N_2064,In_2849,In_1635);
or U2065 (N_2065,In_2376,In_290);
xor U2066 (N_2066,In_918,In_1161);
or U2067 (N_2067,In_767,In_2775);
and U2068 (N_2068,In_2008,In_701);
or U2069 (N_2069,In_1977,In_1832);
and U2070 (N_2070,In_888,In_1648);
or U2071 (N_2071,In_2635,In_2642);
nand U2072 (N_2072,In_2566,In_494);
or U2073 (N_2073,In_1212,In_2561);
and U2074 (N_2074,In_145,In_1323);
nor U2075 (N_2075,In_392,In_2081);
or U2076 (N_2076,In_845,In_2202);
nand U2077 (N_2077,In_1527,In_2435);
nand U2078 (N_2078,In_906,In_651);
nor U2079 (N_2079,In_1599,In_2123);
nand U2080 (N_2080,In_1563,In_1283);
nand U2081 (N_2081,In_1041,In_652);
or U2082 (N_2082,In_2332,In_918);
nor U2083 (N_2083,In_4,In_1612);
and U2084 (N_2084,In_2731,In_446);
xor U2085 (N_2085,In_183,In_2549);
nand U2086 (N_2086,In_2378,In_757);
xnor U2087 (N_2087,In_1270,In_2045);
xor U2088 (N_2088,In_1864,In_2902);
nor U2089 (N_2089,In_2963,In_2263);
or U2090 (N_2090,In_568,In_270);
and U2091 (N_2091,In_216,In_157);
xnor U2092 (N_2092,In_1692,In_692);
xor U2093 (N_2093,In_2188,In_2447);
xnor U2094 (N_2094,In_2925,In_1532);
and U2095 (N_2095,In_1487,In_2215);
or U2096 (N_2096,In_1402,In_2819);
and U2097 (N_2097,In_1058,In_2034);
nor U2098 (N_2098,In_1934,In_2575);
nor U2099 (N_2099,In_1760,In_1341);
nand U2100 (N_2100,In_1478,In_1650);
or U2101 (N_2101,In_95,In_462);
and U2102 (N_2102,In_1732,In_1433);
nor U2103 (N_2103,In_2437,In_335);
xor U2104 (N_2104,In_994,In_2322);
nor U2105 (N_2105,In_439,In_2161);
nand U2106 (N_2106,In_535,In_977);
xor U2107 (N_2107,In_159,In_2514);
nor U2108 (N_2108,In_1809,In_161);
and U2109 (N_2109,In_1607,In_1338);
or U2110 (N_2110,In_1684,In_526);
nand U2111 (N_2111,In_1124,In_831);
nor U2112 (N_2112,In_2928,In_1233);
nand U2113 (N_2113,In_645,In_544);
nor U2114 (N_2114,In_1682,In_792);
and U2115 (N_2115,In_1221,In_2329);
and U2116 (N_2116,In_1609,In_758);
or U2117 (N_2117,In_2369,In_216);
or U2118 (N_2118,In_1764,In_410);
xor U2119 (N_2119,In_757,In_572);
nor U2120 (N_2120,In_2709,In_2107);
nor U2121 (N_2121,In_1982,In_2901);
nor U2122 (N_2122,In_1184,In_2364);
or U2123 (N_2123,In_1829,In_2087);
xnor U2124 (N_2124,In_2609,In_73);
xor U2125 (N_2125,In_2128,In_2688);
or U2126 (N_2126,In_159,In_335);
or U2127 (N_2127,In_1494,In_2234);
or U2128 (N_2128,In_2629,In_665);
and U2129 (N_2129,In_2703,In_2076);
and U2130 (N_2130,In_2967,In_2061);
nor U2131 (N_2131,In_241,In_2844);
or U2132 (N_2132,In_956,In_1960);
and U2133 (N_2133,In_2182,In_516);
and U2134 (N_2134,In_2330,In_1518);
or U2135 (N_2135,In_1099,In_2703);
and U2136 (N_2136,In_2337,In_1352);
nor U2137 (N_2137,In_747,In_288);
xor U2138 (N_2138,In_2900,In_2925);
xnor U2139 (N_2139,In_950,In_2207);
or U2140 (N_2140,In_464,In_1319);
or U2141 (N_2141,In_2282,In_1719);
and U2142 (N_2142,In_346,In_767);
nand U2143 (N_2143,In_1715,In_874);
xor U2144 (N_2144,In_134,In_103);
and U2145 (N_2145,In_2104,In_1778);
xnor U2146 (N_2146,In_2810,In_2850);
xor U2147 (N_2147,In_2775,In_2719);
and U2148 (N_2148,In_1364,In_2418);
or U2149 (N_2149,In_123,In_2313);
and U2150 (N_2150,In_2166,In_1683);
or U2151 (N_2151,In_1347,In_1213);
xnor U2152 (N_2152,In_1928,In_535);
xor U2153 (N_2153,In_151,In_30);
or U2154 (N_2154,In_1952,In_2128);
nor U2155 (N_2155,In_1231,In_2199);
xnor U2156 (N_2156,In_678,In_1359);
xnor U2157 (N_2157,In_1141,In_1190);
xnor U2158 (N_2158,In_1121,In_1412);
or U2159 (N_2159,In_2606,In_1097);
or U2160 (N_2160,In_2188,In_1701);
and U2161 (N_2161,In_1081,In_2850);
and U2162 (N_2162,In_1123,In_1172);
xor U2163 (N_2163,In_1084,In_2173);
nor U2164 (N_2164,In_90,In_1638);
nand U2165 (N_2165,In_558,In_26);
and U2166 (N_2166,In_2035,In_2127);
nand U2167 (N_2167,In_835,In_2467);
or U2168 (N_2168,In_452,In_2691);
nor U2169 (N_2169,In_1320,In_1805);
or U2170 (N_2170,In_2046,In_2072);
and U2171 (N_2171,In_1394,In_580);
nand U2172 (N_2172,In_1448,In_2992);
nand U2173 (N_2173,In_2420,In_790);
or U2174 (N_2174,In_41,In_929);
and U2175 (N_2175,In_1426,In_156);
or U2176 (N_2176,In_2761,In_2778);
or U2177 (N_2177,In_559,In_2425);
nor U2178 (N_2178,In_1791,In_1289);
and U2179 (N_2179,In_1850,In_1570);
nor U2180 (N_2180,In_2403,In_1851);
or U2181 (N_2181,In_1083,In_1872);
xnor U2182 (N_2182,In_2620,In_1361);
nor U2183 (N_2183,In_526,In_985);
or U2184 (N_2184,In_1283,In_2052);
xnor U2185 (N_2185,In_617,In_1779);
xnor U2186 (N_2186,In_737,In_2683);
and U2187 (N_2187,In_2411,In_1919);
and U2188 (N_2188,In_412,In_215);
and U2189 (N_2189,In_955,In_11);
xor U2190 (N_2190,In_2760,In_78);
xor U2191 (N_2191,In_2116,In_2720);
nor U2192 (N_2192,In_2937,In_1626);
xor U2193 (N_2193,In_884,In_1477);
nand U2194 (N_2194,In_975,In_2217);
or U2195 (N_2195,In_975,In_345);
nor U2196 (N_2196,In_965,In_2917);
nor U2197 (N_2197,In_1809,In_134);
nor U2198 (N_2198,In_1099,In_1443);
nand U2199 (N_2199,In_2967,In_2067);
nand U2200 (N_2200,In_395,In_1106);
and U2201 (N_2201,In_1725,In_2762);
nor U2202 (N_2202,In_861,In_20);
or U2203 (N_2203,In_679,In_1962);
and U2204 (N_2204,In_1477,In_1744);
and U2205 (N_2205,In_1048,In_1578);
nor U2206 (N_2206,In_2563,In_1279);
xnor U2207 (N_2207,In_1760,In_2642);
and U2208 (N_2208,In_358,In_1345);
or U2209 (N_2209,In_2742,In_2686);
nand U2210 (N_2210,In_2073,In_1577);
xnor U2211 (N_2211,In_419,In_1602);
nor U2212 (N_2212,In_2371,In_1661);
or U2213 (N_2213,In_241,In_124);
and U2214 (N_2214,In_1433,In_2900);
nand U2215 (N_2215,In_1390,In_714);
nor U2216 (N_2216,In_156,In_2805);
nand U2217 (N_2217,In_2604,In_2293);
and U2218 (N_2218,In_806,In_2490);
xor U2219 (N_2219,In_2766,In_2824);
and U2220 (N_2220,In_400,In_30);
or U2221 (N_2221,In_1957,In_400);
nor U2222 (N_2222,In_107,In_833);
xnor U2223 (N_2223,In_1107,In_2051);
nand U2224 (N_2224,In_1666,In_552);
or U2225 (N_2225,In_741,In_298);
xnor U2226 (N_2226,In_82,In_2456);
xor U2227 (N_2227,In_1478,In_1389);
or U2228 (N_2228,In_2601,In_1207);
nand U2229 (N_2229,In_2107,In_1829);
or U2230 (N_2230,In_2406,In_568);
nand U2231 (N_2231,In_1917,In_2329);
or U2232 (N_2232,In_1253,In_2615);
and U2233 (N_2233,In_2271,In_251);
nor U2234 (N_2234,In_1645,In_2699);
or U2235 (N_2235,In_2620,In_820);
or U2236 (N_2236,In_1738,In_2948);
or U2237 (N_2237,In_1153,In_2972);
nand U2238 (N_2238,In_1307,In_941);
nor U2239 (N_2239,In_952,In_1524);
or U2240 (N_2240,In_2648,In_1156);
xor U2241 (N_2241,In_382,In_1270);
nand U2242 (N_2242,In_923,In_651);
and U2243 (N_2243,In_2479,In_302);
or U2244 (N_2244,In_2129,In_1103);
nor U2245 (N_2245,In_560,In_335);
nor U2246 (N_2246,In_652,In_287);
nor U2247 (N_2247,In_1828,In_615);
nand U2248 (N_2248,In_624,In_1065);
or U2249 (N_2249,In_20,In_498);
nand U2250 (N_2250,In_1522,In_2896);
xnor U2251 (N_2251,In_495,In_2837);
nand U2252 (N_2252,In_755,In_843);
nor U2253 (N_2253,In_2159,In_680);
and U2254 (N_2254,In_2524,In_519);
xnor U2255 (N_2255,In_536,In_121);
and U2256 (N_2256,In_406,In_1751);
xnor U2257 (N_2257,In_1376,In_2949);
or U2258 (N_2258,In_2885,In_1119);
and U2259 (N_2259,In_825,In_2610);
xnor U2260 (N_2260,In_2085,In_2490);
xor U2261 (N_2261,In_2795,In_2776);
or U2262 (N_2262,In_1081,In_2656);
or U2263 (N_2263,In_2334,In_55);
and U2264 (N_2264,In_697,In_2148);
xnor U2265 (N_2265,In_2053,In_2627);
and U2266 (N_2266,In_1997,In_284);
xor U2267 (N_2267,In_1355,In_291);
nor U2268 (N_2268,In_184,In_820);
nand U2269 (N_2269,In_727,In_2787);
and U2270 (N_2270,In_198,In_2358);
and U2271 (N_2271,In_495,In_417);
and U2272 (N_2272,In_22,In_755);
or U2273 (N_2273,In_1131,In_667);
or U2274 (N_2274,In_878,In_40);
or U2275 (N_2275,In_2421,In_664);
and U2276 (N_2276,In_953,In_2965);
xor U2277 (N_2277,In_1189,In_1813);
and U2278 (N_2278,In_542,In_354);
nor U2279 (N_2279,In_2741,In_184);
nor U2280 (N_2280,In_1415,In_810);
or U2281 (N_2281,In_2206,In_667);
xnor U2282 (N_2282,In_1883,In_2287);
xnor U2283 (N_2283,In_2545,In_932);
or U2284 (N_2284,In_420,In_1329);
nor U2285 (N_2285,In_2681,In_462);
or U2286 (N_2286,In_945,In_2945);
and U2287 (N_2287,In_2906,In_462);
nand U2288 (N_2288,In_1543,In_2190);
nand U2289 (N_2289,In_543,In_2423);
and U2290 (N_2290,In_387,In_201);
xnor U2291 (N_2291,In_961,In_24);
xor U2292 (N_2292,In_1379,In_725);
and U2293 (N_2293,In_2815,In_1072);
nor U2294 (N_2294,In_312,In_1059);
xnor U2295 (N_2295,In_598,In_1384);
and U2296 (N_2296,In_655,In_891);
or U2297 (N_2297,In_252,In_498);
or U2298 (N_2298,In_181,In_486);
nand U2299 (N_2299,In_105,In_619);
nand U2300 (N_2300,In_1315,In_2930);
nand U2301 (N_2301,In_1132,In_2266);
nor U2302 (N_2302,In_367,In_14);
nor U2303 (N_2303,In_1306,In_1998);
or U2304 (N_2304,In_2642,In_2424);
nand U2305 (N_2305,In_1186,In_257);
xnor U2306 (N_2306,In_2413,In_851);
or U2307 (N_2307,In_661,In_2018);
and U2308 (N_2308,In_1778,In_563);
and U2309 (N_2309,In_240,In_1882);
or U2310 (N_2310,In_2585,In_1555);
nand U2311 (N_2311,In_2194,In_1803);
nor U2312 (N_2312,In_1998,In_778);
nand U2313 (N_2313,In_2822,In_734);
and U2314 (N_2314,In_1772,In_2279);
xor U2315 (N_2315,In_1100,In_2886);
nand U2316 (N_2316,In_965,In_2974);
xnor U2317 (N_2317,In_1693,In_2229);
nor U2318 (N_2318,In_2350,In_399);
xnor U2319 (N_2319,In_2517,In_1872);
nor U2320 (N_2320,In_1639,In_2035);
and U2321 (N_2321,In_2670,In_311);
nor U2322 (N_2322,In_1649,In_347);
nor U2323 (N_2323,In_1028,In_79);
xor U2324 (N_2324,In_44,In_779);
and U2325 (N_2325,In_679,In_2090);
xnor U2326 (N_2326,In_2710,In_1450);
nor U2327 (N_2327,In_2404,In_1368);
xor U2328 (N_2328,In_2162,In_168);
or U2329 (N_2329,In_2348,In_286);
nor U2330 (N_2330,In_1748,In_802);
nor U2331 (N_2331,In_231,In_1907);
xnor U2332 (N_2332,In_2767,In_653);
or U2333 (N_2333,In_2974,In_1335);
or U2334 (N_2334,In_2639,In_1790);
nand U2335 (N_2335,In_657,In_2522);
xnor U2336 (N_2336,In_465,In_2564);
or U2337 (N_2337,In_2604,In_1746);
or U2338 (N_2338,In_1870,In_2941);
or U2339 (N_2339,In_2237,In_1998);
xor U2340 (N_2340,In_2562,In_1066);
or U2341 (N_2341,In_747,In_1555);
and U2342 (N_2342,In_952,In_2588);
and U2343 (N_2343,In_565,In_983);
and U2344 (N_2344,In_10,In_755);
nand U2345 (N_2345,In_755,In_938);
and U2346 (N_2346,In_2426,In_204);
and U2347 (N_2347,In_285,In_52);
xnor U2348 (N_2348,In_2767,In_156);
xnor U2349 (N_2349,In_1002,In_2462);
xor U2350 (N_2350,In_2457,In_553);
nand U2351 (N_2351,In_119,In_1592);
nor U2352 (N_2352,In_221,In_2020);
or U2353 (N_2353,In_2789,In_487);
nor U2354 (N_2354,In_2629,In_1417);
nand U2355 (N_2355,In_744,In_2482);
nor U2356 (N_2356,In_694,In_1202);
and U2357 (N_2357,In_2676,In_1478);
and U2358 (N_2358,In_904,In_2985);
or U2359 (N_2359,In_1045,In_228);
nand U2360 (N_2360,In_2210,In_764);
nor U2361 (N_2361,In_2576,In_2637);
nor U2362 (N_2362,In_2935,In_2683);
nand U2363 (N_2363,In_2882,In_1490);
xnor U2364 (N_2364,In_1520,In_2162);
xnor U2365 (N_2365,In_2629,In_1326);
or U2366 (N_2366,In_428,In_2480);
xnor U2367 (N_2367,In_1965,In_1603);
nor U2368 (N_2368,In_25,In_470);
nand U2369 (N_2369,In_1340,In_101);
and U2370 (N_2370,In_472,In_1826);
and U2371 (N_2371,In_1580,In_245);
nand U2372 (N_2372,In_2408,In_1693);
or U2373 (N_2373,In_1027,In_811);
or U2374 (N_2374,In_2125,In_584);
nor U2375 (N_2375,In_753,In_85);
and U2376 (N_2376,In_1741,In_1510);
xor U2377 (N_2377,In_1273,In_2359);
xor U2378 (N_2378,In_689,In_1961);
or U2379 (N_2379,In_12,In_405);
nor U2380 (N_2380,In_1985,In_1316);
and U2381 (N_2381,In_193,In_1742);
nor U2382 (N_2382,In_1902,In_776);
nor U2383 (N_2383,In_2354,In_14);
or U2384 (N_2384,In_1021,In_1163);
or U2385 (N_2385,In_658,In_598);
nor U2386 (N_2386,In_1402,In_459);
nor U2387 (N_2387,In_2335,In_502);
and U2388 (N_2388,In_1832,In_953);
or U2389 (N_2389,In_2630,In_1312);
nor U2390 (N_2390,In_2240,In_801);
and U2391 (N_2391,In_2443,In_1099);
or U2392 (N_2392,In_805,In_742);
xor U2393 (N_2393,In_1725,In_2991);
and U2394 (N_2394,In_1241,In_2796);
xor U2395 (N_2395,In_1931,In_209);
nor U2396 (N_2396,In_652,In_2724);
nand U2397 (N_2397,In_1038,In_2316);
and U2398 (N_2398,In_639,In_691);
or U2399 (N_2399,In_1032,In_2596);
and U2400 (N_2400,In_2613,In_689);
nor U2401 (N_2401,In_361,In_2465);
nor U2402 (N_2402,In_1805,In_2494);
xnor U2403 (N_2403,In_126,In_1590);
or U2404 (N_2404,In_2001,In_2210);
or U2405 (N_2405,In_873,In_2805);
or U2406 (N_2406,In_2425,In_2786);
xnor U2407 (N_2407,In_252,In_1479);
and U2408 (N_2408,In_1342,In_2265);
xor U2409 (N_2409,In_2284,In_395);
or U2410 (N_2410,In_339,In_2578);
nor U2411 (N_2411,In_2599,In_2116);
xnor U2412 (N_2412,In_1827,In_1009);
xnor U2413 (N_2413,In_115,In_1180);
nor U2414 (N_2414,In_1787,In_1617);
and U2415 (N_2415,In_333,In_1980);
nor U2416 (N_2416,In_1323,In_580);
or U2417 (N_2417,In_2935,In_1816);
nor U2418 (N_2418,In_765,In_1938);
or U2419 (N_2419,In_968,In_355);
and U2420 (N_2420,In_2681,In_1074);
and U2421 (N_2421,In_1639,In_2093);
xor U2422 (N_2422,In_29,In_2083);
or U2423 (N_2423,In_758,In_2429);
nor U2424 (N_2424,In_1248,In_2137);
xor U2425 (N_2425,In_179,In_2528);
nand U2426 (N_2426,In_2229,In_2254);
nand U2427 (N_2427,In_726,In_776);
nor U2428 (N_2428,In_396,In_1757);
nor U2429 (N_2429,In_351,In_2418);
xor U2430 (N_2430,In_2003,In_297);
and U2431 (N_2431,In_362,In_194);
nand U2432 (N_2432,In_1223,In_2456);
or U2433 (N_2433,In_2204,In_1006);
or U2434 (N_2434,In_1791,In_2359);
nand U2435 (N_2435,In_1238,In_1756);
and U2436 (N_2436,In_678,In_1176);
and U2437 (N_2437,In_1327,In_1331);
and U2438 (N_2438,In_10,In_2559);
xnor U2439 (N_2439,In_1853,In_2663);
and U2440 (N_2440,In_1356,In_1188);
nor U2441 (N_2441,In_661,In_121);
or U2442 (N_2442,In_554,In_534);
xnor U2443 (N_2443,In_2814,In_1830);
or U2444 (N_2444,In_520,In_2062);
xor U2445 (N_2445,In_2510,In_1102);
xor U2446 (N_2446,In_2090,In_2001);
and U2447 (N_2447,In_1843,In_2921);
xnor U2448 (N_2448,In_1114,In_1016);
or U2449 (N_2449,In_929,In_70);
and U2450 (N_2450,In_1288,In_1041);
xor U2451 (N_2451,In_2685,In_2024);
xor U2452 (N_2452,In_2744,In_279);
nor U2453 (N_2453,In_1859,In_722);
and U2454 (N_2454,In_2577,In_1638);
nand U2455 (N_2455,In_2456,In_1687);
nand U2456 (N_2456,In_2132,In_2441);
nor U2457 (N_2457,In_1796,In_2021);
xnor U2458 (N_2458,In_1739,In_653);
nand U2459 (N_2459,In_2791,In_2053);
nand U2460 (N_2460,In_1376,In_257);
nand U2461 (N_2461,In_2501,In_1985);
and U2462 (N_2462,In_730,In_377);
and U2463 (N_2463,In_963,In_110);
or U2464 (N_2464,In_1319,In_2098);
or U2465 (N_2465,In_1946,In_2919);
or U2466 (N_2466,In_2561,In_2696);
nor U2467 (N_2467,In_1780,In_143);
nor U2468 (N_2468,In_1893,In_326);
or U2469 (N_2469,In_70,In_1423);
or U2470 (N_2470,In_2818,In_2266);
xnor U2471 (N_2471,In_1302,In_2519);
nand U2472 (N_2472,In_292,In_615);
or U2473 (N_2473,In_2844,In_2868);
or U2474 (N_2474,In_56,In_294);
nor U2475 (N_2475,In_382,In_2533);
and U2476 (N_2476,In_2344,In_1674);
or U2477 (N_2477,In_66,In_1058);
nand U2478 (N_2478,In_2601,In_257);
xnor U2479 (N_2479,In_1411,In_465);
xor U2480 (N_2480,In_2656,In_131);
xor U2481 (N_2481,In_1937,In_1038);
nand U2482 (N_2482,In_1265,In_2765);
xnor U2483 (N_2483,In_23,In_275);
and U2484 (N_2484,In_2111,In_2839);
nor U2485 (N_2485,In_43,In_1898);
xor U2486 (N_2486,In_2400,In_1212);
and U2487 (N_2487,In_1984,In_1243);
nand U2488 (N_2488,In_413,In_2590);
nand U2489 (N_2489,In_1114,In_115);
xor U2490 (N_2490,In_997,In_1058);
and U2491 (N_2491,In_2375,In_245);
xnor U2492 (N_2492,In_1013,In_1574);
nand U2493 (N_2493,In_2021,In_2883);
nor U2494 (N_2494,In_2038,In_496);
nand U2495 (N_2495,In_747,In_49);
xnor U2496 (N_2496,In_1664,In_1337);
or U2497 (N_2497,In_592,In_1247);
or U2498 (N_2498,In_696,In_1568);
nand U2499 (N_2499,In_1928,In_918);
nand U2500 (N_2500,In_2876,In_1189);
or U2501 (N_2501,In_670,In_1661);
or U2502 (N_2502,In_1567,In_279);
and U2503 (N_2503,In_2414,In_707);
and U2504 (N_2504,In_622,In_2349);
nand U2505 (N_2505,In_602,In_2062);
xnor U2506 (N_2506,In_2164,In_1381);
xnor U2507 (N_2507,In_882,In_1270);
xnor U2508 (N_2508,In_2589,In_99);
xnor U2509 (N_2509,In_1371,In_271);
nand U2510 (N_2510,In_436,In_57);
nor U2511 (N_2511,In_320,In_2805);
or U2512 (N_2512,In_2615,In_160);
nor U2513 (N_2513,In_1401,In_373);
xnor U2514 (N_2514,In_2810,In_1704);
xor U2515 (N_2515,In_632,In_2426);
nand U2516 (N_2516,In_2729,In_1680);
and U2517 (N_2517,In_354,In_1494);
or U2518 (N_2518,In_995,In_70);
xnor U2519 (N_2519,In_1853,In_1811);
nor U2520 (N_2520,In_471,In_1822);
or U2521 (N_2521,In_2522,In_2846);
and U2522 (N_2522,In_1859,In_2238);
xor U2523 (N_2523,In_425,In_797);
nor U2524 (N_2524,In_2863,In_614);
xor U2525 (N_2525,In_1352,In_2483);
nand U2526 (N_2526,In_2074,In_970);
nand U2527 (N_2527,In_2224,In_1806);
nor U2528 (N_2528,In_2720,In_517);
and U2529 (N_2529,In_2214,In_434);
nand U2530 (N_2530,In_502,In_2388);
or U2531 (N_2531,In_2300,In_400);
xor U2532 (N_2532,In_552,In_1927);
nand U2533 (N_2533,In_1278,In_2957);
xnor U2534 (N_2534,In_642,In_2888);
nand U2535 (N_2535,In_1328,In_1995);
or U2536 (N_2536,In_678,In_1501);
xnor U2537 (N_2537,In_2246,In_1518);
nand U2538 (N_2538,In_1929,In_2996);
xor U2539 (N_2539,In_854,In_307);
and U2540 (N_2540,In_2261,In_2066);
xor U2541 (N_2541,In_1943,In_137);
and U2542 (N_2542,In_451,In_2830);
nor U2543 (N_2543,In_1949,In_1706);
nor U2544 (N_2544,In_2744,In_226);
xor U2545 (N_2545,In_1729,In_1291);
or U2546 (N_2546,In_771,In_59);
or U2547 (N_2547,In_365,In_326);
nor U2548 (N_2548,In_1927,In_63);
or U2549 (N_2549,In_604,In_2109);
nor U2550 (N_2550,In_240,In_1613);
and U2551 (N_2551,In_494,In_793);
xor U2552 (N_2552,In_131,In_2505);
nor U2553 (N_2553,In_2780,In_158);
and U2554 (N_2554,In_1249,In_357);
and U2555 (N_2555,In_2973,In_331);
xnor U2556 (N_2556,In_819,In_1461);
nor U2557 (N_2557,In_1443,In_1853);
and U2558 (N_2558,In_1766,In_1170);
and U2559 (N_2559,In_824,In_2455);
and U2560 (N_2560,In_1894,In_1929);
or U2561 (N_2561,In_435,In_846);
nand U2562 (N_2562,In_2964,In_258);
xnor U2563 (N_2563,In_2938,In_2607);
and U2564 (N_2564,In_1646,In_2337);
xor U2565 (N_2565,In_452,In_65);
nor U2566 (N_2566,In_2086,In_1233);
xnor U2567 (N_2567,In_1741,In_1894);
nand U2568 (N_2568,In_2659,In_1161);
nor U2569 (N_2569,In_2878,In_2450);
xnor U2570 (N_2570,In_80,In_2827);
or U2571 (N_2571,In_936,In_2690);
xnor U2572 (N_2572,In_836,In_2027);
or U2573 (N_2573,In_1546,In_2721);
nand U2574 (N_2574,In_1463,In_2031);
xor U2575 (N_2575,In_1016,In_511);
xor U2576 (N_2576,In_1681,In_2139);
or U2577 (N_2577,In_1629,In_764);
xnor U2578 (N_2578,In_1738,In_537);
or U2579 (N_2579,In_1624,In_1898);
nor U2580 (N_2580,In_1695,In_853);
and U2581 (N_2581,In_1045,In_2587);
and U2582 (N_2582,In_2059,In_2073);
xor U2583 (N_2583,In_1019,In_197);
nor U2584 (N_2584,In_2582,In_1489);
nand U2585 (N_2585,In_43,In_2080);
or U2586 (N_2586,In_2772,In_1327);
or U2587 (N_2587,In_1843,In_2217);
xor U2588 (N_2588,In_523,In_2036);
nor U2589 (N_2589,In_482,In_2756);
nor U2590 (N_2590,In_126,In_2325);
or U2591 (N_2591,In_1488,In_1997);
and U2592 (N_2592,In_1117,In_2869);
or U2593 (N_2593,In_2262,In_2864);
and U2594 (N_2594,In_686,In_547);
nor U2595 (N_2595,In_601,In_2482);
nand U2596 (N_2596,In_2228,In_198);
or U2597 (N_2597,In_2305,In_782);
and U2598 (N_2598,In_1166,In_616);
or U2599 (N_2599,In_56,In_1524);
and U2600 (N_2600,In_1317,In_1264);
nor U2601 (N_2601,In_2229,In_299);
nor U2602 (N_2602,In_340,In_1168);
nand U2603 (N_2603,In_2091,In_2959);
nor U2604 (N_2604,In_605,In_1523);
and U2605 (N_2605,In_821,In_1813);
nand U2606 (N_2606,In_1036,In_2612);
xor U2607 (N_2607,In_1995,In_2079);
or U2608 (N_2608,In_309,In_147);
nor U2609 (N_2609,In_1094,In_1344);
nor U2610 (N_2610,In_1386,In_2581);
nor U2611 (N_2611,In_303,In_1624);
nand U2612 (N_2612,In_2459,In_1952);
and U2613 (N_2613,In_2386,In_1345);
or U2614 (N_2614,In_386,In_622);
or U2615 (N_2615,In_1673,In_960);
xnor U2616 (N_2616,In_1193,In_2941);
nand U2617 (N_2617,In_2399,In_2921);
xnor U2618 (N_2618,In_2430,In_229);
and U2619 (N_2619,In_1505,In_564);
and U2620 (N_2620,In_1792,In_1866);
nand U2621 (N_2621,In_222,In_797);
or U2622 (N_2622,In_401,In_1889);
nand U2623 (N_2623,In_1389,In_2500);
and U2624 (N_2624,In_755,In_1628);
nor U2625 (N_2625,In_1325,In_1835);
and U2626 (N_2626,In_678,In_1441);
or U2627 (N_2627,In_118,In_116);
nor U2628 (N_2628,In_2934,In_2049);
nor U2629 (N_2629,In_609,In_1293);
xor U2630 (N_2630,In_1989,In_849);
nand U2631 (N_2631,In_2727,In_752);
nand U2632 (N_2632,In_1687,In_2173);
nor U2633 (N_2633,In_1877,In_2776);
nor U2634 (N_2634,In_806,In_443);
nand U2635 (N_2635,In_1539,In_718);
nor U2636 (N_2636,In_663,In_2431);
nand U2637 (N_2637,In_654,In_298);
nor U2638 (N_2638,In_2748,In_2129);
and U2639 (N_2639,In_2326,In_745);
or U2640 (N_2640,In_2230,In_807);
xor U2641 (N_2641,In_1839,In_1872);
nand U2642 (N_2642,In_1252,In_2294);
nor U2643 (N_2643,In_651,In_1204);
or U2644 (N_2644,In_1903,In_1524);
nor U2645 (N_2645,In_1473,In_2124);
nor U2646 (N_2646,In_1913,In_1150);
or U2647 (N_2647,In_2129,In_787);
nor U2648 (N_2648,In_1063,In_967);
or U2649 (N_2649,In_1874,In_2619);
and U2650 (N_2650,In_1774,In_2603);
nor U2651 (N_2651,In_596,In_2488);
and U2652 (N_2652,In_706,In_1945);
xnor U2653 (N_2653,In_2557,In_2172);
xnor U2654 (N_2654,In_443,In_2754);
xnor U2655 (N_2655,In_900,In_2542);
nor U2656 (N_2656,In_2961,In_2439);
nand U2657 (N_2657,In_2552,In_2713);
or U2658 (N_2658,In_2510,In_362);
nand U2659 (N_2659,In_187,In_1940);
or U2660 (N_2660,In_2747,In_1446);
nor U2661 (N_2661,In_2540,In_336);
nor U2662 (N_2662,In_402,In_1059);
xor U2663 (N_2663,In_1914,In_1310);
nor U2664 (N_2664,In_926,In_1609);
nand U2665 (N_2665,In_2493,In_501);
nand U2666 (N_2666,In_585,In_202);
or U2667 (N_2667,In_2087,In_1034);
xnor U2668 (N_2668,In_2391,In_1920);
or U2669 (N_2669,In_2715,In_1285);
nor U2670 (N_2670,In_2354,In_1738);
xor U2671 (N_2671,In_2462,In_2352);
or U2672 (N_2672,In_476,In_728);
nor U2673 (N_2673,In_160,In_1651);
and U2674 (N_2674,In_418,In_1896);
nor U2675 (N_2675,In_2320,In_992);
nor U2676 (N_2676,In_975,In_2324);
nor U2677 (N_2677,In_2612,In_1617);
or U2678 (N_2678,In_885,In_911);
xnor U2679 (N_2679,In_2027,In_1477);
and U2680 (N_2680,In_649,In_156);
nand U2681 (N_2681,In_589,In_542);
or U2682 (N_2682,In_216,In_2013);
and U2683 (N_2683,In_1817,In_1331);
nand U2684 (N_2684,In_2335,In_560);
and U2685 (N_2685,In_1288,In_1598);
nand U2686 (N_2686,In_2580,In_2117);
nor U2687 (N_2687,In_1794,In_424);
nand U2688 (N_2688,In_1406,In_1515);
and U2689 (N_2689,In_1441,In_1088);
and U2690 (N_2690,In_312,In_1092);
xnor U2691 (N_2691,In_2704,In_2031);
xnor U2692 (N_2692,In_2799,In_2128);
xor U2693 (N_2693,In_2785,In_1633);
nor U2694 (N_2694,In_422,In_2496);
or U2695 (N_2695,In_2335,In_2388);
nor U2696 (N_2696,In_1924,In_869);
nor U2697 (N_2697,In_1700,In_2724);
nand U2698 (N_2698,In_1537,In_359);
or U2699 (N_2699,In_796,In_1443);
nand U2700 (N_2700,In_579,In_148);
nor U2701 (N_2701,In_1583,In_2533);
and U2702 (N_2702,In_2678,In_272);
or U2703 (N_2703,In_884,In_593);
and U2704 (N_2704,In_2771,In_570);
nor U2705 (N_2705,In_670,In_2250);
and U2706 (N_2706,In_1441,In_1287);
nor U2707 (N_2707,In_366,In_2704);
and U2708 (N_2708,In_1910,In_1755);
xnor U2709 (N_2709,In_1373,In_1519);
xnor U2710 (N_2710,In_2597,In_57);
nand U2711 (N_2711,In_1386,In_2517);
and U2712 (N_2712,In_2999,In_1083);
xor U2713 (N_2713,In_2438,In_1272);
xor U2714 (N_2714,In_1981,In_1391);
or U2715 (N_2715,In_2436,In_1019);
or U2716 (N_2716,In_895,In_535);
nand U2717 (N_2717,In_2912,In_1279);
nor U2718 (N_2718,In_2035,In_2562);
nor U2719 (N_2719,In_1781,In_2088);
nor U2720 (N_2720,In_611,In_784);
or U2721 (N_2721,In_2731,In_45);
nand U2722 (N_2722,In_2870,In_1841);
and U2723 (N_2723,In_2979,In_1978);
and U2724 (N_2724,In_2196,In_617);
or U2725 (N_2725,In_2395,In_2706);
or U2726 (N_2726,In_2206,In_1924);
nand U2727 (N_2727,In_2130,In_837);
or U2728 (N_2728,In_1439,In_2276);
or U2729 (N_2729,In_2937,In_1635);
or U2730 (N_2730,In_1002,In_1148);
nor U2731 (N_2731,In_2887,In_1602);
or U2732 (N_2732,In_66,In_1815);
nand U2733 (N_2733,In_1183,In_2493);
nor U2734 (N_2734,In_2734,In_299);
or U2735 (N_2735,In_2153,In_2399);
xor U2736 (N_2736,In_1911,In_1740);
nand U2737 (N_2737,In_2215,In_1217);
xnor U2738 (N_2738,In_594,In_2815);
xor U2739 (N_2739,In_1856,In_2113);
and U2740 (N_2740,In_2975,In_2887);
xnor U2741 (N_2741,In_1875,In_1572);
xor U2742 (N_2742,In_2568,In_2722);
nand U2743 (N_2743,In_2219,In_1601);
nor U2744 (N_2744,In_975,In_2935);
and U2745 (N_2745,In_1498,In_493);
xnor U2746 (N_2746,In_1355,In_298);
and U2747 (N_2747,In_513,In_1489);
or U2748 (N_2748,In_1669,In_1972);
nor U2749 (N_2749,In_2357,In_1938);
or U2750 (N_2750,In_1807,In_967);
nand U2751 (N_2751,In_2527,In_2481);
nand U2752 (N_2752,In_47,In_1616);
nor U2753 (N_2753,In_2426,In_2215);
xnor U2754 (N_2754,In_2393,In_505);
nand U2755 (N_2755,In_2557,In_1685);
nand U2756 (N_2756,In_1107,In_2867);
xnor U2757 (N_2757,In_2662,In_946);
nor U2758 (N_2758,In_1480,In_2418);
nor U2759 (N_2759,In_2862,In_853);
or U2760 (N_2760,In_2063,In_1450);
and U2761 (N_2761,In_2719,In_2334);
xnor U2762 (N_2762,In_1152,In_333);
nor U2763 (N_2763,In_2755,In_2841);
or U2764 (N_2764,In_2241,In_1782);
nand U2765 (N_2765,In_650,In_2012);
nor U2766 (N_2766,In_1696,In_1947);
and U2767 (N_2767,In_2648,In_257);
nor U2768 (N_2768,In_1949,In_1355);
and U2769 (N_2769,In_2294,In_2020);
nand U2770 (N_2770,In_239,In_1021);
xor U2771 (N_2771,In_864,In_812);
or U2772 (N_2772,In_2460,In_227);
or U2773 (N_2773,In_519,In_2732);
or U2774 (N_2774,In_535,In_1229);
nand U2775 (N_2775,In_1223,In_20);
nand U2776 (N_2776,In_1643,In_1858);
nor U2777 (N_2777,In_2486,In_643);
nand U2778 (N_2778,In_444,In_2648);
nor U2779 (N_2779,In_690,In_2311);
and U2780 (N_2780,In_555,In_1147);
and U2781 (N_2781,In_2966,In_2656);
nor U2782 (N_2782,In_2866,In_1452);
and U2783 (N_2783,In_655,In_451);
and U2784 (N_2784,In_2442,In_2972);
or U2785 (N_2785,In_1227,In_1760);
and U2786 (N_2786,In_1049,In_2975);
xor U2787 (N_2787,In_399,In_1023);
nand U2788 (N_2788,In_2644,In_286);
nand U2789 (N_2789,In_1233,In_1138);
xor U2790 (N_2790,In_2663,In_2661);
and U2791 (N_2791,In_1147,In_859);
nor U2792 (N_2792,In_1836,In_2111);
and U2793 (N_2793,In_2833,In_1578);
and U2794 (N_2794,In_1053,In_87);
or U2795 (N_2795,In_1986,In_1860);
or U2796 (N_2796,In_1482,In_114);
nand U2797 (N_2797,In_751,In_789);
xnor U2798 (N_2798,In_1323,In_1093);
nor U2799 (N_2799,In_1929,In_2964);
xor U2800 (N_2800,In_2052,In_568);
and U2801 (N_2801,In_2764,In_936);
nor U2802 (N_2802,In_603,In_1347);
and U2803 (N_2803,In_290,In_413);
and U2804 (N_2804,In_2621,In_1876);
and U2805 (N_2805,In_2790,In_2087);
nor U2806 (N_2806,In_1943,In_1571);
and U2807 (N_2807,In_179,In_2634);
and U2808 (N_2808,In_1737,In_593);
xor U2809 (N_2809,In_667,In_2223);
nor U2810 (N_2810,In_750,In_557);
xor U2811 (N_2811,In_927,In_1167);
xor U2812 (N_2812,In_218,In_1467);
xor U2813 (N_2813,In_2160,In_610);
nor U2814 (N_2814,In_2843,In_866);
nor U2815 (N_2815,In_1655,In_2015);
and U2816 (N_2816,In_295,In_148);
nor U2817 (N_2817,In_1264,In_2333);
xor U2818 (N_2818,In_778,In_1618);
xnor U2819 (N_2819,In_2062,In_696);
or U2820 (N_2820,In_1781,In_1889);
or U2821 (N_2821,In_966,In_777);
xor U2822 (N_2822,In_2197,In_1898);
or U2823 (N_2823,In_2122,In_37);
nand U2824 (N_2824,In_2245,In_825);
or U2825 (N_2825,In_1629,In_673);
nand U2826 (N_2826,In_2542,In_40);
or U2827 (N_2827,In_1975,In_1266);
and U2828 (N_2828,In_2481,In_1115);
nand U2829 (N_2829,In_2115,In_437);
nor U2830 (N_2830,In_2442,In_2610);
xnor U2831 (N_2831,In_694,In_2125);
nor U2832 (N_2832,In_2389,In_439);
nor U2833 (N_2833,In_1730,In_1381);
or U2834 (N_2834,In_2005,In_2616);
and U2835 (N_2835,In_2844,In_2891);
and U2836 (N_2836,In_1417,In_2809);
or U2837 (N_2837,In_1896,In_1893);
and U2838 (N_2838,In_482,In_2586);
nor U2839 (N_2839,In_1343,In_1505);
xor U2840 (N_2840,In_1660,In_1015);
nand U2841 (N_2841,In_1254,In_1620);
xor U2842 (N_2842,In_2341,In_1133);
or U2843 (N_2843,In_1124,In_78);
nor U2844 (N_2844,In_2086,In_1884);
xor U2845 (N_2845,In_619,In_2604);
xnor U2846 (N_2846,In_439,In_377);
or U2847 (N_2847,In_992,In_1726);
nor U2848 (N_2848,In_1388,In_2924);
xor U2849 (N_2849,In_548,In_1251);
nand U2850 (N_2850,In_1584,In_1901);
or U2851 (N_2851,In_2232,In_448);
and U2852 (N_2852,In_2581,In_422);
nand U2853 (N_2853,In_37,In_1028);
nor U2854 (N_2854,In_86,In_2374);
nor U2855 (N_2855,In_511,In_848);
or U2856 (N_2856,In_1685,In_1922);
nor U2857 (N_2857,In_1583,In_2331);
nor U2858 (N_2858,In_2050,In_2696);
or U2859 (N_2859,In_1775,In_1434);
xor U2860 (N_2860,In_1728,In_2823);
nand U2861 (N_2861,In_1270,In_2794);
nor U2862 (N_2862,In_2495,In_787);
nor U2863 (N_2863,In_1378,In_2406);
nor U2864 (N_2864,In_1799,In_86);
or U2865 (N_2865,In_302,In_2786);
xor U2866 (N_2866,In_642,In_2991);
nor U2867 (N_2867,In_1832,In_2231);
nand U2868 (N_2868,In_576,In_1462);
or U2869 (N_2869,In_2123,In_1825);
nand U2870 (N_2870,In_836,In_1903);
or U2871 (N_2871,In_1861,In_1242);
nor U2872 (N_2872,In_2602,In_1664);
nor U2873 (N_2873,In_1190,In_759);
xor U2874 (N_2874,In_2678,In_781);
xor U2875 (N_2875,In_507,In_836);
nand U2876 (N_2876,In_2572,In_2021);
nand U2877 (N_2877,In_1941,In_2129);
xor U2878 (N_2878,In_2855,In_699);
or U2879 (N_2879,In_485,In_2494);
and U2880 (N_2880,In_2517,In_22);
and U2881 (N_2881,In_959,In_620);
and U2882 (N_2882,In_1983,In_740);
nor U2883 (N_2883,In_2715,In_2897);
or U2884 (N_2884,In_79,In_1059);
nor U2885 (N_2885,In_488,In_2781);
nand U2886 (N_2886,In_2767,In_67);
or U2887 (N_2887,In_2467,In_817);
nor U2888 (N_2888,In_518,In_1710);
and U2889 (N_2889,In_495,In_2598);
nand U2890 (N_2890,In_674,In_1201);
or U2891 (N_2891,In_197,In_55);
nor U2892 (N_2892,In_2162,In_216);
xnor U2893 (N_2893,In_1201,In_1090);
or U2894 (N_2894,In_834,In_1931);
xor U2895 (N_2895,In_2994,In_1138);
or U2896 (N_2896,In_2841,In_2722);
nor U2897 (N_2897,In_2731,In_1565);
or U2898 (N_2898,In_1503,In_689);
xor U2899 (N_2899,In_955,In_657);
nand U2900 (N_2900,In_2168,In_2111);
xnor U2901 (N_2901,In_2423,In_2369);
nor U2902 (N_2902,In_863,In_597);
nand U2903 (N_2903,In_1519,In_2140);
nor U2904 (N_2904,In_44,In_1179);
xnor U2905 (N_2905,In_1011,In_584);
nor U2906 (N_2906,In_2163,In_2282);
or U2907 (N_2907,In_153,In_69);
nand U2908 (N_2908,In_551,In_192);
xor U2909 (N_2909,In_1214,In_1399);
and U2910 (N_2910,In_2467,In_1896);
nor U2911 (N_2911,In_872,In_639);
nand U2912 (N_2912,In_693,In_1106);
and U2913 (N_2913,In_0,In_1424);
nand U2914 (N_2914,In_2468,In_1921);
or U2915 (N_2915,In_2874,In_11);
nand U2916 (N_2916,In_824,In_997);
nand U2917 (N_2917,In_1539,In_408);
nand U2918 (N_2918,In_1954,In_2265);
or U2919 (N_2919,In_2854,In_2884);
nor U2920 (N_2920,In_1215,In_1569);
or U2921 (N_2921,In_2859,In_339);
or U2922 (N_2922,In_2444,In_860);
or U2923 (N_2923,In_2907,In_2335);
nand U2924 (N_2924,In_2697,In_1175);
xnor U2925 (N_2925,In_1107,In_1120);
and U2926 (N_2926,In_852,In_871);
xor U2927 (N_2927,In_1143,In_2764);
or U2928 (N_2928,In_323,In_2280);
xnor U2929 (N_2929,In_1164,In_721);
xor U2930 (N_2930,In_444,In_729);
and U2931 (N_2931,In_1668,In_1697);
or U2932 (N_2932,In_2275,In_490);
and U2933 (N_2933,In_302,In_458);
nand U2934 (N_2934,In_2040,In_2159);
or U2935 (N_2935,In_2521,In_2966);
nand U2936 (N_2936,In_2142,In_1891);
nor U2937 (N_2937,In_540,In_1581);
xnor U2938 (N_2938,In_2289,In_305);
nand U2939 (N_2939,In_553,In_1130);
or U2940 (N_2940,In_1153,In_1095);
or U2941 (N_2941,In_1056,In_1450);
nor U2942 (N_2942,In_48,In_696);
nor U2943 (N_2943,In_2543,In_2012);
xor U2944 (N_2944,In_1415,In_1894);
nand U2945 (N_2945,In_2267,In_483);
or U2946 (N_2946,In_612,In_571);
nor U2947 (N_2947,In_411,In_2393);
nand U2948 (N_2948,In_2603,In_2371);
or U2949 (N_2949,In_2376,In_1613);
or U2950 (N_2950,In_1481,In_2479);
nand U2951 (N_2951,In_203,In_221);
nor U2952 (N_2952,In_1603,In_1766);
nand U2953 (N_2953,In_149,In_2430);
nor U2954 (N_2954,In_563,In_2334);
or U2955 (N_2955,In_1966,In_1804);
nor U2956 (N_2956,In_66,In_2268);
nand U2957 (N_2957,In_1986,In_306);
xor U2958 (N_2958,In_1678,In_1889);
nand U2959 (N_2959,In_2074,In_1297);
xnor U2960 (N_2960,In_2638,In_1689);
nand U2961 (N_2961,In_1215,In_453);
and U2962 (N_2962,In_1296,In_1509);
nor U2963 (N_2963,In_1178,In_2827);
or U2964 (N_2964,In_1966,In_1935);
xor U2965 (N_2965,In_1692,In_449);
and U2966 (N_2966,In_2538,In_2286);
or U2967 (N_2967,In_237,In_2396);
or U2968 (N_2968,In_1095,In_1733);
and U2969 (N_2969,In_2921,In_1920);
nor U2970 (N_2970,In_176,In_1952);
xor U2971 (N_2971,In_1313,In_2598);
or U2972 (N_2972,In_128,In_765);
and U2973 (N_2973,In_1441,In_1264);
or U2974 (N_2974,In_1466,In_2152);
and U2975 (N_2975,In_2304,In_2259);
nand U2976 (N_2976,In_2126,In_1364);
nor U2977 (N_2977,In_2797,In_2967);
nor U2978 (N_2978,In_1075,In_1232);
nand U2979 (N_2979,In_1721,In_1520);
nand U2980 (N_2980,In_1371,In_229);
nand U2981 (N_2981,In_383,In_150);
xnor U2982 (N_2982,In_2842,In_1329);
nand U2983 (N_2983,In_2430,In_283);
or U2984 (N_2984,In_1010,In_527);
nand U2985 (N_2985,In_1841,In_1624);
nand U2986 (N_2986,In_2279,In_1046);
nor U2987 (N_2987,In_2293,In_1304);
nor U2988 (N_2988,In_976,In_1211);
and U2989 (N_2989,In_177,In_1136);
nand U2990 (N_2990,In_1700,In_2931);
and U2991 (N_2991,In_2479,In_775);
and U2992 (N_2992,In_2988,In_1119);
xnor U2993 (N_2993,In_2691,In_1122);
xor U2994 (N_2994,In_1187,In_2902);
and U2995 (N_2995,In_1331,In_2012);
nor U2996 (N_2996,In_1408,In_2330);
nand U2997 (N_2997,In_1617,In_2175);
and U2998 (N_2998,In_2192,In_1880);
nand U2999 (N_2999,In_1609,In_904);
nand U3000 (N_3000,In_2666,In_556);
nor U3001 (N_3001,In_1072,In_401);
xnor U3002 (N_3002,In_71,In_2386);
nand U3003 (N_3003,In_2543,In_2298);
and U3004 (N_3004,In_1637,In_428);
nand U3005 (N_3005,In_2048,In_260);
or U3006 (N_3006,In_2641,In_44);
and U3007 (N_3007,In_1763,In_1502);
xor U3008 (N_3008,In_2314,In_358);
and U3009 (N_3009,In_162,In_481);
nand U3010 (N_3010,In_777,In_587);
xor U3011 (N_3011,In_351,In_884);
nor U3012 (N_3012,In_2128,In_2588);
xnor U3013 (N_3013,In_450,In_1969);
nor U3014 (N_3014,In_1868,In_1551);
xnor U3015 (N_3015,In_2538,In_1665);
and U3016 (N_3016,In_172,In_2841);
xnor U3017 (N_3017,In_674,In_2526);
nor U3018 (N_3018,In_2107,In_1018);
xor U3019 (N_3019,In_2642,In_2813);
and U3020 (N_3020,In_2347,In_2166);
and U3021 (N_3021,In_350,In_861);
nand U3022 (N_3022,In_1927,In_240);
and U3023 (N_3023,In_1823,In_684);
and U3024 (N_3024,In_2788,In_1188);
or U3025 (N_3025,In_1340,In_255);
nor U3026 (N_3026,In_1252,In_1159);
and U3027 (N_3027,In_1008,In_2018);
xnor U3028 (N_3028,In_1892,In_467);
nor U3029 (N_3029,In_1812,In_2769);
xnor U3030 (N_3030,In_1226,In_2125);
or U3031 (N_3031,In_277,In_599);
xnor U3032 (N_3032,In_812,In_2234);
or U3033 (N_3033,In_739,In_2974);
and U3034 (N_3034,In_2561,In_227);
and U3035 (N_3035,In_794,In_1277);
or U3036 (N_3036,In_2220,In_2715);
and U3037 (N_3037,In_2536,In_1314);
or U3038 (N_3038,In_1498,In_2202);
or U3039 (N_3039,In_1267,In_753);
or U3040 (N_3040,In_2415,In_1176);
nor U3041 (N_3041,In_2906,In_209);
nor U3042 (N_3042,In_2999,In_2944);
and U3043 (N_3043,In_1242,In_2240);
nor U3044 (N_3044,In_870,In_1950);
and U3045 (N_3045,In_1546,In_2299);
and U3046 (N_3046,In_2551,In_1048);
nand U3047 (N_3047,In_1646,In_653);
nor U3048 (N_3048,In_612,In_359);
xnor U3049 (N_3049,In_571,In_2096);
and U3050 (N_3050,In_1113,In_879);
or U3051 (N_3051,In_2758,In_2901);
nand U3052 (N_3052,In_1825,In_368);
nor U3053 (N_3053,In_936,In_68);
nand U3054 (N_3054,In_1997,In_1436);
nand U3055 (N_3055,In_487,In_2780);
nand U3056 (N_3056,In_671,In_2266);
nand U3057 (N_3057,In_1481,In_491);
or U3058 (N_3058,In_2032,In_2425);
and U3059 (N_3059,In_1014,In_2361);
and U3060 (N_3060,In_1094,In_1022);
nor U3061 (N_3061,In_1731,In_184);
nor U3062 (N_3062,In_420,In_1838);
nand U3063 (N_3063,In_2859,In_2714);
and U3064 (N_3064,In_1466,In_2508);
or U3065 (N_3065,In_1647,In_834);
nor U3066 (N_3066,In_1239,In_2038);
or U3067 (N_3067,In_820,In_1430);
or U3068 (N_3068,In_1032,In_769);
nor U3069 (N_3069,In_2923,In_2984);
or U3070 (N_3070,In_2516,In_1954);
or U3071 (N_3071,In_2508,In_2990);
nand U3072 (N_3072,In_2649,In_1730);
xor U3073 (N_3073,In_1157,In_1277);
nor U3074 (N_3074,In_2185,In_701);
or U3075 (N_3075,In_544,In_1302);
nand U3076 (N_3076,In_1250,In_1163);
xor U3077 (N_3077,In_1992,In_2711);
and U3078 (N_3078,In_1173,In_344);
and U3079 (N_3079,In_1749,In_1372);
or U3080 (N_3080,In_749,In_2990);
and U3081 (N_3081,In_2825,In_2031);
xnor U3082 (N_3082,In_933,In_2300);
xor U3083 (N_3083,In_102,In_82);
or U3084 (N_3084,In_1958,In_1648);
nor U3085 (N_3085,In_1476,In_337);
nor U3086 (N_3086,In_71,In_2164);
nor U3087 (N_3087,In_680,In_1131);
or U3088 (N_3088,In_187,In_2248);
xnor U3089 (N_3089,In_2393,In_1042);
xor U3090 (N_3090,In_1145,In_1289);
nand U3091 (N_3091,In_2034,In_1246);
or U3092 (N_3092,In_842,In_2135);
nor U3093 (N_3093,In_1398,In_1030);
xnor U3094 (N_3094,In_1247,In_912);
or U3095 (N_3095,In_1737,In_1568);
and U3096 (N_3096,In_111,In_2831);
nor U3097 (N_3097,In_1187,In_1516);
and U3098 (N_3098,In_1925,In_439);
xor U3099 (N_3099,In_2114,In_1403);
and U3100 (N_3100,In_227,In_1045);
xnor U3101 (N_3101,In_129,In_277);
nand U3102 (N_3102,In_1639,In_1073);
nand U3103 (N_3103,In_128,In_241);
or U3104 (N_3104,In_1214,In_1228);
nand U3105 (N_3105,In_2965,In_220);
nand U3106 (N_3106,In_2155,In_1365);
and U3107 (N_3107,In_937,In_711);
and U3108 (N_3108,In_872,In_2680);
and U3109 (N_3109,In_1923,In_811);
xnor U3110 (N_3110,In_1222,In_1492);
or U3111 (N_3111,In_660,In_1390);
or U3112 (N_3112,In_2631,In_437);
and U3113 (N_3113,In_1106,In_2130);
and U3114 (N_3114,In_1367,In_703);
and U3115 (N_3115,In_78,In_977);
or U3116 (N_3116,In_740,In_792);
xor U3117 (N_3117,In_2830,In_2518);
and U3118 (N_3118,In_2897,In_2476);
nand U3119 (N_3119,In_2369,In_14);
xnor U3120 (N_3120,In_1252,In_2187);
xnor U3121 (N_3121,In_862,In_1356);
and U3122 (N_3122,In_128,In_2571);
nand U3123 (N_3123,In_2978,In_2968);
or U3124 (N_3124,In_1038,In_706);
nor U3125 (N_3125,In_86,In_457);
or U3126 (N_3126,In_667,In_1144);
or U3127 (N_3127,In_2131,In_1476);
xnor U3128 (N_3128,In_634,In_505);
nand U3129 (N_3129,In_1856,In_2409);
or U3130 (N_3130,In_913,In_930);
xnor U3131 (N_3131,In_292,In_1826);
nand U3132 (N_3132,In_754,In_565);
nor U3133 (N_3133,In_1867,In_280);
nor U3134 (N_3134,In_2781,In_1862);
nand U3135 (N_3135,In_1776,In_846);
nand U3136 (N_3136,In_1619,In_1579);
nor U3137 (N_3137,In_2067,In_2877);
nor U3138 (N_3138,In_728,In_2768);
and U3139 (N_3139,In_601,In_1858);
and U3140 (N_3140,In_2846,In_674);
nand U3141 (N_3141,In_2778,In_2419);
xnor U3142 (N_3142,In_2503,In_192);
or U3143 (N_3143,In_375,In_2413);
or U3144 (N_3144,In_333,In_365);
and U3145 (N_3145,In_514,In_2059);
xor U3146 (N_3146,In_2343,In_363);
xor U3147 (N_3147,In_1248,In_2428);
nor U3148 (N_3148,In_13,In_1884);
nor U3149 (N_3149,In_1421,In_1630);
nand U3150 (N_3150,In_2946,In_990);
nor U3151 (N_3151,In_1173,In_1276);
nand U3152 (N_3152,In_1817,In_137);
xor U3153 (N_3153,In_2808,In_2351);
nor U3154 (N_3154,In_1685,In_776);
xor U3155 (N_3155,In_2940,In_850);
nor U3156 (N_3156,In_303,In_108);
xnor U3157 (N_3157,In_830,In_351);
xor U3158 (N_3158,In_645,In_371);
and U3159 (N_3159,In_1466,In_2630);
xnor U3160 (N_3160,In_936,In_1017);
nand U3161 (N_3161,In_2678,In_1294);
nor U3162 (N_3162,In_341,In_1064);
xor U3163 (N_3163,In_2988,In_1283);
nand U3164 (N_3164,In_2906,In_1443);
and U3165 (N_3165,In_88,In_1785);
nand U3166 (N_3166,In_2351,In_562);
nor U3167 (N_3167,In_160,In_546);
or U3168 (N_3168,In_615,In_2985);
and U3169 (N_3169,In_2463,In_1818);
and U3170 (N_3170,In_341,In_1866);
xnor U3171 (N_3171,In_2527,In_392);
nand U3172 (N_3172,In_2568,In_1898);
nand U3173 (N_3173,In_417,In_2848);
nand U3174 (N_3174,In_1040,In_1167);
or U3175 (N_3175,In_2313,In_1895);
or U3176 (N_3176,In_2145,In_401);
or U3177 (N_3177,In_1679,In_2225);
and U3178 (N_3178,In_2104,In_1892);
or U3179 (N_3179,In_639,In_2903);
nand U3180 (N_3180,In_1056,In_2958);
or U3181 (N_3181,In_2869,In_1894);
nand U3182 (N_3182,In_2334,In_1010);
nand U3183 (N_3183,In_458,In_117);
or U3184 (N_3184,In_1275,In_2126);
nor U3185 (N_3185,In_1679,In_1223);
or U3186 (N_3186,In_28,In_2057);
nor U3187 (N_3187,In_2606,In_2811);
or U3188 (N_3188,In_496,In_2117);
nor U3189 (N_3189,In_452,In_551);
nor U3190 (N_3190,In_1865,In_1228);
and U3191 (N_3191,In_2744,In_2246);
and U3192 (N_3192,In_120,In_2141);
nor U3193 (N_3193,In_1674,In_2050);
nor U3194 (N_3194,In_2409,In_1062);
and U3195 (N_3195,In_879,In_1664);
nor U3196 (N_3196,In_2401,In_2156);
and U3197 (N_3197,In_2956,In_426);
or U3198 (N_3198,In_1024,In_2208);
xnor U3199 (N_3199,In_2762,In_458);
nand U3200 (N_3200,In_2351,In_93);
nand U3201 (N_3201,In_1830,In_906);
nand U3202 (N_3202,In_2814,In_78);
and U3203 (N_3203,In_469,In_1100);
or U3204 (N_3204,In_2639,In_2833);
or U3205 (N_3205,In_1700,In_262);
nor U3206 (N_3206,In_1320,In_410);
or U3207 (N_3207,In_2957,In_1147);
and U3208 (N_3208,In_2292,In_381);
nand U3209 (N_3209,In_2626,In_2693);
and U3210 (N_3210,In_33,In_1919);
or U3211 (N_3211,In_238,In_558);
or U3212 (N_3212,In_14,In_1963);
xor U3213 (N_3213,In_1552,In_2221);
or U3214 (N_3214,In_416,In_2749);
nand U3215 (N_3215,In_1618,In_1162);
nor U3216 (N_3216,In_60,In_2189);
nor U3217 (N_3217,In_119,In_2651);
nand U3218 (N_3218,In_1120,In_72);
xor U3219 (N_3219,In_2162,In_1278);
or U3220 (N_3220,In_2832,In_2784);
and U3221 (N_3221,In_2988,In_1295);
and U3222 (N_3222,In_1290,In_266);
and U3223 (N_3223,In_66,In_1526);
nand U3224 (N_3224,In_497,In_1340);
and U3225 (N_3225,In_199,In_1765);
or U3226 (N_3226,In_2672,In_1287);
and U3227 (N_3227,In_223,In_359);
nand U3228 (N_3228,In_1002,In_2002);
xnor U3229 (N_3229,In_1617,In_1055);
xor U3230 (N_3230,In_1243,In_550);
xor U3231 (N_3231,In_2727,In_616);
and U3232 (N_3232,In_1948,In_1046);
xor U3233 (N_3233,In_2536,In_2719);
nor U3234 (N_3234,In_1899,In_1920);
and U3235 (N_3235,In_1683,In_160);
nor U3236 (N_3236,In_2764,In_2342);
xor U3237 (N_3237,In_1209,In_2844);
or U3238 (N_3238,In_1553,In_1495);
nand U3239 (N_3239,In_2904,In_2642);
nand U3240 (N_3240,In_2107,In_1156);
nor U3241 (N_3241,In_1498,In_1400);
and U3242 (N_3242,In_2101,In_2284);
nor U3243 (N_3243,In_726,In_1077);
or U3244 (N_3244,In_2625,In_1446);
xnor U3245 (N_3245,In_1982,In_116);
nand U3246 (N_3246,In_2309,In_2212);
nor U3247 (N_3247,In_568,In_1719);
xor U3248 (N_3248,In_2791,In_1394);
or U3249 (N_3249,In_514,In_205);
nand U3250 (N_3250,In_436,In_2150);
nand U3251 (N_3251,In_50,In_2645);
and U3252 (N_3252,In_2475,In_1059);
nand U3253 (N_3253,In_2449,In_23);
nand U3254 (N_3254,In_2009,In_290);
or U3255 (N_3255,In_68,In_778);
nor U3256 (N_3256,In_1288,In_1764);
or U3257 (N_3257,In_690,In_2610);
nand U3258 (N_3258,In_1879,In_1855);
nor U3259 (N_3259,In_2352,In_1392);
nor U3260 (N_3260,In_2412,In_674);
or U3261 (N_3261,In_195,In_1588);
nand U3262 (N_3262,In_696,In_1270);
nor U3263 (N_3263,In_2734,In_2689);
or U3264 (N_3264,In_2283,In_1935);
and U3265 (N_3265,In_207,In_1389);
xnor U3266 (N_3266,In_2512,In_132);
nand U3267 (N_3267,In_2049,In_2267);
nand U3268 (N_3268,In_171,In_14);
nor U3269 (N_3269,In_2515,In_1042);
nand U3270 (N_3270,In_1299,In_366);
and U3271 (N_3271,In_1583,In_820);
nand U3272 (N_3272,In_862,In_776);
or U3273 (N_3273,In_1581,In_2299);
nor U3274 (N_3274,In_2947,In_2166);
nand U3275 (N_3275,In_2080,In_1430);
nor U3276 (N_3276,In_1894,In_2212);
and U3277 (N_3277,In_2859,In_1900);
nor U3278 (N_3278,In_2975,In_489);
xor U3279 (N_3279,In_162,In_215);
nand U3280 (N_3280,In_2667,In_430);
and U3281 (N_3281,In_812,In_1199);
and U3282 (N_3282,In_1120,In_1077);
or U3283 (N_3283,In_899,In_671);
nor U3284 (N_3284,In_1548,In_2350);
nand U3285 (N_3285,In_788,In_665);
and U3286 (N_3286,In_579,In_1587);
xor U3287 (N_3287,In_2515,In_1944);
nand U3288 (N_3288,In_1915,In_513);
nor U3289 (N_3289,In_307,In_2216);
or U3290 (N_3290,In_1234,In_591);
nand U3291 (N_3291,In_2370,In_2838);
or U3292 (N_3292,In_1886,In_1674);
nor U3293 (N_3293,In_2165,In_616);
nand U3294 (N_3294,In_2768,In_1644);
xnor U3295 (N_3295,In_2554,In_1958);
and U3296 (N_3296,In_2581,In_2738);
or U3297 (N_3297,In_2407,In_1326);
xnor U3298 (N_3298,In_476,In_257);
nand U3299 (N_3299,In_2191,In_1739);
nand U3300 (N_3300,In_2993,In_2269);
or U3301 (N_3301,In_2368,In_1683);
and U3302 (N_3302,In_2091,In_2736);
nand U3303 (N_3303,In_88,In_460);
nand U3304 (N_3304,In_2994,In_1546);
nand U3305 (N_3305,In_1487,In_1453);
or U3306 (N_3306,In_1381,In_2362);
and U3307 (N_3307,In_1851,In_699);
xnor U3308 (N_3308,In_2183,In_115);
nor U3309 (N_3309,In_425,In_2755);
xor U3310 (N_3310,In_285,In_406);
or U3311 (N_3311,In_1302,In_2056);
and U3312 (N_3312,In_1289,In_1974);
nand U3313 (N_3313,In_1095,In_1313);
xnor U3314 (N_3314,In_405,In_2477);
nor U3315 (N_3315,In_1146,In_2084);
and U3316 (N_3316,In_2745,In_1684);
or U3317 (N_3317,In_83,In_1218);
or U3318 (N_3318,In_1437,In_2075);
nor U3319 (N_3319,In_2109,In_2505);
nand U3320 (N_3320,In_990,In_2032);
nand U3321 (N_3321,In_1370,In_2109);
xor U3322 (N_3322,In_738,In_342);
xor U3323 (N_3323,In_1635,In_871);
nand U3324 (N_3324,In_1916,In_1177);
or U3325 (N_3325,In_902,In_1056);
and U3326 (N_3326,In_1776,In_2795);
xnor U3327 (N_3327,In_1742,In_2098);
xor U3328 (N_3328,In_2497,In_2796);
and U3329 (N_3329,In_696,In_2138);
xor U3330 (N_3330,In_916,In_1957);
and U3331 (N_3331,In_2506,In_763);
xnor U3332 (N_3332,In_444,In_2383);
xor U3333 (N_3333,In_130,In_1273);
or U3334 (N_3334,In_1206,In_2686);
xor U3335 (N_3335,In_2837,In_1032);
nor U3336 (N_3336,In_418,In_1782);
and U3337 (N_3337,In_1850,In_85);
nand U3338 (N_3338,In_2200,In_1461);
nand U3339 (N_3339,In_2710,In_2318);
xor U3340 (N_3340,In_2587,In_2467);
or U3341 (N_3341,In_1015,In_1503);
nand U3342 (N_3342,In_292,In_1334);
or U3343 (N_3343,In_2081,In_1770);
and U3344 (N_3344,In_320,In_1014);
nand U3345 (N_3345,In_2464,In_2584);
or U3346 (N_3346,In_766,In_1742);
nor U3347 (N_3347,In_1828,In_708);
and U3348 (N_3348,In_2323,In_1638);
nand U3349 (N_3349,In_2309,In_496);
nand U3350 (N_3350,In_1857,In_1032);
and U3351 (N_3351,In_1837,In_2870);
xnor U3352 (N_3352,In_1203,In_209);
nand U3353 (N_3353,In_1249,In_2372);
xor U3354 (N_3354,In_1427,In_2515);
xnor U3355 (N_3355,In_1319,In_72);
or U3356 (N_3356,In_2404,In_1961);
nand U3357 (N_3357,In_2224,In_2132);
nand U3358 (N_3358,In_1508,In_1502);
and U3359 (N_3359,In_727,In_457);
or U3360 (N_3360,In_2710,In_185);
nor U3361 (N_3361,In_817,In_1461);
or U3362 (N_3362,In_1585,In_2950);
and U3363 (N_3363,In_249,In_839);
nand U3364 (N_3364,In_2364,In_2566);
nand U3365 (N_3365,In_2277,In_922);
nand U3366 (N_3366,In_2662,In_2396);
or U3367 (N_3367,In_774,In_2223);
or U3368 (N_3368,In_2792,In_1997);
or U3369 (N_3369,In_2392,In_1134);
nor U3370 (N_3370,In_1477,In_1593);
or U3371 (N_3371,In_1260,In_856);
nand U3372 (N_3372,In_2880,In_117);
nand U3373 (N_3373,In_604,In_2790);
xnor U3374 (N_3374,In_814,In_1733);
or U3375 (N_3375,In_1731,In_738);
xor U3376 (N_3376,In_2602,In_83);
nor U3377 (N_3377,In_1840,In_522);
nand U3378 (N_3378,In_942,In_220);
xor U3379 (N_3379,In_892,In_543);
xnor U3380 (N_3380,In_2967,In_65);
xor U3381 (N_3381,In_2689,In_2445);
xnor U3382 (N_3382,In_2269,In_1532);
nor U3383 (N_3383,In_2314,In_509);
and U3384 (N_3384,In_2931,In_248);
and U3385 (N_3385,In_2374,In_1962);
and U3386 (N_3386,In_2092,In_336);
and U3387 (N_3387,In_2749,In_2110);
nand U3388 (N_3388,In_2477,In_111);
nand U3389 (N_3389,In_2361,In_1866);
or U3390 (N_3390,In_2958,In_138);
nand U3391 (N_3391,In_2132,In_1445);
xor U3392 (N_3392,In_925,In_2136);
nand U3393 (N_3393,In_835,In_2200);
nor U3394 (N_3394,In_1505,In_179);
and U3395 (N_3395,In_42,In_16);
or U3396 (N_3396,In_2704,In_1754);
nor U3397 (N_3397,In_1639,In_1574);
nand U3398 (N_3398,In_515,In_1027);
or U3399 (N_3399,In_903,In_733);
xor U3400 (N_3400,In_1949,In_786);
xor U3401 (N_3401,In_1301,In_1623);
or U3402 (N_3402,In_578,In_32);
nor U3403 (N_3403,In_2666,In_2399);
xnor U3404 (N_3404,In_840,In_2119);
or U3405 (N_3405,In_1854,In_922);
nor U3406 (N_3406,In_1565,In_2297);
nand U3407 (N_3407,In_1224,In_2704);
and U3408 (N_3408,In_2860,In_2103);
or U3409 (N_3409,In_1756,In_816);
xnor U3410 (N_3410,In_2606,In_1808);
or U3411 (N_3411,In_1904,In_59);
and U3412 (N_3412,In_2333,In_2161);
or U3413 (N_3413,In_590,In_1509);
and U3414 (N_3414,In_2645,In_879);
xnor U3415 (N_3415,In_68,In_770);
or U3416 (N_3416,In_2137,In_2052);
nand U3417 (N_3417,In_426,In_467);
nor U3418 (N_3418,In_1310,In_1039);
and U3419 (N_3419,In_694,In_2265);
xnor U3420 (N_3420,In_2334,In_2216);
or U3421 (N_3421,In_2132,In_231);
xor U3422 (N_3422,In_711,In_2310);
xor U3423 (N_3423,In_2535,In_2436);
nand U3424 (N_3424,In_613,In_77);
xor U3425 (N_3425,In_185,In_887);
or U3426 (N_3426,In_1929,In_2369);
xor U3427 (N_3427,In_2512,In_2579);
or U3428 (N_3428,In_229,In_1148);
nor U3429 (N_3429,In_423,In_2475);
nand U3430 (N_3430,In_2596,In_214);
or U3431 (N_3431,In_789,In_819);
xor U3432 (N_3432,In_560,In_1188);
xor U3433 (N_3433,In_1158,In_1744);
xor U3434 (N_3434,In_2102,In_449);
or U3435 (N_3435,In_2672,In_370);
nor U3436 (N_3436,In_2814,In_973);
nand U3437 (N_3437,In_901,In_965);
and U3438 (N_3438,In_885,In_146);
or U3439 (N_3439,In_2298,In_870);
xnor U3440 (N_3440,In_915,In_1630);
xor U3441 (N_3441,In_2026,In_354);
or U3442 (N_3442,In_2930,In_2973);
nor U3443 (N_3443,In_2302,In_2753);
or U3444 (N_3444,In_2025,In_678);
xnor U3445 (N_3445,In_2942,In_2364);
or U3446 (N_3446,In_1059,In_2344);
nor U3447 (N_3447,In_2347,In_1050);
nand U3448 (N_3448,In_2980,In_80);
nand U3449 (N_3449,In_1122,In_732);
nor U3450 (N_3450,In_2650,In_1071);
nand U3451 (N_3451,In_1938,In_2478);
nor U3452 (N_3452,In_1838,In_773);
or U3453 (N_3453,In_927,In_865);
and U3454 (N_3454,In_46,In_2418);
nand U3455 (N_3455,In_1659,In_1805);
nand U3456 (N_3456,In_1494,In_1024);
xor U3457 (N_3457,In_483,In_1030);
or U3458 (N_3458,In_23,In_652);
nor U3459 (N_3459,In_525,In_1191);
or U3460 (N_3460,In_1474,In_887);
nand U3461 (N_3461,In_1564,In_245);
nor U3462 (N_3462,In_474,In_1821);
or U3463 (N_3463,In_1842,In_1498);
nand U3464 (N_3464,In_1982,In_2238);
or U3465 (N_3465,In_2392,In_657);
xor U3466 (N_3466,In_2129,In_923);
nor U3467 (N_3467,In_2415,In_2629);
and U3468 (N_3468,In_1619,In_1763);
and U3469 (N_3469,In_2842,In_1548);
and U3470 (N_3470,In_540,In_2996);
or U3471 (N_3471,In_705,In_767);
and U3472 (N_3472,In_349,In_235);
and U3473 (N_3473,In_1402,In_2015);
nand U3474 (N_3474,In_2976,In_1556);
nor U3475 (N_3475,In_1755,In_508);
nor U3476 (N_3476,In_2467,In_2488);
xnor U3477 (N_3477,In_364,In_1741);
xor U3478 (N_3478,In_106,In_2126);
nand U3479 (N_3479,In_1494,In_2761);
nand U3480 (N_3480,In_593,In_292);
and U3481 (N_3481,In_1663,In_2340);
xor U3482 (N_3482,In_2200,In_451);
nand U3483 (N_3483,In_2408,In_1519);
nand U3484 (N_3484,In_1613,In_813);
nor U3485 (N_3485,In_1719,In_1357);
nand U3486 (N_3486,In_1158,In_2674);
nor U3487 (N_3487,In_2910,In_451);
nand U3488 (N_3488,In_2059,In_12);
xnor U3489 (N_3489,In_1089,In_1539);
or U3490 (N_3490,In_2087,In_1721);
and U3491 (N_3491,In_659,In_388);
xor U3492 (N_3492,In_129,In_1096);
xor U3493 (N_3493,In_2471,In_2769);
or U3494 (N_3494,In_2326,In_2953);
nand U3495 (N_3495,In_578,In_1589);
or U3496 (N_3496,In_981,In_1177);
and U3497 (N_3497,In_2966,In_648);
nor U3498 (N_3498,In_2405,In_2004);
nand U3499 (N_3499,In_1377,In_429);
nor U3500 (N_3500,In_2156,In_2172);
or U3501 (N_3501,In_2963,In_1889);
and U3502 (N_3502,In_1714,In_1693);
or U3503 (N_3503,In_2108,In_2796);
nor U3504 (N_3504,In_1393,In_1845);
xor U3505 (N_3505,In_391,In_2667);
nand U3506 (N_3506,In_2287,In_2115);
nor U3507 (N_3507,In_1620,In_1726);
nand U3508 (N_3508,In_1276,In_2497);
and U3509 (N_3509,In_2339,In_1845);
nor U3510 (N_3510,In_1508,In_2678);
and U3511 (N_3511,In_2992,In_1395);
xor U3512 (N_3512,In_1861,In_1899);
xor U3513 (N_3513,In_403,In_818);
and U3514 (N_3514,In_2940,In_134);
and U3515 (N_3515,In_1314,In_773);
nand U3516 (N_3516,In_1065,In_2372);
and U3517 (N_3517,In_1839,In_2637);
or U3518 (N_3518,In_1579,In_1449);
and U3519 (N_3519,In_2862,In_477);
xor U3520 (N_3520,In_296,In_853);
or U3521 (N_3521,In_2883,In_901);
or U3522 (N_3522,In_555,In_283);
xnor U3523 (N_3523,In_2566,In_1596);
and U3524 (N_3524,In_748,In_2698);
nand U3525 (N_3525,In_632,In_590);
and U3526 (N_3526,In_730,In_204);
nand U3527 (N_3527,In_1355,In_473);
or U3528 (N_3528,In_1955,In_1798);
or U3529 (N_3529,In_819,In_1736);
nand U3530 (N_3530,In_1048,In_932);
nand U3531 (N_3531,In_1952,In_216);
and U3532 (N_3532,In_2157,In_2601);
or U3533 (N_3533,In_2482,In_1630);
nand U3534 (N_3534,In_670,In_246);
and U3535 (N_3535,In_1771,In_1089);
or U3536 (N_3536,In_472,In_1490);
xnor U3537 (N_3537,In_1036,In_2375);
xnor U3538 (N_3538,In_1012,In_833);
and U3539 (N_3539,In_1134,In_37);
and U3540 (N_3540,In_986,In_99);
or U3541 (N_3541,In_2545,In_1521);
xor U3542 (N_3542,In_2492,In_1679);
or U3543 (N_3543,In_1709,In_1725);
xor U3544 (N_3544,In_1911,In_2526);
nand U3545 (N_3545,In_1872,In_2261);
nor U3546 (N_3546,In_2835,In_2416);
nor U3547 (N_3547,In_1557,In_2872);
or U3548 (N_3548,In_481,In_1321);
nor U3549 (N_3549,In_1216,In_664);
nand U3550 (N_3550,In_2830,In_1034);
nor U3551 (N_3551,In_2510,In_882);
nor U3552 (N_3552,In_1190,In_2060);
and U3553 (N_3553,In_2558,In_231);
xor U3554 (N_3554,In_936,In_2129);
xor U3555 (N_3555,In_2460,In_1725);
nor U3556 (N_3556,In_348,In_2897);
xor U3557 (N_3557,In_1369,In_225);
xor U3558 (N_3558,In_2974,In_2466);
nand U3559 (N_3559,In_2897,In_1383);
nand U3560 (N_3560,In_2730,In_754);
xnor U3561 (N_3561,In_2692,In_2909);
or U3562 (N_3562,In_1888,In_2173);
nor U3563 (N_3563,In_2847,In_1901);
xnor U3564 (N_3564,In_1150,In_1730);
nor U3565 (N_3565,In_1842,In_1297);
and U3566 (N_3566,In_2201,In_1571);
or U3567 (N_3567,In_2032,In_1859);
nor U3568 (N_3568,In_2792,In_2433);
nand U3569 (N_3569,In_371,In_2921);
nor U3570 (N_3570,In_2291,In_1558);
nand U3571 (N_3571,In_1435,In_1107);
xnor U3572 (N_3572,In_492,In_840);
nand U3573 (N_3573,In_1990,In_2514);
xor U3574 (N_3574,In_1117,In_287);
xnor U3575 (N_3575,In_1452,In_988);
nand U3576 (N_3576,In_1418,In_1268);
nor U3577 (N_3577,In_947,In_2870);
and U3578 (N_3578,In_1873,In_2927);
or U3579 (N_3579,In_1215,In_1148);
nand U3580 (N_3580,In_1919,In_2501);
nand U3581 (N_3581,In_51,In_1671);
nor U3582 (N_3582,In_2271,In_267);
and U3583 (N_3583,In_2259,In_2429);
or U3584 (N_3584,In_1265,In_2265);
nor U3585 (N_3585,In_2781,In_461);
nand U3586 (N_3586,In_64,In_2314);
xor U3587 (N_3587,In_2373,In_2343);
nor U3588 (N_3588,In_946,In_532);
or U3589 (N_3589,In_2594,In_2842);
or U3590 (N_3590,In_2380,In_2421);
nor U3591 (N_3591,In_876,In_158);
nor U3592 (N_3592,In_513,In_2166);
nand U3593 (N_3593,In_302,In_560);
nor U3594 (N_3594,In_1277,In_1017);
xnor U3595 (N_3595,In_1285,In_476);
nor U3596 (N_3596,In_834,In_301);
nor U3597 (N_3597,In_2647,In_2076);
or U3598 (N_3598,In_1782,In_1453);
and U3599 (N_3599,In_2982,In_474);
and U3600 (N_3600,In_751,In_11);
xor U3601 (N_3601,In_269,In_1775);
xor U3602 (N_3602,In_1316,In_2992);
nand U3603 (N_3603,In_2471,In_1958);
xor U3604 (N_3604,In_581,In_2961);
and U3605 (N_3605,In_1434,In_1886);
or U3606 (N_3606,In_1804,In_1354);
nor U3607 (N_3607,In_1357,In_1636);
nand U3608 (N_3608,In_1904,In_462);
and U3609 (N_3609,In_2890,In_538);
and U3610 (N_3610,In_1858,In_2041);
nor U3611 (N_3611,In_1270,In_2249);
xnor U3612 (N_3612,In_716,In_1948);
nor U3613 (N_3613,In_829,In_1999);
xnor U3614 (N_3614,In_790,In_53);
and U3615 (N_3615,In_216,In_594);
nor U3616 (N_3616,In_1381,In_120);
xnor U3617 (N_3617,In_2911,In_1992);
or U3618 (N_3618,In_1437,In_381);
xor U3619 (N_3619,In_1388,In_234);
nand U3620 (N_3620,In_1995,In_1163);
xnor U3621 (N_3621,In_1340,In_1948);
or U3622 (N_3622,In_227,In_605);
nor U3623 (N_3623,In_2713,In_2534);
nor U3624 (N_3624,In_700,In_184);
nand U3625 (N_3625,In_2878,In_549);
xor U3626 (N_3626,In_2672,In_970);
xnor U3627 (N_3627,In_2072,In_1725);
nand U3628 (N_3628,In_1394,In_2472);
and U3629 (N_3629,In_2404,In_158);
nor U3630 (N_3630,In_1274,In_438);
and U3631 (N_3631,In_2081,In_2031);
xnor U3632 (N_3632,In_2693,In_1669);
xor U3633 (N_3633,In_1936,In_1310);
and U3634 (N_3634,In_1326,In_1943);
and U3635 (N_3635,In_402,In_635);
nand U3636 (N_3636,In_290,In_1404);
nand U3637 (N_3637,In_2954,In_2838);
nand U3638 (N_3638,In_930,In_2614);
xor U3639 (N_3639,In_1597,In_883);
nand U3640 (N_3640,In_399,In_1497);
xnor U3641 (N_3641,In_2767,In_2122);
or U3642 (N_3642,In_358,In_445);
xnor U3643 (N_3643,In_1972,In_839);
or U3644 (N_3644,In_2225,In_2271);
or U3645 (N_3645,In_1897,In_2652);
xor U3646 (N_3646,In_921,In_1096);
and U3647 (N_3647,In_2342,In_1561);
nor U3648 (N_3648,In_1468,In_2312);
nor U3649 (N_3649,In_2040,In_625);
xor U3650 (N_3650,In_1326,In_555);
and U3651 (N_3651,In_1287,In_2770);
or U3652 (N_3652,In_2870,In_2431);
nor U3653 (N_3653,In_1019,In_759);
or U3654 (N_3654,In_328,In_1426);
nor U3655 (N_3655,In_1455,In_2193);
and U3656 (N_3656,In_2482,In_2290);
and U3657 (N_3657,In_570,In_1167);
or U3658 (N_3658,In_2579,In_2618);
or U3659 (N_3659,In_1362,In_263);
xnor U3660 (N_3660,In_2663,In_1091);
and U3661 (N_3661,In_2496,In_2730);
nand U3662 (N_3662,In_1784,In_1798);
and U3663 (N_3663,In_2080,In_2555);
nand U3664 (N_3664,In_2849,In_359);
nand U3665 (N_3665,In_1706,In_1674);
and U3666 (N_3666,In_499,In_718);
xor U3667 (N_3667,In_647,In_273);
nand U3668 (N_3668,In_2852,In_454);
xor U3669 (N_3669,In_1717,In_2881);
xnor U3670 (N_3670,In_243,In_1953);
and U3671 (N_3671,In_2744,In_1290);
and U3672 (N_3672,In_956,In_1404);
nor U3673 (N_3673,In_1420,In_1887);
nand U3674 (N_3674,In_1138,In_422);
nor U3675 (N_3675,In_1734,In_1984);
nor U3676 (N_3676,In_2205,In_2085);
and U3677 (N_3677,In_2346,In_80);
nand U3678 (N_3678,In_605,In_2574);
and U3679 (N_3679,In_540,In_804);
xnor U3680 (N_3680,In_1981,In_408);
nor U3681 (N_3681,In_2330,In_1659);
or U3682 (N_3682,In_2730,In_66);
nor U3683 (N_3683,In_1053,In_2014);
or U3684 (N_3684,In_1087,In_2406);
nand U3685 (N_3685,In_2247,In_527);
or U3686 (N_3686,In_2330,In_1423);
or U3687 (N_3687,In_2821,In_1614);
xor U3688 (N_3688,In_674,In_591);
and U3689 (N_3689,In_2854,In_2141);
nand U3690 (N_3690,In_978,In_1538);
nand U3691 (N_3691,In_2896,In_1451);
or U3692 (N_3692,In_2973,In_1508);
nand U3693 (N_3693,In_601,In_1915);
nand U3694 (N_3694,In_2625,In_952);
nand U3695 (N_3695,In_88,In_564);
xnor U3696 (N_3696,In_1783,In_1271);
nor U3697 (N_3697,In_992,In_2121);
nand U3698 (N_3698,In_2096,In_15);
or U3699 (N_3699,In_2865,In_1162);
xnor U3700 (N_3700,In_237,In_2758);
or U3701 (N_3701,In_2755,In_2788);
nand U3702 (N_3702,In_1899,In_124);
nor U3703 (N_3703,In_2675,In_627);
nand U3704 (N_3704,In_2713,In_2807);
or U3705 (N_3705,In_1922,In_1429);
or U3706 (N_3706,In_1521,In_2474);
nand U3707 (N_3707,In_621,In_1594);
xnor U3708 (N_3708,In_765,In_2347);
and U3709 (N_3709,In_2319,In_426);
nor U3710 (N_3710,In_2375,In_373);
xor U3711 (N_3711,In_1921,In_1719);
nand U3712 (N_3712,In_2873,In_146);
or U3713 (N_3713,In_1967,In_2187);
nand U3714 (N_3714,In_334,In_1959);
nor U3715 (N_3715,In_1267,In_2586);
and U3716 (N_3716,In_719,In_1334);
and U3717 (N_3717,In_1356,In_1222);
or U3718 (N_3718,In_1399,In_657);
nand U3719 (N_3719,In_2069,In_2329);
nor U3720 (N_3720,In_252,In_2927);
nor U3721 (N_3721,In_316,In_51);
and U3722 (N_3722,In_2491,In_312);
nor U3723 (N_3723,In_2650,In_986);
nor U3724 (N_3724,In_2862,In_1596);
or U3725 (N_3725,In_695,In_478);
and U3726 (N_3726,In_1073,In_2830);
or U3727 (N_3727,In_2240,In_1755);
xor U3728 (N_3728,In_2548,In_2095);
nand U3729 (N_3729,In_1607,In_1190);
or U3730 (N_3730,In_1420,In_1666);
nor U3731 (N_3731,In_2228,In_1310);
and U3732 (N_3732,In_1118,In_369);
and U3733 (N_3733,In_1008,In_752);
nand U3734 (N_3734,In_798,In_2567);
or U3735 (N_3735,In_1149,In_722);
or U3736 (N_3736,In_2457,In_593);
nand U3737 (N_3737,In_2927,In_827);
xnor U3738 (N_3738,In_2631,In_1608);
xnor U3739 (N_3739,In_1995,In_2766);
or U3740 (N_3740,In_36,In_1065);
or U3741 (N_3741,In_2102,In_1852);
nand U3742 (N_3742,In_2928,In_1570);
and U3743 (N_3743,In_2056,In_1194);
and U3744 (N_3744,In_2345,In_1406);
xnor U3745 (N_3745,In_1182,In_2643);
or U3746 (N_3746,In_90,In_473);
nand U3747 (N_3747,In_2014,In_1197);
and U3748 (N_3748,In_120,In_911);
nor U3749 (N_3749,In_2181,In_884);
xnor U3750 (N_3750,In_2591,In_790);
xor U3751 (N_3751,In_1644,In_1338);
nand U3752 (N_3752,In_2146,In_1912);
nor U3753 (N_3753,In_2059,In_484);
xor U3754 (N_3754,In_509,In_505);
nand U3755 (N_3755,In_1633,In_1218);
and U3756 (N_3756,In_1591,In_32);
nor U3757 (N_3757,In_515,In_1432);
nand U3758 (N_3758,In_623,In_2064);
and U3759 (N_3759,In_2808,In_1867);
or U3760 (N_3760,In_1244,In_1182);
nor U3761 (N_3761,In_529,In_2120);
xnor U3762 (N_3762,In_2544,In_425);
and U3763 (N_3763,In_1236,In_1863);
or U3764 (N_3764,In_800,In_2417);
or U3765 (N_3765,In_1263,In_2996);
or U3766 (N_3766,In_539,In_430);
or U3767 (N_3767,In_166,In_604);
nand U3768 (N_3768,In_384,In_1836);
or U3769 (N_3769,In_2625,In_2775);
nor U3770 (N_3770,In_239,In_1188);
xnor U3771 (N_3771,In_2810,In_2758);
xnor U3772 (N_3772,In_2702,In_795);
and U3773 (N_3773,In_2671,In_376);
nand U3774 (N_3774,In_2905,In_642);
xnor U3775 (N_3775,In_1746,In_394);
nor U3776 (N_3776,In_1852,In_1396);
and U3777 (N_3777,In_1639,In_628);
nor U3778 (N_3778,In_288,In_2463);
or U3779 (N_3779,In_1174,In_1491);
nor U3780 (N_3780,In_305,In_585);
xnor U3781 (N_3781,In_1829,In_857);
or U3782 (N_3782,In_1303,In_1077);
xnor U3783 (N_3783,In_1369,In_2139);
xnor U3784 (N_3784,In_1845,In_2982);
and U3785 (N_3785,In_2673,In_201);
xnor U3786 (N_3786,In_2432,In_2088);
xor U3787 (N_3787,In_1210,In_1907);
nor U3788 (N_3788,In_1849,In_1021);
xnor U3789 (N_3789,In_2604,In_2301);
xor U3790 (N_3790,In_2773,In_93);
xor U3791 (N_3791,In_2484,In_2300);
nor U3792 (N_3792,In_182,In_417);
nand U3793 (N_3793,In_2811,In_1596);
or U3794 (N_3794,In_2134,In_534);
and U3795 (N_3795,In_2840,In_394);
or U3796 (N_3796,In_1626,In_2612);
nor U3797 (N_3797,In_1123,In_2044);
and U3798 (N_3798,In_1773,In_99);
or U3799 (N_3799,In_462,In_86);
nor U3800 (N_3800,In_515,In_1610);
nand U3801 (N_3801,In_100,In_1391);
and U3802 (N_3802,In_2516,In_2134);
xnor U3803 (N_3803,In_2542,In_2744);
nand U3804 (N_3804,In_108,In_262);
and U3805 (N_3805,In_623,In_611);
nand U3806 (N_3806,In_1107,In_2657);
nor U3807 (N_3807,In_1908,In_2596);
or U3808 (N_3808,In_2280,In_438);
nor U3809 (N_3809,In_2739,In_487);
nor U3810 (N_3810,In_1602,In_2584);
and U3811 (N_3811,In_2160,In_693);
and U3812 (N_3812,In_430,In_2456);
nor U3813 (N_3813,In_1181,In_1603);
or U3814 (N_3814,In_196,In_1835);
nand U3815 (N_3815,In_2530,In_2020);
xor U3816 (N_3816,In_1434,In_1752);
and U3817 (N_3817,In_19,In_2739);
or U3818 (N_3818,In_1060,In_2843);
or U3819 (N_3819,In_2517,In_2872);
nand U3820 (N_3820,In_2635,In_1144);
xnor U3821 (N_3821,In_137,In_851);
or U3822 (N_3822,In_1007,In_2389);
and U3823 (N_3823,In_954,In_232);
nand U3824 (N_3824,In_1357,In_580);
nor U3825 (N_3825,In_730,In_809);
and U3826 (N_3826,In_876,In_616);
xnor U3827 (N_3827,In_1039,In_740);
and U3828 (N_3828,In_1897,In_2414);
nor U3829 (N_3829,In_2506,In_1428);
and U3830 (N_3830,In_2538,In_2336);
or U3831 (N_3831,In_2621,In_1649);
nand U3832 (N_3832,In_1083,In_2260);
nand U3833 (N_3833,In_2033,In_1264);
and U3834 (N_3834,In_2001,In_1027);
and U3835 (N_3835,In_2563,In_1493);
and U3836 (N_3836,In_898,In_1788);
nand U3837 (N_3837,In_2701,In_456);
xnor U3838 (N_3838,In_2082,In_2577);
or U3839 (N_3839,In_1241,In_2886);
or U3840 (N_3840,In_344,In_332);
nand U3841 (N_3841,In_514,In_273);
xor U3842 (N_3842,In_2274,In_1553);
nand U3843 (N_3843,In_1520,In_1703);
xnor U3844 (N_3844,In_1092,In_288);
or U3845 (N_3845,In_1009,In_1686);
or U3846 (N_3846,In_1576,In_113);
nand U3847 (N_3847,In_682,In_2080);
nor U3848 (N_3848,In_1965,In_2176);
or U3849 (N_3849,In_2511,In_878);
xnor U3850 (N_3850,In_1399,In_219);
nor U3851 (N_3851,In_2659,In_1834);
xor U3852 (N_3852,In_900,In_1502);
nand U3853 (N_3853,In_821,In_500);
and U3854 (N_3854,In_562,In_2191);
nor U3855 (N_3855,In_1898,In_1699);
or U3856 (N_3856,In_937,In_285);
and U3857 (N_3857,In_1069,In_198);
or U3858 (N_3858,In_2134,In_290);
nand U3859 (N_3859,In_816,In_463);
xor U3860 (N_3860,In_2938,In_1818);
xnor U3861 (N_3861,In_2841,In_707);
nand U3862 (N_3862,In_1846,In_375);
nor U3863 (N_3863,In_1940,In_9);
xnor U3864 (N_3864,In_1698,In_2349);
nor U3865 (N_3865,In_1239,In_2072);
and U3866 (N_3866,In_1118,In_1724);
nor U3867 (N_3867,In_20,In_226);
and U3868 (N_3868,In_1763,In_254);
nor U3869 (N_3869,In_2910,In_231);
nand U3870 (N_3870,In_1328,In_2620);
nand U3871 (N_3871,In_819,In_2987);
or U3872 (N_3872,In_2030,In_2281);
xnor U3873 (N_3873,In_1063,In_2877);
nor U3874 (N_3874,In_971,In_2344);
nor U3875 (N_3875,In_1105,In_1910);
and U3876 (N_3876,In_2979,In_321);
and U3877 (N_3877,In_1928,In_1633);
nor U3878 (N_3878,In_2382,In_291);
or U3879 (N_3879,In_989,In_1672);
nand U3880 (N_3880,In_2717,In_1587);
and U3881 (N_3881,In_2417,In_603);
xor U3882 (N_3882,In_147,In_123);
nand U3883 (N_3883,In_2404,In_1136);
and U3884 (N_3884,In_195,In_138);
or U3885 (N_3885,In_1100,In_919);
and U3886 (N_3886,In_896,In_24);
xor U3887 (N_3887,In_1815,In_1640);
nor U3888 (N_3888,In_2834,In_884);
or U3889 (N_3889,In_917,In_756);
xnor U3890 (N_3890,In_2648,In_2052);
nor U3891 (N_3891,In_271,In_2617);
nor U3892 (N_3892,In_2469,In_2556);
and U3893 (N_3893,In_4,In_655);
nand U3894 (N_3894,In_1557,In_1743);
xor U3895 (N_3895,In_1581,In_2284);
xor U3896 (N_3896,In_2522,In_1383);
nand U3897 (N_3897,In_1468,In_2159);
nor U3898 (N_3898,In_841,In_2883);
nand U3899 (N_3899,In_1142,In_2341);
nand U3900 (N_3900,In_2668,In_1364);
and U3901 (N_3901,In_195,In_2244);
and U3902 (N_3902,In_1144,In_803);
nor U3903 (N_3903,In_230,In_1856);
nand U3904 (N_3904,In_2555,In_1917);
or U3905 (N_3905,In_1328,In_2654);
xor U3906 (N_3906,In_695,In_2708);
nand U3907 (N_3907,In_2514,In_2802);
nand U3908 (N_3908,In_2304,In_846);
nor U3909 (N_3909,In_4,In_2390);
nand U3910 (N_3910,In_1115,In_2568);
and U3911 (N_3911,In_388,In_1810);
and U3912 (N_3912,In_2428,In_2785);
and U3913 (N_3913,In_2359,In_55);
xnor U3914 (N_3914,In_2149,In_2014);
xnor U3915 (N_3915,In_214,In_662);
nor U3916 (N_3916,In_303,In_367);
nor U3917 (N_3917,In_1122,In_1377);
or U3918 (N_3918,In_2794,In_2930);
nor U3919 (N_3919,In_2226,In_1399);
nor U3920 (N_3920,In_2884,In_838);
and U3921 (N_3921,In_2666,In_811);
and U3922 (N_3922,In_2783,In_1947);
nand U3923 (N_3923,In_1992,In_620);
or U3924 (N_3924,In_1789,In_1861);
nor U3925 (N_3925,In_1218,In_2247);
and U3926 (N_3926,In_2407,In_562);
or U3927 (N_3927,In_577,In_2726);
nand U3928 (N_3928,In_1047,In_2270);
and U3929 (N_3929,In_2096,In_646);
and U3930 (N_3930,In_1008,In_1678);
nand U3931 (N_3931,In_1033,In_2895);
nand U3932 (N_3932,In_1322,In_1057);
nor U3933 (N_3933,In_106,In_881);
and U3934 (N_3934,In_2931,In_1871);
nor U3935 (N_3935,In_442,In_872);
nor U3936 (N_3936,In_1061,In_1646);
and U3937 (N_3937,In_675,In_796);
nor U3938 (N_3938,In_1022,In_322);
xor U3939 (N_3939,In_58,In_1437);
or U3940 (N_3940,In_2328,In_2519);
or U3941 (N_3941,In_2731,In_609);
xnor U3942 (N_3942,In_1804,In_252);
xor U3943 (N_3943,In_884,In_2439);
or U3944 (N_3944,In_2283,In_2330);
or U3945 (N_3945,In_2691,In_2319);
or U3946 (N_3946,In_1386,In_1168);
nor U3947 (N_3947,In_2,In_1224);
and U3948 (N_3948,In_2229,In_1285);
nand U3949 (N_3949,In_1308,In_1333);
and U3950 (N_3950,In_1960,In_2075);
or U3951 (N_3951,In_2029,In_512);
nor U3952 (N_3952,In_1221,In_1262);
xor U3953 (N_3953,In_2953,In_89);
nor U3954 (N_3954,In_2217,In_1744);
and U3955 (N_3955,In_1624,In_199);
or U3956 (N_3956,In_2072,In_248);
xnor U3957 (N_3957,In_805,In_2323);
nand U3958 (N_3958,In_1976,In_1479);
xnor U3959 (N_3959,In_2401,In_2404);
nor U3960 (N_3960,In_484,In_2691);
xor U3961 (N_3961,In_2565,In_854);
or U3962 (N_3962,In_2827,In_2565);
xor U3963 (N_3963,In_493,In_2831);
and U3964 (N_3964,In_157,In_2383);
nand U3965 (N_3965,In_820,In_1886);
xor U3966 (N_3966,In_1289,In_1490);
nand U3967 (N_3967,In_1279,In_2898);
or U3968 (N_3968,In_1022,In_1116);
xor U3969 (N_3969,In_2555,In_1686);
and U3970 (N_3970,In_1076,In_169);
and U3971 (N_3971,In_1686,In_2524);
xor U3972 (N_3972,In_1643,In_1075);
or U3973 (N_3973,In_720,In_2709);
and U3974 (N_3974,In_2488,In_2840);
nor U3975 (N_3975,In_348,In_1523);
nor U3976 (N_3976,In_39,In_1458);
nor U3977 (N_3977,In_1100,In_2359);
and U3978 (N_3978,In_2160,In_1827);
nor U3979 (N_3979,In_2310,In_2462);
xor U3980 (N_3980,In_2588,In_1748);
nor U3981 (N_3981,In_2661,In_2583);
and U3982 (N_3982,In_2525,In_2767);
and U3983 (N_3983,In_1025,In_770);
or U3984 (N_3984,In_1893,In_2676);
xor U3985 (N_3985,In_2950,In_1629);
xor U3986 (N_3986,In_444,In_2896);
and U3987 (N_3987,In_446,In_2920);
and U3988 (N_3988,In_2506,In_2330);
or U3989 (N_3989,In_583,In_1448);
xor U3990 (N_3990,In_859,In_1059);
nor U3991 (N_3991,In_454,In_2875);
or U3992 (N_3992,In_794,In_2921);
or U3993 (N_3993,In_1664,In_858);
xor U3994 (N_3994,In_1324,In_2025);
xnor U3995 (N_3995,In_836,In_2858);
xor U3996 (N_3996,In_827,In_2885);
xor U3997 (N_3997,In_2850,In_1454);
xor U3998 (N_3998,In_2316,In_786);
and U3999 (N_3999,In_2556,In_2767);
xnor U4000 (N_4000,In_1442,In_341);
and U4001 (N_4001,In_472,In_908);
xnor U4002 (N_4002,In_1159,In_1932);
or U4003 (N_4003,In_2830,In_1120);
nor U4004 (N_4004,In_2447,In_2003);
nor U4005 (N_4005,In_30,In_2628);
or U4006 (N_4006,In_1891,In_1685);
xor U4007 (N_4007,In_895,In_1818);
or U4008 (N_4008,In_1011,In_1414);
or U4009 (N_4009,In_1183,In_1282);
nor U4010 (N_4010,In_1375,In_2411);
and U4011 (N_4011,In_1233,In_2841);
xnor U4012 (N_4012,In_1609,In_2995);
or U4013 (N_4013,In_1771,In_1990);
or U4014 (N_4014,In_2051,In_1426);
or U4015 (N_4015,In_658,In_2411);
xnor U4016 (N_4016,In_1278,In_1901);
nor U4017 (N_4017,In_2842,In_584);
and U4018 (N_4018,In_2373,In_101);
or U4019 (N_4019,In_2373,In_885);
xnor U4020 (N_4020,In_1149,In_1010);
nor U4021 (N_4021,In_2414,In_1952);
or U4022 (N_4022,In_997,In_2435);
xor U4023 (N_4023,In_21,In_1829);
nand U4024 (N_4024,In_1845,In_2322);
or U4025 (N_4025,In_889,In_1344);
nor U4026 (N_4026,In_1902,In_1814);
or U4027 (N_4027,In_700,In_1689);
or U4028 (N_4028,In_2942,In_2419);
and U4029 (N_4029,In_1024,In_2268);
xnor U4030 (N_4030,In_1344,In_2795);
xnor U4031 (N_4031,In_1715,In_172);
or U4032 (N_4032,In_64,In_2127);
nor U4033 (N_4033,In_2955,In_282);
or U4034 (N_4034,In_215,In_1755);
xor U4035 (N_4035,In_1681,In_157);
nor U4036 (N_4036,In_1879,In_1649);
and U4037 (N_4037,In_2797,In_732);
nand U4038 (N_4038,In_1639,In_2534);
xnor U4039 (N_4039,In_1040,In_2919);
nand U4040 (N_4040,In_120,In_876);
nand U4041 (N_4041,In_1549,In_1606);
nand U4042 (N_4042,In_571,In_2714);
xor U4043 (N_4043,In_61,In_2529);
and U4044 (N_4044,In_1252,In_2285);
and U4045 (N_4045,In_914,In_2109);
xnor U4046 (N_4046,In_23,In_2192);
nor U4047 (N_4047,In_1121,In_1292);
and U4048 (N_4048,In_2971,In_1107);
and U4049 (N_4049,In_1477,In_37);
or U4050 (N_4050,In_253,In_2952);
xnor U4051 (N_4051,In_2102,In_2587);
xnor U4052 (N_4052,In_503,In_1347);
nand U4053 (N_4053,In_1082,In_2813);
and U4054 (N_4054,In_2411,In_115);
nor U4055 (N_4055,In_1923,In_2556);
nand U4056 (N_4056,In_452,In_2913);
nand U4057 (N_4057,In_2070,In_10);
xor U4058 (N_4058,In_1259,In_1478);
nor U4059 (N_4059,In_1413,In_1353);
or U4060 (N_4060,In_108,In_525);
nor U4061 (N_4061,In_2676,In_447);
nor U4062 (N_4062,In_912,In_2556);
or U4063 (N_4063,In_2983,In_34);
and U4064 (N_4064,In_1797,In_2978);
xnor U4065 (N_4065,In_890,In_35);
nor U4066 (N_4066,In_2838,In_2826);
nor U4067 (N_4067,In_110,In_2674);
nand U4068 (N_4068,In_2321,In_879);
or U4069 (N_4069,In_1098,In_893);
and U4070 (N_4070,In_162,In_1634);
nand U4071 (N_4071,In_628,In_2907);
and U4072 (N_4072,In_1754,In_2431);
or U4073 (N_4073,In_1785,In_2432);
nand U4074 (N_4074,In_67,In_954);
nor U4075 (N_4075,In_2949,In_2128);
nand U4076 (N_4076,In_1657,In_2065);
or U4077 (N_4077,In_2331,In_1325);
xor U4078 (N_4078,In_500,In_2893);
and U4079 (N_4079,In_2564,In_2039);
nand U4080 (N_4080,In_2751,In_1610);
or U4081 (N_4081,In_1755,In_1516);
and U4082 (N_4082,In_2400,In_1482);
nor U4083 (N_4083,In_2025,In_2265);
nor U4084 (N_4084,In_1057,In_1814);
nand U4085 (N_4085,In_1385,In_2331);
xor U4086 (N_4086,In_114,In_2916);
and U4087 (N_4087,In_1217,In_1132);
and U4088 (N_4088,In_687,In_1548);
and U4089 (N_4089,In_1729,In_2855);
nor U4090 (N_4090,In_65,In_2376);
nor U4091 (N_4091,In_2947,In_2857);
and U4092 (N_4092,In_2608,In_181);
or U4093 (N_4093,In_1417,In_2024);
and U4094 (N_4094,In_1107,In_2189);
nor U4095 (N_4095,In_62,In_16);
and U4096 (N_4096,In_2014,In_483);
or U4097 (N_4097,In_2846,In_2422);
nand U4098 (N_4098,In_2833,In_1878);
nand U4099 (N_4099,In_1871,In_2943);
nand U4100 (N_4100,In_1647,In_1735);
and U4101 (N_4101,In_2691,In_120);
xnor U4102 (N_4102,In_1030,In_277);
nor U4103 (N_4103,In_2889,In_1782);
nand U4104 (N_4104,In_1761,In_2107);
or U4105 (N_4105,In_2136,In_2754);
or U4106 (N_4106,In_2942,In_946);
xor U4107 (N_4107,In_1449,In_2517);
and U4108 (N_4108,In_1436,In_1974);
xor U4109 (N_4109,In_885,In_26);
and U4110 (N_4110,In_2951,In_276);
and U4111 (N_4111,In_552,In_1212);
nand U4112 (N_4112,In_232,In_821);
nor U4113 (N_4113,In_1552,In_1257);
or U4114 (N_4114,In_2038,In_2617);
xnor U4115 (N_4115,In_1173,In_696);
xnor U4116 (N_4116,In_2605,In_40);
nor U4117 (N_4117,In_902,In_978);
or U4118 (N_4118,In_9,In_320);
nor U4119 (N_4119,In_1396,In_251);
xor U4120 (N_4120,In_1146,In_234);
nor U4121 (N_4121,In_2291,In_2420);
and U4122 (N_4122,In_2133,In_1263);
xor U4123 (N_4123,In_1998,In_2987);
nor U4124 (N_4124,In_428,In_481);
nor U4125 (N_4125,In_239,In_2951);
xor U4126 (N_4126,In_1802,In_2134);
nand U4127 (N_4127,In_1370,In_1973);
nor U4128 (N_4128,In_1397,In_1033);
nor U4129 (N_4129,In_794,In_2121);
nor U4130 (N_4130,In_56,In_395);
nor U4131 (N_4131,In_2605,In_2822);
nand U4132 (N_4132,In_79,In_369);
nand U4133 (N_4133,In_2362,In_1616);
nor U4134 (N_4134,In_1210,In_2022);
xor U4135 (N_4135,In_1866,In_2322);
and U4136 (N_4136,In_140,In_2867);
nor U4137 (N_4137,In_2064,In_211);
xnor U4138 (N_4138,In_2305,In_2646);
xnor U4139 (N_4139,In_1849,In_2391);
nand U4140 (N_4140,In_2088,In_472);
nor U4141 (N_4141,In_1947,In_2806);
xnor U4142 (N_4142,In_758,In_2593);
nor U4143 (N_4143,In_996,In_1246);
nand U4144 (N_4144,In_1344,In_2601);
nand U4145 (N_4145,In_1533,In_789);
nand U4146 (N_4146,In_1548,In_25);
xnor U4147 (N_4147,In_1592,In_2994);
xor U4148 (N_4148,In_997,In_2208);
xor U4149 (N_4149,In_1120,In_214);
and U4150 (N_4150,In_2969,In_2218);
nor U4151 (N_4151,In_1462,In_1501);
xor U4152 (N_4152,In_2691,In_542);
and U4153 (N_4153,In_501,In_1358);
and U4154 (N_4154,In_2980,In_123);
xnor U4155 (N_4155,In_192,In_2848);
xnor U4156 (N_4156,In_965,In_377);
nor U4157 (N_4157,In_862,In_1996);
or U4158 (N_4158,In_569,In_2738);
and U4159 (N_4159,In_1564,In_762);
nor U4160 (N_4160,In_2907,In_619);
or U4161 (N_4161,In_610,In_123);
nand U4162 (N_4162,In_1289,In_138);
nor U4163 (N_4163,In_2351,In_1495);
and U4164 (N_4164,In_1630,In_2206);
xnor U4165 (N_4165,In_129,In_2189);
or U4166 (N_4166,In_1116,In_1602);
or U4167 (N_4167,In_2307,In_2722);
and U4168 (N_4168,In_572,In_544);
or U4169 (N_4169,In_393,In_1469);
nor U4170 (N_4170,In_793,In_2);
nand U4171 (N_4171,In_2855,In_727);
nor U4172 (N_4172,In_1500,In_994);
or U4173 (N_4173,In_1552,In_2174);
or U4174 (N_4174,In_1150,In_2937);
and U4175 (N_4175,In_1197,In_1300);
nand U4176 (N_4176,In_857,In_2582);
nand U4177 (N_4177,In_1585,In_1201);
nand U4178 (N_4178,In_2474,In_117);
nor U4179 (N_4179,In_63,In_620);
and U4180 (N_4180,In_2551,In_2055);
nor U4181 (N_4181,In_695,In_2043);
or U4182 (N_4182,In_760,In_655);
xor U4183 (N_4183,In_682,In_2885);
nor U4184 (N_4184,In_812,In_205);
nor U4185 (N_4185,In_971,In_1700);
nand U4186 (N_4186,In_1609,In_1683);
or U4187 (N_4187,In_809,In_811);
xor U4188 (N_4188,In_2320,In_2293);
or U4189 (N_4189,In_1863,In_2706);
and U4190 (N_4190,In_1305,In_988);
or U4191 (N_4191,In_398,In_556);
xor U4192 (N_4192,In_396,In_2710);
or U4193 (N_4193,In_1571,In_887);
and U4194 (N_4194,In_1676,In_1922);
nor U4195 (N_4195,In_2378,In_2995);
or U4196 (N_4196,In_1536,In_1402);
or U4197 (N_4197,In_2740,In_1293);
nand U4198 (N_4198,In_1666,In_1687);
xnor U4199 (N_4199,In_1441,In_2158);
nor U4200 (N_4200,In_673,In_2173);
nand U4201 (N_4201,In_7,In_501);
or U4202 (N_4202,In_519,In_5);
nand U4203 (N_4203,In_879,In_969);
nand U4204 (N_4204,In_2207,In_2262);
nand U4205 (N_4205,In_2986,In_325);
and U4206 (N_4206,In_1296,In_459);
and U4207 (N_4207,In_1823,In_291);
and U4208 (N_4208,In_436,In_789);
nor U4209 (N_4209,In_128,In_1365);
nor U4210 (N_4210,In_2950,In_1612);
and U4211 (N_4211,In_2592,In_573);
or U4212 (N_4212,In_109,In_2106);
and U4213 (N_4213,In_649,In_1988);
nor U4214 (N_4214,In_1493,In_2207);
nand U4215 (N_4215,In_2834,In_2243);
or U4216 (N_4216,In_1049,In_2730);
xor U4217 (N_4217,In_1570,In_1265);
and U4218 (N_4218,In_1036,In_1226);
and U4219 (N_4219,In_358,In_1530);
xor U4220 (N_4220,In_451,In_1129);
and U4221 (N_4221,In_2677,In_73);
nand U4222 (N_4222,In_958,In_2714);
nor U4223 (N_4223,In_410,In_774);
xor U4224 (N_4224,In_1226,In_1580);
and U4225 (N_4225,In_2480,In_1835);
xor U4226 (N_4226,In_2230,In_131);
or U4227 (N_4227,In_1022,In_2952);
or U4228 (N_4228,In_1635,In_753);
nand U4229 (N_4229,In_2126,In_2846);
xor U4230 (N_4230,In_2939,In_2911);
or U4231 (N_4231,In_2604,In_1870);
nand U4232 (N_4232,In_2532,In_1813);
or U4233 (N_4233,In_955,In_2448);
or U4234 (N_4234,In_207,In_1490);
nor U4235 (N_4235,In_1952,In_375);
or U4236 (N_4236,In_2596,In_372);
nand U4237 (N_4237,In_629,In_1049);
and U4238 (N_4238,In_544,In_1294);
nor U4239 (N_4239,In_2437,In_2270);
nand U4240 (N_4240,In_763,In_2472);
nor U4241 (N_4241,In_2588,In_2038);
nor U4242 (N_4242,In_2602,In_359);
xor U4243 (N_4243,In_2390,In_984);
and U4244 (N_4244,In_178,In_1604);
or U4245 (N_4245,In_2259,In_339);
and U4246 (N_4246,In_1015,In_952);
or U4247 (N_4247,In_2007,In_1923);
xor U4248 (N_4248,In_2188,In_625);
or U4249 (N_4249,In_1262,In_1544);
or U4250 (N_4250,In_2246,In_701);
xnor U4251 (N_4251,In_717,In_2496);
xor U4252 (N_4252,In_129,In_1258);
or U4253 (N_4253,In_2089,In_269);
nor U4254 (N_4254,In_2004,In_2932);
nor U4255 (N_4255,In_2687,In_2060);
nand U4256 (N_4256,In_1413,In_466);
and U4257 (N_4257,In_2332,In_74);
or U4258 (N_4258,In_970,In_409);
xor U4259 (N_4259,In_1741,In_60);
or U4260 (N_4260,In_1722,In_566);
xor U4261 (N_4261,In_1544,In_136);
nor U4262 (N_4262,In_1212,In_1899);
or U4263 (N_4263,In_1421,In_1265);
nor U4264 (N_4264,In_1774,In_2977);
or U4265 (N_4265,In_2519,In_2247);
xor U4266 (N_4266,In_2162,In_1849);
or U4267 (N_4267,In_2133,In_1681);
or U4268 (N_4268,In_1248,In_1475);
nand U4269 (N_4269,In_1935,In_2650);
or U4270 (N_4270,In_297,In_348);
and U4271 (N_4271,In_2209,In_2674);
or U4272 (N_4272,In_220,In_2390);
xnor U4273 (N_4273,In_1319,In_799);
xor U4274 (N_4274,In_1801,In_1403);
and U4275 (N_4275,In_933,In_1397);
and U4276 (N_4276,In_127,In_2290);
nand U4277 (N_4277,In_2851,In_15);
or U4278 (N_4278,In_2464,In_1119);
nand U4279 (N_4279,In_2118,In_2278);
nor U4280 (N_4280,In_40,In_1170);
or U4281 (N_4281,In_1935,In_826);
nor U4282 (N_4282,In_1327,In_390);
or U4283 (N_4283,In_2806,In_2861);
nand U4284 (N_4284,In_685,In_1481);
or U4285 (N_4285,In_894,In_725);
xor U4286 (N_4286,In_784,In_2785);
nor U4287 (N_4287,In_1677,In_184);
or U4288 (N_4288,In_892,In_2260);
nand U4289 (N_4289,In_2582,In_2979);
nand U4290 (N_4290,In_1257,In_2503);
xnor U4291 (N_4291,In_437,In_2982);
nand U4292 (N_4292,In_408,In_2357);
or U4293 (N_4293,In_1972,In_14);
or U4294 (N_4294,In_959,In_531);
xor U4295 (N_4295,In_1432,In_1425);
and U4296 (N_4296,In_595,In_319);
xor U4297 (N_4297,In_2770,In_2292);
xor U4298 (N_4298,In_597,In_861);
xnor U4299 (N_4299,In_1031,In_2975);
xor U4300 (N_4300,In_410,In_1677);
or U4301 (N_4301,In_1865,In_9);
or U4302 (N_4302,In_211,In_575);
nor U4303 (N_4303,In_2558,In_2141);
nand U4304 (N_4304,In_1875,In_2805);
nor U4305 (N_4305,In_2325,In_1426);
xnor U4306 (N_4306,In_833,In_1304);
or U4307 (N_4307,In_1040,In_2009);
xor U4308 (N_4308,In_2222,In_2517);
or U4309 (N_4309,In_1207,In_2696);
and U4310 (N_4310,In_1874,In_2258);
nor U4311 (N_4311,In_2126,In_474);
xor U4312 (N_4312,In_679,In_993);
and U4313 (N_4313,In_513,In_652);
xor U4314 (N_4314,In_857,In_528);
or U4315 (N_4315,In_2313,In_1309);
nor U4316 (N_4316,In_858,In_1238);
nand U4317 (N_4317,In_1271,In_1796);
nand U4318 (N_4318,In_2713,In_1898);
and U4319 (N_4319,In_84,In_45);
nand U4320 (N_4320,In_1914,In_2961);
nor U4321 (N_4321,In_401,In_2105);
or U4322 (N_4322,In_155,In_517);
xnor U4323 (N_4323,In_2850,In_1126);
xor U4324 (N_4324,In_1629,In_1985);
nor U4325 (N_4325,In_2790,In_2968);
and U4326 (N_4326,In_2467,In_504);
xnor U4327 (N_4327,In_869,In_1894);
nand U4328 (N_4328,In_1682,In_742);
nor U4329 (N_4329,In_2464,In_408);
or U4330 (N_4330,In_2855,In_1862);
or U4331 (N_4331,In_518,In_2630);
nor U4332 (N_4332,In_2690,In_337);
nand U4333 (N_4333,In_838,In_649);
xor U4334 (N_4334,In_2293,In_1368);
or U4335 (N_4335,In_266,In_2316);
nand U4336 (N_4336,In_1162,In_838);
xor U4337 (N_4337,In_1082,In_2726);
and U4338 (N_4338,In_930,In_907);
xnor U4339 (N_4339,In_2809,In_819);
or U4340 (N_4340,In_631,In_582);
nand U4341 (N_4341,In_2883,In_2242);
and U4342 (N_4342,In_944,In_1308);
or U4343 (N_4343,In_1503,In_624);
nor U4344 (N_4344,In_1468,In_202);
and U4345 (N_4345,In_2858,In_405);
nand U4346 (N_4346,In_2173,In_2160);
nand U4347 (N_4347,In_2207,In_2539);
nor U4348 (N_4348,In_2479,In_30);
and U4349 (N_4349,In_231,In_679);
xnor U4350 (N_4350,In_1700,In_265);
or U4351 (N_4351,In_2118,In_2293);
and U4352 (N_4352,In_1979,In_945);
and U4353 (N_4353,In_1184,In_630);
xor U4354 (N_4354,In_2169,In_2827);
nor U4355 (N_4355,In_674,In_2098);
and U4356 (N_4356,In_2235,In_549);
and U4357 (N_4357,In_470,In_1181);
xor U4358 (N_4358,In_2489,In_1865);
nor U4359 (N_4359,In_1304,In_2590);
or U4360 (N_4360,In_1881,In_1143);
nor U4361 (N_4361,In_2919,In_2584);
nor U4362 (N_4362,In_1455,In_1526);
nor U4363 (N_4363,In_2114,In_2639);
nor U4364 (N_4364,In_154,In_578);
or U4365 (N_4365,In_2404,In_712);
and U4366 (N_4366,In_367,In_699);
nor U4367 (N_4367,In_706,In_1529);
xnor U4368 (N_4368,In_2114,In_2808);
nand U4369 (N_4369,In_1099,In_2049);
and U4370 (N_4370,In_1031,In_340);
and U4371 (N_4371,In_2637,In_122);
nand U4372 (N_4372,In_1296,In_2550);
and U4373 (N_4373,In_2862,In_243);
nand U4374 (N_4374,In_1082,In_628);
xor U4375 (N_4375,In_1182,In_101);
nand U4376 (N_4376,In_154,In_1704);
and U4377 (N_4377,In_1710,In_2961);
or U4378 (N_4378,In_1947,In_2306);
nand U4379 (N_4379,In_774,In_1533);
nand U4380 (N_4380,In_2928,In_2900);
nand U4381 (N_4381,In_205,In_1915);
and U4382 (N_4382,In_1516,In_2581);
xor U4383 (N_4383,In_71,In_120);
nor U4384 (N_4384,In_2699,In_98);
or U4385 (N_4385,In_418,In_2712);
and U4386 (N_4386,In_229,In_295);
nor U4387 (N_4387,In_742,In_789);
nor U4388 (N_4388,In_565,In_1092);
xor U4389 (N_4389,In_1320,In_1936);
or U4390 (N_4390,In_299,In_1653);
nand U4391 (N_4391,In_1257,In_2983);
and U4392 (N_4392,In_380,In_2381);
or U4393 (N_4393,In_2914,In_2642);
and U4394 (N_4394,In_51,In_2706);
xnor U4395 (N_4395,In_1285,In_2990);
xor U4396 (N_4396,In_2100,In_607);
or U4397 (N_4397,In_36,In_1372);
and U4398 (N_4398,In_1861,In_867);
or U4399 (N_4399,In_592,In_331);
nor U4400 (N_4400,In_1658,In_2255);
nor U4401 (N_4401,In_2323,In_381);
nand U4402 (N_4402,In_2352,In_2153);
nand U4403 (N_4403,In_1285,In_2962);
nand U4404 (N_4404,In_2407,In_368);
and U4405 (N_4405,In_2914,In_984);
xnor U4406 (N_4406,In_178,In_44);
nand U4407 (N_4407,In_1761,In_2199);
nand U4408 (N_4408,In_1892,In_1495);
or U4409 (N_4409,In_506,In_2145);
nor U4410 (N_4410,In_721,In_1021);
and U4411 (N_4411,In_1120,In_1798);
nor U4412 (N_4412,In_651,In_1641);
nand U4413 (N_4413,In_2488,In_2825);
nand U4414 (N_4414,In_1463,In_2813);
and U4415 (N_4415,In_996,In_115);
nand U4416 (N_4416,In_531,In_1788);
nor U4417 (N_4417,In_1626,In_1522);
or U4418 (N_4418,In_1248,In_2434);
or U4419 (N_4419,In_2649,In_1984);
and U4420 (N_4420,In_1406,In_642);
and U4421 (N_4421,In_93,In_1013);
and U4422 (N_4422,In_2919,In_1648);
or U4423 (N_4423,In_2931,In_1505);
xor U4424 (N_4424,In_691,In_550);
nand U4425 (N_4425,In_2635,In_217);
xnor U4426 (N_4426,In_2765,In_86);
and U4427 (N_4427,In_1137,In_2193);
nand U4428 (N_4428,In_2348,In_2981);
xor U4429 (N_4429,In_926,In_227);
or U4430 (N_4430,In_877,In_1936);
or U4431 (N_4431,In_1608,In_2997);
xor U4432 (N_4432,In_478,In_2136);
or U4433 (N_4433,In_2461,In_267);
and U4434 (N_4434,In_2019,In_1443);
or U4435 (N_4435,In_2930,In_199);
and U4436 (N_4436,In_2607,In_1840);
nand U4437 (N_4437,In_745,In_643);
or U4438 (N_4438,In_2886,In_2880);
or U4439 (N_4439,In_2849,In_1079);
and U4440 (N_4440,In_2168,In_1979);
or U4441 (N_4441,In_2442,In_479);
nor U4442 (N_4442,In_556,In_457);
xor U4443 (N_4443,In_2574,In_1105);
nand U4444 (N_4444,In_255,In_1333);
nor U4445 (N_4445,In_491,In_1424);
nand U4446 (N_4446,In_1679,In_95);
and U4447 (N_4447,In_763,In_2735);
or U4448 (N_4448,In_680,In_2228);
nor U4449 (N_4449,In_2520,In_1371);
xor U4450 (N_4450,In_1922,In_548);
and U4451 (N_4451,In_1193,In_1450);
and U4452 (N_4452,In_2685,In_267);
nand U4453 (N_4453,In_1764,In_2728);
xor U4454 (N_4454,In_1510,In_730);
nor U4455 (N_4455,In_753,In_2533);
nor U4456 (N_4456,In_684,In_2034);
nand U4457 (N_4457,In_75,In_2757);
or U4458 (N_4458,In_1250,In_2680);
or U4459 (N_4459,In_2460,In_1294);
nor U4460 (N_4460,In_151,In_1720);
nand U4461 (N_4461,In_1053,In_482);
xnor U4462 (N_4462,In_321,In_406);
xor U4463 (N_4463,In_2610,In_828);
xnor U4464 (N_4464,In_1374,In_2892);
or U4465 (N_4465,In_271,In_1501);
xor U4466 (N_4466,In_940,In_1346);
nand U4467 (N_4467,In_2156,In_1901);
and U4468 (N_4468,In_1694,In_752);
nor U4469 (N_4469,In_1036,In_899);
nor U4470 (N_4470,In_1070,In_229);
nand U4471 (N_4471,In_1460,In_855);
nor U4472 (N_4472,In_2391,In_456);
or U4473 (N_4473,In_1356,In_309);
xor U4474 (N_4474,In_1145,In_524);
nand U4475 (N_4475,In_912,In_2051);
nor U4476 (N_4476,In_1318,In_331);
and U4477 (N_4477,In_2243,In_315);
nand U4478 (N_4478,In_2857,In_2575);
or U4479 (N_4479,In_2389,In_567);
and U4480 (N_4480,In_1672,In_143);
nand U4481 (N_4481,In_2504,In_2818);
xor U4482 (N_4482,In_2027,In_8);
nand U4483 (N_4483,In_43,In_1546);
and U4484 (N_4484,In_127,In_1867);
or U4485 (N_4485,In_244,In_2688);
nor U4486 (N_4486,In_1374,In_2032);
and U4487 (N_4487,In_1977,In_1879);
and U4488 (N_4488,In_1799,In_2374);
or U4489 (N_4489,In_1440,In_1124);
xor U4490 (N_4490,In_1200,In_2687);
nor U4491 (N_4491,In_2630,In_2700);
or U4492 (N_4492,In_2916,In_1333);
nand U4493 (N_4493,In_295,In_1348);
nor U4494 (N_4494,In_1966,In_1726);
nand U4495 (N_4495,In_2152,In_957);
and U4496 (N_4496,In_2730,In_5);
or U4497 (N_4497,In_1808,In_2991);
or U4498 (N_4498,In_1106,In_132);
xnor U4499 (N_4499,In_2444,In_1588);
nand U4500 (N_4500,In_513,In_1250);
or U4501 (N_4501,In_1335,In_2880);
and U4502 (N_4502,In_2077,In_380);
nand U4503 (N_4503,In_1475,In_2688);
or U4504 (N_4504,In_1103,In_965);
nor U4505 (N_4505,In_2032,In_2991);
xnor U4506 (N_4506,In_1340,In_879);
xnor U4507 (N_4507,In_259,In_2778);
nor U4508 (N_4508,In_965,In_1074);
xnor U4509 (N_4509,In_92,In_2871);
or U4510 (N_4510,In_220,In_2532);
nor U4511 (N_4511,In_544,In_2273);
or U4512 (N_4512,In_2923,In_2405);
nor U4513 (N_4513,In_2605,In_508);
and U4514 (N_4514,In_783,In_1675);
nand U4515 (N_4515,In_1140,In_365);
and U4516 (N_4516,In_661,In_722);
xor U4517 (N_4517,In_1697,In_932);
xnor U4518 (N_4518,In_2131,In_1378);
or U4519 (N_4519,In_1954,In_1446);
and U4520 (N_4520,In_186,In_264);
or U4521 (N_4521,In_1973,In_2750);
nor U4522 (N_4522,In_2433,In_583);
or U4523 (N_4523,In_1674,In_1205);
xnor U4524 (N_4524,In_1836,In_1109);
nand U4525 (N_4525,In_2415,In_2739);
and U4526 (N_4526,In_1002,In_2645);
nor U4527 (N_4527,In_2472,In_2908);
nand U4528 (N_4528,In_414,In_125);
nand U4529 (N_4529,In_1297,In_1133);
xnor U4530 (N_4530,In_2812,In_1226);
xnor U4531 (N_4531,In_541,In_1726);
nand U4532 (N_4532,In_2608,In_1061);
and U4533 (N_4533,In_607,In_1174);
and U4534 (N_4534,In_2177,In_1406);
and U4535 (N_4535,In_565,In_2092);
nand U4536 (N_4536,In_1300,In_1088);
nand U4537 (N_4537,In_1496,In_1494);
and U4538 (N_4538,In_567,In_1394);
nor U4539 (N_4539,In_2404,In_1667);
and U4540 (N_4540,In_1989,In_2585);
and U4541 (N_4541,In_1283,In_1971);
or U4542 (N_4542,In_2975,In_946);
or U4543 (N_4543,In_2686,In_1696);
and U4544 (N_4544,In_2601,In_1409);
nand U4545 (N_4545,In_810,In_2017);
nand U4546 (N_4546,In_1044,In_2824);
nor U4547 (N_4547,In_1125,In_2565);
nor U4548 (N_4548,In_482,In_628);
or U4549 (N_4549,In_2807,In_1012);
or U4550 (N_4550,In_1103,In_1390);
nand U4551 (N_4551,In_293,In_2250);
or U4552 (N_4552,In_2721,In_302);
nand U4553 (N_4553,In_66,In_1407);
nor U4554 (N_4554,In_1288,In_2369);
and U4555 (N_4555,In_2601,In_2806);
or U4556 (N_4556,In_1921,In_2142);
and U4557 (N_4557,In_703,In_914);
nor U4558 (N_4558,In_1251,In_36);
or U4559 (N_4559,In_828,In_94);
and U4560 (N_4560,In_532,In_1477);
or U4561 (N_4561,In_1931,In_2295);
xor U4562 (N_4562,In_138,In_992);
or U4563 (N_4563,In_2427,In_1750);
xor U4564 (N_4564,In_2646,In_1888);
nand U4565 (N_4565,In_373,In_1968);
nor U4566 (N_4566,In_2957,In_2411);
nand U4567 (N_4567,In_2337,In_1023);
or U4568 (N_4568,In_1998,In_1355);
nand U4569 (N_4569,In_614,In_954);
nand U4570 (N_4570,In_2791,In_842);
and U4571 (N_4571,In_2964,In_2197);
nand U4572 (N_4572,In_2020,In_2190);
or U4573 (N_4573,In_1177,In_1634);
xnor U4574 (N_4574,In_2688,In_2146);
xnor U4575 (N_4575,In_1261,In_2764);
or U4576 (N_4576,In_2067,In_2951);
nor U4577 (N_4577,In_887,In_1850);
or U4578 (N_4578,In_1159,In_1755);
and U4579 (N_4579,In_719,In_1407);
and U4580 (N_4580,In_290,In_492);
nor U4581 (N_4581,In_2401,In_430);
nand U4582 (N_4582,In_854,In_2669);
xor U4583 (N_4583,In_2163,In_883);
nand U4584 (N_4584,In_2676,In_1043);
and U4585 (N_4585,In_1000,In_1273);
nand U4586 (N_4586,In_77,In_1483);
or U4587 (N_4587,In_2244,In_2966);
and U4588 (N_4588,In_1550,In_2866);
nand U4589 (N_4589,In_1004,In_2807);
nand U4590 (N_4590,In_1644,In_93);
or U4591 (N_4591,In_1960,In_1110);
nor U4592 (N_4592,In_324,In_1323);
nand U4593 (N_4593,In_2183,In_2950);
and U4594 (N_4594,In_508,In_815);
and U4595 (N_4595,In_23,In_1696);
xnor U4596 (N_4596,In_2772,In_1879);
xnor U4597 (N_4597,In_2759,In_256);
nor U4598 (N_4598,In_1267,In_1924);
xor U4599 (N_4599,In_2041,In_2481);
and U4600 (N_4600,In_110,In_821);
or U4601 (N_4601,In_2355,In_2316);
or U4602 (N_4602,In_1562,In_1992);
xnor U4603 (N_4603,In_194,In_658);
nand U4604 (N_4604,In_1388,In_2740);
nand U4605 (N_4605,In_326,In_481);
nand U4606 (N_4606,In_910,In_1289);
nand U4607 (N_4607,In_2137,In_1422);
nor U4608 (N_4608,In_2044,In_2701);
xor U4609 (N_4609,In_2403,In_2248);
and U4610 (N_4610,In_2235,In_439);
and U4611 (N_4611,In_2959,In_835);
nor U4612 (N_4612,In_2712,In_1794);
or U4613 (N_4613,In_427,In_2987);
xor U4614 (N_4614,In_1190,In_471);
or U4615 (N_4615,In_566,In_2354);
nor U4616 (N_4616,In_1837,In_1889);
nand U4617 (N_4617,In_1127,In_2552);
nor U4618 (N_4618,In_403,In_864);
nor U4619 (N_4619,In_714,In_2516);
and U4620 (N_4620,In_1438,In_1417);
and U4621 (N_4621,In_693,In_546);
xor U4622 (N_4622,In_975,In_1026);
and U4623 (N_4623,In_1630,In_2172);
nor U4624 (N_4624,In_2524,In_694);
nand U4625 (N_4625,In_1985,In_512);
and U4626 (N_4626,In_2080,In_1132);
and U4627 (N_4627,In_782,In_396);
and U4628 (N_4628,In_1645,In_434);
or U4629 (N_4629,In_1629,In_2807);
xor U4630 (N_4630,In_30,In_2804);
nor U4631 (N_4631,In_2548,In_2011);
nor U4632 (N_4632,In_2764,In_2915);
nor U4633 (N_4633,In_2122,In_70);
and U4634 (N_4634,In_1263,In_812);
and U4635 (N_4635,In_1761,In_1909);
nor U4636 (N_4636,In_1397,In_1137);
or U4637 (N_4637,In_401,In_653);
and U4638 (N_4638,In_636,In_2802);
and U4639 (N_4639,In_2169,In_1578);
and U4640 (N_4640,In_406,In_2539);
or U4641 (N_4641,In_2551,In_1586);
nor U4642 (N_4642,In_187,In_1837);
nor U4643 (N_4643,In_2004,In_1199);
nand U4644 (N_4644,In_2222,In_876);
or U4645 (N_4645,In_1024,In_1237);
nor U4646 (N_4646,In_2730,In_1507);
xor U4647 (N_4647,In_2283,In_1527);
and U4648 (N_4648,In_933,In_2423);
nand U4649 (N_4649,In_1270,In_486);
and U4650 (N_4650,In_124,In_235);
and U4651 (N_4651,In_638,In_1886);
and U4652 (N_4652,In_1804,In_2444);
or U4653 (N_4653,In_1061,In_226);
xor U4654 (N_4654,In_1838,In_2138);
or U4655 (N_4655,In_1729,In_850);
or U4656 (N_4656,In_2524,In_1310);
or U4657 (N_4657,In_2300,In_399);
or U4658 (N_4658,In_2263,In_1794);
nand U4659 (N_4659,In_1573,In_542);
xnor U4660 (N_4660,In_1376,In_2797);
or U4661 (N_4661,In_2196,In_2727);
and U4662 (N_4662,In_1607,In_2882);
nor U4663 (N_4663,In_1933,In_1428);
or U4664 (N_4664,In_2230,In_2295);
nand U4665 (N_4665,In_1712,In_1482);
or U4666 (N_4666,In_2957,In_317);
or U4667 (N_4667,In_2454,In_2637);
or U4668 (N_4668,In_967,In_1846);
or U4669 (N_4669,In_2074,In_654);
nand U4670 (N_4670,In_148,In_1974);
and U4671 (N_4671,In_651,In_2221);
nand U4672 (N_4672,In_939,In_835);
nand U4673 (N_4673,In_1926,In_2228);
xnor U4674 (N_4674,In_1310,In_246);
and U4675 (N_4675,In_2014,In_1489);
or U4676 (N_4676,In_1007,In_1359);
nor U4677 (N_4677,In_2618,In_1092);
nand U4678 (N_4678,In_1374,In_2611);
nand U4679 (N_4679,In_1766,In_2230);
or U4680 (N_4680,In_1107,In_1825);
and U4681 (N_4681,In_2072,In_1578);
nand U4682 (N_4682,In_1117,In_90);
nor U4683 (N_4683,In_2618,In_1778);
and U4684 (N_4684,In_1099,In_467);
or U4685 (N_4685,In_2907,In_324);
nor U4686 (N_4686,In_2649,In_1837);
or U4687 (N_4687,In_2206,In_1336);
xnor U4688 (N_4688,In_1726,In_2172);
nand U4689 (N_4689,In_1335,In_1397);
nor U4690 (N_4690,In_1365,In_1745);
and U4691 (N_4691,In_1363,In_2275);
nand U4692 (N_4692,In_118,In_8);
nand U4693 (N_4693,In_582,In_884);
xnor U4694 (N_4694,In_1678,In_521);
and U4695 (N_4695,In_1998,In_2097);
and U4696 (N_4696,In_463,In_1693);
or U4697 (N_4697,In_2327,In_1350);
nor U4698 (N_4698,In_2764,In_262);
nand U4699 (N_4699,In_1578,In_1315);
nand U4700 (N_4700,In_2551,In_16);
nand U4701 (N_4701,In_1121,In_1574);
and U4702 (N_4702,In_1305,In_282);
nor U4703 (N_4703,In_2630,In_537);
nor U4704 (N_4704,In_2363,In_1668);
xnor U4705 (N_4705,In_1598,In_1966);
nand U4706 (N_4706,In_2656,In_1489);
nor U4707 (N_4707,In_2989,In_2560);
nor U4708 (N_4708,In_332,In_1778);
and U4709 (N_4709,In_1282,In_1915);
and U4710 (N_4710,In_1843,In_206);
nand U4711 (N_4711,In_1919,In_1549);
nand U4712 (N_4712,In_2911,In_2783);
nand U4713 (N_4713,In_1766,In_1869);
and U4714 (N_4714,In_1672,In_1101);
xnor U4715 (N_4715,In_168,In_1182);
xor U4716 (N_4716,In_2864,In_2597);
nor U4717 (N_4717,In_2208,In_1664);
or U4718 (N_4718,In_703,In_839);
xnor U4719 (N_4719,In_2060,In_1733);
xor U4720 (N_4720,In_1141,In_2546);
xnor U4721 (N_4721,In_606,In_1502);
and U4722 (N_4722,In_1628,In_2894);
nor U4723 (N_4723,In_1277,In_1700);
or U4724 (N_4724,In_2725,In_782);
xnor U4725 (N_4725,In_1987,In_425);
nand U4726 (N_4726,In_2538,In_2612);
nor U4727 (N_4727,In_1723,In_1900);
nor U4728 (N_4728,In_647,In_2590);
or U4729 (N_4729,In_767,In_1646);
nand U4730 (N_4730,In_90,In_486);
or U4731 (N_4731,In_1259,In_1661);
nor U4732 (N_4732,In_775,In_418);
nand U4733 (N_4733,In_1927,In_1096);
nor U4734 (N_4734,In_752,In_699);
nor U4735 (N_4735,In_419,In_2791);
xnor U4736 (N_4736,In_1051,In_277);
and U4737 (N_4737,In_1041,In_2124);
xor U4738 (N_4738,In_1696,In_615);
nor U4739 (N_4739,In_2578,In_1592);
nor U4740 (N_4740,In_1548,In_2853);
nor U4741 (N_4741,In_513,In_946);
nand U4742 (N_4742,In_2447,In_1706);
and U4743 (N_4743,In_925,In_2217);
and U4744 (N_4744,In_1434,In_1131);
or U4745 (N_4745,In_1947,In_1137);
xnor U4746 (N_4746,In_756,In_2908);
nand U4747 (N_4747,In_2343,In_499);
xnor U4748 (N_4748,In_1445,In_2292);
nand U4749 (N_4749,In_113,In_273);
nor U4750 (N_4750,In_2952,In_2945);
or U4751 (N_4751,In_2506,In_2309);
xor U4752 (N_4752,In_1769,In_2409);
and U4753 (N_4753,In_456,In_1503);
nand U4754 (N_4754,In_687,In_51);
nor U4755 (N_4755,In_2728,In_270);
and U4756 (N_4756,In_433,In_2069);
xnor U4757 (N_4757,In_940,In_572);
or U4758 (N_4758,In_1685,In_545);
or U4759 (N_4759,In_2211,In_337);
and U4760 (N_4760,In_2008,In_1765);
nand U4761 (N_4761,In_2349,In_409);
nand U4762 (N_4762,In_1736,In_2402);
or U4763 (N_4763,In_175,In_2899);
nor U4764 (N_4764,In_915,In_2937);
nor U4765 (N_4765,In_73,In_1224);
nor U4766 (N_4766,In_217,In_2600);
xor U4767 (N_4767,In_32,In_2448);
nand U4768 (N_4768,In_372,In_761);
nor U4769 (N_4769,In_2656,In_1010);
nand U4770 (N_4770,In_1529,In_2054);
nand U4771 (N_4771,In_1792,In_1916);
xnor U4772 (N_4772,In_1903,In_556);
or U4773 (N_4773,In_2324,In_578);
xor U4774 (N_4774,In_1412,In_1232);
xnor U4775 (N_4775,In_908,In_1539);
xnor U4776 (N_4776,In_1584,In_1368);
nand U4777 (N_4777,In_220,In_164);
nor U4778 (N_4778,In_2872,In_1673);
nand U4779 (N_4779,In_340,In_762);
and U4780 (N_4780,In_2018,In_1428);
nor U4781 (N_4781,In_2120,In_1038);
xor U4782 (N_4782,In_688,In_2630);
xnor U4783 (N_4783,In_98,In_2765);
nand U4784 (N_4784,In_673,In_374);
nor U4785 (N_4785,In_2929,In_2265);
and U4786 (N_4786,In_2112,In_2267);
xor U4787 (N_4787,In_2419,In_475);
nand U4788 (N_4788,In_153,In_1191);
or U4789 (N_4789,In_542,In_1397);
xor U4790 (N_4790,In_118,In_229);
and U4791 (N_4791,In_847,In_1781);
xnor U4792 (N_4792,In_1977,In_2091);
nand U4793 (N_4793,In_2559,In_1548);
nor U4794 (N_4794,In_2528,In_543);
or U4795 (N_4795,In_2267,In_712);
nand U4796 (N_4796,In_222,In_2866);
and U4797 (N_4797,In_805,In_1918);
nor U4798 (N_4798,In_2989,In_649);
nand U4799 (N_4799,In_2585,In_2913);
and U4800 (N_4800,In_1958,In_2937);
nand U4801 (N_4801,In_2173,In_1210);
nor U4802 (N_4802,In_1816,In_322);
nand U4803 (N_4803,In_2123,In_1915);
nand U4804 (N_4804,In_2934,In_2472);
xor U4805 (N_4805,In_1728,In_556);
nand U4806 (N_4806,In_1723,In_382);
xnor U4807 (N_4807,In_2841,In_1930);
xor U4808 (N_4808,In_1664,In_2476);
nand U4809 (N_4809,In_1075,In_2732);
and U4810 (N_4810,In_2210,In_30);
nor U4811 (N_4811,In_200,In_2902);
nand U4812 (N_4812,In_2714,In_600);
and U4813 (N_4813,In_1015,In_502);
xnor U4814 (N_4814,In_479,In_319);
or U4815 (N_4815,In_2371,In_1272);
xor U4816 (N_4816,In_2760,In_2142);
xor U4817 (N_4817,In_1815,In_874);
or U4818 (N_4818,In_2653,In_1495);
and U4819 (N_4819,In_1499,In_406);
and U4820 (N_4820,In_1399,In_1417);
or U4821 (N_4821,In_1891,In_2143);
or U4822 (N_4822,In_146,In_104);
nor U4823 (N_4823,In_26,In_2418);
nor U4824 (N_4824,In_531,In_2024);
nand U4825 (N_4825,In_2796,In_237);
xnor U4826 (N_4826,In_1811,In_2367);
or U4827 (N_4827,In_9,In_862);
xnor U4828 (N_4828,In_1678,In_2090);
or U4829 (N_4829,In_2537,In_1850);
nand U4830 (N_4830,In_1699,In_2990);
nand U4831 (N_4831,In_2593,In_1929);
and U4832 (N_4832,In_863,In_2509);
nor U4833 (N_4833,In_2662,In_17);
nor U4834 (N_4834,In_1348,In_2291);
xor U4835 (N_4835,In_311,In_753);
nor U4836 (N_4836,In_1659,In_1268);
and U4837 (N_4837,In_903,In_284);
or U4838 (N_4838,In_1792,In_1511);
or U4839 (N_4839,In_1670,In_638);
xnor U4840 (N_4840,In_1933,In_2894);
nand U4841 (N_4841,In_1027,In_1638);
xor U4842 (N_4842,In_1478,In_2013);
nor U4843 (N_4843,In_1321,In_2231);
or U4844 (N_4844,In_2682,In_49);
and U4845 (N_4845,In_2821,In_1749);
and U4846 (N_4846,In_784,In_1708);
and U4847 (N_4847,In_422,In_2198);
nor U4848 (N_4848,In_538,In_2305);
nor U4849 (N_4849,In_2532,In_2104);
and U4850 (N_4850,In_2462,In_2795);
and U4851 (N_4851,In_2506,In_2692);
xnor U4852 (N_4852,In_1530,In_311);
nor U4853 (N_4853,In_1795,In_2644);
nand U4854 (N_4854,In_520,In_1009);
and U4855 (N_4855,In_1306,In_135);
and U4856 (N_4856,In_553,In_1504);
and U4857 (N_4857,In_181,In_1764);
or U4858 (N_4858,In_70,In_883);
and U4859 (N_4859,In_774,In_2151);
nor U4860 (N_4860,In_2161,In_2135);
nor U4861 (N_4861,In_1136,In_1842);
nor U4862 (N_4862,In_2493,In_1512);
nor U4863 (N_4863,In_2604,In_944);
nor U4864 (N_4864,In_191,In_710);
and U4865 (N_4865,In_832,In_2793);
or U4866 (N_4866,In_2792,In_163);
and U4867 (N_4867,In_1681,In_1036);
nand U4868 (N_4868,In_2152,In_1851);
xor U4869 (N_4869,In_448,In_17);
or U4870 (N_4870,In_2460,In_1435);
nand U4871 (N_4871,In_610,In_2655);
xnor U4872 (N_4872,In_1495,In_1043);
or U4873 (N_4873,In_628,In_1364);
nor U4874 (N_4874,In_268,In_990);
nor U4875 (N_4875,In_2528,In_497);
and U4876 (N_4876,In_137,In_1502);
and U4877 (N_4877,In_2273,In_560);
nor U4878 (N_4878,In_536,In_1667);
nor U4879 (N_4879,In_1768,In_1359);
xor U4880 (N_4880,In_2413,In_1465);
and U4881 (N_4881,In_2380,In_2097);
xor U4882 (N_4882,In_1254,In_2428);
xor U4883 (N_4883,In_2031,In_1529);
nor U4884 (N_4884,In_298,In_2165);
nor U4885 (N_4885,In_1014,In_1845);
nor U4886 (N_4886,In_1521,In_1674);
xor U4887 (N_4887,In_2878,In_2710);
nand U4888 (N_4888,In_1197,In_2659);
nor U4889 (N_4889,In_1159,In_355);
xnor U4890 (N_4890,In_108,In_1982);
xnor U4891 (N_4891,In_1538,In_646);
nand U4892 (N_4892,In_1644,In_2571);
nor U4893 (N_4893,In_2391,In_399);
nor U4894 (N_4894,In_1173,In_2390);
nand U4895 (N_4895,In_175,In_2874);
xor U4896 (N_4896,In_852,In_2361);
nand U4897 (N_4897,In_1030,In_2212);
nand U4898 (N_4898,In_109,In_2150);
xnor U4899 (N_4899,In_622,In_2085);
xnor U4900 (N_4900,In_2755,In_1982);
nand U4901 (N_4901,In_681,In_2904);
or U4902 (N_4902,In_41,In_17);
and U4903 (N_4903,In_204,In_1309);
or U4904 (N_4904,In_1112,In_2764);
or U4905 (N_4905,In_2562,In_308);
and U4906 (N_4906,In_232,In_1546);
nand U4907 (N_4907,In_1479,In_1450);
nand U4908 (N_4908,In_773,In_2364);
xor U4909 (N_4909,In_2040,In_1474);
xor U4910 (N_4910,In_2590,In_1551);
xnor U4911 (N_4911,In_1155,In_2508);
xor U4912 (N_4912,In_952,In_2443);
or U4913 (N_4913,In_215,In_2707);
nor U4914 (N_4914,In_2467,In_1322);
or U4915 (N_4915,In_2329,In_865);
and U4916 (N_4916,In_1434,In_2955);
xor U4917 (N_4917,In_388,In_1493);
and U4918 (N_4918,In_2729,In_929);
or U4919 (N_4919,In_899,In_410);
and U4920 (N_4920,In_1987,In_2817);
and U4921 (N_4921,In_1500,In_970);
xnor U4922 (N_4922,In_2430,In_738);
and U4923 (N_4923,In_2432,In_1939);
and U4924 (N_4924,In_1736,In_2418);
or U4925 (N_4925,In_391,In_371);
and U4926 (N_4926,In_1212,In_299);
xor U4927 (N_4927,In_640,In_2456);
nand U4928 (N_4928,In_2231,In_581);
xnor U4929 (N_4929,In_2780,In_2628);
nor U4930 (N_4930,In_1316,In_1848);
nor U4931 (N_4931,In_2550,In_397);
nor U4932 (N_4932,In_351,In_932);
nor U4933 (N_4933,In_1802,In_917);
or U4934 (N_4934,In_2041,In_1680);
nand U4935 (N_4935,In_1311,In_2123);
nor U4936 (N_4936,In_106,In_1836);
and U4937 (N_4937,In_2710,In_2182);
and U4938 (N_4938,In_345,In_270);
or U4939 (N_4939,In_2095,In_1514);
nor U4940 (N_4940,In_1779,In_721);
nor U4941 (N_4941,In_1110,In_1268);
nor U4942 (N_4942,In_194,In_1009);
nor U4943 (N_4943,In_198,In_676);
xnor U4944 (N_4944,In_862,In_815);
and U4945 (N_4945,In_385,In_2684);
and U4946 (N_4946,In_2008,In_228);
nand U4947 (N_4947,In_569,In_159);
nand U4948 (N_4948,In_1185,In_1830);
or U4949 (N_4949,In_464,In_2472);
xor U4950 (N_4950,In_1697,In_2999);
and U4951 (N_4951,In_2489,In_594);
xor U4952 (N_4952,In_371,In_1444);
nand U4953 (N_4953,In_2191,In_29);
or U4954 (N_4954,In_421,In_1752);
or U4955 (N_4955,In_970,In_1060);
nand U4956 (N_4956,In_2949,In_1562);
and U4957 (N_4957,In_2539,In_466);
nor U4958 (N_4958,In_1162,In_499);
xor U4959 (N_4959,In_731,In_2914);
nor U4960 (N_4960,In_284,In_1776);
nor U4961 (N_4961,In_2352,In_2928);
or U4962 (N_4962,In_1147,In_785);
nand U4963 (N_4963,In_2995,In_1427);
and U4964 (N_4964,In_2407,In_556);
xnor U4965 (N_4965,In_861,In_1631);
and U4966 (N_4966,In_2452,In_81);
xnor U4967 (N_4967,In_2375,In_1527);
or U4968 (N_4968,In_2115,In_219);
or U4969 (N_4969,In_2529,In_767);
nor U4970 (N_4970,In_355,In_1919);
xnor U4971 (N_4971,In_1784,In_639);
or U4972 (N_4972,In_2517,In_701);
and U4973 (N_4973,In_86,In_1001);
or U4974 (N_4974,In_2495,In_1625);
or U4975 (N_4975,In_1505,In_488);
or U4976 (N_4976,In_2237,In_2065);
or U4977 (N_4977,In_2007,In_2774);
xnor U4978 (N_4978,In_476,In_1888);
nor U4979 (N_4979,In_2519,In_2453);
and U4980 (N_4980,In_2076,In_520);
nand U4981 (N_4981,In_133,In_219);
nor U4982 (N_4982,In_2338,In_110);
nand U4983 (N_4983,In_2443,In_2249);
xnor U4984 (N_4984,In_940,In_1887);
nor U4985 (N_4985,In_710,In_1769);
and U4986 (N_4986,In_1309,In_1292);
nor U4987 (N_4987,In_1609,In_1617);
xor U4988 (N_4988,In_2715,In_1745);
xor U4989 (N_4989,In_2788,In_538);
nor U4990 (N_4990,In_1078,In_2865);
or U4991 (N_4991,In_981,In_881);
or U4992 (N_4992,In_1836,In_2043);
nor U4993 (N_4993,In_794,In_1270);
nor U4994 (N_4994,In_995,In_459);
and U4995 (N_4995,In_2189,In_1976);
nor U4996 (N_4996,In_1703,In_2789);
and U4997 (N_4997,In_821,In_2689);
nor U4998 (N_4998,In_1290,In_2391);
xnor U4999 (N_4999,In_656,In_1594);
xnor U5000 (N_5000,In_2986,In_282);
xor U5001 (N_5001,In_377,In_51);
nand U5002 (N_5002,In_35,In_749);
nor U5003 (N_5003,In_611,In_923);
and U5004 (N_5004,In_17,In_2402);
nand U5005 (N_5005,In_1330,In_558);
nor U5006 (N_5006,In_1951,In_2137);
nand U5007 (N_5007,In_2395,In_275);
or U5008 (N_5008,In_2262,In_378);
nor U5009 (N_5009,In_493,In_1353);
nand U5010 (N_5010,In_1012,In_1021);
or U5011 (N_5011,In_1790,In_2659);
or U5012 (N_5012,In_2841,In_2930);
xnor U5013 (N_5013,In_2184,In_2978);
xnor U5014 (N_5014,In_267,In_893);
nand U5015 (N_5015,In_937,In_2490);
and U5016 (N_5016,In_2775,In_1710);
nor U5017 (N_5017,In_225,In_2273);
xnor U5018 (N_5018,In_1734,In_2155);
nor U5019 (N_5019,In_405,In_2225);
and U5020 (N_5020,In_168,In_140);
xor U5021 (N_5021,In_1025,In_593);
nand U5022 (N_5022,In_1216,In_237);
nand U5023 (N_5023,In_1415,In_1223);
or U5024 (N_5024,In_1208,In_1893);
xnor U5025 (N_5025,In_858,In_2610);
or U5026 (N_5026,In_2288,In_1047);
and U5027 (N_5027,In_2454,In_2213);
nor U5028 (N_5028,In_2810,In_1577);
or U5029 (N_5029,In_2117,In_2426);
and U5030 (N_5030,In_1935,In_888);
and U5031 (N_5031,In_2292,In_1024);
or U5032 (N_5032,In_684,In_2428);
or U5033 (N_5033,In_1308,In_2732);
and U5034 (N_5034,In_705,In_1807);
and U5035 (N_5035,In_515,In_1278);
nor U5036 (N_5036,In_836,In_665);
nand U5037 (N_5037,In_1213,In_1718);
nor U5038 (N_5038,In_2104,In_259);
nor U5039 (N_5039,In_2224,In_670);
nand U5040 (N_5040,In_2697,In_1050);
nor U5041 (N_5041,In_871,In_625);
nand U5042 (N_5042,In_481,In_2268);
and U5043 (N_5043,In_1453,In_2166);
and U5044 (N_5044,In_2071,In_2097);
xnor U5045 (N_5045,In_2525,In_792);
nor U5046 (N_5046,In_2725,In_1296);
and U5047 (N_5047,In_1512,In_1769);
and U5048 (N_5048,In_2640,In_2535);
nor U5049 (N_5049,In_738,In_731);
xnor U5050 (N_5050,In_739,In_542);
xor U5051 (N_5051,In_378,In_940);
xnor U5052 (N_5052,In_359,In_832);
and U5053 (N_5053,In_1610,In_824);
or U5054 (N_5054,In_1145,In_2698);
xor U5055 (N_5055,In_1119,In_1091);
xor U5056 (N_5056,In_360,In_2914);
nor U5057 (N_5057,In_2794,In_2192);
xnor U5058 (N_5058,In_2815,In_646);
nand U5059 (N_5059,In_153,In_1428);
nand U5060 (N_5060,In_912,In_607);
nor U5061 (N_5061,In_1390,In_2167);
nand U5062 (N_5062,In_2754,In_2330);
nand U5063 (N_5063,In_490,In_2784);
nor U5064 (N_5064,In_1321,In_2966);
and U5065 (N_5065,In_790,In_762);
nand U5066 (N_5066,In_1339,In_812);
nor U5067 (N_5067,In_121,In_1947);
or U5068 (N_5068,In_1591,In_921);
xnor U5069 (N_5069,In_2146,In_913);
xor U5070 (N_5070,In_2144,In_457);
nand U5071 (N_5071,In_129,In_2311);
and U5072 (N_5072,In_1791,In_2475);
or U5073 (N_5073,In_629,In_2910);
or U5074 (N_5074,In_1194,In_2694);
and U5075 (N_5075,In_2654,In_85);
nor U5076 (N_5076,In_2393,In_1744);
or U5077 (N_5077,In_525,In_853);
xnor U5078 (N_5078,In_1251,In_162);
nand U5079 (N_5079,In_1135,In_2218);
xnor U5080 (N_5080,In_1568,In_2441);
and U5081 (N_5081,In_317,In_998);
or U5082 (N_5082,In_956,In_1187);
nand U5083 (N_5083,In_1582,In_1649);
nor U5084 (N_5084,In_1503,In_825);
xnor U5085 (N_5085,In_2344,In_2671);
and U5086 (N_5086,In_2234,In_1652);
nand U5087 (N_5087,In_2467,In_2737);
or U5088 (N_5088,In_1303,In_2690);
and U5089 (N_5089,In_2859,In_2242);
nand U5090 (N_5090,In_590,In_2982);
or U5091 (N_5091,In_2837,In_2440);
or U5092 (N_5092,In_208,In_1792);
xnor U5093 (N_5093,In_1221,In_1651);
nand U5094 (N_5094,In_1653,In_1906);
and U5095 (N_5095,In_703,In_446);
or U5096 (N_5096,In_395,In_1598);
nor U5097 (N_5097,In_490,In_2042);
xor U5098 (N_5098,In_1496,In_2326);
or U5099 (N_5099,In_2432,In_2170);
nor U5100 (N_5100,In_1847,In_1039);
and U5101 (N_5101,In_1924,In_1607);
or U5102 (N_5102,In_2709,In_2324);
xor U5103 (N_5103,In_557,In_2349);
or U5104 (N_5104,In_1108,In_2059);
nor U5105 (N_5105,In_710,In_91);
xnor U5106 (N_5106,In_2469,In_601);
nand U5107 (N_5107,In_217,In_2172);
or U5108 (N_5108,In_1111,In_2849);
and U5109 (N_5109,In_2127,In_1741);
and U5110 (N_5110,In_2125,In_1280);
and U5111 (N_5111,In_1761,In_90);
xnor U5112 (N_5112,In_2714,In_2559);
xnor U5113 (N_5113,In_1322,In_2555);
xor U5114 (N_5114,In_1505,In_1994);
xnor U5115 (N_5115,In_481,In_869);
xnor U5116 (N_5116,In_2408,In_2004);
or U5117 (N_5117,In_636,In_594);
xor U5118 (N_5118,In_1021,In_513);
or U5119 (N_5119,In_1931,In_1338);
or U5120 (N_5120,In_2751,In_1669);
nand U5121 (N_5121,In_1437,In_1925);
nand U5122 (N_5122,In_1022,In_2960);
nand U5123 (N_5123,In_1759,In_2939);
nor U5124 (N_5124,In_1402,In_2596);
nor U5125 (N_5125,In_2782,In_640);
nor U5126 (N_5126,In_2707,In_2316);
nor U5127 (N_5127,In_1457,In_1404);
xnor U5128 (N_5128,In_2192,In_2530);
or U5129 (N_5129,In_549,In_133);
nand U5130 (N_5130,In_410,In_1459);
or U5131 (N_5131,In_2761,In_1430);
nand U5132 (N_5132,In_729,In_1859);
nor U5133 (N_5133,In_717,In_2605);
nand U5134 (N_5134,In_2005,In_2827);
nand U5135 (N_5135,In_1424,In_2429);
nor U5136 (N_5136,In_1050,In_1888);
or U5137 (N_5137,In_315,In_1628);
and U5138 (N_5138,In_2743,In_1812);
or U5139 (N_5139,In_1004,In_2259);
and U5140 (N_5140,In_2929,In_1685);
and U5141 (N_5141,In_2710,In_2551);
nand U5142 (N_5142,In_2753,In_1262);
or U5143 (N_5143,In_2442,In_105);
or U5144 (N_5144,In_480,In_2963);
and U5145 (N_5145,In_2120,In_834);
or U5146 (N_5146,In_623,In_2718);
or U5147 (N_5147,In_2397,In_2224);
nand U5148 (N_5148,In_1824,In_984);
or U5149 (N_5149,In_2262,In_466);
xnor U5150 (N_5150,In_1522,In_1670);
and U5151 (N_5151,In_174,In_405);
xor U5152 (N_5152,In_260,In_321);
and U5153 (N_5153,In_1781,In_1992);
nand U5154 (N_5154,In_1996,In_1092);
nand U5155 (N_5155,In_2677,In_2916);
or U5156 (N_5156,In_463,In_1671);
nand U5157 (N_5157,In_1506,In_1878);
nor U5158 (N_5158,In_1435,In_810);
xnor U5159 (N_5159,In_401,In_1843);
nand U5160 (N_5160,In_829,In_688);
nor U5161 (N_5161,In_887,In_1688);
nor U5162 (N_5162,In_532,In_906);
nor U5163 (N_5163,In_1587,In_1324);
and U5164 (N_5164,In_2192,In_1204);
and U5165 (N_5165,In_2563,In_262);
xnor U5166 (N_5166,In_803,In_1612);
nand U5167 (N_5167,In_1288,In_784);
and U5168 (N_5168,In_783,In_1016);
nor U5169 (N_5169,In_675,In_2932);
nor U5170 (N_5170,In_1365,In_2942);
nand U5171 (N_5171,In_404,In_1757);
nand U5172 (N_5172,In_777,In_2527);
and U5173 (N_5173,In_888,In_1068);
xor U5174 (N_5174,In_849,In_2214);
or U5175 (N_5175,In_2310,In_2828);
xor U5176 (N_5176,In_2413,In_837);
xor U5177 (N_5177,In_1768,In_2479);
xor U5178 (N_5178,In_1009,In_2217);
nor U5179 (N_5179,In_987,In_1648);
or U5180 (N_5180,In_2502,In_803);
and U5181 (N_5181,In_1411,In_2348);
xor U5182 (N_5182,In_479,In_23);
nand U5183 (N_5183,In_2161,In_2325);
nand U5184 (N_5184,In_1896,In_2472);
nand U5185 (N_5185,In_2514,In_1797);
and U5186 (N_5186,In_1765,In_1848);
nand U5187 (N_5187,In_336,In_2665);
nor U5188 (N_5188,In_1394,In_2956);
nor U5189 (N_5189,In_203,In_555);
or U5190 (N_5190,In_499,In_2631);
and U5191 (N_5191,In_1321,In_2652);
or U5192 (N_5192,In_1976,In_232);
or U5193 (N_5193,In_89,In_518);
or U5194 (N_5194,In_479,In_830);
nand U5195 (N_5195,In_1442,In_1260);
nor U5196 (N_5196,In_1975,In_55);
and U5197 (N_5197,In_85,In_956);
nand U5198 (N_5198,In_1418,In_1100);
nand U5199 (N_5199,In_2276,In_1050);
xor U5200 (N_5200,In_2720,In_1063);
nor U5201 (N_5201,In_1041,In_1937);
nand U5202 (N_5202,In_1669,In_2755);
and U5203 (N_5203,In_165,In_63);
xnor U5204 (N_5204,In_1127,In_2762);
and U5205 (N_5205,In_12,In_371);
nor U5206 (N_5206,In_1100,In_492);
and U5207 (N_5207,In_100,In_1219);
nand U5208 (N_5208,In_1570,In_1108);
xnor U5209 (N_5209,In_2535,In_1267);
xor U5210 (N_5210,In_1481,In_592);
nand U5211 (N_5211,In_2737,In_2709);
or U5212 (N_5212,In_1574,In_2912);
xnor U5213 (N_5213,In_386,In_1264);
nor U5214 (N_5214,In_59,In_277);
xor U5215 (N_5215,In_2585,In_509);
xnor U5216 (N_5216,In_1764,In_1544);
xor U5217 (N_5217,In_1374,In_951);
nand U5218 (N_5218,In_850,In_2237);
nand U5219 (N_5219,In_1275,In_2931);
xnor U5220 (N_5220,In_1005,In_2403);
and U5221 (N_5221,In_2880,In_1508);
xnor U5222 (N_5222,In_1605,In_1932);
and U5223 (N_5223,In_2831,In_1415);
and U5224 (N_5224,In_2970,In_2109);
xnor U5225 (N_5225,In_2130,In_2221);
nor U5226 (N_5226,In_1232,In_2784);
nand U5227 (N_5227,In_1729,In_562);
nor U5228 (N_5228,In_241,In_1751);
or U5229 (N_5229,In_2313,In_2314);
nand U5230 (N_5230,In_2539,In_97);
xnor U5231 (N_5231,In_215,In_1899);
nor U5232 (N_5232,In_2448,In_2657);
xor U5233 (N_5233,In_2809,In_1449);
nand U5234 (N_5234,In_1098,In_1374);
nor U5235 (N_5235,In_1264,In_1368);
nor U5236 (N_5236,In_2116,In_1338);
and U5237 (N_5237,In_2026,In_2454);
xnor U5238 (N_5238,In_1510,In_781);
nand U5239 (N_5239,In_482,In_1075);
and U5240 (N_5240,In_2237,In_601);
and U5241 (N_5241,In_2354,In_2930);
xnor U5242 (N_5242,In_756,In_300);
and U5243 (N_5243,In_1078,In_1696);
xor U5244 (N_5244,In_1813,In_2221);
and U5245 (N_5245,In_408,In_46);
nor U5246 (N_5246,In_1693,In_818);
and U5247 (N_5247,In_1869,In_1568);
xnor U5248 (N_5248,In_820,In_139);
or U5249 (N_5249,In_1550,In_2007);
or U5250 (N_5250,In_555,In_235);
nor U5251 (N_5251,In_2481,In_1221);
and U5252 (N_5252,In_411,In_2233);
xor U5253 (N_5253,In_1856,In_1224);
or U5254 (N_5254,In_64,In_1967);
nor U5255 (N_5255,In_871,In_564);
and U5256 (N_5256,In_1403,In_2404);
or U5257 (N_5257,In_2058,In_2864);
and U5258 (N_5258,In_927,In_2761);
or U5259 (N_5259,In_1281,In_2117);
nand U5260 (N_5260,In_1390,In_785);
nand U5261 (N_5261,In_1858,In_2894);
and U5262 (N_5262,In_1743,In_2917);
nor U5263 (N_5263,In_618,In_280);
nand U5264 (N_5264,In_1241,In_930);
or U5265 (N_5265,In_302,In_2673);
or U5266 (N_5266,In_1343,In_2055);
nand U5267 (N_5267,In_1988,In_917);
xor U5268 (N_5268,In_2226,In_1517);
nand U5269 (N_5269,In_2348,In_1093);
or U5270 (N_5270,In_653,In_907);
nor U5271 (N_5271,In_873,In_206);
nand U5272 (N_5272,In_2649,In_1815);
nand U5273 (N_5273,In_1191,In_1698);
or U5274 (N_5274,In_660,In_1855);
or U5275 (N_5275,In_646,In_2967);
nor U5276 (N_5276,In_1874,In_2703);
or U5277 (N_5277,In_2893,In_1389);
and U5278 (N_5278,In_806,In_935);
or U5279 (N_5279,In_2323,In_1955);
or U5280 (N_5280,In_1421,In_1550);
or U5281 (N_5281,In_626,In_2601);
or U5282 (N_5282,In_1378,In_2207);
and U5283 (N_5283,In_1168,In_118);
nor U5284 (N_5284,In_173,In_2729);
nand U5285 (N_5285,In_1416,In_1486);
and U5286 (N_5286,In_222,In_448);
nor U5287 (N_5287,In_170,In_2984);
nor U5288 (N_5288,In_349,In_467);
and U5289 (N_5289,In_1334,In_961);
or U5290 (N_5290,In_2958,In_1521);
nor U5291 (N_5291,In_277,In_618);
and U5292 (N_5292,In_2039,In_1660);
nand U5293 (N_5293,In_1073,In_1671);
nand U5294 (N_5294,In_2302,In_1993);
nor U5295 (N_5295,In_1939,In_2675);
or U5296 (N_5296,In_769,In_558);
nor U5297 (N_5297,In_1199,In_1340);
xnor U5298 (N_5298,In_556,In_1600);
nor U5299 (N_5299,In_19,In_2054);
or U5300 (N_5300,In_2784,In_1943);
nor U5301 (N_5301,In_440,In_2148);
or U5302 (N_5302,In_2303,In_2219);
nand U5303 (N_5303,In_298,In_1880);
nor U5304 (N_5304,In_2049,In_587);
nand U5305 (N_5305,In_467,In_712);
xnor U5306 (N_5306,In_2518,In_572);
nand U5307 (N_5307,In_1108,In_1305);
xnor U5308 (N_5308,In_1332,In_1080);
nor U5309 (N_5309,In_1433,In_1776);
or U5310 (N_5310,In_2519,In_894);
or U5311 (N_5311,In_2149,In_2365);
or U5312 (N_5312,In_1910,In_1029);
xor U5313 (N_5313,In_876,In_828);
or U5314 (N_5314,In_246,In_82);
xnor U5315 (N_5315,In_1791,In_1695);
or U5316 (N_5316,In_2255,In_1495);
nand U5317 (N_5317,In_578,In_2848);
nand U5318 (N_5318,In_2654,In_487);
and U5319 (N_5319,In_2828,In_1905);
and U5320 (N_5320,In_2902,In_29);
and U5321 (N_5321,In_2572,In_1400);
xor U5322 (N_5322,In_538,In_1000);
and U5323 (N_5323,In_830,In_1240);
xnor U5324 (N_5324,In_606,In_864);
xnor U5325 (N_5325,In_1485,In_805);
nand U5326 (N_5326,In_1004,In_2785);
xnor U5327 (N_5327,In_1884,In_18);
and U5328 (N_5328,In_923,In_1622);
or U5329 (N_5329,In_161,In_1937);
nor U5330 (N_5330,In_446,In_1562);
nand U5331 (N_5331,In_2142,In_154);
nor U5332 (N_5332,In_511,In_2639);
and U5333 (N_5333,In_359,In_2981);
xnor U5334 (N_5334,In_1772,In_1002);
or U5335 (N_5335,In_1605,In_218);
nor U5336 (N_5336,In_1856,In_2168);
nor U5337 (N_5337,In_2341,In_2239);
nor U5338 (N_5338,In_965,In_950);
nand U5339 (N_5339,In_2344,In_737);
and U5340 (N_5340,In_462,In_2298);
xor U5341 (N_5341,In_730,In_1321);
nand U5342 (N_5342,In_366,In_2452);
and U5343 (N_5343,In_80,In_915);
nor U5344 (N_5344,In_2565,In_1624);
nand U5345 (N_5345,In_325,In_1411);
or U5346 (N_5346,In_654,In_520);
and U5347 (N_5347,In_343,In_1299);
or U5348 (N_5348,In_2987,In_729);
xnor U5349 (N_5349,In_1145,In_535);
nor U5350 (N_5350,In_1924,In_992);
nor U5351 (N_5351,In_273,In_914);
xor U5352 (N_5352,In_2995,In_868);
or U5353 (N_5353,In_1477,In_1843);
or U5354 (N_5354,In_265,In_2583);
xnor U5355 (N_5355,In_2415,In_1738);
or U5356 (N_5356,In_31,In_2987);
nor U5357 (N_5357,In_2258,In_37);
and U5358 (N_5358,In_974,In_2058);
nor U5359 (N_5359,In_625,In_2454);
and U5360 (N_5360,In_715,In_2024);
nor U5361 (N_5361,In_2576,In_416);
and U5362 (N_5362,In_2617,In_2628);
or U5363 (N_5363,In_1382,In_2901);
or U5364 (N_5364,In_175,In_2046);
or U5365 (N_5365,In_2897,In_1620);
and U5366 (N_5366,In_239,In_430);
or U5367 (N_5367,In_2565,In_1233);
xnor U5368 (N_5368,In_2223,In_1143);
xor U5369 (N_5369,In_1357,In_2354);
nor U5370 (N_5370,In_2510,In_1404);
and U5371 (N_5371,In_2831,In_104);
nor U5372 (N_5372,In_2787,In_2784);
nand U5373 (N_5373,In_921,In_372);
nand U5374 (N_5374,In_2134,In_2421);
and U5375 (N_5375,In_658,In_1213);
nor U5376 (N_5376,In_522,In_232);
and U5377 (N_5377,In_418,In_2805);
and U5378 (N_5378,In_2128,In_2928);
xor U5379 (N_5379,In_2519,In_2072);
xnor U5380 (N_5380,In_2618,In_1523);
xnor U5381 (N_5381,In_2503,In_2352);
or U5382 (N_5382,In_268,In_2633);
xnor U5383 (N_5383,In_2036,In_1348);
nor U5384 (N_5384,In_5,In_926);
and U5385 (N_5385,In_1974,In_2113);
xnor U5386 (N_5386,In_1183,In_2352);
or U5387 (N_5387,In_1653,In_1724);
xor U5388 (N_5388,In_1410,In_466);
xnor U5389 (N_5389,In_120,In_386);
nand U5390 (N_5390,In_1772,In_2105);
or U5391 (N_5391,In_1476,In_2397);
and U5392 (N_5392,In_1779,In_1392);
and U5393 (N_5393,In_216,In_1554);
nand U5394 (N_5394,In_2815,In_600);
nand U5395 (N_5395,In_2905,In_1133);
xor U5396 (N_5396,In_1293,In_387);
nand U5397 (N_5397,In_2304,In_1046);
nor U5398 (N_5398,In_2110,In_2101);
xnor U5399 (N_5399,In_2754,In_2097);
and U5400 (N_5400,In_2357,In_789);
and U5401 (N_5401,In_198,In_1759);
nand U5402 (N_5402,In_845,In_425);
or U5403 (N_5403,In_925,In_858);
and U5404 (N_5404,In_2122,In_2148);
and U5405 (N_5405,In_2562,In_2167);
nor U5406 (N_5406,In_2055,In_746);
nand U5407 (N_5407,In_114,In_1065);
xnor U5408 (N_5408,In_1637,In_790);
or U5409 (N_5409,In_1452,In_1601);
or U5410 (N_5410,In_877,In_1260);
or U5411 (N_5411,In_378,In_1649);
and U5412 (N_5412,In_1583,In_1669);
nor U5413 (N_5413,In_2903,In_1378);
xnor U5414 (N_5414,In_46,In_822);
or U5415 (N_5415,In_2442,In_1423);
nor U5416 (N_5416,In_1551,In_2341);
xor U5417 (N_5417,In_2421,In_440);
and U5418 (N_5418,In_905,In_86);
xnor U5419 (N_5419,In_1181,In_141);
and U5420 (N_5420,In_2375,In_1754);
nand U5421 (N_5421,In_2561,In_529);
and U5422 (N_5422,In_809,In_2673);
or U5423 (N_5423,In_2600,In_139);
xor U5424 (N_5424,In_207,In_1296);
nand U5425 (N_5425,In_1358,In_2696);
nand U5426 (N_5426,In_801,In_2035);
nor U5427 (N_5427,In_940,In_1303);
and U5428 (N_5428,In_1633,In_790);
and U5429 (N_5429,In_2183,In_1670);
nor U5430 (N_5430,In_567,In_1681);
nand U5431 (N_5431,In_1888,In_1488);
nor U5432 (N_5432,In_2048,In_2200);
nand U5433 (N_5433,In_2093,In_2036);
nand U5434 (N_5434,In_369,In_461);
and U5435 (N_5435,In_1933,In_517);
or U5436 (N_5436,In_2541,In_2217);
nand U5437 (N_5437,In_2873,In_1259);
or U5438 (N_5438,In_2730,In_2856);
nand U5439 (N_5439,In_1868,In_16);
nand U5440 (N_5440,In_1174,In_824);
xnor U5441 (N_5441,In_2359,In_1694);
nor U5442 (N_5442,In_2860,In_597);
nand U5443 (N_5443,In_1635,In_961);
nand U5444 (N_5444,In_47,In_539);
nor U5445 (N_5445,In_2977,In_2755);
nand U5446 (N_5446,In_688,In_2205);
or U5447 (N_5447,In_898,In_517);
xnor U5448 (N_5448,In_700,In_647);
nor U5449 (N_5449,In_166,In_2958);
and U5450 (N_5450,In_1376,In_2739);
nor U5451 (N_5451,In_2162,In_1097);
or U5452 (N_5452,In_1979,In_722);
nor U5453 (N_5453,In_637,In_1304);
and U5454 (N_5454,In_1943,In_2772);
xor U5455 (N_5455,In_86,In_2952);
nor U5456 (N_5456,In_2011,In_1091);
nand U5457 (N_5457,In_2657,In_188);
and U5458 (N_5458,In_1167,In_2135);
nor U5459 (N_5459,In_745,In_2661);
or U5460 (N_5460,In_2770,In_806);
and U5461 (N_5461,In_2591,In_2123);
nor U5462 (N_5462,In_73,In_1192);
xor U5463 (N_5463,In_627,In_1370);
nor U5464 (N_5464,In_2873,In_1082);
xor U5465 (N_5465,In_456,In_2508);
nand U5466 (N_5466,In_2619,In_1791);
nand U5467 (N_5467,In_2825,In_351);
or U5468 (N_5468,In_828,In_1682);
nand U5469 (N_5469,In_2332,In_1053);
or U5470 (N_5470,In_805,In_1211);
nand U5471 (N_5471,In_41,In_701);
nor U5472 (N_5472,In_2761,In_198);
and U5473 (N_5473,In_2678,In_2960);
nand U5474 (N_5474,In_2973,In_2968);
and U5475 (N_5475,In_2602,In_1137);
and U5476 (N_5476,In_2209,In_2190);
or U5477 (N_5477,In_850,In_2008);
nor U5478 (N_5478,In_1273,In_725);
and U5479 (N_5479,In_1958,In_333);
and U5480 (N_5480,In_2100,In_981);
and U5481 (N_5481,In_1834,In_2437);
nor U5482 (N_5482,In_2422,In_1720);
xor U5483 (N_5483,In_229,In_1754);
and U5484 (N_5484,In_2594,In_1146);
and U5485 (N_5485,In_1364,In_525);
nand U5486 (N_5486,In_191,In_1703);
and U5487 (N_5487,In_978,In_358);
xor U5488 (N_5488,In_501,In_950);
and U5489 (N_5489,In_2482,In_2847);
or U5490 (N_5490,In_2081,In_1633);
xnor U5491 (N_5491,In_646,In_2431);
or U5492 (N_5492,In_825,In_1924);
xnor U5493 (N_5493,In_1087,In_1715);
nand U5494 (N_5494,In_289,In_585);
or U5495 (N_5495,In_861,In_1365);
xor U5496 (N_5496,In_1342,In_2327);
xnor U5497 (N_5497,In_866,In_1236);
xnor U5498 (N_5498,In_358,In_801);
xor U5499 (N_5499,In_1087,In_215);
nor U5500 (N_5500,In_2974,In_2157);
xor U5501 (N_5501,In_1362,In_2389);
xor U5502 (N_5502,In_405,In_391);
and U5503 (N_5503,In_544,In_2243);
xnor U5504 (N_5504,In_1546,In_2149);
nor U5505 (N_5505,In_734,In_2990);
nand U5506 (N_5506,In_1120,In_6);
nor U5507 (N_5507,In_2940,In_2253);
and U5508 (N_5508,In_2805,In_481);
or U5509 (N_5509,In_1441,In_2499);
and U5510 (N_5510,In_2107,In_790);
or U5511 (N_5511,In_1088,In_2808);
and U5512 (N_5512,In_1773,In_1302);
nor U5513 (N_5513,In_1188,In_1580);
xor U5514 (N_5514,In_1233,In_2277);
nand U5515 (N_5515,In_754,In_2524);
and U5516 (N_5516,In_187,In_2073);
and U5517 (N_5517,In_1574,In_2091);
or U5518 (N_5518,In_161,In_737);
or U5519 (N_5519,In_840,In_2219);
and U5520 (N_5520,In_1433,In_470);
and U5521 (N_5521,In_540,In_749);
and U5522 (N_5522,In_1618,In_755);
or U5523 (N_5523,In_1403,In_2106);
or U5524 (N_5524,In_20,In_961);
or U5525 (N_5525,In_2456,In_527);
nor U5526 (N_5526,In_2927,In_977);
nor U5527 (N_5527,In_915,In_636);
nand U5528 (N_5528,In_1313,In_1179);
xor U5529 (N_5529,In_2353,In_112);
xnor U5530 (N_5530,In_1573,In_2314);
and U5531 (N_5531,In_205,In_44);
nand U5532 (N_5532,In_1321,In_134);
nand U5533 (N_5533,In_2043,In_2190);
nand U5534 (N_5534,In_1102,In_2482);
nand U5535 (N_5535,In_2440,In_30);
and U5536 (N_5536,In_1658,In_1095);
and U5537 (N_5537,In_323,In_43);
and U5538 (N_5538,In_1306,In_1496);
nand U5539 (N_5539,In_975,In_2404);
nor U5540 (N_5540,In_1277,In_2498);
and U5541 (N_5541,In_364,In_2327);
or U5542 (N_5542,In_211,In_1482);
and U5543 (N_5543,In_2094,In_1075);
xor U5544 (N_5544,In_2882,In_15);
xor U5545 (N_5545,In_1764,In_379);
nand U5546 (N_5546,In_2057,In_1681);
and U5547 (N_5547,In_452,In_1343);
nand U5548 (N_5548,In_1210,In_640);
or U5549 (N_5549,In_2630,In_548);
nand U5550 (N_5550,In_335,In_1544);
or U5551 (N_5551,In_176,In_243);
nor U5552 (N_5552,In_329,In_1065);
nand U5553 (N_5553,In_1471,In_82);
xor U5554 (N_5554,In_2707,In_2);
nand U5555 (N_5555,In_844,In_2478);
nand U5556 (N_5556,In_1149,In_1607);
and U5557 (N_5557,In_1579,In_1285);
or U5558 (N_5558,In_164,In_349);
nor U5559 (N_5559,In_995,In_2222);
nand U5560 (N_5560,In_1294,In_1571);
nor U5561 (N_5561,In_2389,In_2773);
nor U5562 (N_5562,In_1115,In_2837);
nor U5563 (N_5563,In_1279,In_271);
and U5564 (N_5564,In_500,In_775);
nor U5565 (N_5565,In_733,In_569);
nor U5566 (N_5566,In_2169,In_1486);
and U5567 (N_5567,In_1167,In_1892);
nand U5568 (N_5568,In_2928,In_1175);
or U5569 (N_5569,In_2063,In_84);
nor U5570 (N_5570,In_922,In_657);
nor U5571 (N_5571,In_923,In_1021);
and U5572 (N_5572,In_543,In_157);
nor U5573 (N_5573,In_1507,In_2566);
and U5574 (N_5574,In_2149,In_2148);
nor U5575 (N_5575,In_2019,In_2645);
or U5576 (N_5576,In_2709,In_1467);
nor U5577 (N_5577,In_336,In_633);
or U5578 (N_5578,In_1786,In_2392);
and U5579 (N_5579,In_2066,In_2799);
nand U5580 (N_5580,In_1394,In_2123);
xor U5581 (N_5581,In_999,In_2609);
xnor U5582 (N_5582,In_170,In_2225);
nand U5583 (N_5583,In_1953,In_343);
and U5584 (N_5584,In_2382,In_1365);
and U5585 (N_5585,In_365,In_2048);
xor U5586 (N_5586,In_237,In_3);
or U5587 (N_5587,In_1508,In_1525);
and U5588 (N_5588,In_2364,In_2905);
xnor U5589 (N_5589,In_2601,In_2505);
nor U5590 (N_5590,In_2990,In_2373);
and U5591 (N_5591,In_2807,In_1784);
nand U5592 (N_5592,In_987,In_2401);
xnor U5593 (N_5593,In_176,In_1945);
xnor U5594 (N_5594,In_1511,In_1666);
xnor U5595 (N_5595,In_1403,In_1949);
nor U5596 (N_5596,In_1364,In_1632);
nand U5597 (N_5597,In_157,In_2697);
or U5598 (N_5598,In_1889,In_234);
xor U5599 (N_5599,In_2023,In_369);
nand U5600 (N_5600,In_2519,In_350);
nor U5601 (N_5601,In_1894,In_686);
nor U5602 (N_5602,In_876,In_1729);
nor U5603 (N_5603,In_153,In_1048);
nor U5604 (N_5604,In_195,In_2276);
nor U5605 (N_5605,In_2878,In_1075);
nand U5606 (N_5606,In_1195,In_16);
and U5607 (N_5607,In_2220,In_1810);
or U5608 (N_5608,In_1714,In_2775);
nor U5609 (N_5609,In_167,In_259);
or U5610 (N_5610,In_1393,In_2004);
or U5611 (N_5611,In_2733,In_2894);
or U5612 (N_5612,In_1494,In_1116);
nor U5613 (N_5613,In_2910,In_2816);
nand U5614 (N_5614,In_1167,In_2531);
and U5615 (N_5615,In_1780,In_897);
nand U5616 (N_5616,In_1642,In_1005);
nand U5617 (N_5617,In_944,In_2957);
nor U5618 (N_5618,In_427,In_1803);
or U5619 (N_5619,In_1139,In_2177);
xnor U5620 (N_5620,In_1316,In_1449);
or U5621 (N_5621,In_389,In_1524);
or U5622 (N_5622,In_1251,In_808);
nor U5623 (N_5623,In_1558,In_1603);
nor U5624 (N_5624,In_846,In_1406);
nor U5625 (N_5625,In_1012,In_2968);
or U5626 (N_5626,In_194,In_1380);
nor U5627 (N_5627,In_620,In_2930);
nand U5628 (N_5628,In_1525,In_2411);
nand U5629 (N_5629,In_1887,In_1981);
nand U5630 (N_5630,In_1905,In_270);
or U5631 (N_5631,In_651,In_2916);
and U5632 (N_5632,In_655,In_361);
and U5633 (N_5633,In_1013,In_1704);
xor U5634 (N_5634,In_614,In_1646);
and U5635 (N_5635,In_2034,In_1540);
nor U5636 (N_5636,In_2485,In_2068);
xor U5637 (N_5637,In_106,In_1199);
nand U5638 (N_5638,In_2973,In_853);
nand U5639 (N_5639,In_1998,In_2591);
and U5640 (N_5640,In_1887,In_1685);
or U5641 (N_5641,In_1917,In_2863);
nand U5642 (N_5642,In_2722,In_908);
xnor U5643 (N_5643,In_1534,In_1799);
or U5644 (N_5644,In_1396,In_1355);
xnor U5645 (N_5645,In_2120,In_1199);
and U5646 (N_5646,In_1671,In_1737);
xnor U5647 (N_5647,In_1095,In_491);
nand U5648 (N_5648,In_1172,In_1548);
or U5649 (N_5649,In_2795,In_1083);
or U5650 (N_5650,In_1483,In_937);
nor U5651 (N_5651,In_2356,In_2440);
and U5652 (N_5652,In_2314,In_1801);
nand U5653 (N_5653,In_998,In_1527);
or U5654 (N_5654,In_1549,In_1011);
xnor U5655 (N_5655,In_2351,In_1040);
nand U5656 (N_5656,In_2127,In_2470);
xnor U5657 (N_5657,In_73,In_2027);
nor U5658 (N_5658,In_1506,In_1146);
nand U5659 (N_5659,In_1233,In_1456);
or U5660 (N_5660,In_1654,In_2640);
nand U5661 (N_5661,In_1082,In_1793);
and U5662 (N_5662,In_2471,In_798);
nor U5663 (N_5663,In_2159,In_1333);
nor U5664 (N_5664,In_2861,In_566);
or U5665 (N_5665,In_618,In_2925);
nand U5666 (N_5666,In_871,In_2709);
or U5667 (N_5667,In_2581,In_1337);
and U5668 (N_5668,In_2720,In_87);
xor U5669 (N_5669,In_579,In_1698);
nor U5670 (N_5670,In_1358,In_300);
xnor U5671 (N_5671,In_2609,In_2143);
and U5672 (N_5672,In_2780,In_2042);
and U5673 (N_5673,In_1009,In_2654);
nor U5674 (N_5674,In_1904,In_2001);
xor U5675 (N_5675,In_1533,In_857);
nand U5676 (N_5676,In_1896,In_979);
xor U5677 (N_5677,In_28,In_1570);
nor U5678 (N_5678,In_405,In_817);
nor U5679 (N_5679,In_961,In_1687);
nor U5680 (N_5680,In_20,In_1003);
nor U5681 (N_5681,In_1679,In_947);
nand U5682 (N_5682,In_51,In_121);
nand U5683 (N_5683,In_1484,In_210);
and U5684 (N_5684,In_2469,In_2333);
and U5685 (N_5685,In_1432,In_1486);
nand U5686 (N_5686,In_2129,In_2691);
xnor U5687 (N_5687,In_1479,In_381);
nand U5688 (N_5688,In_524,In_285);
nand U5689 (N_5689,In_141,In_2007);
nor U5690 (N_5690,In_1354,In_509);
and U5691 (N_5691,In_720,In_652);
xor U5692 (N_5692,In_1113,In_1376);
nor U5693 (N_5693,In_2338,In_303);
nand U5694 (N_5694,In_671,In_1554);
xnor U5695 (N_5695,In_203,In_465);
nor U5696 (N_5696,In_959,In_1965);
or U5697 (N_5697,In_936,In_2003);
and U5698 (N_5698,In_450,In_2643);
nor U5699 (N_5699,In_2269,In_331);
nand U5700 (N_5700,In_1055,In_2564);
nand U5701 (N_5701,In_1124,In_2212);
nor U5702 (N_5702,In_459,In_1300);
nor U5703 (N_5703,In_238,In_1903);
nand U5704 (N_5704,In_1017,In_2533);
or U5705 (N_5705,In_1838,In_2865);
nand U5706 (N_5706,In_1209,In_2208);
or U5707 (N_5707,In_191,In_1190);
or U5708 (N_5708,In_2350,In_649);
and U5709 (N_5709,In_1888,In_1212);
or U5710 (N_5710,In_664,In_1237);
nor U5711 (N_5711,In_2786,In_2788);
nand U5712 (N_5712,In_2417,In_972);
or U5713 (N_5713,In_544,In_652);
or U5714 (N_5714,In_1641,In_2797);
and U5715 (N_5715,In_2558,In_2157);
and U5716 (N_5716,In_7,In_2635);
nand U5717 (N_5717,In_1652,In_389);
xor U5718 (N_5718,In_2329,In_669);
nand U5719 (N_5719,In_1845,In_99);
and U5720 (N_5720,In_2613,In_2848);
or U5721 (N_5721,In_2107,In_283);
xor U5722 (N_5722,In_1660,In_642);
xnor U5723 (N_5723,In_2955,In_1143);
nor U5724 (N_5724,In_551,In_2706);
xor U5725 (N_5725,In_2686,In_2104);
or U5726 (N_5726,In_1355,In_1622);
or U5727 (N_5727,In_155,In_2561);
and U5728 (N_5728,In_1326,In_56);
nor U5729 (N_5729,In_2559,In_1451);
and U5730 (N_5730,In_252,In_2401);
nand U5731 (N_5731,In_758,In_43);
xnor U5732 (N_5732,In_2924,In_517);
nor U5733 (N_5733,In_1797,In_291);
or U5734 (N_5734,In_2906,In_1157);
nand U5735 (N_5735,In_2408,In_803);
or U5736 (N_5736,In_2393,In_1836);
or U5737 (N_5737,In_2435,In_2980);
xnor U5738 (N_5738,In_842,In_338);
and U5739 (N_5739,In_818,In_531);
or U5740 (N_5740,In_1629,In_483);
or U5741 (N_5741,In_461,In_336);
or U5742 (N_5742,In_1310,In_1572);
nand U5743 (N_5743,In_2978,In_639);
or U5744 (N_5744,In_2521,In_1867);
nor U5745 (N_5745,In_1262,In_992);
nand U5746 (N_5746,In_1054,In_117);
and U5747 (N_5747,In_825,In_2934);
or U5748 (N_5748,In_2107,In_2976);
xor U5749 (N_5749,In_2556,In_27);
or U5750 (N_5750,In_1916,In_376);
nor U5751 (N_5751,In_623,In_510);
xnor U5752 (N_5752,In_1233,In_844);
or U5753 (N_5753,In_2781,In_1345);
and U5754 (N_5754,In_2685,In_778);
nor U5755 (N_5755,In_1823,In_142);
and U5756 (N_5756,In_471,In_2368);
and U5757 (N_5757,In_2541,In_2827);
nor U5758 (N_5758,In_2302,In_1636);
nand U5759 (N_5759,In_1427,In_1839);
xor U5760 (N_5760,In_21,In_1270);
or U5761 (N_5761,In_1359,In_1666);
nor U5762 (N_5762,In_176,In_832);
nand U5763 (N_5763,In_425,In_944);
xnor U5764 (N_5764,In_2159,In_2351);
nand U5765 (N_5765,In_256,In_1125);
nand U5766 (N_5766,In_2322,In_2);
xnor U5767 (N_5767,In_2223,In_1511);
and U5768 (N_5768,In_41,In_1880);
nor U5769 (N_5769,In_1688,In_2850);
nor U5770 (N_5770,In_1429,In_2749);
or U5771 (N_5771,In_29,In_1883);
nand U5772 (N_5772,In_68,In_163);
and U5773 (N_5773,In_1702,In_2958);
and U5774 (N_5774,In_2831,In_2600);
nand U5775 (N_5775,In_1537,In_1472);
and U5776 (N_5776,In_2832,In_234);
and U5777 (N_5777,In_2591,In_538);
nor U5778 (N_5778,In_144,In_1459);
nor U5779 (N_5779,In_336,In_2152);
nor U5780 (N_5780,In_2089,In_141);
xnor U5781 (N_5781,In_2559,In_802);
xnor U5782 (N_5782,In_30,In_417);
and U5783 (N_5783,In_2004,In_2597);
nand U5784 (N_5784,In_1435,In_1035);
xor U5785 (N_5785,In_54,In_2038);
xor U5786 (N_5786,In_2606,In_2349);
nor U5787 (N_5787,In_1438,In_1046);
or U5788 (N_5788,In_2504,In_2090);
or U5789 (N_5789,In_818,In_745);
xnor U5790 (N_5790,In_1206,In_2910);
and U5791 (N_5791,In_72,In_1691);
xnor U5792 (N_5792,In_1448,In_418);
xor U5793 (N_5793,In_2024,In_2200);
nand U5794 (N_5794,In_429,In_1741);
nor U5795 (N_5795,In_615,In_1349);
nor U5796 (N_5796,In_851,In_2412);
nand U5797 (N_5797,In_2026,In_2407);
or U5798 (N_5798,In_826,In_1777);
and U5799 (N_5799,In_1290,In_274);
xor U5800 (N_5800,In_1101,In_2490);
nor U5801 (N_5801,In_1940,In_2343);
nor U5802 (N_5802,In_658,In_897);
xnor U5803 (N_5803,In_1825,In_2939);
nor U5804 (N_5804,In_2453,In_918);
xor U5805 (N_5805,In_1477,In_226);
nor U5806 (N_5806,In_790,In_2810);
nor U5807 (N_5807,In_2820,In_2662);
or U5808 (N_5808,In_909,In_26);
and U5809 (N_5809,In_12,In_1110);
or U5810 (N_5810,In_338,In_2875);
and U5811 (N_5811,In_1984,In_1971);
and U5812 (N_5812,In_396,In_124);
or U5813 (N_5813,In_2872,In_1458);
nor U5814 (N_5814,In_679,In_18);
and U5815 (N_5815,In_199,In_2504);
xnor U5816 (N_5816,In_713,In_2487);
nand U5817 (N_5817,In_2707,In_1585);
xnor U5818 (N_5818,In_2699,In_2465);
xor U5819 (N_5819,In_2726,In_379);
and U5820 (N_5820,In_2372,In_2482);
xor U5821 (N_5821,In_731,In_437);
nand U5822 (N_5822,In_2368,In_620);
nand U5823 (N_5823,In_776,In_903);
xor U5824 (N_5824,In_2313,In_763);
nand U5825 (N_5825,In_1562,In_622);
nand U5826 (N_5826,In_2666,In_810);
and U5827 (N_5827,In_2829,In_1633);
xnor U5828 (N_5828,In_496,In_1427);
or U5829 (N_5829,In_1470,In_1922);
and U5830 (N_5830,In_2913,In_1733);
and U5831 (N_5831,In_1873,In_174);
and U5832 (N_5832,In_1990,In_1898);
or U5833 (N_5833,In_654,In_2972);
or U5834 (N_5834,In_2633,In_145);
or U5835 (N_5835,In_2225,In_1);
xnor U5836 (N_5836,In_345,In_1569);
or U5837 (N_5837,In_2580,In_470);
nor U5838 (N_5838,In_602,In_2985);
and U5839 (N_5839,In_816,In_2515);
xnor U5840 (N_5840,In_294,In_1363);
and U5841 (N_5841,In_1664,In_1857);
nor U5842 (N_5842,In_1599,In_402);
xnor U5843 (N_5843,In_900,In_147);
and U5844 (N_5844,In_1752,In_1616);
xor U5845 (N_5845,In_446,In_454);
xnor U5846 (N_5846,In_1678,In_2010);
nor U5847 (N_5847,In_2168,In_34);
nand U5848 (N_5848,In_2552,In_2602);
nor U5849 (N_5849,In_890,In_754);
xnor U5850 (N_5850,In_1748,In_2030);
and U5851 (N_5851,In_589,In_2602);
and U5852 (N_5852,In_2110,In_2979);
xor U5853 (N_5853,In_2940,In_2004);
and U5854 (N_5854,In_1942,In_1693);
or U5855 (N_5855,In_48,In_1972);
xor U5856 (N_5856,In_2141,In_2134);
nand U5857 (N_5857,In_1777,In_2276);
nor U5858 (N_5858,In_799,In_1949);
nor U5859 (N_5859,In_1287,In_2174);
and U5860 (N_5860,In_116,In_1498);
or U5861 (N_5861,In_1740,In_2352);
nor U5862 (N_5862,In_2164,In_2509);
and U5863 (N_5863,In_954,In_1134);
or U5864 (N_5864,In_1117,In_1333);
nor U5865 (N_5865,In_2205,In_2027);
nand U5866 (N_5866,In_1374,In_676);
or U5867 (N_5867,In_2160,In_1699);
nor U5868 (N_5868,In_102,In_1721);
or U5869 (N_5869,In_2955,In_398);
nor U5870 (N_5870,In_1787,In_14);
nor U5871 (N_5871,In_1433,In_2878);
or U5872 (N_5872,In_2262,In_2733);
xor U5873 (N_5873,In_2953,In_1529);
nor U5874 (N_5874,In_1966,In_2498);
nor U5875 (N_5875,In_1236,In_2105);
or U5876 (N_5876,In_2895,In_587);
nor U5877 (N_5877,In_875,In_1487);
nor U5878 (N_5878,In_75,In_2129);
nand U5879 (N_5879,In_249,In_427);
nand U5880 (N_5880,In_1927,In_48);
xor U5881 (N_5881,In_1481,In_2947);
or U5882 (N_5882,In_2993,In_1039);
nand U5883 (N_5883,In_368,In_54);
or U5884 (N_5884,In_2193,In_2322);
nor U5885 (N_5885,In_430,In_2104);
nand U5886 (N_5886,In_2845,In_344);
nand U5887 (N_5887,In_1844,In_600);
xnor U5888 (N_5888,In_412,In_2333);
and U5889 (N_5889,In_1553,In_2054);
xnor U5890 (N_5890,In_2456,In_2880);
and U5891 (N_5891,In_1660,In_1411);
xor U5892 (N_5892,In_2406,In_1641);
xnor U5893 (N_5893,In_2999,In_1406);
xnor U5894 (N_5894,In_2988,In_520);
and U5895 (N_5895,In_2833,In_2852);
nand U5896 (N_5896,In_306,In_2804);
xor U5897 (N_5897,In_641,In_167);
nand U5898 (N_5898,In_363,In_1104);
xnor U5899 (N_5899,In_896,In_1540);
or U5900 (N_5900,In_175,In_2812);
xor U5901 (N_5901,In_17,In_1575);
and U5902 (N_5902,In_2181,In_1255);
xor U5903 (N_5903,In_1093,In_2967);
and U5904 (N_5904,In_329,In_602);
nand U5905 (N_5905,In_574,In_767);
or U5906 (N_5906,In_2255,In_2356);
and U5907 (N_5907,In_2020,In_2663);
xnor U5908 (N_5908,In_2117,In_1280);
or U5909 (N_5909,In_1946,In_1661);
or U5910 (N_5910,In_260,In_1464);
and U5911 (N_5911,In_727,In_525);
and U5912 (N_5912,In_793,In_1803);
and U5913 (N_5913,In_1229,In_2640);
xor U5914 (N_5914,In_2316,In_2259);
and U5915 (N_5915,In_2009,In_1519);
nor U5916 (N_5916,In_908,In_170);
nand U5917 (N_5917,In_1508,In_967);
nand U5918 (N_5918,In_501,In_128);
nor U5919 (N_5919,In_2960,In_4);
nand U5920 (N_5920,In_2039,In_68);
nand U5921 (N_5921,In_375,In_713);
xnor U5922 (N_5922,In_2979,In_1939);
or U5923 (N_5923,In_44,In_247);
nor U5924 (N_5924,In_2519,In_2767);
nor U5925 (N_5925,In_638,In_1840);
or U5926 (N_5926,In_2372,In_218);
or U5927 (N_5927,In_735,In_2111);
nor U5928 (N_5928,In_2170,In_141);
nand U5929 (N_5929,In_325,In_355);
or U5930 (N_5930,In_1969,In_699);
nor U5931 (N_5931,In_1242,In_332);
and U5932 (N_5932,In_1104,In_2);
nor U5933 (N_5933,In_2654,In_772);
and U5934 (N_5934,In_1841,In_241);
nor U5935 (N_5935,In_2431,In_128);
and U5936 (N_5936,In_776,In_2325);
xor U5937 (N_5937,In_1118,In_1028);
and U5938 (N_5938,In_1489,In_2719);
nand U5939 (N_5939,In_927,In_1681);
nand U5940 (N_5940,In_1814,In_917);
nor U5941 (N_5941,In_10,In_1337);
nand U5942 (N_5942,In_367,In_1048);
nor U5943 (N_5943,In_515,In_800);
nand U5944 (N_5944,In_1698,In_2987);
nor U5945 (N_5945,In_2991,In_879);
or U5946 (N_5946,In_189,In_545);
xnor U5947 (N_5947,In_563,In_1709);
and U5948 (N_5948,In_1520,In_2470);
and U5949 (N_5949,In_71,In_431);
xnor U5950 (N_5950,In_2258,In_942);
xnor U5951 (N_5951,In_2090,In_761);
or U5952 (N_5952,In_1985,In_28);
nand U5953 (N_5953,In_325,In_1518);
and U5954 (N_5954,In_1009,In_2704);
or U5955 (N_5955,In_1324,In_2859);
nor U5956 (N_5956,In_1601,In_792);
nand U5957 (N_5957,In_614,In_2096);
xor U5958 (N_5958,In_1269,In_1604);
xor U5959 (N_5959,In_2623,In_1923);
or U5960 (N_5960,In_2238,In_2163);
nand U5961 (N_5961,In_889,In_2005);
nand U5962 (N_5962,In_1496,In_408);
and U5963 (N_5963,In_2879,In_111);
nand U5964 (N_5964,In_2741,In_2114);
nor U5965 (N_5965,In_683,In_2658);
nand U5966 (N_5966,In_2344,In_915);
and U5967 (N_5967,In_200,In_1623);
xnor U5968 (N_5968,In_1416,In_1832);
nor U5969 (N_5969,In_2190,In_1280);
and U5970 (N_5970,In_2867,In_1540);
nor U5971 (N_5971,In_1405,In_1644);
and U5972 (N_5972,In_2683,In_2885);
xnor U5973 (N_5973,In_721,In_1538);
nand U5974 (N_5974,In_638,In_2497);
or U5975 (N_5975,In_180,In_1794);
nor U5976 (N_5976,In_1547,In_1356);
or U5977 (N_5977,In_1932,In_2187);
xor U5978 (N_5978,In_951,In_1407);
and U5979 (N_5979,In_205,In_672);
nor U5980 (N_5980,In_2477,In_2658);
nor U5981 (N_5981,In_715,In_2809);
nor U5982 (N_5982,In_831,In_2818);
and U5983 (N_5983,In_1973,In_2085);
nor U5984 (N_5984,In_2111,In_37);
or U5985 (N_5985,In_1905,In_767);
nor U5986 (N_5986,In_392,In_623);
nand U5987 (N_5987,In_77,In_1359);
xnor U5988 (N_5988,In_40,In_585);
and U5989 (N_5989,In_881,In_2492);
and U5990 (N_5990,In_2701,In_1172);
or U5991 (N_5991,In_1778,In_2576);
nor U5992 (N_5992,In_924,In_236);
or U5993 (N_5993,In_724,In_2358);
and U5994 (N_5994,In_415,In_1809);
nor U5995 (N_5995,In_706,In_560);
xnor U5996 (N_5996,In_2050,In_1083);
nor U5997 (N_5997,In_1944,In_90);
nand U5998 (N_5998,In_1822,In_1115);
nor U5999 (N_5999,In_333,In_256);
xor U6000 (N_6000,N_1981,N_830);
or U6001 (N_6001,N_1587,N_2478);
xnor U6002 (N_6002,N_931,N_921);
nor U6003 (N_6003,N_2625,N_1711);
and U6004 (N_6004,N_4859,N_0);
and U6005 (N_6005,N_1624,N_982);
or U6006 (N_6006,N_4076,N_486);
and U6007 (N_6007,N_3262,N_2409);
nand U6008 (N_6008,N_3434,N_1382);
or U6009 (N_6009,N_1143,N_5518);
or U6010 (N_6010,N_1815,N_5758);
nand U6011 (N_6011,N_1511,N_2814);
or U6012 (N_6012,N_4569,N_4712);
nor U6013 (N_6013,N_1034,N_5702);
or U6014 (N_6014,N_5210,N_5485);
and U6015 (N_6015,N_4243,N_3244);
and U6016 (N_6016,N_5155,N_3046);
nand U6017 (N_6017,N_2595,N_5587);
nor U6018 (N_6018,N_799,N_1144);
or U6019 (N_6019,N_29,N_2944);
xnor U6020 (N_6020,N_579,N_540);
and U6021 (N_6021,N_4265,N_1375);
and U6022 (N_6022,N_151,N_3934);
xor U6023 (N_6023,N_2018,N_1770);
nand U6024 (N_6024,N_1854,N_1191);
nand U6025 (N_6025,N_2060,N_1162);
nand U6026 (N_6026,N_5270,N_136);
xor U6027 (N_6027,N_3087,N_1556);
and U6028 (N_6028,N_4677,N_2330);
nand U6029 (N_6029,N_4074,N_4193);
xnor U6030 (N_6030,N_2370,N_4507);
nor U6031 (N_6031,N_3560,N_5173);
nor U6032 (N_6032,N_5068,N_108);
xor U6033 (N_6033,N_582,N_3701);
and U6034 (N_6034,N_5509,N_1812);
xnor U6035 (N_6035,N_2017,N_5062);
xnor U6036 (N_6036,N_1,N_2314);
nor U6037 (N_6037,N_1181,N_3731);
or U6038 (N_6038,N_3698,N_976);
nand U6039 (N_6039,N_5868,N_301);
nor U6040 (N_6040,N_1160,N_3117);
nand U6041 (N_6041,N_5902,N_2177);
or U6042 (N_6042,N_1709,N_490);
xor U6043 (N_6043,N_1544,N_2526);
and U6044 (N_6044,N_2262,N_2118);
nor U6045 (N_6045,N_1048,N_4828);
or U6046 (N_6046,N_1581,N_2766);
nand U6047 (N_6047,N_731,N_5054);
and U6048 (N_6048,N_1080,N_5601);
xor U6049 (N_6049,N_5424,N_4278);
xor U6050 (N_6050,N_5033,N_219);
nand U6051 (N_6051,N_4440,N_5167);
or U6052 (N_6052,N_1005,N_2214);
and U6053 (N_6053,N_5462,N_1203);
and U6054 (N_6054,N_891,N_5126);
nand U6055 (N_6055,N_4536,N_1920);
and U6056 (N_6056,N_3332,N_4852);
nor U6057 (N_6057,N_1280,N_4112);
nand U6058 (N_6058,N_1427,N_3660);
nor U6059 (N_6059,N_3475,N_1677);
and U6060 (N_6060,N_5002,N_1500);
or U6061 (N_6061,N_1007,N_2890);
or U6062 (N_6062,N_1460,N_3221);
nand U6063 (N_6063,N_3488,N_5675);
nor U6064 (N_6064,N_3596,N_1670);
xor U6065 (N_6065,N_824,N_3872);
or U6066 (N_6066,N_2534,N_2139);
nor U6067 (N_6067,N_558,N_4368);
nor U6068 (N_6068,N_4523,N_1692);
nand U6069 (N_6069,N_1602,N_2319);
nand U6070 (N_6070,N_1769,N_554);
nor U6071 (N_6071,N_1728,N_4558);
nor U6072 (N_6072,N_77,N_5076);
or U6073 (N_6073,N_2775,N_5171);
nand U6074 (N_6074,N_2398,N_3818);
nor U6075 (N_6075,N_1623,N_3792);
nand U6076 (N_6076,N_4402,N_5153);
or U6077 (N_6077,N_4079,N_5281);
or U6078 (N_6078,N_1644,N_2929);
xnor U6079 (N_6079,N_4018,N_5562);
and U6080 (N_6080,N_259,N_567);
xor U6081 (N_6081,N_60,N_1345);
or U6082 (N_6082,N_4660,N_362);
or U6083 (N_6083,N_263,N_648);
nand U6084 (N_6084,N_1618,N_2758);
or U6085 (N_6085,N_386,N_13);
nand U6086 (N_6086,N_1953,N_4474);
or U6087 (N_6087,N_2326,N_4101);
and U6088 (N_6088,N_2436,N_851);
xnor U6089 (N_6089,N_4605,N_2673);
and U6090 (N_6090,N_1204,N_2987);
nor U6091 (N_6091,N_4547,N_4966);
and U6092 (N_6092,N_389,N_1469);
nand U6093 (N_6093,N_2129,N_5012);
nor U6094 (N_6094,N_5266,N_1254);
xnor U6095 (N_6095,N_2980,N_3567);
nand U6096 (N_6096,N_5089,N_2873);
and U6097 (N_6097,N_1138,N_3176);
xnor U6098 (N_6098,N_3606,N_237);
xor U6099 (N_6099,N_2747,N_2298);
or U6100 (N_6100,N_1503,N_5788);
xor U6101 (N_6101,N_2631,N_1946);
and U6102 (N_6102,N_4465,N_5093);
or U6103 (N_6103,N_294,N_4103);
or U6104 (N_6104,N_5719,N_30);
nor U6105 (N_6105,N_2267,N_3507);
and U6106 (N_6106,N_4810,N_2296);
nor U6107 (N_6107,N_2040,N_5605);
nand U6108 (N_6108,N_1560,N_5347);
nand U6109 (N_6109,N_1439,N_1262);
nand U6110 (N_6110,N_5956,N_4630);
and U6111 (N_6111,N_1290,N_785);
or U6112 (N_6112,N_1908,N_2406);
nand U6113 (N_6113,N_2215,N_5236);
or U6114 (N_6114,N_3291,N_5638);
nand U6115 (N_6115,N_5559,N_4108);
and U6116 (N_6116,N_5438,N_1242);
or U6117 (N_6117,N_1317,N_1459);
and U6118 (N_6118,N_9,N_2710);
or U6119 (N_6119,N_680,N_875);
and U6120 (N_6120,N_5394,N_3530);
xnor U6121 (N_6121,N_5763,N_5691);
or U6122 (N_6122,N_5976,N_4053);
nor U6123 (N_6123,N_2049,N_804);
xnor U6124 (N_6124,N_2057,N_5551);
nand U6125 (N_6125,N_2071,N_4464);
nand U6126 (N_6126,N_491,N_5050);
nor U6127 (N_6127,N_3636,N_4177);
nand U6128 (N_6128,N_3785,N_5814);
and U6129 (N_6129,N_2759,N_2141);
nor U6130 (N_6130,N_1661,N_2044);
nand U6131 (N_6131,N_1348,N_2169);
and U6132 (N_6132,N_3398,N_5696);
or U6133 (N_6133,N_1287,N_4351);
or U6134 (N_6134,N_3566,N_275);
or U6135 (N_6135,N_3017,N_3749);
xor U6136 (N_6136,N_4151,N_4671);
or U6137 (N_6137,N_1286,N_3941);
and U6138 (N_6138,N_1790,N_3180);
nand U6139 (N_6139,N_723,N_171);
xor U6140 (N_6140,N_5795,N_2554);
nor U6141 (N_6141,N_2772,N_3406);
or U6142 (N_6142,N_2800,N_4403);
xor U6143 (N_6143,N_5287,N_250);
and U6144 (N_6144,N_3473,N_5538);
and U6145 (N_6145,N_285,N_4977);
or U6146 (N_6146,N_966,N_1111);
or U6147 (N_6147,N_2431,N_3524);
nand U6148 (N_6148,N_1893,N_1279);
or U6149 (N_6149,N_4651,N_3094);
nor U6150 (N_6150,N_334,N_3420);
xor U6151 (N_6151,N_5244,N_3597);
nand U6152 (N_6152,N_5196,N_3761);
nor U6153 (N_6153,N_4941,N_2425);
nand U6154 (N_6154,N_3718,N_69);
nor U6155 (N_6155,N_3512,N_3284);
nor U6156 (N_6156,N_2977,N_5824);
nand U6157 (N_6157,N_5521,N_5781);
or U6158 (N_6158,N_1697,N_4503);
or U6159 (N_6159,N_46,N_1185);
or U6160 (N_6160,N_699,N_2531);
nand U6161 (N_6161,N_4843,N_5880);
and U6162 (N_6162,N_2277,N_1918);
xnor U6163 (N_6163,N_5109,N_2972);
and U6164 (N_6164,N_4663,N_5860);
nand U6165 (N_6165,N_5930,N_5722);
and U6166 (N_6166,N_4531,N_4750);
nor U6167 (N_6167,N_172,N_5177);
nand U6168 (N_6168,N_1519,N_1258);
nor U6169 (N_6169,N_1473,N_462);
xnor U6170 (N_6170,N_1738,N_4580);
and U6171 (N_6171,N_188,N_3938);
and U6172 (N_6172,N_2206,N_1821);
and U6173 (N_6173,N_5227,N_5289);
nand U6174 (N_6174,N_194,N_2790);
and U6175 (N_6175,N_2802,N_3357);
nor U6176 (N_6176,N_4357,N_2995);
nand U6177 (N_6177,N_3447,N_2774);
nor U6178 (N_6178,N_3839,N_4428);
or U6179 (N_6179,N_4805,N_3353);
or U6180 (N_6180,N_5015,N_4506);
xor U6181 (N_6181,N_3271,N_1608);
xor U6182 (N_6182,N_1848,N_2811);
or U6183 (N_6183,N_1649,N_1452);
nand U6184 (N_6184,N_5871,N_3345);
xor U6185 (N_6185,N_1081,N_3364);
nand U6186 (N_6186,N_64,N_1958);
xor U6187 (N_6187,N_4945,N_3550);
or U6188 (N_6188,N_1320,N_4266);
or U6189 (N_6189,N_3769,N_5513);
and U6190 (N_6190,N_2852,N_1910);
and U6191 (N_6191,N_5494,N_4504);
nor U6192 (N_6192,N_2839,N_995);
nor U6193 (N_6193,N_2429,N_1036);
xnor U6194 (N_6194,N_2446,N_1593);
nand U6195 (N_6195,N_4946,N_434);
nor U6196 (N_6196,N_3456,N_1360);
and U6197 (N_6197,N_2463,N_873);
nand U6198 (N_6198,N_3562,N_459);
or U6199 (N_6199,N_1247,N_2764);
and U6200 (N_6200,N_4980,N_5129);
and U6201 (N_6201,N_4490,N_2809);
or U6202 (N_6202,N_305,N_3953);
nand U6203 (N_6203,N_1532,N_1078);
and U6204 (N_6204,N_3011,N_3181);
nand U6205 (N_6205,N_198,N_3788);
and U6206 (N_6206,N_2316,N_5903);
and U6207 (N_6207,N_2282,N_5712);
and U6208 (N_6208,N_4857,N_2638);
nand U6209 (N_6209,N_1917,N_5892);
nor U6210 (N_6210,N_1293,N_4114);
and U6211 (N_6211,N_2116,N_5476);
nor U6212 (N_6212,N_4466,N_4848);
nand U6213 (N_6213,N_779,N_1380);
nor U6214 (N_6214,N_2646,N_2936);
and U6215 (N_6215,N_4785,N_4856);
nor U6216 (N_6216,N_2850,N_5931);
or U6217 (N_6217,N_1391,N_414);
xor U6218 (N_6218,N_729,N_5773);
nor U6219 (N_6219,N_3754,N_5686);
and U6220 (N_6220,N_3423,N_1488);
nand U6221 (N_6221,N_5460,N_4756);
nor U6222 (N_6222,N_3464,N_3499);
and U6223 (N_6223,N_4839,N_2506);
xor U6224 (N_6224,N_4920,N_5957);
xor U6225 (N_6225,N_5853,N_4137);
and U6226 (N_6226,N_4253,N_3266);
xnor U6227 (N_6227,N_2942,N_1079);
or U6228 (N_6228,N_92,N_1495);
or U6229 (N_6229,N_569,N_4110);
or U6230 (N_6230,N_1625,N_4261);
nor U6231 (N_6231,N_4049,N_4325);
xor U6232 (N_6232,N_5350,N_1050);
xor U6233 (N_6233,N_979,N_1533);
nor U6234 (N_6234,N_3984,N_2097);
nand U6235 (N_6235,N_4821,N_913);
nor U6236 (N_6236,N_808,N_176);
xnor U6237 (N_6237,N_1827,N_3976);
xnor U6238 (N_6238,N_5046,N_3168);
or U6239 (N_6239,N_2461,N_2170);
or U6240 (N_6240,N_4827,N_4444);
nand U6241 (N_6241,N_5051,N_5679);
nand U6242 (N_6242,N_5664,N_1565);
nand U6243 (N_6243,N_2487,N_1127);
or U6244 (N_6244,N_4228,N_5900);
or U6245 (N_6245,N_2492,N_4701);
xor U6246 (N_6246,N_920,N_1850);
or U6247 (N_6247,N_4923,N_2163);
or U6248 (N_6248,N_5870,N_4426);
nor U6249 (N_6249,N_4885,N_159);
and U6250 (N_6250,N_3959,N_656);
and U6251 (N_6251,N_3838,N_2697);
nor U6252 (N_6252,N_812,N_3809);
or U6253 (N_6253,N_2223,N_694);
xnor U6254 (N_6254,N_2430,N_495);
xnor U6255 (N_6255,N_5962,N_3916);
or U6256 (N_6256,N_404,N_542);
nor U6257 (N_6257,N_1259,N_5989);
nor U6258 (N_6258,N_2975,N_5876);
and U6259 (N_6259,N_5571,N_2404);
nand U6260 (N_6260,N_1730,N_4284);
and U6261 (N_6261,N_872,N_1338);
and U6262 (N_6262,N_42,N_512);
xnor U6263 (N_6263,N_1870,N_3366);
or U6264 (N_6264,N_3091,N_1903);
nor U6265 (N_6265,N_955,N_4858);
and U6266 (N_6266,N_5934,N_4779);
and U6267 (N_6267,N_235,N_5443);
or U6268 (N_6268,N_4525,N_3051);
xnor U6269 (N_6269,N_4924,N_4639);
xnor U6270 (N_6270,N_3328,N_3449);
xor U6271 (N_6271,N_2469,N_1426);
xor U6272 (N_6272,N_3191,N_1887);
nand U6273 (N_6273,N_2205,N_3654);
xnor U6274 (N_6274,N_2901,N_2149);
xor U6275 (N_6275,N_5274,N_280);
xnor U6276 (N_6276,N_3248,N_4673);
or U6277 (N_6277,N_1582,N_3990);
nand U6278 (N_6278,N_911,N_2866);
xor U6279 (N_6279,N_4321,N_2145);
nor U6280 (N_6280,N_5854,N_1083);
and U6281 (N_6281,N_2922,N_3723);
or U6282 (N_6282,N_2034,N_5835);
or U6283 (N_6283,N_4005,N_3721);
or U6284 (N_6284,N_475,N_3173);
and U6285 (N_6285,N_820,N_2113);
or U6286 (N_6286,N_3707,N_5316);
nand U6287 (N_6287,N_5708,N_5831);
or U6288 (N_6288,N_701,N_4405);
xor U6289 (N_6289,N_3556,N_7);
xnor U6290 (N_6290,N_519,N_1970);
xnor U6291 (N_6291,N_4165,N_4058);
nor U6292 (N_6292,N_5657,N_3807);
and U6293 (N_6293,N_1808,N_4794);
or U6294 (N_6294,N_2843,N_2159);
and U6295 (N_6295,N_2609,N_4694);
nand U6296 (N_6296,N_5291,N_2066);
or U6297 (N_6297,N_5042,N_4290);
and U6298 (N_6298,N_5447,N_5586);
nand U6299 (N_6299,N_111,N_5604);
nor U6300 (N_6300,N_4851,N_4275);
and U6301 (N_6301,N_4086,N_1358);
and U6302 (N_6302,N_3012,N_4089);
and U6303 (N_6303,N_2791,N_5720);
xnor U6304 (N_6304,N_5371,N_719);
nand U6305 (N_6305,N_584,N_2105);
and U6306 (N_6306,N_1312,N_818);
or U6307 (N_6307,N_4695,N_2745);
nor U6308 (N_6308,N_2954,N_2119);
xor U6309 (N_6309,N_5410,N_2355);
and U6310 (N_6310,N_1678,N_1658);
xor U6311 (N_6311,N_1417,N_4755);
nand U6312 (N_6312,N_884,N_3431);
nand U6313 (N_6313,N_71,N_2310);
or U6314 (N_6314,N_1632,N_999);
xnor U6315 (N_6315,N_3511,N_114);
xnor U6316 (N_6316,N_959,N_2109);
and U6317 (N_6317,N_1629,N_3145);
and U6318 (N_6318,N_2700,N_3495);
nor U6319 (N_6319,N_4971,N_5417);
and U6320 (N_6320,N_737,N_3000);
xnor U6321 (N_6321,N_517,N_4668);
and U6322 (N_6322,N_187,N_591);
nand U6323 (N_6323,N_967,N_994);
nor U6324 (N_6324,N_1679,N_2629);
or U6325 (N_6325,N_315,N_4144);
xor U6326 (N_6326,N_4052,N_1039);
and U6327 (N_6327,N_5366,N_5941);
nor U6328 (N_6328,N_3160,N_5439);
and U6329 (N_6329,N_2108,N_2914);
or U6330 (N_6330,N_1789,N_2730);
nand U6331 (N_6331,N_541,N_397);
nor U6332 (N_6332,N_4667,N_1173);
and U6333 (N_6333,N_855,N_2668);
nand U6334 (N_6334,N_2965,N_5985);
nand U6335 (N_6335,N_5887,N_2252);
nand U6336 (N_6336,N_1364,N_5058);
or U6337 (N_6337,N_2867,N_261);
nor U6338 (N_6338,N_3622,N_5817);
xnor U6339 (N_6339,N_732,N_347);
or U6340 (N_6340,N_5631,N_2336);
nor U6341 (N_6341,N_1273,N_4907);
and U6342 (N_6342,N_2196,N_1156);
nor U6343 (N_6343,N_5241,N_321);
xor U6344 (N_6344,N_2473,N_3786);
or U6345 (N_6345,N_2880,N_1889);
xor U6346 (N_6346,N_5114,N_2447);
and U6347 (N_6347,N_3483,N_3368);
or U6348 (N_6348,N_1306,N_1218);
xnor U6349 (N_6349,N_2058,N_968);
or U6350 (N_6350,N_3086,N_2162);
and U6351 (N_6351,N_1357,N_3367);
nand U6352 (N_6352,N_1211,N_2333);
or U6353 (N_6353,N_5507,N_3529);
nand U6354 (N_6354,N_4943,N_2645);
and U6355 (N_6355,N_2357,N_2385);
xor U6356 (N_6356,N_5116,N_4831);
nand U6357 (N_6357,N_5212,N_2460);
nor U6358 (N_6358,N_721,N_2112);
nor U6359 (N_6359,N_1707,N_1121);
and U6360 (N_6360,N_2931,N_3480);
nand U6361 (N_6361,N_2517,N_2689);
and U6362 (N_6362,N_3847,N_599);
nand U6363 (N_6363,N_856,N_1455);
nand U6364 (N_6364,N_2382,N_5649);
xnor U6365 (N_6365,N_2321,N_2281);
nor U6366 (N_6366,N_3365,N_5841);
xnor U6367 (N_6367,N_2714,N_5425);
and U6368 (N_6368,N_3129,N_726);
nand U6369 (N_6369,N_5336,N_1101);
xnor U6370 (N_6370,N_4850,N_2648);
nor U6371 (N_6371,N_3477,N_3967);
or U6372 (N_6372,N_5774,N_496);
nor U6373 (N_6373,N_5967,N_12);
and U6374 (N_6374,N_2665,N_5181);
nor U6375 (N_6375,N_3664,N_3192);
or U6376 (N_6376,N_311,N_5437);
and U6377 (N_6377,N_4960,N_4216);
or U6378 (N_6378,N_2746,N_3358);
nor U6379 (N_6379,N_5688,N_3233);
nand U6380 (N_6380,N_4308,N_2172);
nand U6381 (N_6381,N_3432,N_2209);
and U6382 (N_6382,N_270,N_2219);
or U6383 (N_6383,N_5536,N_1368);
nand U6384 (N_6384,N_2821,N_3570);
or U6385 (N_6385,N_5827,N_4727);
nand U6386 (N_6386,N_2832,N_2426);
nand U6387 (N_6387,N_5749,N_381);
xor U6388 (N_6388,N_245,N_3049);
and U6389 (N_6389,N_21,N_3392);
or U6390 (N_6390,N_3092,N_2115);
and U6391 (N_6391,N_4925,N_5189);
nand U6392 (N_6392,N_5247,N_866);
nand U6393 (N_6393,N_4819,N_3790);
xnor U6394 (N_6394,N_4641,N_2982);
nor U6395 (N_6395,N_2963,N_3607);
nand U6396 (N_6396,N_2293,N_725);
nand U6397 (N_6397,N_2851,N_2588);
or U6398 (N_6398,N_3451,N_1952);
and U6399 (N_6399,N_1553,N_3558);
nand U6400 (N_6400,N_2846,N_3772);
nor U6401 (N_6401,N_2256,N_3155);
or U6402 (N_6402,N_122,N_2618);
or U6403 (N_6403,N_2120,N_1653);
and U6404 (N_6404,N_5359,N_3929);
nand U6405 (N_6405,N_5666,N_5319);
and U6406 (N_6406,N_2723,N_1001);
nor U6407 (N_6407,N_4397,N_1355);
nor U6408 (N_6408,N_3508,N_1588);
xor U6409 (N_6409,N_3819,N_536);
nor U6410 (N_6410,N_3068,N_438);
nand U6411 (N_6411,N_2073,N_3796);
and U6412 (N_6412,N_4807,N_1405);
and U6413 (N_6413,N_1209,N_593);
or U6414 (N_6414,N_1044,N_5807);
nor U6415 (N_6415,N_734,N_1786);
nand U6416 (N_6416,N_1841,N_2362);
or U6417 (N_6417,N_5678,N_5829);
nand U6418 (N_6418,N_1186,N_3797);
and U6419 (N_6419,N_2918,N_1717);
or U6420 (N_6420,N_877,N_1328);
and U6421 (N_6421,N_142,N_5326);
and U6422 (N_6422,N_4042,N_2221);
nor U6423 (N_6423,N_3513,N_1552);
nand U6424 (N_6424,N_1824,N_3459);
xor U6425 (N_6425,N_3518,N_4627);
nand U6426 (N_6426,N_4921,N_5743);
and U6427 (N_6427,N_1183,N_3982);
or U6428 (N_6428,N_5648,N_291);
nand U6429 (N_6429,N_402,N_3494);
nand U6430 (N_6430,N_3055,N_2713);
xnor U6431 (N_6431,N_4762,N_1929);
or U6432 (N_6432,N_70,N_248);
nor U6433 (N_6433,N_4524,N_2862);
nand U6434 (N_6434,N_3065,N_3167);
and U6435 (N_6435,N_174,N_5499);
or U6436 (N_6436,N_1112,N_5211);
or U6437 (N_6437,N_5305,N_3);
nor U6438 (N_6438,N_2468,N_3631);
xnor U6439 (N_6439,N_1558,N_276);
xor U6440 (N_6440,N_1289,N_786);
or U6441 (N_6441,N_303,N_1535);
xnor U6442 (N_6442,N_4720,N_5851);
and U6443 (N_6443,N_4272,N_2189);
nand U6444 (N_6444,N_3661,N_5088);
xor U6445 (N_6445,N_325,N_2284);
xnor U6446 (N_6446,N_5435,N_914);
nor U6447 (N_6447,N_2416,N_50);
nand U6448 (N_6448,N_4908,N_3439);
and U6449 (N_6449,N_4430,N_4407);
or U6450 (N_6450,N_4883,N_411);
or U6451 (N_6451,N_2919,N_1134);
xnor U6452 (N_6452,N_5428,N_5393);
xor U6453 (N_6453,N_4733,N_5919);
nor U6454 (N_6454,N_524,N_4961);
and U6455 (N_6455,N_5580,N_2796);
xnor U6456 (N_6456,N_346,N_1414);
nand U6457 (N_6457,N_5778,N_4223);
nor U6458 (N_6458,N_4586,N_2672);
and U6459 (N_6459,N_5409,N_5579);
xor U6460 (N_6460,N_5377,N_1818);
nor U6461 (N_6461,N_1806,N_5262);
nor U6462 (N_6462,N_3409,N_1170);
or U6463 (N_6463,N_484,N_2064);
and U6464 (N_6464,N_2892,N_2403);
xnor U6465 (N_6465,N_342,N_4860);
nand U6466 (N_6466,N_1626,N_2380);
and U6467 (N_6467,N_1387,N_1527);
and U6468 (N_6468,N_183,N_2444);
or U6469 (N_6469,N_4167,N_4476);
xor U6470 (N_6470,N_1294,N_4552);
nand U6471 (N_6471,N_2334,N_1187);
xor U6472 (N_6472,N_5429,N_2056);
xor U6473 (N_6473,N_2967,N_838);
and U6474 (N_6474,N_1480,N_5037);
or U6475 (N_6475,N_2653,N_3894);
nand U6476 (N_6476,N_868,N_146);
or U6477 (N_6477,N_4059,N_5195);
and U6478 (N_6478,N_2372,N_3540);
nor U6479 (N_6479,N_3583,N_1525);
or U6480 (N_6480,N_5286,N_278);
xor U6481 (N_6481,N_91,N_3768);
xnor U6482 (N_6482,N_4777,N_2146);
nor U6483 (N_6483,N_659,N_2973);
and U6484 (N_6484,N_5235,N_130);
or U6485 (N_6485,N_4502,N_1773);
and U6486 (N_6486,N_746,N_3214);
or U6487 (N_6487,N_1662,N_2369);
nand U6488 (N_6488,N_1809,N_5199);
nand U6489 (N_6489,N_4400,N_4380);
or U6490 (N_6490,N_4739,N_987);
and U6491 (N_6491,N_4539,N_3762);
and U6492 (N_6492,N_5971,N_367);
or U6493 (N_6493,N_4655,N_3725);
nand U6494 (N_6494,N_1190,N_750);
xnor U6495 (N_6495,N_697,N_4719);
and U6496 (N_6496,N_5498,N_3895);
or U6497 (N_6497,N_3289,N_223);
nand U6498 (N_6498,N_2715,N_5395);
nand U6499 (N_6499,N_240,N_4209);
nor U6500 (N_6500,N_1136,N_4543);
nand U6501 (N_6501,N_4152,N_1508);
nand U6502 (N_6502,N_73,N_3727);
xnor U6503 (N_6503,N_1515,N_3858);
nor U6504 (N_6504,N_3330,N_5908);
nor U6505 (N_6505,N_2573,N_1740);
and U6506 (N_6506,N_249,N_3165);
nor U6507 (N_6507,N_5246,N_5535);
or U6508 (N_6508,N_5353,N_4201);
nor U6509 (N_6509,N_2486,N_3962);
nor U6510 (N_6510,N_478,N_933);
nor U6511 (N_6511,N_3446,N_3997);
and U6512 (N_6512,N_3777,N_3919);
xnor U6513 (N_6513,N_4344,N_912);
nand U6514 (N_6514,N_56,N_3854);
xor U6515 (N_6515,N_2400,N_2613);
nor U6516 (N_6516,N_3604,N_5798);
nor U6517 (N_6517,N_2611,N_3356);
xor U6518 (N_6518,N_5935,N_4323);
or U6519 (N_6519,N_4889,N_1762);
nand U6520 (N_6520,N_23,N_3071);
and U6521 (N_6521,N_3073,N_5261);
and U6522 (N_6522,N_2164,N_2649);
and U6523 (N_6523,N_4330,N_5312);
nand U6524 (N_6524,N_2509,N_2010);
nand U6525 (N_6525,N_2489,N_5440);
or U6526 (N_6526,N_5802,N_4302);
nand U6527 (N_6527,N_2886,N_422);
nor U6528 (N_6528,N_428,N_4538);
or U6529 (N_6529,N_3314,N_3361);
nand U6530 (N_6530,N_390,N_3076);
and U6531 (N_6531,N_4808,N_3082);
and U6532 (N_6532,N_760,N_826);
or U6533 (N_6533,N_2020,N_370);
or U6534 (N_6534,N_2456,N_1399);
xor U6535 (N_6535,N_3712,N_1664);
and U6536 (N_6536,N_1526,N_2464);
and U6537 (N_6537,N_3323,N_4700);
nand U6538 (N_6538,N_2530,N_1778);
and U6539 (N_6539,N_5514,N_3052);
xnor U6540 (N_6540,N_2346,N_2889);
and U6541 (N_6541,N_1142,N_412);
nor U6542 (N_6542,N_4642,N_1992);
xor U6543 (N_6543,N_2352,N_1330);
or U6544 (N_6544,N_1340,N_5889);
or U6545 (N_6545,N_3993,N_5924);
or U6546 (N_6546,N_450,N_1126);
or U6547 (N_6547,N_3084,N_836);
nand U6548 (N_6548,N_420,N_421);
xor U6549 (N_6549,N_255,N_1443);
xor U6550 (N_6550,N_2636,N_1716);
and U6551 (N_6551,N_5304,N_3106);
xor U6552 (N_6552,N_1329,N_2732);
nor U6553 (N_6553,N_1379,N_5936);
nand U6554 (N_6554,N_5228,N_1643);
and U6555 (N_6555,N_236,N_5556);
and U6556 (N_6556,N_5006,N_4320);
nor U6557 (N_6557,N_1575,N_658);
nor U6558 (N_6558,N_1047,N_3671);
and U6559 (N_6559,N_3471,N_112);
nor U6560 (N_6560,N_1152,N_4431);
nor U6561 (N_6561,N_2667,N_3975);
nor U6562 (N_6562,N_4553,N_1976);
or U6563 (N_6563,N_1310,N_80);
xnor U6564 (N_6564,N_767,N_4953);
or U6565 (N_6565,N_4371,N_145);
nor U6566 (N_6566,N_1363,N_5768);
nand U6567 (N_6567,N_4429,N_2903);
nand U6568 (N_6568,N_5804,N_3978);
and U6569 (N_6569,N_4307,N_1695);
nor U6570 (N_6570,N_969,N_2448);
and U6571 (N_6571,N_539,N_1339);
nand U6572 (N_6572,N_2439,N_672);
nand U6573 (N_6573,N_4123,N_2864);
nand U6574 (N_6574,N_22,N_5893);
xor U6575 (N_6575,N_1836,N_2801);
xor U6576 (N_6576,N_5527,N_1070);
nand U6577 (N_6577,N_4205,N_1141);
nor U6578 (N_6578,N_2349,N_3756);
and U6579 (N_6579,N_2742,N_1145);
nand U6580 (N_6580,N_4749,N_2082);
nand U6581 (N_6581,N_4281,N_4597);
nor U6582 (N_6582,N_2960,N_5208);
or U6583 (N_6583,N_3948,N_1755);
nand U6584 (N_6584,N_2959,N_5540);
nand U6585 (N_6585,N_1940,N_4686);
xnor U6586 (N_6586,N_5271,N_4625);
nand U6587 (N_6587,N_4067,N_2095);
or U6588 (N_6588,N_3150,N_338);
xnor U6589 (N_6589,N_3824,N_3584);
nor U6590 (N_6590,N_1336,N_4117);
and U6591 (N_6591,N_1255,N_5998);
xnor U6592 (N_6592,N_2525,N_794);
nor U6593 (N_6593,N_5629,N_2229);
nor U6594 (N_6594,N_3034,N_5441);
nand U6595 (N_6595,N_1436,N_3733);
xor U6596 (N_6596,N_5585,N_1767);
and U6597 (N_6597,N_5386,N_951);
or U6598 (N_6598,N_3569,N_661);
nand U6599 (N_6599,N_326,N_5233);
or U6600 (N_6600,N_1243,N_5145);
and U6601 (N_6601,N_265,N_520);
or U6602 (N_6602,N_2694,N_4002);
and U6603 (N_6603,N_4258,N_1652);
nand U6604 (N_6604,N_741,N_1820);
or U6605 (N_6605,N_418,N_4743);
xnor U6606 (N_6606,N_5388,N_4149);
or U6607 (N_6607,N_5687,N_1223);
nor U6608 (N_6608,N_1043,N_2842);
nor U6609 (N_6609,N_1640,N_5730);
nor U6610 (N_6610,N_2485,N_1215);
xor U6611 (N_6611,N_1901,N_5090);
and U6612 (N_6612,N_678,N_3845);
nand U6613 (N_6613,N_160,N_2168);
xor U6614 (N_6614,N_427,N_2780);
and U6615 (N_6615,N_3913,N_5565);
nor U6616 (N_6616,N_4761,N_5007);
nor U6617 (N_6617,N_1683,N_989);
or U6618 (N_6618,N_5360,N_1720);
or U6619 (N_6619,N_576,N_1943);
and U6620 (N_6620,N_807,N_4845);
nor U6621 (N_6621,N_3227,N_4632);
nor U6622 (N_6622,N_413,N_596);
xnor U6623 (N_6623,N_3196,N_2716);
or U6624 (N_6624,N_2476,N_1549);
nand U6625 (N_6625,N_1975,N_4315);
or U6626 (N_6626,N_4958,N_1063);
xor U6627 (N_6627,N_5321,N_2291);
xor U6628 (N_6628,N_3140,N_3344);
and U6629 (N_6629,N_4458,N_3515);
nand U6630 (N_6630,N_5009,N_4496);
xnor U6631 (N_6631,N_4352,N_3188);
nor U6632 (N_6632,N_1384,N_3205);
or U6633 (N_6633,N_5330,N_1261);
nand U6634 (N_6634,N_1014,N_345);
nand U6635 (N_6635,N_5133,N_3137);
and U6636 (N_6636,N_5256,N_2528);
or U6637 (N_6637,N_4721,N_148);
or U6638 (N_6638,N_1299,N_216);
xor U6639 (N_6639,N_4225,N_1563);
nor U6640 (N_6640,N_3413,N_4023);
and U6641 (N_6641,N_2235,N_4637);
nand U6642 (N_6642,N_5981,N_2777);
and U6643 (N_6643,N_2033,N_3917);
xor U6644 (N_6644,N_1471,N_2008);
and U6645 (N_6645,N_3573,N_2484);
and U6646 (N_6646,N_547,N_643);
nor U6647 (N_6647,N_4905,N_3380);
and U6648 (N_6648,N_2104,N_3637);
and U6649 (N_6649,N_5789,N_889);
and U6650 (N_6650,N_2111,N_5610);
nand U6651 (N_6651,N_4954,N_4066);
nor U6652 (N_6652,N_2688,N_3774);
xnor U6653 (N_6653,N_3555,N_369);
nor U6654 (N_6654,N_5332,N_399);
nor U6655 (N_6655,N_197,N_5392);
nand U6656 (N_6656,N_568,N_4334);
nand U6657 (N_6657,N_3755,N_2654);
xor U6658 (N_6658,N_1628,N_698);
nor U6659 (N_6659,N_2475,N_5483);
nor U6660 (N_6660,N_143,N_98);
nor U6661 (N_6661,N_1482,N_544);
and U6662 (N_6662,N_5863,N_4951);
or U6663 (N_6663,N_5769,N_4999);
or U6664 (N_6664,N_2974,N_4868);
nor U6665 (N_6665,N_3444,N_1578);
or U6666 (N_6666,N_1221,N_1479);
nor U6667 (N_6667,N_4835,N_4636);
xnor U6668 (N_6668,N_2244,N_5620);
xnor U6669 (N_6669,N_2883,N_5407);
and U6670 (N_6670,N_950,N_5555);
nand U6671 (N_6671,N_4994,N_3478);
and U6672 (N_6672,N_388,N_5665);
nand U6673 (N_6673,N_2368,N_1963);
xor U6674 (N_6674,N_4998,N_3226);
and U6675 (N_6675,N_1419,N_3269);
nor U6676 (N_6676,N_4220,N_3516);
and U6677 (N_6677,N_2575,N_638);
and U6678 (N_6678,N_4595,N_1655);
xnor U6679 (N_6679,N_2663,N_4659);
nor U6680 (N_6680,N_5929,N_3612);
xor U6681 (N_6681,N_762,N_1059);
or U6682 (N_6682,N_3635,N_4121);
nand U6683 (N_6683,N_3490,N_1863);
or U6684 (N_6684,N_2174,N_3442);
or U6685 (N_6685,N_59,N_4008);
and U6686 (N_6686,N_1494,N_3911);
xnor U6687 (N_6687,N_5677,N_5103);
or U6688 (N_6688,N_580,N_3683);
nor U6689 (N_6689,N_2418,N_4598);
and U6690 (N_6690,N_2749,N_917);
or U6691 (N_6691,N_3108,N_2970);
nand U6692 (N_6692,N_2581,N_3537);
nor U6693 (N_6693,N_508,N_260);
or U6694 (N_6694,N_5980,N_5999);
nor U6695 (N_6695,N_2424,N_1377);
and U6696 (N_6696,N_3319,N_3259);
nor U6697 (N_6697,N_2493,N_4221);
or U6698 (N_6698,N_1574,N_2160);
and U6699 (N_6699,N_1065,N_5973);
and U6700 (N_6700,N_4242,N_2810);
or U6701 (N_6701,N_5695,N_2292);
xnor U6702 (N_6702,N_1109,N_25);
and U6703 (N_6703,N_4034,N_2098);
xor U6704 (N_6704,N_1916,N_1275);
and U6705 (N_6705,N_570,N_2156);
or U6706 (N_6706,N_2571,N_5432);
or U6707 (N_6707,N_1053,N_5081);
and U6708 (N_6708,N_1008,N_3536);
or U6709 (N_6709,N_3321,N_90);
and U6710 (N_6710,N_553,N_2988);
nand U6711 (N_6711,N_4432,N_4838);
or U6712 (N_6712,N_2505,N_3868);
and U6713 (N_6713,N_384,N_161);
or U6714 (N_6714,N_3424,N_5119);
and U6715 (N_6715,N_193,N_5458);
nand U6716 (N_6716,N_2664,N_1486);
or U6717 (N_6717,N_168,N_881);
xor U6718 (N_6718,N_1125,N_2147);
xnor U6719 (N_6719,N_2195,N_2641);
nand U6720 (N_6720,N_635,N_2661);
xnor U6721 (N_6721,N_3599,N_1398);
and U6722 (N_6722,N_273,N_2590);
nand U6723 (N_6723,N_2304,N_1365);
or U6724 (N_6724,N_5035,N_258);
or U6725 (N_6725,N_3374,N_4599);
or U6726 (N_6726,N_4728,N_4319);
xor U6727 (N_6727,N_1163,N_571);
nand U6728 (N_6728,N_3901,N_1968);
nand U6729 (N_6729,N_4650,N_1555);
and U6730 (N_6730,N_1091,N_970);
or U6731 (N_6731,N_1092,N_1431);
or U6732 (N_6732,N_227,N_4210);
and U6733 (N_6733,N_1027,N_2812);
nor U6734 (N_6734,N_2757,N_3971);
nand U6735 (N_6735,N_150,N_5451);
nand U6736 (N_6736,N_1729,N_3242);
nor U6737 (N_6737,N_1107,N_3220);
nand U6738 (N_6738,N_1219,N_1834);
nor U6739 (N_6739,N_4304,N_3659);
and U6740 (N_6740,N_4247,N_5372);
and U6741 (N_6741,N_1086,N_778);
xor U6742 (N_6742,N_769,N_738);
nand U6743 (N_6743,N_2939,N_2197);
or U6744 (N_6744,N_3977,N_2187);
and U6745 (N_6745,N_4949,N_297);
xor U6746 (N_6746,N_4296,N_2662);
and U6747 (N_6747,N_5859,N_3641);
nor U6748 (N_6748,N_487,N_2806);
and U6749 (N_6749,N_154,N_1990);
xor U6750 (N_6750,N_1856,N_5408);
nand U6751 (N_6751,N_101,N_2392);
nor U6752 (N_6752,N_4704,N_5775);
and U6753 (N_6753,N_2043,N_3088);
or U6754 (N_6754,N_1745,N_2940);
or U6755 (N_6755,N_2729,N_4792);
xnor U6756 (N_6756,N_1906,N_3161);
xor U6757 (N_6757,N_4025,N_1230);
nand U6758 (N_6758,N_1458,N_5322);
nor U6759 (N_6759,N_3618,N_4237);
xnor U6760 (N_6760,N_4834,N_3169);
nand U6761 (N_6761,N_4372,N_644);
nand U6762 (N_6762,N_3122,N_313);
nand U6763 (N_6763,N_5782,N_1094);
or U6764 (N_6764,N_257,N_349);
nor U6765 (N_6765,N_971,N_3359);
xor U6766 (N_6766,N_1595,N_2592);
nand U6767 (N_6767,N_3888,N_2186);
nand U6768 (N_6768,N_631,N_527);
nor U6769 (N_6769,N_4765,N_1325);
or U6770 (N_6770,N_3010,N_1252);
nor U6771 (N_6771,N_2826,N_1268);
and U6772 (N_6772,N_4195,N_5295);
nor U6773 (N_6773,N_2089,N_4235);
nand U6774 (N_6774,N_2756,N_1857);
or U6775 (N_6775,N_4895,N_355);
and U6776 (N_6776,N_3066,N_4741);
xnor U6777 (N_6777,N_3784,N_4965);
xnor U6778 (N_6778,N_1038,N_2761);
nor U6779 (N_6779,N_4537,N_5943);
and U6780 (N_6780,N_1719,N_5008);
xnor U6781 (N_6781,N_383,N_4396);
or U6782 (N_6782,N_5647,N_2069);
nor U6783 (N_6783,N_5086,N_5715);
and U6784 (N_6784,N_5421,N_5770);
nand U6785 (N_6785,N_268,N_3143);
nand U6786 (N_6786,N_5385,N_5823);
and U6787 (N_6787,N_961,N_218);
nor U6788 (N_6788,N_1301,N_2467);
and U6789 (N_6789,N_1305,N_1571);
nand U6790 (N_6790,N_610,N_5744);
nor U6791 (N_6791,N_3737,N_2032);
nor U6792 (N_6792,N_320,N_3889);
or U6793 (N_6793,N_3870,N_1924);
and U6794 (N_6794,N_4491,N_4976);
xor U6795 (N_6795,N_3770,N_4984);
nand U6796 (N_6796,N_3219,N_1499);
nor U6797 (N_6797,N_4786,N_232);
nor U6798 (N_6798,N_5740,N_5329);
nor U6799 (N_6799,N_3891,N_4196);
nor U6800 (N_6800,N_3862,N_4661);
nor U6801 (N_6801,N_814,N_5115);
nor U6802 (N_6802,N_2072,N_2213);
and U6803 (N_6803,N_3458,N_451);
nand U6804 (N_6804,N_1478,N_1932);
or U6805 (N_6805,N_4722,N_4068);
xnor U6806 (N_6806,N_39,N_2541);
or U6807 (N_6807,N_2041,N_560);
nor U6808 (N_6808,N_4989,N_844);
nor U6809 (N_6809,N_4335,N_2309);
nand U6810 (N_6810,N_3744,N_2952);
nor U6811 (N_6811,N_5224,N_5954);
xnor U6812 (N_6812,N_5275,N_3179);
xor U6813 (N_6813,N_1172,N_5301);
or U6814 (N_6814,N_4780,N_2853);
xor U6815 (N_6815,N_1057,N_1612);
or U6816 (N_6816,N_5165,N_1037);
or U6817 (N_6817,N_1104,N_5668);
nor U6818 (N_6818,N_1931,N_3950);
nor U6819 (N_6819,N_1651,N_1539);
and U6820 (N_6820,N_1114,N_1311);
or U6821 (N_6821,N_3158,N_2707);
or U6822 (N_6822,N_87,N_3469);
xnor U6823 (N_6823,N_1260,N_2254);
or U6824 (N_6824,N_612,N_4891);
and U6825 (N_6825,N_5290,N_1938);
nor U6826 (N_6826,N_5318,N_310);
nand U6827 (N_6827,N_1184,N_5577);
and U6828 (N_6828,N_5121,N_5693);
or U6829 (N_6829,N_271,N_5010);
nand U6830 (N_6830,N_2720,N_3944);
xnor U6831 (N_6831,N_5234,N_48);
xnor U6832 (N_6832,N_4493,N_2258);
nand U6833 (N_6833,N_2234,N_665);
nand U6834 (N_6834,N_4781,N_3617);
or U6835 (N_6835,N_210,N_5519);
or U6836 (N_6836,N_131,N_1052);
nor U6837 (N_6837,N_4187,N_5107);
and U6838 (N_6838,N_51,N_1023);
or U6839 (N_6839,N_1964,N_5311);
nand U6840 (N_6840,N_1922,N_4609);
and U6841 (N_6841,N_4732,N_963);
nor U6842 (N_6842,N_5005,N_4904);
xor U6843 (N_6843,N_489,N_3794);
nand U6844 (N_6844,N_4199,N_5944);
or U6845 (N_6845,N_5812,N_2763);
nor U6846 (N_6846,N_5144,N_1421);
nand U6847 (N_6847,N_1256,N_2106);
xor U6848 (N_6848,N_4029,N_2305);
nand U6849 (N_6849,N_5627,N_3253);
nor U6850 (N_6850,N_5803,N_4870);
xnor U6851 (N_6851,N_181,N_1196);
and U6852 (N_6852,N_4740,N_4688);
xnor U6853 (N_6853,N_1674,N_352);
or U6854 (N_6854,N_3646,N_5020);
nor U6855 (N_6855,N_406,N_2823);
nand U6856 (N_6856,N_1022,N_2323);
xor U6857 (N_6857,N_745,N_1984);
or U6858 (N_6858,N_5049,N_2226);
nand U6859 (N_6859,N_5589,N_1236);
and U6860 (N_6860,N_243,N_2006);
nand U6861 (N_6861,N_4494,N_5237);
xor U6862 (N_6862,N_5576,N_1746);
or U6863 (N_6863,N_3381,N_4421);
and U6864 (N_6864,N_2928,N_4666);
and U6865 (N_6865,N_4929,N_5490);
nor U6866 (N_6866,N_4326,N_2443);
and U6867 (N_6867,N_2036,N_1140);
or U6868 (N_6868,N_1669,N_811);
nor U6869 (N_6869,N_4855,N_5656);
and U6870 (N_6870,N_1276,N_4800);
and U6871 (N_6871,N_104,N_2634);
or U6872 (N_6872,N_4437,N_5862);
nor U6873 (N_6873,N_4603,N_2992);
nor U6874 (N_6874,N_5331,N_2307);
and U6875 (N_6875,N_4584,N_135);
or U6876 (N_6876,N_5747,N_3964);
and U6877 (N_6877,N_5718,N_4484);
or U6878 (N_6878,N_4950,N_2676);
or U6879 (N_6879,N_2863,N_3299);
nand U6880 (N_6880,N_5180,N_5127);
or U6881 (N_6881,N_1957,N_2178);
or U6882 (N_6882,N_137,N_4896);
nor U6883 (N_6883,N_2927,N_1410);
nor U6884 (N_6884,N_4231,N_204);
xor U6885 (N_6885,N_3625,N_5406);
xor U6886 (N_6886,N_1939,N_5752);
nand U6887 (N_6887,N_1446,N_1700);
xor U6888 (N_6888,N_5108,N_217);
xnor U6889 (N_6889,N_5742,N_2127);
or U6890 (N_6890,N_4236,N_1886);
or U6891 (N_6891,N_4702,N_5222);
xnor U6892 (N_6892,N_5434,N_4770);
and U6893 (N_6893,N_1179,N_1376);
nor U6894 (N_6894,N_5135,N_4427);
nand U6895 (N_6895,N_4146,N_4901);
xnor U6896 (N_6896,N_474,N_5810);
xnor U6897 (N_6897,N_3382,N_4798);
nor U6898 (N_6898,N_646,N_4693);
nand U6899 (N_6899,N_4338,N_322);
nand U6900 (N_6900,N_3639,N_3834);
nand U6901 (N_6901,N_4037,N_5299);
xor U6902 (N_6902,N_5075,N_5);
nand U6903 (N_6903,N_40,N_4081);
nand U6904 (N_6904,N_3746,N_5206);
xor U6905 (N_6905,N_4975,N_2591);
nand U6906 (N_6906,N_3930,N_2228);
or U6907 (N_6907,N_3987,N_4417);
and U6908 (N_6908,N_3608,N_1313);
and U6909 (N_6909,N_375,N_5578);
or U6910 (N_6910,N_3097,N_2088);
nand U6911 (N_6911,N_4297,N_4027);
nand U6912 (N_6912,N_319,N_2402);
xnor U6913 (N_6913,N_4568,N_2516);
nor U6914 (N_6914,N_2311,N_2123);
or U6915 (N_6915,N_3994,N_453);
or U6916 (N_6916,N_4825,N_716);
nor U6917 (N_6917,N_5961,N_1885);
nand U6918 (N_6918,N_2962,N_2388);
xnor U6919 (N_6919,N_4535,N_614);
xor U6920 (N_6920,N_2520,N_1839);
nand U6921 (N_6921,N_1694,N_290);
and U6922 (N_6922,N_3496,N_2550);
or U6923 (N_6923,N_3254,N_2612);
and U6924 (N_6924,N_3936,N_4972);
or U6925 (N_6925,N_4515,N_3902);
or U6926 (N_6926,N_5412,N_1253);
nand U6927 (N_6927,N_1352,N_1441);
nand U6928 (N_6928,N_34,N_2200);
xor U6929 (N_6929,N_626,N_4212);
nand U6930 (N_6930,N_2837,N_4388);
nand U6931 (N_6931,N_3500,N_5765);
and U6932 (N_6932,N_5654,N_5726);
xor U6933 (N_6933,N_781,N_2513);
xor U6934 (N_6934,N_3825,N_2976);
and U6935 (N_6935,N_926,N_4422);
xnor U6936 (N_6936,N_607,N_2619);
xnor U6937 (N_6937,N_4381,N_5138);
or U6938 (N_6938,N_852,N_3510);
xor U6939 (N_6939,N_2847,N_1009);
xor U6940 (N_6940,N_2583,N_2440);
nand U6941 (N_6941,N_528,N_4753);
or U6942 (N_6942,N_1538,N_1613);
or U6943 (N_6943,N_5309,N_1282);
xor U6944 (N_6944,N_359,N_1566);
nor U6945 (N_6945,N_4419,N_3811);
and U6946 (N_6946,N_4514,N_4548);
nor U6947 (N_6947,N_3102,N_5223);
nor U6948 (N_6948,N_2943,N_4240);
and U6949 (N_6949,N_4030,N_687);
nor U6950 (N_6950,N_531,N_3387);
xnor U6951 (N_6951,N_5615,N_4299);
nor U6952 (N_6952,N_75,N_409);
xnor U6953 (N_6953,N_5684,N_4287);
nor U6954 (N_6954,N_505,N_879);
and U6955 (N_6955,N_79,N_2397);
nor U6956 (N_6956,N_5048,N_4044);
nor U6957 (N_6957,N_1088,N_2572);
xnor U6958 (N_6958,N_5898,N_4178);
and U6959 (N_6959,N_3633,N_683);
or U6960 (N_6960,N_2558,N_4181);
xor U6961 (N_6961,N_2602,N_1461);
nor U6962 (N_6962,N_3803,N_2133);
xor U6963 (N_6963,N_981,N_1472);
nor U6964 (N_6964,N_391,N_5640);
nand U6965 (N_6965,N_4241,N_4656);
xnor U6966 (N_6966,N_993,N_95);
and U6967 (N_6967,N_1161,N_5294);
nor U6968 (N_6968,N_5716,N_3229);
nand U6969 (N_6969,N_2755,N_2290);
and U6970 (N_6970,N_2705,N_3448);
nor U6971 (N_6971,N_2627,N_4631);
or U6972 (N_6972,N_3985,N_965);
or U6973 (N_6973,N_504,N_3470);
xor U6974 (N_6974,N_4171,N_2421);
nand U6975 (N_6975,N_5239,N_3023);
and U6976 (N_6976,N_5611,N_3096);
or U6977 (N_6977,N_5265,N_1481);
and U6978 (N_6978,N_2083,N_1084);
nand U6979 (N_6979,N_1337,N_3293);
and U6980 (N_6980,N_1645,N_590);
nand U6981 (N_6981,N_5820,N_289);
nand U6982 (N_6982,N_3648,N_3371);
nor U6983 (N_6983,N_5461,N_4256);
and U6984 (N_6984,N_2014,N_2225);
nor U6985 (N_6985,N_1326,N_458);
nand U6986 (N_6986,N_5567,N_5197);
xor U6987 (N_6987,N_4618,N_5504);
nor U6988 (N_6988,N_2556,N_1671);
xor U6989 (N_6989,N_669,N_252);
or U6990 (N_6990,N_5599,N_3695);
nand U6991 (N_6991,N_783,N_4955);
and U6992 (N_6992,N_892,N_3170);
or U6993 (N_6993,N_5027,N_3408);
nor U6994 (N_6994,N_4270,N_4197);
nor U6995 (N_6995,N_2577,N_3224);
xor U6996 (N_6996,N_5156,N_4401);
nand U6997 (N_6997,N_492,N_1741);
nand U6998 (N_6998,N_2738,N_615);
or U6999 (N_6999,N_155,N_972);
nand U7000 (N_7000,N_1832,N_2844);
and U7001 (N_7001,N_2438,N_4892);
nand U7002 (N_7002,N_2275,N_739);
or U7003 (N_7003,N_3572,N_3417);
nand U7004 (N_7004,N_3216,N_3937);
or U7005 (N_7005,N_916,N_3235);
and U7006 (N_7006,N_1288,N_66);
xor U7007 (N_7007,N_4813,N_2427);
nand U7008 (N_7008,N_461,N_2045);
nor U7009 (N_7009,N_2158,N_3611);
and U7010 (N_7010,N_3144,N_538);
and U7011 (N_7011,N_1568,N_329);
nor U7012 (N_7012,N_964,N_1332);
nor U7013 (N_7013,N_3798,N_3722);
nor U7014 (N_7014,N_4633,N_5949);
nand U7015 (N_7015,N_5314,N_2567);
or U7016 (N_7016,N_2607,N_2308);
nor U7017 (N_7017,N_208,N_816);
and U7018 (N_7018,N_4988,N_5215);
xor U7019 (N_7019,N_5543,N_2371);
xnor U7020 (N_7020,N_2872,N_4992);
nor U7021 (N_7021,N_3307,N_4269);
nand U7022 (N_7022,N_1082,N_53);
and U7023 (N_7023,N_4423,N_4349);
nor U7024 (N_7024,N_3491,N_600);
and U7025 (N_7025,N_5800,N_3687);
or U7026 (N_7026,N_586,N_1702);
xor U7027 (N_7027,N_936,N_4658);
nand U7028 (N_7028,N_3013,N_944);
or U7029 (N_7029,N_2035,N_1122);
and U7030 (N_7030,N_4711,N_5120);
nand U7031 (N_7031,N_880,N_4416);
xnor U7032 (N_7032,N_4439,N_682);
nand U7033 (N_7033,N_5091,N_3133);
nor U7034 (N_7034,N_354,N_3545);
nor U7035 (N_7035,N_1524,N_332);
xnor U7036 (N_7036,N_1826,N_761);
and U7037 (N_7037,N_4488,N_2542);
and U7038 (N_7038,N_2029,N_339);
and U7039 (N_7039,N_5865,N_5221);
or U7040 (N_7040,N_5024,N_4717);
nand U7041 (N_7041,N_922,N_562);
nand U7042 (N_7042,N_4847,N_1004);
nor U7043 (N_7043,N_1504,N_1167);
nor U7044 (N_7044,N_3757,N_3062);
or U7045 (N_7045,N_894,N_4602);
or U7046 (N_7046,N_5642,N_4500);
nor U7047 (N_7047,N_3280,N_3085);
nor U7048 (N_7048,N_4160,N_1936);
xnor U7049 (N_7049,N_431,N_5229);
nor U7050 (N_7050,N_5583,N_4305);
and U7051 (N_7051,N_4601,N_1876);
or U7052 (N_7052,N_1457,N_3095);
or U7053 (N_7053,N_3123,N_3153);
and U7054 (N_7054,N_763,N_1987);
and U7055 (N_7055,N_5324,N_1807);
nand U7056 (N_7056,N_1342,N_1099);
nor U7057 (N_7057,N_5284,N_4107);
or U7058 (N_7058,N_106,N_4708);
nor U7059 (N_7059,N_2331,N_5403);
or U7060 (N_7060,N_775,N_2562);
nand U7061 (N_7061,N_771,N_18);
xnor U7062 (N_7062,N_3841,N_1631);
nand U7063 (N_7063,N_5508,N_3559);
or U7064 (N_7064,N_850,N_400);
nor U7065 (N_7065,N_1941,N_3325);
nand U7066 (N_7066,N_5674,N_3019);
or U7067 (N_7067,N_744,N_1062);
nor U7068 (N_7068,N_4937,N_1307);
nor U7069 (N_7069,N_4365,N_1120);
nor U7070 (N_7070,N_2719,N_3028);
nor U7071 (N_7071,N_4085,N_2690);
nand U7072 (N_7072,N_5021,N_3400);
xor U7073 (N_7073,N_3057,N_3876);
and U7074 (N_7074,N_1706,N_3193);
or U7075 (N_7075,N_2264,N_5055);
nand U7076 (N_7076,N_3793,N_1822);
or U7077 (N_7077,N_1991,N_1768);
or U7078 (N_7078,N_3487,N_5313);
nor U7079 (N_7079,N_1962,N_2937);
xnor U7080 (N_7080,N_1225,N_3270);
nor U7081 (N_7081,N_2608,N_4303);
xnor U7082 (N_7082,N_3195,N_664);
nand U7083 (N_7083,N_5636,N_4162);
and U7084 (N_7084,N_1010,N_3301);
or U7085 (N_7085,N_3175,N_5644);
nor U7086 (N_7086,N_3112,N_4760);
xor U7087 (N_7087,N_5469,N_5391);
xor U7088 (N_7088,N_3680,N_4166);
nor U7089 (N_7089,N_2647,N_1791);
nand U7090 (N_7090,N_3893,N_1980);
xnor U7091 (N_7091,N_973,N_4271);
nor U7092 (N_7092,N_841,N_1998);
nand U7093 (N_7093,N_3308,N_5056);
or U7094 (N_7094,N_2983,N_2462);
xor U7095 (N_7095,N_2080,N_4118);
nor U7096 (N_7096,N_5455,N_138);
nor U7097 (N_7097,N_3776,N_5659);
and U7098 (N_7098,N_5901,N_3656);
nand U7099 (N_7099,N_4613,N_727);
and U7100 (N_7100,N_3586,N_4190);
and U7101 (N_7101,N_4017,N_1752);
and U7102 (N_7102,N_3799,N_3670);
and U7103 (N_7103,N_3174,N_3054);
xor U7104 (N_7104,N_3905,N_1814);
or U7105 (N_7105,N_1601,N_2785);
xnor U7106 (N_7106,N_4823,N_5057);
and U7107 (N_7107,N_5272,N_768);
or U7108 (N_7108,N_1966,N_3890);
nand U7109 (N_7109,N_1117,N_3047);
and U7110 (N_7110,N_81,N_577);
xor U7111 (N_7111,N_953,N_1217);
or U7112 (N_7112,N_2859,N_2359);
xnor U7113 (N_7113,N_4788,N_4674);
or U7114 (N_7114,N_5003,N_4653);
xor U7115 (N_7115,N_4940,N_5760);
nand U7116 (N_7116,N_5094,N_2549);
xnor U7117 (N_7117,N_3812,N_792);
xnor U7118 (N_7118,N_1772,N_3867);
nor U7119 (N_7119,N_3067,N_1165);
or U7120 (N_7120,N_3072,N_1234);
nand U7121 (N_7121,N_4763,N_3004);
nand U7122 (N_7122,N_286,N_4342);
and U7123 (N_7123,N_2496,N_842);
nor U7124 (N_7124,N_4829,N_1753);
xor U7125 (N_7125,N_4145,N_4664);
xnor U7126 (N_7126,N_1638,N_1194);
or U7127 (N_7127,N_2320,N_632);
nor U7128 (N_7128,N_2656,N_5184);
nand U7129 (N_7129,N_1366,N_2287);
nand U7130 (N_7130,N_1487,N_2260);
or U7131 (N_7131,N_2411,N_251);
or U7132 (N_7132,N_4608,N_2926);
xnor U7133 (N_7133,N_3672,N_498);
nand U7134 (N_7134,N_3020,N_5877);
or U7135 (N_7135,N_3326,N_1604);
nor U7136 (N_7136,N_5232,N_1577);
nor U7137 (N_7137,N_2412,N_2899);
nor U7138 (N_7138,N_5658,N_1823);
or U7139 (N_7139,N_565,N_4313);
nand U7140 (N_7140,N_3410,N_3025);
nand U7141 (N_7141,N_1263,N_3402);
or U7142 (N_7142,N_1245,N_3800);
xnor U7143 (N_7143,N_4218,N_681);
nor U7144 (N_7144,N_1971,N_1703);
nand U7145 (N_7145,N_685,N_3272);
and U7146 (N_7146,N_3241,N_2586);
or U7147 (N_7147,N_1606,N_3623);
nand U7148 (N_7148,N_4075,N_1547);
or U7149 (N_7149,N_1731,N_1988);
or U7150 (N_7150,N_4119,N_1071);
or U7151 (N_7151,N_4369,N_4267);
xnor U7152 (N_7152,N_3880,N_3503);
or U7153 (N_7153,N_304,N_5164);
nor U7154 (N_7154,N_5982,N_5193);
nand U7155 (N_7155,N_5082,N_4147);
xor U7156 (N_7156,N_5947,N_4995);
nor U7157 (N_7157,N_1054,N_1316);
nand U7158 (N_7158,N_1110,N_2);
xor U7159 (N_7159,N_393,N_1845);
nor U7160 (N_7160,N_231,N_4936);
nand U7161 (N_7161,N_1641,N_1130);
and U7162 (N_7162,N_5570,N_2861);
and U7163 (N_7163,N_3422,N_4832);
xor U7164 (N_7164,N_4350,N_4944);
xnor U7165 (N_7165,N_5984,N_2680);
xnor U7166 (N_7166,N_5036,N_634);
or U7167 (N_7167,N_5022,N_5097);
nand U7168 (N_7168,N_361,N_455);
xnor U7169 (N_7169,N_4408,N_3763);
and U7170 (N_7170,N_4692,N_3802);
nand U7171 (N_7171,N_5471,N_5204);
nor U7172 (N_7172,N_3758,N_5729);
xnor U7173 (N_7173,N_3030,N_5905);
or U7174 (N_7174,N_2068,N_4129);
xor U7175 (N_7175,N_4758,N_5515);
or U7176 (N_7176,N_372,N_1733);
or U7177 (N_7177,N_4967,N_3871);
or U7178 (N_7178,N_1228,N_4917);
and U7179 (N_7179,N_3544,N_4696);
nand U7180 (N_7180,N_5542,N_3125);
nor U7181 (N_7181,N_595,N_4731);
xor U7182 (N_7182,N_689,N_5297);
and U7183 (N_7183,N_3542,N_5939);
or U7184 (N_7184,N_5252,N_1634);
or U7185 (N_7185,N_5118,N_4096);
and U7186 (N_7186,N_3005,N_3651);
or U7187 (N_7187,N_4963,N_5151);
or U7188 (N_7188,N_1220,N_3951);
nor U7189 (N_7189,N_3697,N_2803);
xnor U7190 (N_7190,N_1955,N_5069);
or U7191 (N_7191,N_1859,N_460);
or U7192 (N_7192,N_5662,N_5468);
or U7193 (N_7193,N_2840,N_4064);
and U7194 (N_7194,N_3640,N_3699);
nor U7195 (N_7195,N_5095,N_4772);
and U7196 (N_7196,N_5754,N_1146);
nor U7197 (N_7197,N_5572,N_4377);
nand U7198 (N_7198,N_3859,N_5292);
nand U7199 (N_7199,N_5484,N_1766);
nand U7200 (N_7200,N_711,N_2503);
nor U7201 (N_7201,N_4028,N_2783);
xnor U7202 (N_7202,N_1873,N_3943);
or U7203 (N_7203,N_513,N_4282);
xor U7204 (N_7204,N_3650,N_633);
and U7205 (N_7205,N_209,N_4128);
or U7206 (N_7206,N_5895,N_2704);
nor U7207 (N_7207,N_1712,N_2019);
or U7208 (N_7208,N_2650,N_2628);
and U7209 (N_7209,N_2770,N_1322);
xor U7210 (N_7210,N_3171,N_2218);
nor U7211 (N_7211,N_429,N_5479);
and U7212 (N_7212,N_1369,N_5532);
or U7213 (N_7213,N_1149,N_2718);
and U7214 (N_7214,N_3388,N_3912);
xor U7215 (N_7215,N_3135,N_627);
nor U7216 (N_7216,N_1838,N_756);
nand U7217 (N_7217,N_2529,N_2459);
xor U7218 (N_7218,N_4803,N_3120);
and U7219 (N_7219,N_3856,N_4624);
nor U7220 (N_7220,N_1137,N_1303);
xor U7221 (N_7221,N_5766,N_833);
xor U7222 (N_7222,N_2941,N_247);
and U7223 (N_7223,N_5453,N_928);
nor U7224 (N_7224,N_1781,N_5786);
xor U7225 (N_7225,N_2731,N_2813);
nand U7226 (N_7226,N_805,N_534);
nor U7227 (N_7227,N_2038,N_2909);
and U7228 (N_7228,N_3547,N_2155);
and U7229 (N_7229,N_2317,N_5596);
xnor U7230 (N_7230,N_1407,N_5380);
or U7231 (N_7231,N_5045,N_4286);
or U7232 (N_7232,N_2171,N_4382);
xnor U7233 (N_7233,N_2820,N_1935);
nor U7234 (N_7234,N_2896,N_5147);
or U7235 (N_7235,N_1592,N_5362);
nand U7236 (N_7236,N_1801,N_4884);
nand U7237 (N_7237,N_4509,N_3260);
nor U7238 (N_7238,N_4822,N_5751);
nand U7239 (N_7239,N_5013,N_6);
or U7240 (N_7240,N_2273,N_2691);
nor U7241 (N_7241,N_859,N_3211);
nand U7242 (N_7242,N_456,N_5624);
xnor U7243 (N_7243,N_78,N_4148);
xor U7244 (N_7244,N_119,N_3141);
nand U7245 (N_7245,N_1550,N_597);
nor U7246 (N_7246,N_772,N_324);
and U7247 (N_7247,N_4384,N_870);
or U7248 (N_7248,N_2345,N_1522);
xor U7249 (N_7249,N_1169,N_5139);
nand U7250 (N_7250,N_3083,N_5592);
or U7251 (N_7251,N_5338,N_5796);
nand U7252 (N_7252,N_5142,N_3275);
nor U7253 (N_7253,N_1505,N_1513);
nand U7254 (N_7254,N_704,N_1688);
or U7255 (N_7255,N_2888,N_4657);
nor U7256 (N_7256,N_4006,N_854);
xor U7257 (N_7257,N_2524,N_1327);
or U7258 (N_7258,N_5834,N_3942);
and U7259 (N_7259,N_295,N_3817);
nand U7260 (N_7260,N_2376,N_3146);
nand U7261 (N_7261,N_3832,N_1198);
xnor U7262 (N_7262,N_281,N_3338);
and U7263 (N_7263,N_3836,N_2968);
or U7264 (N_7264,N_1926,N_2351);
nand U7265 (N_7265,N_509,N_2547);
and U7266 (N_7266,N_246,N_2137);
nor U7267 (N_7267,N_765,N_2490);
nor U7268 (N_7268,N_2678,N_3257);
nand U7269 (N_7269,N_3598,N_3126);
or U7270 (N_7270,N_865,N_348);
and U7271 (N_7271,N_3928,N_585);
xnor U7272 (N_7272,N_2522,N_1408);
nor U7273 (N_7273,N_2771,N_2989);
xnor U7274 (N_7274,N_773,N_1115);
or U7275 (N_7275,N_5669,N_5549);
and U7276 (N_7276,N_4389,N_238);
and U7277 (N_7277,N_1463,N_2134);
or U7278 (N_7278,N_445,N_5201);
xnor U7279 (N_7279,N_1639,N_1453);
xor U7280 (N_7280,N_5650,N_2217);
xnor U7281 (N_7281,N_5794,N_1269);
nand U7282 (N_7282,N_5563,N_266);
xor U7283 (N_7283,N_309,N_1150);
xor U7284 (N_7284,N_2752,N_3910);
nor U7285 (N_7285,N_2793,N_5427);
and U7286 (N_7286,N_5959,N_1543);
xnor U7287 (N_7287,N_2318,N_5721);
or U7288 (N_7288,N_3177,N_1518);
xnor U7289 (N_7289,N_3835,N_125);
and U7290 (N_7290,N_930,N_3290);
or U7291 (N_7291,N_3875,N_1476);
or U7292 (N_7292,N_5162,N_5379);
and U7293 (N_7293,N_588,N_5553);
or U7294 (N_7294,N_5502,N_177);
or U7295 (N_7295,N_5965,N_5374);
and U7296 (N_7296,N_780,N_4591);
and U7297 (N_7297,N_4289,N_5706);
and U7298 (N_7298,N_5283,N_1875);
xor U7299 (N_7299,N_927,N_2191);
and U7300 (N_7300,N_5217,N_4250);
and U7301 (N_7301,N_3969,N_5345);
and U7302 (N_7302,N_4239,N_848);
nor U7303 (N_7303,N_2932,N_2671);
nor U7304 (N_7304,N_5832,N_4939);
nor U7305 (N_7305,N_1239,N_5389);
xor U7306 (N_7306,N_4804,N_5117);
nor U7307 (N_7307,N_1049,N_1507);
nor U7308 (N_7308,N_1030,N_5238);
xor U7309 (N_7309,N_3717,N_898);
and U7310 (N_7310,N_256,N_2224);
or U7311 (N_7311,N_452,N_1747);
or U7312 (N_7312,N_2265,N_4188);
or U7313 (N_7313,N_5472,N_3318);
nand U7314 (N_7314,N_986,N_3682);
xor U7315 (N_7315,N_4499,N_479);
and U7316 (N_7316,N_1177,N_43);
nor U7317 (N_7317,N_3630,N_377);
and U7318 (N_7318,N_942,N_2389);
nor U7319 (N_7319,N_1241,N_3002);
xor U7320 (N_7320,N_5801,N_4615);
nor U7321 (N_7321,N_4996,N_2897);
nand U7322 (N_7322,N_433,N_2564);
and U7323 (N_7323,N_1866,N_3535);
xnor U7324 (N_7324,N_5874,N_3109);
and U7325 (N_7325,N_5588,N_736);
nor U7326 (N_7326,N_5414,N_4363);
nand U7327 (N_7327,N_109,N_4470);
xor U7328 (N_7328,N_494,N_4183);
nor U7329 (N_7329,N_1656,N_2521);
or U7330 (N_7330,N_4489,N_564);
nor U7331 (N_7331,N_1776,N_4158);
or U7332 (N_7332,N_5767,N_2660);
xnor U7333 (N_7333,N_1381,N_2110);
and U7334 (N_7334,N_4862,N_3593);
and U7335 (N_7335,N_4232,N_469);
xor U7336 (N_7336,N_2617,N_679);
nand U7337 (N_7337,N_1334,N_333);
nor U7338 (N_7338,N_985,N_4043);
or U7339 (N_7339,N_2854,N_467);
or U7340 (N_7340,N_2935,N_52);
nand U7341 (N_7341,N_4564,N_3264);
or U7342 (N_7342,N_4039,N_649);
nor U7343 (N_7343,N_2693,N_4341);
xor U7344 (N_7344,N_4024,N_2585);
xnor U7345 (N_7345,N_1739,N_1862);
and U7346 (N_7346,N_5609,N_3814);
and U7347 (N_7347,N_1210,N_1849);
or U7348 (N_7348,N_4219,N_5630);
and U7349 (N_7349,N_4592,N_1599);
nand U7350 (N_7350,N_3806,N_1617);
xnor U7351 (N_7351,N_4587,N_552);
xnor U7352 (N_7352,N_2395,N_1580);
nor U7353 (N_7353,N_4764,N_485);
or U7354 (N_7354,N_4887,N_4268);
xnor U7355 (N_7355,N_1912,N_2337);
nand U7356 (N_7356,N_537,N_5525);
nor U7357 (N_7357,N_514,N_2100);
nor U7358 (N_7358,N_4806,N_4559);
nand U7359 (N_7359,N_4355,N_5001);
or U7360 (N_7360,N_4748,N_5174);
and U7361 (N_7361,N_4714,N_68);
or U7362 (N_7362,N_3662,N_1321);
xor U7363 (N_7363,N_5602,N_5633);
or U7364 (N_7364,N_5317,N_714);
or U7365 (N_7365,N_2423,N_1087);
nor U7366 (N_7366,N_3898,N_340);
nor U7367 (N_7367,N_1139,N_2479);
and U7368 (N_7368,N_957,N_1069);
nor U7369 (N_7369,N_5975,N_3517);
or U7370 (N_7370,N_3232,N_2348);
xnor U7371 (N_7371,N_99,N_5183);
and U7372 (N_7372,N_2379,N_3230);
nand U7373 (N_7373,N_2086,N_5641);
nor U7374 (N_7374,N_3860,N_5968);
xor U7375 (N_7375,N_4826,N_153);
or U7376 (N_7376,N_5137,N_5849);
or U7377 (N_7377,N_3866,N_2878);
nor U7378 (N_7378,N_1620,N_2140);
nor U7379 (N_7379,N_5100,N_5411);
nor U7380 (N_7380,N_2964,N_674);
xor U7381 (N_7381,N_2199,N_5822);
or U7382 (N_7382,N_2474,N_5701);
nand U7383 (N_7383,N_923,N_49);
nand U7384 (N_7384,N_3696,N_4254);
nand U7385 (N_7385,N_1226,N_1758);
xor U7386 (N_7386,N_3156,N_3676);
xor U7387 (N_7387,N_3645,N_3287);
and U7388 (N_7388,N_3703,N_3059);
or U7389 (N_7389,N_3037,N_733);
xnor U7390 (N_7390,N_521,N_3404);
and U7391 (N_7391,N_5838,N_5288);
or U7392 (N_7392,N_3463,N_874);
xor U7393 (N_7393,N_229,N_3909);
xnor U7394 (N_7394,N_4367,N_5545);
or U7395 (N_7395,N_2231,N_1614);
xnor U7396 (N_7396,N_2997,N_201);
xor U7397 (N_7397,N_3968,N_962);
or U7398 (N_7398,N_5735,N_140);
nand U7399 (N_7399,N_287,N_845);
nor U7400 (N_7400,N_5102,N_4836);
and U7401 (N_7401,N_4038,N_2891);
and U7402 (N_7402,N_4698,N_5520);
xnor U7403 (N_7403,N_2744,N_3629);
nand U7404 (N_7404,N_3995,N_1648);
nor U7405 (N_7405,N_5128,N_4047);
xor U7406 (N_7406,N_3949,N_4185);
or U7407 (N_7407,N_2240,N_3843);
xnor U7408 (N_7408,N_5497,N_1096);
or U7409 (N_7409,N_1308,N_2092);
or U7410 (N_7410,N_2350,N_3677);
nor U7411 (N_7411,N_4527,N_3435);
or U7412 (N_7412,N_2167,N_1517);
or U7413 (N_7413,N_4452,N_5692);
and U7414 (N_7414,N_3182,N_660);
nand U7415 (N_7415,N_4638,N_1314);
nor U7416 (N_7416,N_3209,N_1155);
and U7417 (N_7417,N_4062,N_4051);
and U7418 (N_7418,N_3377,N_3668);
nand U7419 (N_7419,N_896,N_1799);
nor U7420 (N_7420,N_1777,N_1003);
xnor U7421 (N_7421,N_1902,N_2815);
nand U7422 (N_7422,N_5869,N_4716);
nand U7423 (N_7423,N_3705,N_4752);
nand U7424 (N_7424,N_800,N_2300);
nand U7425 (N_7425,N_3554,N_5978);
nor U7426 (N_7426,N_598,N_200);
nor U7427 (N_7427,N_1603,N_2515);
nor U7428 (N_7428,N_2482,N_3563);
nand U7429 (N_7429,N_105,N_415);
and U7430 (N_7430,N_1264,N_1396);
or U7431 (N_7431,N_4796,N_2166);
and U7432 (N_7432,N_1106,N_2908);
and U7433 (N_7433,N_5906,N_5634);
or U7434 (N_7434,N_5966,N_3719);
xor U7435 (N_7435,N_2227,N_244);
nor U7436 (N_7436,N_1864,N_2906);
and U7437 (N_7437,N_3479,N_3329);
nand U7438 (N_7438,N_625,N_4073);
or U7439 (N_7439,N_2250,N_3035);
xnor U7440 (N_7440,N_1954,N_5178);
xor U7441 (N_7441,N_4477,N_3614);
and U7442 (N_7442,N_82,N_587);
and U7443 (N_7443,N_1687,N_3653);
and U7444 (N_7444,N_4055,N_2559);
or U7445 (N_7445,N_2415,N_3202);
and U7446 (N_7446,N_1609,N_2488);
nand U7447 (N_7447,N_915,N_2236);
nor U7448 (N_7448,N_4095,N_1858);
and U7449 (N_7449,N_1897,N_4549);
and U7450 (N_7450,N_1636,N_2094);
or U7451 (N_7451,N_1385,N_5591);
or U7452 (N_7452,N_992,N_3679);
and U7453 (N_7453,N_1103,N_2176);
nand U7454 (N_7454,N_5790,N_1267);
xnor U7455 (N_7455,N_5480,N_126);
and U7456 (N_7456,N_1675,N_2957);
nor U7457 (N_7457,N_3857,N_5079);
nand U7458 (N_7458,N_3282,N_974);
and U7459 (N_7459,N_4968,N_35);
xor U7460 (N_7460,N_481,N_5442);
nand U7461 (N_7461,N_2589,N_5367);
nor U7462 (N_7462,N_5492,N_3846);
nand U7463 (N_7463,N_3238,N_620);
or U7464 (N_7464,N_5310,N_4251);
or U7465 (N_7465,N_589,N_3590);
or U7466 (N_7466,N_2514,N_1829);
nand U7467 (N_7467,N_559,N_4447);
and U7468 (N_7468,N_1579,N_3462);
nor U7469 (N_7469,N_2220,N_191);
nor U7470 (N_7470,N_4252,N_3708);
and U7471 (N_7471,N_2626,N_1158);
or U7472 (N_7472,N_5552,N_1779);
xnor U7473 (N_7473,N_709,N_3370);
nor U7474 (N_7474,N_1520,N_3738);
nor U7475 (N_7475,N_493,N_4682);
nor U7476 (N_7476,N_5830,N_447);
nand U7477 (N_7477,N_4288,N_1429);
and U7478 (N_7478,N_5847,N_5653);
nand U7479 (N_7479,N_3925,N_2703);
nor U7480 (N_7480,N_1732,N_4912);
xnor U7481 (N_7481,N_318,N_5753);
xnor U7482 (N_7482,N_703,N_5209);
xnor U7483 (N_7483,N_371,N_3401);
and U7484 (N_7484,N_5157,N_3115);
or U7485 (N_7485,N_190,N_1296);
or U7486 (N_7486,N_3436,N_2934);
nand U7487 (N_7487,N_1684,N_3603);
or U7488 (N_7488,N_5561,N_89);
and U7489 (N_7489,N_4634,N_1557);
nand U7490 (N_7490,N_1750,N_2002);
nor U7491 (N_7491,N_1076,N_1448);
xor U7492 (N_7492,N_134,N_4875);
nor U7493 (N_7493,N_163,N_4957);
or U7494 (N_7494,N_1914,N_3315);
xnor U7495 (N_7495,N_2243,N_317);
nand U7496 (N_7496,N_4974,N_4768);
nand U7497 (N_7497,N_2784,N_5757);
nand U7498 (N_7498,N_5426,N_1833);
nand U7499 (N_7499,N_4644,N_2454);
xnor U7500 (N_7500,N_2085,N_5278);
nor U7501 (N_7501,N_96,N_5500);
or U7502 (N_7502,N_3265,N_506);
and U7503 (N_7503,N_5354,N_5489);
and U7504 (N_7504,N_2533,N_4783);
and U7505 (N_7505,N_5672,N_465);
xor U7506 (N_7506,N_4629,N_2391);
or U7507 (N_7507,N_3250,N_984);
or U7508 (N_7508,N_3716,N_3131);
nand U7509 (N_7509,N_834,N_4579);
nor U7510 (N_7510,N_4479,N_4550);
xnor U7511 (N_7511,N_1409,N_2472);
nand U7512 (N_7512,N_5612,N_581);
nor U7513 (N_7513,N_888,N_4136);
xor U7514 (N_7514,N_1635,N_1090);
nor U7515 (N_7515,N_2597,N_5028);
nor U7516 (N_7516,N_3840,N_2499);
nand U7517 (N_7517,N_1193,N_4230);
nand U7518 (N_7518,N_3333,N_173);
and U7519 (N_7519,N_5550,N_5655);
nor U7520 (N_7520,N_1147,N_5912);
and U7521 (N_7521,N_4522,N_2313);
nor U7522 (N_7522,N_1851,N_1985);
nor U7523 (N_7523,N_3922,N_4283);
and U7524 (N_7524,N_5176,N_4374);
nand U7525 (N_7525,N_4581,N_2767);
nand U7526 (N_7526,N_690,N_5821);
nor U7527 (N_7527,N_5503,N_4516);
and U7528 (N_7528,N_1271,N_1512);
or U7529 (N_7529,N_1780,N_2360);
nor U7530 (N_7530,N_2408,N_3430);
nand U7531 (N_7531,N_2601,N_2978);
or U7532 (N_7532,N_3681,N_4154);
or U7533 (N_7533,N_2180,N_5645);
nor U7534 (N_7534,N_225,N_5700);
or U7535 (N_7535,N_3574,N_4864);
xnor U7536 (N_7536,N_1531,N_3389);
xor U7537 (N_7537,N_3276,N_3736);
or U7538 (N_7538,N_2107,N_2794);
nor U7539 (N_7539,N_1585,N_2182);
or U7540 (N_7540,N_1270,N_621);
nand U7541 (N_7541,N_5031,N_4446);
nor U7542 (N_7542,N_1425,N_3302);
and U7543 (N_7543,N_2565,N_980);
nand U7544 (N_7544,N_1891,N_184);
and U7545 (N_7545,N_1216,N_4346);
nand U7546 (N_7546,N_3999,N_1089);
and U7547 (N_7547,N_4176,N_323);
xnor U7548 (N_7548,N_2358,N_5996);
nor U7549 (N_7549,N_2681,N_4046);
nor U7550 (N_7550,N_4610,N_4699);
xnor U7551 (N_7551,N_3669,N_3460);
or U7552 (N_7552,N_185,N_3042);
nand U7553 (N_7553,N_2884,N_1231);
or U7554 (N_7554,N_3748,N_1000);
or U7555 (N_7555,N_4546,N_5932);
and U7556 (N_7556,N_205,N_5660);
or U7557 (N_7557,N_3956,N_4902);
and U7558 (N_7558,N_3658,N_1093);
or U7559 (N_7559,N_5341,N_63);
and U7560 (N_7560,N_2190,N_4947);
nor U7561 (N_7561,N_2798,N_604);
or U7562 (N_7562,N_179,N_5707);
nand U7563 (N_7563,N_1442,N_4736);
or U7564 (N_7564,N_2991,N_4790);
or U7565 (N_7565,N_2046,N_5914);
or U7566 (N_7566,N_2012,N_2315);
xnor U7567 (N_7567,N_784,N_4041);
xnor U7568 (N_7568,N_4683,N_639);
nand U7569 (N_7569,N_1206,N_945);
or U7570 (N_7570,N_3485,N_622);
xor U7571 (N_7571,N_2184,N_4709);
and U7572 (N_7572,N_960,N_4497);
or U7573 (N_7573,N_5416,N_4469);
nor U7574 (N_7574,N_3394,N_4997);
nand U7575 (N_7575,N_2769,N_752);
and U7576 (N_7576,N_3061,N_4056);
xor U7577 (N_7577,N_4102,N_2449);
nor U7578 (N_7578,N_4645,N_3212);
and U7579 (N_7579,N_4084,N_2675);
or U7580 (N_7580,N_5927,N_4443);
or U7581 (N_7581,N_2450,N_37);
xor U7582 (N_7582,N_1734,N_3412);
nor U7583 (N_7583,N_4113,N_2743);
nand U7584 (N_7584,N_5273,N_1570);
nor U7585 (N_7585,N_608,N_5546);
nand U7586 (N_7586,N_3278,N_3568);
nor U7587 (N_7587,N_425,N_1816);
and U7588 (N_7588,N_1085,N_2458);
and U7589 (N_7589,N_1403,N_357);
nand U7590 (N_7590,N_4910,N_4774);
nand U7591 (N_7591,N_2004,N_4818);
and U7592 (N_7592,N_4604,N_3501);
nand U7593 (N_7593,N_61,N_3313);
xor U7594 (N_7594,N_5303,N_4982);
xor U7595 (N_7595,N_3580,N_510);
or U7596 (N_7596,N_2211,N_1704);
and U7597 (N_7597,N_3787,N_3805);
or U7598 (N_7598,N_3728,N_941);
or U7599 (N_7599,N_4082,N_2741);
xnor U7600 (N_7600,N_4540,N_2470);
and U7601 (N_7601,N_2498,N_905);
nand U7602 (N_7602,N_770,N_3200);
or U7603 (N_7603,N_5792,N_164);
nor U7604 (N_7604,N_3955,N_3764);
and U7605 (N_7605,N_1784,N_4347);
nor U7606 (N_7606,N_5172,N_1947);
nand U7607 (N_7607,N_5182,N_3850);
or U7608 (N_7608,N_3429,N_3621);
or U7609 (N_7609,N_4391,N_4574);
nor U7610 (N_7610,N_5016,N_5680);
xor U7611 (N_7611,N_5257,N_3715);
xor U7612 (N_7612,N_1277,N_4611);
and U7613 (N_7613,N_1237,N_4092);
or U7614 (N_7614,N_3354,N_3589);
nor U7615 (N_7615,N_2386,N_5072);
or U7616 (N_7616,N_1698,N_4164);
nor U7617 (N_7617,N_5398,N_777);
nor U7618 (N_7618,N_5839,N_4678);
nand U7619 (N_7619,N_224,N_424);
nand U7620 (N_7620,N_2188,N_946);
nor U7621 (N_7621,N_4420,N_2737);
nand U7622 (N_7622,N_4911,N_2028);
and U7623 (N_7623,N_3773,N_4878);
or U7624 (N_7624,N_5533,N_764);
nand U7625 (N_7625,N_5897,N_3615);
xnor U7626 (N_7626,N_3090,N_906);
xnor U7627 (N_7627,N_2643,N_5092);
or U7628 (N_7628,N_3148,N_4099);
or U7629 (N_7629,N_358,N_2924);
or U7630 (N_7630,N_3667,N_5293);
xor U7631 (N_7631,N_3666,N_1233);
nand U7632 (N_7632,N_1982,N_2532);
nor U7633 (N_7633,N_3771,N_3295);
xnor U7634 (N_7634,N_3886,N_3992);
nand U7635 (N_7635,N_2280,N_5065);
xnor U7636 (N_7636,N_1197,N_2981);
and U7637 (N_7637,N_753,N_211);
xnor U7638 (N_7638,N_1213,N_948);
and U7639 (N_7639,N_1994,N_535);
nand U7640 (N_7640,N_1973,N_1529);
nor U7641 (N_7641,N_457,N_1319);
nor U7642 (N_7642,N_5351,N_1986);
and U7643 (N_7643,N_5066,N_4723);
nand U7644 (N_7644,N_4771,N_1895);
nand U7645 (N_7645,N_330,N_3166);
nor U7646 (N_7646,N_5148,N_2913);
nor U7647 (N_7647,N_5837,N_1607);
nand U7648 (N_7648,N_3081,N_2288);
xnor U7649 (N_7649,N_3958,N_5190);
or U7650 (N_7650,N_3904,N_1449);
nand U7651 (N_7651,N_4675,N_5105);
xnor U7652 (N_7652,N_5534,N_2841);
and U7653 (N_7653,N_1035,N_628);
or U7654 (N_7654,N_4206,N_4399);
or U7655 (N_7655,N_2795,N_4681);
or U7656 (N_7656,N_2099,N_663);
and U7657 (N_7657,N_605,N_2500);
or U7658 (N_7658,N_1266,N_4567);
nand U7659 (N_7659,N_3228,N_796);
and U7660 (N_7660,N_3486,N_3602);
nor U7661 (N_7661,N_515,N_1415);
or U7662 (N_7662,N_3369,N_5878);
xor U7663 (N_7663,N_1440,N_4526);
nor U7664 (N_7664,N_3390,N_5858);
or U7665 (N_7665,N_2027,N_2070);
and U7666 (N_7666,N_2143,N_1423);
or U7667 (N_7667,N_2131,N_4669);
xor U7668 (N_7668,N_5840,N_4358);
or U7669 (N_7669,N_1412,N_5809);
or U7670 (N_7670,N_4927,N_2998);
nand U7671 (N_7671,N_4551,N_4886);
xnor U7672 (N_7672,N_2750,N_2898);
and U7673 (N_7673,N_3760,N_653);
xor U7674 (N_7674,N_2445,N_4035);
nor U7675 (N_7675,N_5748,N_3685);
or U7676 (N_7676,N_1015,N_2894);
or U7677 (N_7677,N_337,N_5594);
nand U7678 (N_7678,N_2151,N_1961);
nor U7679 (N_7679,N_822,N_4457);
or U7680 (N_7680,N_2945,N_5112);
nand U7681 (N_7681,N_272,N_3546);
nand U7682 (N_7682,N_488,N_932);
xnor U7683 (N_7683,N_3527,N_3914);
nor U7684 (N_7684,N_2121,N_4366);
xnor U7685 (N_7685,N_3638,N_4570);
nand U7686 (N_7686,N_1811,N_2030);
xor U7687 (N_7687,N_4156,N_867);
nor U7688 (N_7688,N_2699,N_2299);
nand U7689 (N_7689,N_4450,N_407);
or U7690 (N_7690,N_5784,N_1665);
or U7691 (N_7691,N_5628,N_3218);
nand U7692 (N_7692,N_578,N_1915);
xnor U7693 (N_7693,N_2657,N_940);
or U7694 (N_7694,N_3433,N_3399);
nand U7695 (N_7695,N_3283,N_4487);
nand U7696 (N_7696,N_115,N_651);
xor U7697 (N_7697,N_883,N_2413);
and U7698 (N_7698,N_3136,N_4097);
or U7699 (N_7699,N_2659,N_4541);
nor U7700 (N_7700,N_5420,N_5539);
or U7701 (N_7701,N_1331,N_2297);
nand U7702 (N_7702,N_300,N_3157);
and U7703 (N_7703,N_5166,N_5501);
and U7704 (N_7704,N_2538,N_1997);
and U7705 (N_7705,N_4310,N_5004);
nand U7706 (N_7706,N_262,N_3541);
and U7707 (N_7707,N_4359,N_1977);
and U7708 (N_7708,N_4376,N_3058);
nor U7709 (N_7709,N_5140,N_4643);
nor U7710 (N_7710,N_1666,N_54);
nand U7711 (N_7711,N_5342,N_4115);
xnor U7712 (N_7712,N_4782,N_2994);
and U7713 (N_7713,N_2725,N_4563);
xor U7714 (N_7714,N_2865,N_1545);
nand U7715 (N_7715,N_5524,N_908);
xor U7716 (N_7716,N_2765,N_3519);
nor U7717 (N_7717,N_2546,N_1434);
and U7718 (N_7718,N_477,N_3724);
or U7719 (N_7719,N_1489,N_2799);
xnor U7720 (N_7720,N_1393,N_5937);
nor U7721 (N_7721,N_3750,N_4528);
and U7722 (N_7722,N_523,N_4456);
nand U7723 (N_7723,N_871,N_2052);
xnor U7724 (N_7724,N_416,N_110);
xor U7725 (N_7725,N_1880,N_167);
nor U7726 (N_7726,N_267,N_3509);
nand U7727 (N_7727,N_691,N_2183);
nor U7728 (N_7728,N_2587,N_532);
xnor U7729 (N_7729,N_4294,N_1483);
or U7730 (N_7730,N_3075,N_4415);
nand U7731 (N_7731,N_2466,N_3739);
and U7732 (N_7732,N_5320,N_637);
and U7733 (N_7733,N_1713,N_5907);
nor U7734 (N_7734,N_1708,N_207);
xor U7735 (N_7735,N_2701,N_5160);
nor U7736 (N_7736,N_2063,N_306);
or U7737 (N_7737,N_3864,N_990);
and U7738 (N_7738,N_949,N_2605);
or U7739 (N_7739,N_4019,N_1911);
nor U7740 (N_7740,N_1335,N_1804);
nand U7741 (N_7741,N_4713,N_471);
or U7742 (N_7742,N_5891,N_3957);
nand U7743 (N_7743,N_551,N_3726);
or U7744 (N_7744,N_1108,N_5600);
nor U7745 (N_7745,N_1540,N_1723);
nor U7746 (N_7746,N_3467,N_2696);
nand U7747 (N_7747,N_1356,N_2833);
nor U7748 (N_7748,N_1591,N_2135);
nand U7749 (N_7749,N_860,N_1594);
xor U7750 (N_7750,N_3643,N_19);
xor U7751 (N_7751,N_328,N_2245);
nor U7752 (N_7752,N_4198,N_5974);
nand U7753 (N_7753,N_676,N_4573);
and U7754 (N_7754,N_5382,N_2390);
and U7755 (N_7755,N_3210,N_5067);
nand U7756 (N_7756,N_4409,N_526);
and U7757 (N_7757,N_890,N_3691);
xor U7758 (N_7758,N_5836,N_616);
or U7759 (N_7759,N_4654,N_5368);
xor U7760 (N_7760,N_776,N_3947);
nor U7761 (N_7761,N_2893,N_2600);
or U7762 (N_7762,N_5450,N_5243);
or U7763 (N_7763,N_3553,N_316);
or U7764 (N_7764,N_684,N_3231);
or U7765 (N_7765,N_5154,N_3147);
or U7766 (N_7766,N_4264,N_3644);
nand U7767 (N_7767,N_5818,N_4640);
nand U7768 (N_7768,N_4109,N_1905);
nand U7769 (N_7769,N_2686,N_5745);
nor U7770 (N_7770,N_228,N_5014);
xor U7771 (N_7771,N_1095,N_4510);
or U7772 (N_7772,N_5141,N_5637);
nand U7773 (N_7773,N_1097,N_4814);
nand U7774 (N_7774,N_3217,N_5074);
or U7775 (N_7775,N_730,N_4511);
and U7776 (N_7776,N_2669,N_292);
nand U7777 (N_7777,N_363,N_2877);
nor U7778 (N_7778,N_4425,N_1359);
nand U7779 (N_7779,N_2887,N_1913);
and U7780 (N_7780,N_4312,N_5207);
and U7781 (N_7781,N_41,N_1642);
or U7782 (N_7782,N_3609,N_1257);
and U7783 (N_7783,N_2838,N_2246);
nor U7784 (N_7784,N_3878,N_2702);
or U7785 (N_7785,N_1892,N_4411);
xnor U7786 (N_7786,N_2222,N_1615);
nand U7787 (N_7787,N_4393,N_702);
and U7788 (N_7788,N_1246,N_2950);
and U7789 (N_7789,N_1128,N_1274);
nand U7790 (N_7790,N_5225,N_1567);
xnor U7791 (N_7791,N_5104,N_4956);
nor U7792 (N_7792,N_1590,N_5864);
or U7793 (N_7793,N_5573,N_3983);
xor U7794 (N_7794,N_2338,N_1796);
nor U7795 (N_7795,N_3255,N_1969);
nor U7796 (N_7796,N_2212,N_3989);
nor U7797 (N_7797,N_398,N_3601);
xnor U7798 (N_7798,N_4590,N_4462);
nand U7799 (N_7799,N_4130,N_5488);
nand U7800 (N_7800,N_2979,N_2381);
nor U7801 (N_7801,N_3351,N_3678);
xnor U7802 (N_7802,N_430,N_797);
xnor U7803 (N_7803,N_1433,N_1042);
or U7804 (N_7804,N_1536,N_1761);
nor U7805 (N_7805,N_1224,N_1944);
or U7806 (N_7806,N_4285,N_2067);
and U7807 (N_7807,N_886,N_2857);
xor U7808 (N_7808,N_3063,N_5988);
xor U7809 (N_7809,N_327,N_3743);
xnor U7810 (N_7810,N_1584,N_828);
or U7811 (N_7811,N_5419,N_4328);
and U7812 (N_7812,N_436,N_2335);
xor U7813 (N_7813,N_5071,N_1551);
nand U7814 (N_7814,N_3626,N_5704);
nand U7815 (N_7815,N_5073,N_3828);
or U7816 (N_7816,N_4505,N_1468);
xnor U7817 (N_7817,N_3383,N_1240);
nor U7818 (N_7818,N_3808,N_2933);
and U7819 (N_7819,N_1681,N_837);
xnor U7820 (N_7820,N_4277,N_5101);
nand U7821 (N_7821,N_4263,N_1361);
nand U7822 (N_7822,N_4899,N_31);
xor U7823 (N_7823,N_156,N_3592);
and U7824 (N_7824,N_3274,N_4824);
and U7825 (N_7825,N_3285,N_4436);
or U7826 (N_7826,N_127,N_4354);
and U7827 (N_7827,N_2827,N_3585);
nor U7828 (N_7828,N_3729,N_1124);
nand U7829 (N_7829,N_1942,N_4116);
xnor U7830 (N_7830,N_522,N_5689);
nand U7831 (N_7831,N_3694,N_4649);
nor U7832 (N_7832,N_4292,N_117);
and U7833 (N_7833,N_5080,N_566);
or U7834 (N_7834,N_817,N_5993);
xnor U7835 (N_7835,N_2084,N_4141);
nor U7836 (N_7836,N_5344,N_5263);
nor U7837 (N_7837,N_501,N_5446);
and U7838 (N_7838,N_5179,N_640);
xor U7839 (N_7839,N_3327,N_2779);
xor U7840 (N_7840,N_2062,N_4245);
or U7841 (N_7841,N_2938,N_3201);
nor U7842 (N_7842,N_5910,N_1742);
or U7843 (N_7843,N_5739,N_2644);
or U7844 (N_7844,N_5626,N_2535);
nor U7845 (N_7845,N_4274,N_4784);
xor U7846 (N_7846,N_819,N_2923);
xor U7847 (N_7847,N_2009,N_1646);
and U7848 (N_7848,N_2077,N_5951);
and U7849 (N_7849,N_1722,N_3873);
nor U7850 (N_7850,N_3154,N_4142);
and U7851 (N_7851,N_1691,N_5000);
nand U7852 (N_7852,N_3528,N_5017);
and U7853 (N_7853,N_3340,N_3074);
or U7854 (N_7854,N_419,N_4993);
and U7855 (N_7855,N_2128,N_3316);
nor U7856 (N_7856,N_5911,N_3281);
or U7857 (N_7857,N_4919,N_3113);
nor U7858 (N_7858,N_5248,N_717);
or U7859 (N_7859,N_846,N_3552);
or U7860 (N_7860,N_2835,N_4517);
and U7861 (N_7861,N_1466,N_133);
or U7862 (N_7862,N_212,N_1100);
nor U7863 (N_7863,N_5885,N_293);
xor U7864 (N_7864,N_4952,N_380);
nand U7865 (N_7865,N_5842,N_1056);
and U7866 (N_7866,N_4913,N_2216);
nor U7867 (N_7867,N_4202,N_4533);
and U7868 (N_7868,N_827,N_5369);
or U7869 (N_7869,N_943,N_2198);
nand U7870 (N_7870,N_1995,N_1562);
nor U7871 (N_7871,N_4718,N_5566);
nand U7872 (N_7872,N_5713,N_4459);
and U7873 (N_7873,N_2969,N_308);
nor U7874 (N_7874,N_4932,N_4246);
and U7875 (N_7875,N_5799,N_3132);
xor U7876 (N_7876,N_5433,N_939);
nor U7877 (N_7877,N_3752,N_4585);
or U7878 (N_7878,N_2419,N_3657);
nand U7879 (N_7879,N_5356,N_3373);
nand U7880 (N_7880,N_1374,N_3243);
nor U7881 (N_7881,N_5132,N_3309);
or U7882 (N_7882,N_1882,N_5214);
nor U7883 (N_7883,N_4050,N_5791);
xnor U7884 (N_7884,N_657,N_4337);
and U7885 (N_7885,N_3245,N_5723);
and U7886 (N_7886,N_107,N_2302);
and U7887 (N_7887,N_4175,N_5890);
nand U7888 (N_7888,N_751,N_4379);
or U7889 (N_7889,N_869,N_4744);
nand U7890 (N_7890,N_2059,N_4897);
nand U7891 (N_7891,N_5131,N_5673);
nor U7892 (N_7892,N_934,N_102);
nand U7893 (N_7893,N_1072,N_395);
or U7894 (N_7894,N_3720,N_5608);
or U7895 (N_7895,N_2808,N_3414);
nand U7896 (N_7896,N_4125,N_1297);
nor U7897 (N_7897,N_740,N_3306);
nand U7898 (N_7898,N_2401,N_5059);
xnor U7899 (N_7899,N_3974,N_5040);
or U7900 (N_7900,N_5826,N_882);
and U7901 (N_7901,N_4614,N_2807);
nor U7902 (N_7902,N_5632,N_2871);
nand U7903 (N_7903,N_2344,N_4922);
or U7904 (N_7904,N_5463,N_5340);
nor U7905 (N_7905,N_74,N_3268);
nor U7906 (N_7906,N_757,N_3709);
nand U7907 (N_7907,N_1805,N_2289);
nand U7908 (N_7908,N_4080,N_2604);
or U7909 (N_7909,N_2721,N_3674);
or U7910 (N_7910,N_2874,N_5676);
or U7911 (N_7911,N_5705,N_3869);
and U7912 (N_7912,N_432,N_269);
or U7913 (N_7913,N_5593,N_4385);
nand U7914 (N_7914,N_448,N_4745);
nand U7915 (N_7915,N_3441,N_3421);
nor U7916 (N_7916,N_2624,N_5616);
xnor U7917 (N_7917,N_5970,N_4482);
or U7918 (N_7918,N_1159,N_3098);
xor U7919 (N_7919,N_695,N_5737);
nor U7920 (N_7920,N_3502,N_3372);
nor U7921 (N_7921,N_4617,N_2301);
or U7922 (N_7922,N_4032,N_4593);
or U7923 (N_7923,N_3505,N_396);
xor U7924 (N_7924,N_5663,N_2870);
and U7925 (N_7925,N_4127,N_4356);
nor U7926 (N_7926,N_5736,N_4161);
and U7927 (N_7927,N_1751,N_4706);
and U7928 (N_7928,N_825,N_2778);
xnor U7929 (N_7929,N_1576,N_1930);
or U7930 (N_7930,N_4619,N_2130);
and U7931 (N_7931,N_5896,N_4588);
nand U7932 (N_7932,N_5308,N_4959);
xor U7933 (N_7933,N_900,N_2582);
nor U7934 (N_7934,N_602,N_5879);
nor U7935 (N_7935,N_2930,N_1371);
nand U7936 (N_7936,N_277,N_4442);
xnor U7937 (N_7937,N_241,N_4213);
and U7938 (N_7938,N_4348,N_561);
xnor U7939 (N_7939,N_4106,N_3945);
xor U7940 (N_7940,N_284,N_5724);
and U7941 (N_7941,N_1718,N_5646);
nor U7942 (N_7942,N_5423,N_1810);
and U7943 (N_7943,N_2502,N_1373);
nor U7944 (N_7944,N_1432,N_2727);
or U7945 (N_7945,N_4565,N_4088);
and U7946 (N_7946,N_3906,N_1354);
nor U7947 (N_7947,N_4909,N_5383);
nand U7948 (N_7948,N_603,N_1148);
nor U7949 (N_7949,N_84,N_5603);
or U7950 (N_7950,N_1444,N_3581);
nor U7951 (N_7951,N_1129,N_885);
xnor U7952 (N_7952,N_2635,N_3920);
or U7953 (N_7953,N_3504,N_1474);
and U7954 (N_7954,N_5952,N_5969);
and U7955 (N_7955,N_3472,N_4260);
and U7956 (N_7956,N_3915,N_2876);
nor U7957 (N_7957,N_356,N_5597);
nand U7958 (N_7958,N_314,N_3753);
or U7959 (N_7959,N_858,N_4003);
or U7960 (N_7960,N_2666,N_4455);
nor U7961 (N_7961,N_3093,N_5431);
xor U7962 (N_7962,N_1227,N_5717);
and U7963 (N_7963,N_1846,N_1541);
xnor U7964 (N_7964,N_1454,N_3362);
nand U7965 (N_7965,N_3665,N_4273);
or U7966 (N_7966,N_157,N_466);
nor U7967 (N_7967,N_1663,N_4453);
and U7968 (N_7968,N_2375,N_2024);
nor U7969 (N_7969,N_2552,N_3543);
nor U7970 (N_7970,N_1825,N_5560);
nand U7971 (N_7971,N_3907,N_2452);
and U7972 (N_7972,N_720,N_5759);
xnor U7973 (N_7973,N_2061,N_1105);
and U7974 (N_7974,N_3506,N_1283);
nand U7975 (N_7975,N_1690,N_1878);
or U7976 (N_7976,N_1785,N_675);
nor U7977 (N_7977,N_3783,N_2136);
or U7978 (N_7978,N_619,N_3346);
or U7979 (N_7979,N_1600,N_5375);
and U7980 (N_7980,N_4690,N_3303);
or U7981 (N_7981,N_5772,N_4316);
nand U7982 (N_7982,N_3223,N_2428);
nor U7983 (N_7983,N_3734,N_861);
nor U7984 (N_7984,N_5964,N_5761);
xnor U7985 (N_7985,N_4809,N_5819);
nor U7986 (N_7986,N_712,N_563);
nor U7987 (N_7987,N_4757,N_1844);
nor U7988 (N_7988,N_4211,N_4485);
nand U7989 (N_7989,N_3740,N_5953);
nand U7990 (N_7990,N_4463,N_1689);
xor U7991 (N_7991,N_3972,N_32);
and U7992 (N_7992,N_3921,N_1616);
or U7993 (N_7993,N_5625,N_4295);
nand U7994 (N_7994,N_1537,N_1569);
nand U7995 (N_7995,N_2773,N_3522);
and U7996 (N_7996,N_5728,N_5264);
nand U7997 (N_7997,N_2956,N_5349);
xnor U7998 (N_7998,N_1660,N_2483);
nand U7999 (N_7999,N_5875,N_3571);
and U8000 (N_8000,N_3438,N_116);
and U8001 (N_8001,N_5328,N_3114);
xnor U8002 (N_8002,N_1420,N_5255);
nand U8003 (N_8003,N_3693,N_5240);
nand U8004 (N_8004,N_2544,N_5267);
and U8005 (N_8005,N_2782,N_5405);
xor U8006 (N_8006,N_2831,N_4454);
or U8007 (N_8007,N_3183,N_2817);
and U8008 (N_8008,N_3349,N_3029);
nor U8009 (N_8009,N_4300,N_5475);
nor U8010 (N_8010,N_4833,N_4373);
nand U8011 (N_8011,N_4877,N_1205);
nor U8012 (N_8012,N_4200,N_3162);
and U8013 (N_8013,N_3521,N_4001);
nand U8014 (N_8014,N_3710,N_3747);
nand U8015 (N_8015,N_1222,N_5850);
nor U8016 (N_8016,N_5884,N_3822);
nand U8017 (N_8017,N_1123,N_1881);
and U8018 (N_8018,N_1041,N_2576);
xnor U8019 (N_8019,N_350,N_2882);
or U8020 (N_8020,N_3525,N_2907);
xor U8021 (N_8021,N_5083,N_480);
nand U8022 (N_8022,N_222,N_647);
or U8023 (N_8023,N_2632,N_239);
or U8024 (N_8024,N_1993,N_5617);
xnor U8025 (N_8025,N_1596,N_2393);
xnor U8026 (N_8026,N_1428,N_688);
xnor U8027 (N_8027,N_307,N_335);
xor U8028 (N_8028,N_4394,N_3855);
or U8029 (N_8029,N_5487,N_1774);
nor U8030 (N_8030,N_4045,N_2555);
nand U8031 (N_8031,N_1346,N_3610);
nand U8032 (N_8032,N_2377,N_1046);
and U8033 (N_8033,N_3045,N_5523);
nand U8034 (N_8034,N_1682,N_5661);
nor U8035 (N_8035,N_4233,N_2340);
and U8036 (N_8036,N_180,N_4844);
nand U8037 (N_8037,N_705,N_4561);
or U8038 (N_8038,N_5541,N_667);
xnor U8039 (N_8039,N_1928,N_5061);
nor U8040 (N_8040,N_4545,N_3766);
and U8041 (N_8041,N_2946,N_2410);
xnor U8042 (N_8042,N_4894,N_2366);
nand U8043 (N_8043,N_696,N_1509);
or U8044 (N_8044,N_2278,N_4413);
xnor U8045 (N_8045,N_902,N_2717);
and U8046 (N_8046,N_5478,N_2674);
nor U8047 (N_8047,N_5078,N_1817);
nor U8048 (N_8048,N_3341,N_1855);
nand U8049 (N_8049,N_4986,N_2836);
and U8050 (N_8050,N_4301,N_5130);
nor U8051 (N_8051,N_5134,N_630);
and U8052 (N_8052,N_166,N_5699);
xnor U8053 (N_8053,N_3582,N_5124);
nor U8054 (N_8054,N_3688,N_5113);
or U8055 (N_8055,N_3324,N_5064);
nor U8056 (N_8056,N_3415,N_5454);
xor U8057 (N_8057,N_1573,N_3514);
xnor U8058 (N_8058,N_4612,N_3142);
or U8059 (N_8059,N_4361,N_3675);
or U8060 (N_8060,N_4715,N_1033);
xor U8061 (N_8061,N_3996,N_2683);
xor U8062 (N_8062,N_718,N_2365);
and U8063 (N_8063,N_937,N_1113);
or U8064 (N_8064,N_3963,N_1904);
xnor U8065 (N_8065,N_3751,N_1743);
xor U8066 (N_8066,N_2441,N_4012);
nor U8067 (N_8067,N_1024,N_2603);
nand U8068 (N_8068,N_283,N_4224);
nand U8069 (N_8069,N_4009,N_4189);
nor U8070 (N_8070,N_3450,N_2207);
or U8071 (N_8071,N_2568,N_1378);
nand U8072 (N_8072,N_4276,N_788);
and U8073 (N_8073,N_472,N_3903);
nand U8074 (N_8074,N_483,N_5709);
nand U8075 (N_8075,N_4016,N_5298);
nand U8076 (N_8076,N_5805,N_5710);
xor U8077 (N_8077,N_1386,N_1771);
nor U8078 (N_8078,N_2684,N_2414);
xnor U8079 (N_8079,N_5436,N_5575);
nor U8080 (N_8080,N_1406,N_1341);
or U8081 (N_8081,N_2422,N_1333);
xnor U8082 (N_8082,N_650,N_4767);
nor U8083 (N_8083,N_5370,N_5815);
nor U8084 (N_8084,N_5023,N_3207);
nand U8085 (N_8085,N_3128,N_175);
nor U8086 (N_8086,N_4797,N_1392);
or U8087 (N_8087,N_2829,N_4830);
nand U8088 (N_8088,N_4026,N_910);
or U8089 (N_8089,N_5169,N_878);
and U8090 (N_8090,N_4670,N_2797);
nor U8091 (N_8091,N_58,N_3704);
and U8092 (N_8092,N_230,N_1151);
and U8093 (N_8093,N_2101,N_3980);
or U8094 (N_8094,N_708,N_3741);
and U8095 (N_8095,N_2373,N_2405);
or U8096 (N_8096,N_4471,N_550);
nand U8097 (N_8097,N_3064,N_4392);
xnor U8098 (N_8098,N_3363,N_2047);
nand U8099 (N_8099,N_5415,N_4133);
nand U8100 (N_8100,N_5926,N_1546);
xnor U8101 (N_8101,N_3425,N_4257);
nand U8102 (N_8102,N_2580,N_2332);
nor U8103 (N_8103,N_3457,N_4775);
xor U8104 (N_8104,N_3187,N_4647);
xnor U8105 (N_8105,N_5307,N_3107);
or U8106 (N_8106,N_5381,N_4560);
xnor U8107 (N_8107,N_4882,N_4293);
or U8108 (N_8108,N_3965,N_5335);
nand U8109 (N_8109,N_1979,N_706);
xnor U8110 (N_8110,N_3016,N_4726);
nand U8111 (N_8111,N_3881,N_4438);
nor U8112 (N_8112,N_5670,N_4483);
or U8113 (N_8113,N_5904,N_2735);
xnor U8114 (N_8114,N_4872,N_1787);
nand U8115 (N_8115,N_3164,N_5084);
xor U8116 (N_8116,N_2399,N_5226);
xnor U8117 (N_8117,N_2076,N_1506);
nor U8118 (N_8118,N_5909,N_2453);
xnor U8119 (N_8119,N_2327,N_5152);
xor U8120 (N_8120,N_1894,N_3492);
and U8121 (N_8121,N_652,N_2537);
nand U8122 (N_8122,N_3628,N_1657);
nor U8123 (N_8123,N_5671,N_803);
and U8124 (N_8124,N_113,N_5785);
xnor U8125 (N_8125,N_947,N_364);
nand U8126 (N_8126,N_2734,N_3440);
nand U8127 (N_8127,N_749,N_1589);
nand U8128 (N_8128,N_2578,N_3190);
nand U8129 (N_8129,N_787,N_4979);
xor U8130 (N_8130,N_2022,N_5787);
nand U8131 (N_8131,N_724,N_5098);
or U8132 (N_8132,N_4248,N_3532);
xor U8133 (N_8133,N_1619,N_3014);
or U8134 (N_8134,N_1212,N_5491);
and U8135 (N_8135,N_3690,N_5950);
and U8136 (N_8136,N_4778,N_2050);
xor U8137 (N_8137,N_3587,N_2563);
nor U8138 (N_8138,N_3613,N_4157);
and U8139 (N_8139,N_1102,N_673);
nand U8140 (N_8140,N_5467,N_4626);
and U8141 (N_8141,N_5652,N_5052);
and U8142 (N_8142,N_4036,N_4410);
nor U8143 (N_8143,N_5916,N_3813);
nor U8144 (N_8144,N_2545,N_1318);
or U8145 (N_8145,N_2610,N_4697);
nand U8146 (N_8146,N_2548,N_2037);
and U8147 (N_8147,N_382,N_4513);
and U8148 (N_8148,N_4451,N_5921);
xnor U8149 (N_8149,N_1235,N_3443);
or U8150 (N_8150,N_4105,N_2132);
xor U8151 (N_8151,N_4345,N_5750);
xor U8152 (N_8152,N_4707,N_573);
nand U8153 (N_8153,N_952,N_2442);
and U8154 (N_8154,N_186,N_5282);
and U8155 (N_8155,N_935,N_2748);
xor U8156 (N_8156,N_693,N_5219);
nand U8157 (N_8157,N_3924,N_1869);
or U8158 (N_8158,N_2996,N_641);
nor U8159 (N_8159,N_3053,N_5945);
nand U8160 (N_8160,N_4898,N_4020);
xor U8161 (N_8161,N_403,N_3642);
and U8162 (N_8162,N_5811,N_1477);
nand U8163 (N_8163,N_4498,N_2768);
nand U8164 (N_8164,N_1559,N_4742);
xnor U8165 (N_8165,N_2251,N_3821);
nor U8166 (N_8166,N_4222,N_1180);
or U8167 (N_8167,N_3865,N_1031);
nand U8168 (N_8168,N_226,N_747);
nand U8169 (N_8169,N_497,N_5779);
or U8170 (N_8170,N_5276,N_4873);
or U8171 (N_8171,N_801,N_1847);
or U8172 (N_8172,N_5203,N_4766);
or U8173 (N_8173,N_4094,N_5643);
or U8174 (N_8174,N_2096,N_3445);
nand U8175 (N_8175,N_4812,N_2232);
and U8176 (N_8176,N_1272,N_3198);
and U8177 (N_8177,N_1175,N_4475);
xor U8178 (N_8178,N_2179,N_5529);
or U8179 (N_8179,N_2181,N_3138);
nor U8180 (N_8180,N_798,N_5464);
or U8181 (N_8181,N_3311,N_1383);
nor U8182 (N_8182,N_1760,N_4635);
or U8183 (N_8183,N_2971,N_2274);
xor U8184 (N_8184,N_4942,N_3427);
nand U8185 (N_8185,N_3026,N_2193);
and U8186 (N_8186,N_2736,N_1281);
or U8187 (N_8187,N_1530,N_1842);
nor U8188 (N_8188,N_4204,N_686);
nor U8189 (N_8189,N_3101,N_5495);
xnor U8190 (N_8190,N_5258,N_3476);
nand U8191 (N_8191,N_5470,N_1726);
nor U8192 (N_8192,N_3863,N_2569);
and U8193 (N_8193,N_5979,N_5558);
nand U8194 (N_8194,N_1456,N_1983);
and U8195 (N_8195,N_5861,N_1029);
nand U8196 (N_8196,N_5136,N_3197);
or U8197 (N_8197,N_5977,N_5473);
or U8198 (N_8198,N_3003,N_3044);
nand U8199 (N_8199,N_62,N_5146);
xor U8200 (N_8200,N_3236,N_1192);
or U8201 (N_8201,N_4120,N_473);
nand U8202 (N_8202,N_4122,N_4331);
and U8203 (N_8203,N_5323,N_2818);
and U8204 (N_8204,N_4150,N_925);
xnor U8205 (N_8205,N_2805,N_3335);
nand U8206 (N_8206,N_5496,N_843);
nand U8207 (N_8207,N_5041,N_3056);
xnor U8208 (N_8208,N_4441,N_1040);
or U8209 (N_8209,N_4480,N_774);
nand U8210 (N_8210,N_5334,N_4040);
or U8211 (N_8211,N_4087,N_2760);
and U8212 (N_8212,N_4853,N_3549);
and U8213 (N_8213,N_4534,N_1933);
xor U8214 (N_8214,N_823,N_2255);
nor U8215 (N_8215,N_617,N_2126);
nand U8216 (N_8216,N_4279,N_1411);
nor U8217 (N_8217,N_2192,N_4985);
nor U8218 (N_8218,N_5960,N_4628);
and U8219 (N_8219,N_4048,N_464);
and U8220 (N_8220,N_86,N_20);
xor U8221 (N_8221,N_5681,N_3452);
nor U8222 (N_8222,N_444,N_4386);
nand U8223 (N_8223,N_4090,N_4140);
and U8224 (N_8224,N_1627,N_4529);
nand U8225 (N_8225,N_636,N_4623);
xor U8226 (N_8226,N_938,N_2614);
or U8227 (N_8227,N_5948,N_3988);
and U8228 (N_8228,N_4754,N_2247);
nor U8229 (N_8229,N_2283,N_5725);
and U8230 (N_8230,N_3647,N_2709);
or U8231 (N_8231,N_45,N_2848);
xnor U8232 (N_8232,N_4964,N_2271);
xor U8233 (N_8233,N_2026,N_5746);
xnor U8234 (N_8234,N_4,N_5866);
nand U8235 (N_8235,N_4362,N_4918);
nand U8236 (N_8236,N_1465,N_5522);
nand U8237 (N_8237,N_677,N_4554);
and U8238 (N_8238,N_3627,N_443);
xor U8239 (N_8239,N_214,N_4069);
nand U8240 (N_8240,N_3288,N_530);
and U8241 (N_8241,N_1659,N_919);
and U8242 (N_8242,N_454,N_5997);
nand U8243 (N_8243,N_5547,N_2637);
nor U8244 (N_8244,N_3578,N_4208);
nor U8245 (N_8245,N_728,N_254);
xor U8246 (N_8246,N_1068,N_1680);
and U8247 (N_8247,N_3163,N_2920);
nand U8248 (N_8248,N_121,N_4710);
and U8249 (N_8249,N_5845,N_1058);
nor U8250 (N_8250,N_3194,N_5694);
or U8251 (N_8251,N_1898,N_3151);
nor U8252 (N_8252,N_3206,N_2354);
nand U8253 (N_8253,N_1877,N_3247);
xnor U8254 (N_8254,N_1250,N_4104);
nand U8255 (N_8255,N_2912,N_4238);
or U8256 (N_8256,N_2055,N_3337);
or U8257 (N_8257,N_904,N_5808);
or U8258 (N_8258,N_1676,N_2384);
and U8259 (N_8259,N_76,N_1424);
nand U8260 (N_8260,N_3124,N_1800);
nand U8261 (N_8261,N_4013,N_3887);
xnor U8262 (N_8262,N_5277,N_3043);
or U8263 (N_8263,N_5873,N_296);
or U8264 (N_8264,N_2630,N_5486);
or U8265 (N_8265,N_3979,N_754);
nor U8266 (N_8266,N_748,N_1696);
xor U8267 (N_8267,N_549,N_5928);
or U8268 (N_8268,N_5882,N_642);
nor U8269 (N_8269,N_1793,N_789);
and U8270 (N_8270,N_5185,N_4837);
xnor U8271 (N_8271,N_2173,N_5194);
nand U8272 (N_8272,N_2263,N_5806);
nor U8273 (N_8273,N_1757,N_360);
or U8274 (N_8274,N_1951,N_5205);
xnor U8275 (N_8275,N_233,N_1672);
xor U8276 (N_8276,N_118,N_4255);
nor U8277 (N_8277,N_4072,N_5096);
and U8278 (N_8278,N_3899,N_3900);
xor U8279 (N_8279,N_4174,N_3391);
nand U8280 (N_8280,N_1868,N_312);
xnor U8281 (N_8281,N_2175,N_857);
nand U8282 (N_8282,N_3827,N_3339);
nor U8283 (N_8283,N_4329,N_4934);
nand U8284 (N_8284,N_5384,N_2993);
and U8285 (N_8285,N_1011,N_2792);
nand U8286 (N_8286,N_3816,N_3428);
nor U8287 (N_8287,N_5302,N_3304);
xnor U8288 (N_8288,N_5639,N_5361);
and U8289 (N_8289,N_4769,N_3700);
nor U8290 (N_8290,N_4280,N_918);
nand U8291 (N_8291,N_5564,N_3203);
or U8292 (N_8292,N_3927,N_5333);
and U8293 (N_8293,N_3926,N_5339);
or U8294 (N_8294,N_4970,N_2201);
and U8295 (N_8295,N_2724,N_3455);
nand U8296 (N_8296,N_4801,N_609);
or U8297 (N_8297,N_1896,N_3347);
and U8298 (N_8298,N_2090,N_94);
xnor U8299 (N_8299,N_4555,N_3384);
and U8300 (N_8300,N_1006,N_3465);
or U8301 (N_8301,N_192,N_3159);
and U8302 (N_8302,N_1447,N_4311);
or U8303 (N_8303,N_5619,N_3032);
xor U8304 (N_8304,N_10,N_4435);
nor U8305 (N_8305,N_2093,N_4521);
nand U8306 (N_8306,N_4434,N_5198);
and U8307 (N_8307,N_782,N_5477);
nor U8308 (N_8308,N_3620,N_5296);
xnor U8309 (N_8309,N_654,N_624);
nand U8310 (N_8310,N_802,N_2574);
nand U8311 (N_8311,N_149,N_5606);
xnor U8312 (N_8312,N_2708,N_3184);
or U8313 (N_8313,N_2958,N_2363);
or U8314 (N_8314,N_373,N_2144);
nor U8315 (N_8315,N_1860,N_3551);
or U8316 (N_8316,N_4747,N_4931);
or U8317 (N_8317,N_3702,N_2622);
or U8318 (N_8318,N_5306,N_4556);
nor U8319 (N_8319,N_1118,N_4724);
or U8320 (N_8320,N_4449,N_3577);
nand U8321 (N_8321,N_1367,N_2339);
and U8322 (N_8322,N_5505,N_4881);
nand U8323 (N_8323,N_5727,N_2204);
nand U8324 (N_8324,N_5994,N_4170);
nand U8325 (N_8325,N_26,N_1831);
or U8326 (N_8326,N_4578,N_1232);
nor U8327 (N_8327,N_1300,N_1667);
nand U8328 (N_8328,N_5070,N_4406);
nand U8329 (N_8329,N_2640,N_2949);
and U8330 (N_8330,N_4817,N_5047);
xor U8331 (N_8331,N_4014,N_1323);
or U8332 (N_8332,N_3189,N_5548);
or U8333 (N_8333,N_5300,N_4680);
nor U8334 (N_8334,N_3649,N_3331);
nor U8335 (N_8335,N_809,N_4672);
xnor U8336 (N_8336,N_864,N_5202);
nor U8337 (N_8337,N_1949,N_5032);
xnor U8338 (N_8338,N_476,N_2740);
xnor U8339 (N_8339,N_700,N_1561);
xnor U8340 (N_8340,N_5584,N_2364);
xnor U8341 (N_8341,N_5481,N_1045);
nand U8342 (N_8342,N_5883,N_4725);
nor U8343 (N_8343,N_3765,N_5060);
and U8344 (N_8344,N_1501,N_189);
nand U8345 (N_8345,N_4799,N_4738);
nor U8346 (N_8346,N_575,N_1324);
nand U8347 (N_8347,N_2787,N_1788);
xnor U8348 (N_8348,N_4191,N_997);
nor U8349 (N_8349,N_5925,N_1927);
nor U8350 (N_8350,N_5315,N_996);
or U8351 (N_8351,N_1309,N_759);
nor U8352 (N_8352,N_3317,N_2921);
or U8353 (N_8353,N_1622,N_662);
xor U8354 (N_8354,N_3411,N_3033);
or U8355 (N_8355,N_2269,N_2103);
nand U8356 (N_8356,N_2342,N_5466);
and U8357 (N_8357,N_5613,N_3237);
nand U8358 (N_8358,N_5991,N_2900);
and U8359 (N_8359,N_5651,N_2031);
nand U8360 (N_8360,N_298,N_5186);
nand U8361 (N_8361,N_4207,N_4011);
or U8362 (N_8362,N_4532,N_1462);
xnor U8363 (N_8363,N_5990,N_1775);
nor U8364 (N_8364,N_5888,N_2855);
or U8365 (N_8365,N_3484,N_2733);
nor U8366 (N_8366,N_5913,N_1835);
nor U8367 (N_8367,N_4684,N_5346);
and U8368 (N_8368,N_5149,N_1705);
nor U8369 (N_8369,N_1999,N_4582);
or U8370 (N_8370,N_3689,N_2639);
and U8371 (N_8371,N_4322,N_5886);
or U8372 (N_8372,N_2075,N_1251);
nand U8373 (N_8373,N_715,N_4071);
nand U8374 (N_8374,N_3031,N_353);
nand U8375 (N_8375,N_120,N_2471);
xnor U8376 (N_8376,N_5844,N_1168);
nor U8377 (N_8377,N_3892,N_2623);
or U8378 (N_8378,N_2518,N_4057);
nor U8379 (N_8379,N_2917,N_3378);
nor U8380 (N_8380,N_2374,N_2951);
or U8381 (N_8381,N_3121,N_1572);
and U8382 (N_8382,N_57,N_4793);
xnor U8383 (N_8383,N_2208,N_1996);
and U8384 (N_8384,N_1974,N_1548);
and U8385 (N_8385,N_3684,N_3039);
and U8386 (N_8386,N_2356,N_5683);
nor U8387 (N_8387,N_1597,N_2551);
xor U8388 (N_8388,N_3225,N_4333);
or U8389 (N_8389,N_4472,N_4600);
nand U8390 (N_8390,N_1060,N_2407);
or U8391 (N_8391,N_2579,N_2804);
nand U8392 (N_8392,N_3251,N_3348);
nand U8393 (N_8393,N_4583,N_1154);
xor U8394 (N_8394,N_2915,N_5797);
nor U8395 (N_8395,N_440,N_4378);
xnor U8396 (N_8396,N_4987,N_3634);
or U8397 (N_8397,N_4903,N_839);
and U8398 (N_8398,N_545,N_4155);
xnor U8399 (N_8399,N_3320,N_2042);
nor U8400 (N_8400,N_3461,N_3001);
or U8401 (N_8401,N_5857,N_1164);
xnor U8402 (N_8402,N_3286,N_2202);
xnor U8403 (N_8403,N_1018,N_5544);
nor U8404 (N_8404,N_4098,N_668);
xnor U8405 (N_8405,N_3294,N_2507);
nand U8406 (N_8406,N_3981,N_2306);
and U8407 (N_8407,N_5776,N_2881);
or U8408 (N_8408,N_4787,N_1782);
nor U8409 (N_8409,N_3297,N_2786);
or U8410 (N_8410,N_2504,N_2495);
nand U8411 (N_8411,N_55,N_4846);
and U8412 (N_8412,N_1016,N_4867);
nand U8413 (N_8413,N_3322,N_1611);
and U8414 (N_8414,N_623,N_2560);
and U8415 (N_8415,N_893,N_2347);
nand U8416 (N_8416,N_983,N_2420);
or U8417 (N_8417,N_4132,N_4991);
and U8418 (N_8418,N_4928,N_3024);
nand U8419 (N_8419,N_5285,N_5188);
and U8420 (N_8420,N_543,N_1171);
nor U8421 (N_8421,N_3735,N_33);
xor U8422 (N_8422,N_3767,N_4318);
nor U8423 (N_8423,N_3178,N_3801);
xnor U8424 (N_8424,N_1840,N_2712);
nand U8425 (N_8425,N_3208,N_5574);
or U8426 (N_8426,N_5918,N_1304);
and U8427 (N_8427,N_1295,N_3960);
nand U8428 (N_8428,N_4306,N_4861);
or U8429 (N_8429,N_449,N_1315);
and U8430 (N_8430,N_15,N_1884);
nand U8431 (N_8431,N_1372,N_1389);
and U8432 (N_8432,N_4467,N_4572);
xor U8433 (N_8433,N_4481,N_5043);
xor U8434 (N_8434,N_5452,N_2451);
nor U8435 (N_8435,N_2904,N_3970);
and U8436 (N_8436,N_2762,N_5917);
nor U8437 (N_8437,N_2596,N_5422);
xnor U8438 (N_8438,N_2343,N_1201);
or U8439 (N_8439,N_5510,N_439);
nor U8440 (N_8440,N_88,N_2570);
and U8441 (N_8441,N_1736,N_1727);
and U8442 (N_8442,N_1934,N_4703);
xnor U8443 (N_8443,N_5731,N_299);
nand U8444 (N_8444,N_2312,N_3998);
and U8445 (N_8445,N_178,N_3041);
or U8446 (N_8446,N_1394,N_3933);
xnor U8447 (N_8447,N_5242,N_5963);
or U8448 (N_8448,N_1178,N_3334);
and U8449 (N_8449,N_4815,N_2007);
xnor U8450 (N_8450,N_5777,N_1650);
and U8451 (N_8451,N_3222,N_446);
nor U8452 (N_8452,N_5511,N_3006);
xor U8453 (N_8453,N_5191,N_2239);
nor U8454 (N_8454,N_351,N_1200);
and U8455 (N_8455,N_810,N_5915);
or U8456 (N_8456,N_4184,N_2295);
nand U8457 (N_8457,N_67,N_3397);
nor U8458 (N_8458,N_195,N_4445);
nor U8459 (N_8459,N_4492,N_2947);
or U8460 (N_8460,N_2286,N_954);
or U8461 (N_8461,N_4562,N_4869);
or U8462 (N_8462,N_2237,N_1748);
nor U8463 (N_8463,N_1437,N_1737);
nor U8464 (N_8464,N_3261,N_2816);
xor U8465 (N_8465,N_1388,N_4353);
and U8466 (N_8466,N_1967,N_5376);
nor U8467 (N_8467,N_4179,N_4914);
or U8468 (N_8468,N_2955,N_3826);
or U8469 (N_8469,N_1923,N_3759);
nand U8470 (N_8470,N_5771,N_2241);
nand U8471 (N_8471,N_5537,N_2437);
or U8472 (N_8472,N_1647,N_336);
and U8473 (N_8473,N_3523,N_671);
or U8474 (N_8474,N_5387,N_3172);
nor U8475 (N_8475,N_2869,N_1119);
nand U8476 (N_8476,N_4478,N_958);
or U8477 (N_8477,N_1401,N_4691);
nand U8478 (N_8478,N_1395,N_4652);
or U8479 (N_8479,N_3489,N_3355);
nor U8480 (N_8480,N_5618,N_4249);
or U8481 (N_8481,N_3453,N_5364);
nand U8482 (N_8482,N_4544,N_3215);
xnor U8483 (N_8483,N_1344,N_3350);
nand U8484 (N_8484,N_5378,N_5038);
xor U8485 (N_8485,N_4317,N_4557);
nand U8486 (N_8486,N_3273,N_3848);
or U8487 (N_8487,N_5685,N_1989);
nand U8488 (N_8488,N_1872,N_4620);
xnor U8489 (N_8489,N_408,N_594);
and U8490 (N_8490,N_4054,N_4229);
or U8491 (N_8491,N_2670,N_1710);
xor U8492 (N_8492,N_2753,N_1498);
nand U8493 (N_8493,N_4866,N_3576);
nor U8494 (N_8494,N_3775,N_442);
xor U8495 (N_8495,N_5213,N_4021);
nor U8496 (N_8496,N_2885,N_4983);
xor U8497 (N_8497,N_3395,N_5856);
nand U8498 (N_8498,N_831,N_1229);
or U8499 (N_8499,N_4900,N_3594);
and U8500 (N_8500,N_2822,N_1802);
nor U8501 (N_8501,N_2986,N_1166);
xor U8502 (N_8502,N_3711,N_1413);
nand U8503 (N_8503,N_14,N_1132);
and U8504 (N_8504,N_2984,N_2916);
or U8505 (N_8505,N_1067,N_1370);
or U8506 (N_8506,N_2651,N_1907);
or U8507 (N_8507,N_555,N_5123);
nor U8508 (N_8508,N_3831,N_4820);
or U8509 (N_8509,N_4060,N_3305);
and U8510 (N_8510,N_2087,N_1630);
nor U8511 (N_8511,N_2257,N_5449);
and U8512 (N_8512,N_4460,N_3077);
nand U8513 (N_8513,N_832,N_4448);
and U8514 (N_8514,N_17,N_4501);
nand U8515 (N_8515,N_288,N_1724);
nand U8516 (N_8516,N_1701,N_1244);
or U8517 (N_8517,N_3105,N_4616);
nand U8518 (N_8518,N_3588,N_2990);
or U8519 (N_8519,N_5170,N_1075);
or U8520 (N_8520,N_4990,N_2361);
and U8521 (N_8521,N_1586,N_5111);
or U8522 (N_8522,N_546,N_2615);
or U8523 (N_8523,N_3851,N_899);
and U8524 (N_8524,N_2081,N_2455);
nor U8525 (N_8525,N_5528,N_3419);
nand U8526 (N_8526,N_991,N_4876);
or U8527 (N_8527,N_2396,N_4153);
nand U8528 (N_8528,N_3896,N_5531);
and U8529 (N_8529,N_3038,N_3240);
xnor U8530 (N_8530,N_5526,N_5972);
nor U8531 (N_8531,N_93,N_3110);
nor U8532 (N_8532,N_1950,N_2157);
nor U8533 (N_8533,N_1852,N_3991);
nor U8534 (N_8534,N_387,N_2677);
nor U8535 (N_8535,N_4387,N_5516);
xnor U8536 (N_8536,N_556,N_5456);
xnor U8537 (N_8537,N_3256,N_3742);
and U8538 (N_8538,N_4880,N_2726);
nand U8539 (N_8539,N_713,N_1188);
nor U8540 (N_8540,N_368,N_5218);
and U8541 (N_8541,N_3789,N_611);
or U8542 (N_8542,N_1874,N_3557);
or U8543 (N_8543,N_182,N_2117);
xnor U8544 (N_8544,N_4418,N_5357);
nor U8545 (N_8545,N_1721,N_1925);
or U8546 (N_8546,N_1610,N_3375);
and U8547 (N_8547,N_1972,N_4168);
nor U8548 (N_8548,N_4111,N_887);
and U8549 (N_8549,N_1435,N_5200);
nand U8550 (N_8550,N_1521,N_4327);
and U8551 (N_8551,N_4192,N_3277);
and U8552 (N_8552,N_3730,N_3849);
nand U8553 (N_8553,N_3343,N_2011);
xor U8554 (N_8554,N_2434,N_5581);
xor U8555 (N_8555,N_3352,N_3246);
nand U8556 (N_8556,N_4776,N_1871);
and U8557 (N_8557,N_1025,N_2417);
nand U8558 (N_8558,N_1879,N_3952);
nand U8559 (N_8559,N_2378,N_3139);
and U8560 (N_8560,N_853,N_5783);
nand U8561 (N_8561,N_5163,N_5517);
nor U8562 (N_8562,N_3778,N_1017);
nand U8563 (N_8563,N_124,N_5122);
xnor U8564 (N_8564,N_618,N_5399);
xnor U8565 (N_8565,N_2849,N_2494);
nand U8566 (N_8566,N_5373,N_1248);
nor U8567 (N_8567,N_4390,N_583);
and U8568 (N_8568,N_2519,N_3100);
or U8569 (N_8569,N_103,N_2845);
and U8570 (N_8570,N_5459,N_1883);
nand U8571 (N_8571,N_3379,N_2523);
xor U8572 (N_8572,N_2000,N_3815);
or U8573 (N_8573,N_1965,N_3018);
or U8574 (N_8574,N_5568,N_141);
nor U8575 (N_8575,N_3844,N_331);
or U8576 (N_8576,N_2435,N_1828);
nand U8577 (N_8577,N_2341,N_2432);
nor U8578 (N_8578,N_4370,N_1493);
and U8579 (N_8579,N_1116,N_2902);
and U8580 (N_8580,N_5621,N_1853);
nand U8581 (N_8581,N_3595,N_203);
nor U8582 (N_8582,N_5029,N_4978);
and U8583 (N_8583,N_1621,N_557);
xnor U8584 (N_8584,N_1888,N_3935);
or U8585 (N_8585,N_4606,N_1735);
and U8586 (N_8586,N_85,N_3279);
nand U8587 (N_8587,N_1470,N_2259);
xor U8588 (N_8588,N_3853,N_5756);
xor U8589 (N_8589,N_1900,N_2527);
nand U8590 (N_8590,N_4010,N_977);
xnor U8591 (N_8591,N_5482,N_909);
and U8592 (N_8592,N_1764,N_3732);
nand U8593 (N_8593,N_4314,N_1749);
or U8594 (N_8594,N_2594,N_123);
xnor U8595 (N_8595,N_1464,N_2788);
or U8596 (N_8596,N_518,N_4679);
nor U8597 (N_8597,N_16,N_4930);
and U8598 (N_8598,N_3048,N_1803);
xnor U8599 (N_8599,N_97,N_2536);
nand U8600 (N_8600,N_2253,N_862);
xor U8601 (N_8601,N_5813,N_666);
and U8602 (N_8602,N_4227,N_5741);
nand U8603 (N_8603,N_4100,N_196);
nand U8604 (N_8604,N_3396,N_3591);
xnor U8605 (N_8605,N_5249,N_4131);
nand U8606 (N_8606,N_5848,N_1291);
and U8607 (N_8607,N_606,N_821);
nand U8608 (N_8608,N_3482,N_5894);
nand U8609 (N_8609,N_3342,N_4065);
xor U8610 (N_8610,N_3820,N_4662);
nand U8611 (N_8611,N_5077,N_274);
and U8612 (N_8612,N_3897,N_975);
nor U8613 (N_8613,N_3336,N_5732);
and U8614 (N_8614,N_3213,N_5352);
nand U8615 (N_8615,N_2910,N_2165);
and U8616 (N_8616,N_1763,N_4622);
xor U8617 (N_8617,N_5260,N_3782);
nand U8618 (N_8618,N_1715,N_895);
xnor U8619 (N_8619,N_2124,N_1362);
nor U8620 (N_8620,N_139,N_4163);
nand U8621 (N_8621,N_1066,N_3070);
xnor U8622 (N_8622,N_4648,N_5085);
nand U8623 (N_8623,N_1418,N_1390);
or U8624 (N_8624,N_2830,N_1843);
nor U8625 (N_8625,N_5401,N_2303);
xnor U8626 (N_8626,N_3407,N_4737);
and U8627 (N_8627,N_1837,N_5955);
xnor U8628 (N_8628,N_3939,N_4789);
and U8629 (N_8629,N_3810,N_5175);
nand U8630 (N_8630,N_5933,N_4070);
xor U8631 (N_8631,N_1542,N_3152);
and U8632 (N_8632,N_405,N_5396);
nor U8633 (N_8633,N_3539,N_2599);
and U8634 (N_8634,N_4730,N_5855);
nor U8635 (N_8635,N_220,N_302);
nor U8636 (N_8636,N_3416,N_3199);
xor U8637 (N_8637,N_5590,N_5607);
xor U8638 (N_8638,N_5018,N_3118);
nor U8639 (N_8639,N_1699,N_341);
nor U8640 (N_8640,N_5920,N_1564);
nor U8641 (N_8641,N_3564,N_1133);
and U8642 (N_8642,N_4364,N_3249);
or U8643 (N_8643,N_24,N_4879);
or U8644 (N_8644,N_5512,N_5923);
nor U8645 (N_8645,N_2122,N_423);
and U8646 (N_8646,N_4791,N_1061);
nor U8647 (N_8647,N_863,N_4705);
nor U8648 (N_8648,N_5940,N_1956);
or U8649 (N_8649,N_1830,N_5690);
nor U8650 (N_8650,N_5355,N_956);
nor U8651 (N_8651,N_253,N_5992);
and U8652 (N_8652,N_3548,N_876);
nor U8653 (N_8653,N_2858,N_500);
nand U8654 (N_8654,N_2023,N_4061);
nor U8655 (N_8655,N_4169,N_1397);
nor U8656 (N_8656,N_165,N_410);
nor U8657 (N_8657,N_3360,N_4262);
xnor U8658 (N_8658,N_4575,N_1284);
nor U8659 (N_8659,N_5946,N_199);
xor U8660 (N_8660,N_1098,N_3918);
or U8661 (N_8661,N_5063,N_533);
nor U8662 (N_8662,N_2557,N_4871);
nand U8663 (N_8663,N_901,N_426);
and U8664 (N_8664,N_1693,N_806);
xnor U8665 (N_8665,N_4969,N_903);
and U8666 (N_8666,N_4520,N_2606);
nor U8667 (N_8667,N_3292,N_2279);
and U8668 (N_8668,N_1919,N_4840);
xor U8669 (N_8669,N_5030,N_5598);
and U8670 (N_8670,N_3497,N_2539);
nand U8671 (N_8671,N_5833,N_2553);
or U8672 (N_8672,N_3466,N_5530);
xor U8673 (N_8673,N_2003,N_2633);
nand U8674 (N_8674,N_2457,N_4143);
and U8675 (N_8675,N_4139,N_1756);
nor U8676 (N_8676,N_3104,N_435);
and U8677 (N_8677,N_2015,N_2692);
or U8678 (N_8678,N_2655,N_3932);
xor U8679 (N_8679,N_4203,N_3239);
nor U8680 (N_8680,N_147,N_3791);
nor U8681 (N_8681,N_924,N_2150);
nor U8682 (N_8682,N_2065,N_1349);
and U8683 (N_8683,N_4093,N_4842);
nand U8684 (N_8684,N_2013,N_2497);
nand U8685 (N_8685,N_2540,N_5682);
and U8686 (N_8686,N_2754,N_5738);
xnor U8687 (N_8687,N_2739,N_3600);
nor U8688 (N_8688,N_4000,N_4542);
nor U8689 (N_8689,N_2824,N_829);
xnor U8690 (N_8690,N_1583,N_4735);
nand U8691 (N_8691,N_3885,N_735);
nor U8692 (N_8692,N_3008,N_83);
nor U8693 (N_8693,N_2433,N_5698);
nor U8694 (N_8694,N_1960,N_2048);
nor U8695 (N_8695,N_242,N_2905);
nand U8696 (N_8696,N_3258,N_1021);
nor U8697 (N_8697,N_499,N_2698);
xor U8698 (N_8698,N_5938,N_4404);
and U8699 (N_8699,N_4172,N_4646);
and U8700 (N_8700,N_5635,N_1019);
nand U8701 (N_8701,N_2233,N_4217);
and U8702 (N_8702,N_2353,N_2658);
nand U8703 (N_8703,N_793,N_129);
and U8704 (N_8704,N_2152,N_128);
or U8705 (N_8705,N_2272,N_1497);
xnor U8706 (N_8706,N_4865,N_1798);
xnor U8707 (N_8707,N_2249,N_1032);
xor U8708 (N_8708,N_72,N_3842);
nand U8709 (N_8709,N_1554,N_344);
nand U8710 (N_8710,N_2125,N_3940);
nand U8711 (N_8711,N_343,N_2584);
nand U8712 (N_8712,N_998,N_392);
nand U8713 (N_8713,N_5872,N_1978);
nand U8714 (N_8714,N_5034,N_3078);
and U8715 (N_8715,N_3877,N_4126);
nor U8716 (N_8716,N_2387,N_2728);
and U8717 (N_8717,N_4577,N_4926);
and U8718 (N_8718,N_4751,N_441);
nand U8719 (N_8719,N_378,N_5269);
nand U8720 (N_8720,N_470,N_5187);
xor U8721 (N_8721,N_3310,N_3823);
nor U8722 (N_8722,N_2566,N_2966);
and U8723 (N_8723,N_1794,N_4773);
nor U8724 (N_8724,N_36,N_978);
nor U8725 (N_8725,N_1430,N_4324);
xnor U8726 (N_8726,N_1534,N_4360);
and U8727 (N_8727,N_1765,N_5125);
nor U8728 (N_8728,N_2620,N_2860);
and U8729 (N_8729,N_152,N_3386);
xnor U8730 (N_8730,N_4795,N_4676);
nand U8731 (N_8731,N_5733,N_5457);
or U8732 (N_8732,N_1813,N_4186);
and U8733 (N_8733,N_1182,N_1485);
xor U8734 (N_8734,N_5192,N_4915);
nand U8735 (N_8735,N_2005,N_132);
nand U8736 (N_8736,N_2039,N_2051);
xor U8737 (N_8737,N_3079,N_4685);
nor U8738 (N_8738,N_1028,N_766);
xor U8739 (N_8739,N_4759,N_2465);
nor U8740 (N_8740,N_1278,N_158);
and U8741 (N_8741,N_2325,N_1899);
xor U8742 (N_8742,N_1467,N_629);
xnor U8743 (N_8743,N_1285,N_2074);
and U8744 (N_8744,N_366,N_5251);
or U8745 (N_8745,N_5987,N_3561);
nor U8746 (N_8746,N_1795,N_3481);
xor U8747 (N_8747,N_3833,N_4033);
nand U8748 (N_8748,N_2238,N_3663);
nand U8749 (N_8749,N_2543,N_4596);
or U8750 (N_8750,N_3185,N_5400);
xor U8751 (N_8751,N_3961,N_5343);
nor U8752 (N_8752,N_5557,N_3884);
nor U8753 (N_8753,N_2875,N_1959);
and U8754 (N_8754,N_1451,N_3575);
or U8755 (N_8755,N_707,N_1347);
xor U8756 (N_8756,N_790,N_3263);
nand U8757 (N_8757,N_376,N_3036);
nand U8758 (N_8758,N_169,N_144);
nand U8759 (N_8759,N_463,N_4063);
and U8760 (N_8760,N_2695,N_3252);
nor U8761 (N_8761,N_385,N_3393);
or U8762 (N_8762,N_3298,N_3134);
nand U8763 (N_8763,N_5867,N_516);
nor U8764 (N_8764,N_2825,N_1350);
xor U8765 (N_8765,N_5254,N_3119);
xor U8766 (N_8766,N_3385,N_3007);
xor U8767 (N_8767,N_758,N_3130);
or U8768 (N_8768,N_511,N_4890);
or U8769 (N_8769,N_4461,N_3069);
xor U8770 (N_8770,N_3116,N_835);
and U8771 (N_8771,N_847,N_1422);
or U8772 (N_8772,N_5697,N_1937);
nor U8773 (N_8773,N_4571,N_1654);
and U8774 (N_8774,N_897,N_1528);
xor U8775 (N_8775,N_1026,N_5358);
and U8776 (N_8776,N_482,N_2053);
nor U8777 (N_8777,N_3605,N_4687);
and U8778 (N_8778,N_5143,N_2210);
and U8779 (N_8779,N_5714,N_4962);
or U8780 (N_8780,N_592,N_3673);
nor U8781 (N_8781,N_3565,N_5365);
nor U8782 (N_8782,N_3526,N_221);
and U8783 (N_8783,N_2142,N_1502);
nor U8784 (N_8784,N_4124,N_5703);
and U8785 (N_8785,N_692,N_5444);
and U8786 (N_8786,N_4291,N_4938);
or U8787 (N_8787,N_5734,N_5825);
nand U8788 (N_8788,N_5011,N_5846);
xor U8789 (N_8789,N_5268,N_1416);
nor U8790 (N_8790,N_4424,N_3692);
or U8791 (N_8791,N_4863,N_3149);
nor U8792 (N_8792,N_2285,N_5986);
nand U8793 (N_8793,N_3986,N_5493);
nand U8794 (N_8794,N_417,N_1074);
or U8795 (N_8795,N_5780,N_2001);
xnor U8796 (N_8796,N_5363,N_4495);
and U8797 (N_8797,N_2268,N_1153);
nor U8798 (N_8798,N_3267,N_3418);
nor U8799 (N_8799,N_1402,N_4948);
or U8800 (N_8800,N_3533,N_5448);
or U8801 (N_8801,N_722,N_4849);
or U8802 (N_8802,N_2828,N_1668);
nor U8803 (N_8803,N_815,N_38);
and U8804 (N_8804,N_365,N_1214);
xnor U8805 (N_8805,N_4015,N_2491);
or U8806 (N_8806,N_2510,N_2367);
nor U8807 (N_8807,N_2270,N_2153);
nor U8808 (N_8808,N_4729,N_4433);
nand U8809 (N_8809,N_929,N_4078);
and U8810 (N_8810,N_4244,N_3021);
xor U8811 (N_8811,N_2616,N_44);
nor U8812 (N_8812,N_2561,N_1510);
and U8813 (N_8813,N_2148,N_2985);
xor U8814 (N_8814,N_5348,N_5259);
and U8815 (N_8815,N_1523,N_2203);
nor U8816 (N_8816,N_5161,N_3080);
or U8817 (N_8817,N_5958,N_2102);
xnor U8818 (N_8818,N_1450,N_2138);
nor U8819 (N_8819,N_5582,N_3874);
nor U8820 (N_8820,N_3966,N_4468);
and U8821 (N_8821,N_3714,N_3882);
nor U8822 (N_8822,N_4841,N_468);
nor U8823 (N_8823,N_8,N_2324);
nor U8824 (N_8824,N_5168,N_1819);
xor U8825 (N_8825,N_4077,N_2687);
and U8826 (N_8826,N_3655,N_5828);
nor U8827 (N_8827,N_2948,N_1754);
nand U8828 (N_8828,N_548,N_4383);
and U8829 (N_8829,N_2276,N_795);
nor U8830 (N_8830,N_3795,N_65);
and U8831 (N_8831,N_3861,N_4589);
nor U8832 (N_8832,N_1077,N_2329);
xnor U8833 (N_8833,N_4007,N_1135);
and U8834 (N_8834,N_5280,N_613);
nor U8835 (N_8835,N_1445,N_215);
and U8836 (N_8836,N_1867,N_2999);
nor U8837 (N_8837,N_1199,N_4412);
nand U8838 (N_8838,N_2685,N_5253);
xor U8839 (N_8839,N_2856,N_2091);
and U8840 (N_8840,N_1302,N_2230);
nand U8841 (N_8841,N_2480,N_5230);
nand U8842 (N_8842,N_1909,N_213);
nor U8843 (N_8843,N_5150,N_5843);
nor U8844 (N_8844,N_3089,N_3624);
nand U8845 (N_8845,N_3946,N_5159);
and U8846 (N_8846,N_4530,N_3027);
nor U8847 (N_8847,N_3474,N_3616);
or U8848 (N_8848,N_5053,N_1948);
nor U8849 (N_8849,N_2261,N_5216);
xor U8850 (N_8850,N_2652,N_2751);
nand U8851 (N_8851,N_1055,N_4874);
nor U8852 (N_8852,N_5983,N_2706);
and U8853 (N_8853,N_5816,N_3234);
nand U8854 (N_8854,N_1598,N_1685);
nand U8855 (N_8855,N_3437,N_601);
nor U8856 (N_8856,N_813,N_4816);
xnor U8857 (N_8857,N_1921,N_1605);
or U8858 (N_8858,N_1131,N_5474);
nor U8859 (N_8859,N_379,N_4518);
nand U8860 (N_8860,N_2598,N_1945);
nor U8861 (N_8861,N_3022,N_2642);
or U8862 (N_8862,N_4182,N_2621);
or U8863 (N_8863,N_1351,N_5595);
or U8864 (N_8864,N_3619,N_2328);
xor U8865 (N_8865,N_2477,N_1516);
and U8866 (N_8866,N_4935,N_2154);
nand U8867 (N_8867,N_1073,N_3908);
nor U8868 (N_8868,N_3852,N_1343);
and U8869 (N_8869,N_503,N_5025);
nor U8870 (N_8870,N_234,N_279);
or U8871 (N_8871,N_28,N_4981);
nor U8872 (N_8872,N_5337,N_3009);
nor U8873 (N_8873,N_4576,N_2078);
or U8874 (N_8874,N_4594,N_100);
and U8875 (N_8875,N_2194,N_1514);
xnor U8876 (N_8876,N_3204,N_3376);
nand U8877 (N_8877,N_4298,N_529);
nor U8878 (N_8878,N_5506,N_2079);
nand U8879 (N_8879,N_4340,N_3706);
xnor U8880 (N_8880,N_1404,N_4091);
nor U8881 (N_8881,N_840,N_4933);
xnor U8882 (N_8882,N_3713,N_1633);
nand U8883 (N_8883,N_5158,N_5250);
and U8884 (N_8884,N_5667,N_3454);
nor U8885 (N_8885,N_5279,N_4486);
nor U8886 (N_8886,N_4508,N_3973);
nand U8887 (N_8887,N_3468,N_3883);
nor U8888 (N_8888,N_4906,N_907);
nor U8889 (N_8889,N_2185,N_5623);
xor U8890 (N_8890,N_3632,N_4811);
or U8891 (N_8891,N_5026,N_4473);
nand U8892 (N_8892,N_3520,N_4138);
and U8893 (N_8893,N_5430,N_1759);
and U8894 (N_8894,N_5087,N_4746);
or U8895 (N_8895,N_849,N_5614);
nor U8896 (N_8896,N_4621,N_5390);
nand U8897 (N_8897,N_4173,N_3804);
nor U8898 (N_8898,N_3050,N_2776);
or U8899 (N_8899,N_1249,N_5465);
nor U8900 (N_8900,N_507,N_4519);
nor U8901 (N_8901,N_5397,N_2961);
nor U8902 (N_8902,N_5711,N_1484);
or U8903 (N_8903,N_4194,N_5569);
and U8904 (N_8904,N_5110,N_4159);
or U8905 (N_8905,N_1475,N_2711);
xor U8906 (N_8906,N_2054,N_3923);
xor U8907 (N_8907,N_4375,N_1298);
and U8908 (N_8908,N_2114,N_1208);
or U8909 (N_8909,N_5220,N_5231);
and U8910 (N_8910,N_2266,N_1400);
nor U8911 (N_8911,N_1783,N_5622);
xor U8912 (N_8912,N_1064,N_1637);
and U8913 (N_8913,N_5418,N_5413);
nand U8914 (N_8914,N_3186,N_1744);
xnor U8915 (N_8915,N_1195,N_2868);
or U8916 (N_8916,N_1496,N_1020);
nor U8917 (N_8917,N_2781,N_2722);
or U8918 (N_8918,N_3111,N_4888);
or U8919 (N_8919,N_1176,N_1174);
or U8920 (N_8920,N_1292,N_4234);
nand U8921 (N_8921,N_710,N_202);
xnor U8922 (N_8922,N_2508,N_3099);
and U8923 (N_8923,N_5922,N_5099);
nor U8924 (N_8924,N_2925,N_755);
or U8925 (N_8925,N_743,N_374);
or U8926 (N_8926,N_4339,N_1013);
nand U8927 (N_8927,N_2953,N_1491);
and U8928 (N_8928,N_5942,N_2789);
and U8929 (N_8929,N_5762,N_645);
and U8930 (N_8930,N_1157,N_1797);
xnor U8931 (N_8931,N_1189,N_4031);
nand U8932 (N_8932,N_27,N_1686);
or U8933 (N_8933,N_5852,N_4214);
nor U8934 (N_8934,N_4916,N_2016);
or U8935 (N_8935,N_4734,N_1002);
nor U8936 (N_8936,N_4665,N_4395);
and U8937 (N_8937,N_2682,N_394);
or U8938 (N_8938,N_3837,N_3879);
and U8939 (N_8939,N_3538,N_3493);
nor U8940 (N_8940,N_4854,N_502);
nand U8941 (N_8941,N_1673,N_170);
xnor U8942 (N_8942,N_5755,N_2242);
nor U8943 (N_8943,N_3830,N_4607);
or U8944 (N_8944,N_1865,N_655);
nor U8945 (N_8945,N_3405,N_437);
or U8946 (N_8946,N_1202,N_3829);
xnor U8947 (N_8947,N_162,N_4566);
or U8948 (N_8948,N_3579,N_4309);
xor U8949 (N_8949,N_1714,N_11);
nor U8950 (N_8950,N_3015,N_282);
xnor U8951 (N_8951,N_3103,N_742);
nand U8952 (N_8952,N_206,N_3060);
xor U8953 (N_8953,N_3300,N_401);
nand U8954 (N_8954,N_5899,N_3040);
xnor U8955 (N_8955,N_1051,N_4226);
or U8956 (N_8956,N_4343,N_1265);
nor U8957 (N_8957,N_572,N_4180);
nand U8958 (N_8958,N_1207,N_5245);
nand U8959 (N_8959,N_47,N_4135);
or U8960 (N_8960,N_4414,N_2819);
and U8961 (N_8961,N_791,N_4004);
xnor U8962 (N_8962,N_2834,N_5995);
nor U8963 (N_8963,N_3954,N_2025);
nor U8964 (N_8964,N_4893,N_1890);
nor U8965 (N_8965,N_2895,N_2879);
nor U8966 (N_8966,N_3498,N_525);
or U8967 (N_8967,N_4689,N_2294);
and U8968 (N_8968,N_5554,N_2161);
and U8969 (N_8969,N_4083,N_3931);
or U8970 (N_8970,N_2679,N_3127);
or U8971 (N_8971,N_4134,N_2911);
nor U8972 (N_8972,N_4973,N_4332);
xnor U8973 (N_8973,N_5044,N_2501);
nor U8974 (N_8974,N_3780,N_2512);
nand U8975 (N_8975,N_5325,N_1725);
and U8976 (N_8976,N_2481,N_4802);
nor U8977 (N_8977,N_5793,N_3781);
nand U8978 (N_8978,N_1238,N_1353);
nand U8979 (N_8979,N_3531,N_3652);
nand U8980 (N_8980,N_5327,N_5404);
xor U8981 (N_8981,N_1012,N_988);
and U8982 (N_8982,N_1490,N_2021);
nand U8983 (N_8983,N_5039,N_4336);
nor U8984 (N_8984,N_5881,N_3534);
or U8985 (N_8985,N_2322,N_3403);
xor U8986 (N_8986,N_2511,N_2248);
or U8987 (N_8987,N_5019,N_2593);
nand U8988 (N_8988,N_3686,N_4398);
and U8989 (N_8989,N_5106,N_3312);
xnor U8990 (N_8990,N_3296,N_574);
nor U8991 (N_8991,N_3779,N_1792);
and U8992 (N_8992,N_670,N_2383);
nor U8993 (N_8993,N_1438,N_5764);
or U8994 (N_8994,N_3745,N_1492);
nand U8995 (N_8995,N_4215,N_4512);
and U8996 (N_8996,N_5445,N_5402);
and U8997 (N_8997,N_264,N_4259);
or U8998 (N_8998,N_2394,N_1861);
xor U8999 (N_8999,N_4022,N_3426);
or U9000 (N_9000,N_3860,N_3044);
xnor U9001 (N_9001,N_1928,N_328);
nor U9002 (N_9002,N_2080,N_948);
xnor U9003 (N_9003,N_4310,N_5876);
xor U9004 (N_9004,N_16,N_5320);
nor U9005 (N_9005,N_681,N_740);
xnor U9006 (N_9006,N_5140,N_5445);
nand U9007 (N_9007,N_5339,N_5519);
nand U9008 (N_9008,N_4320,N_1164);
and U9009 (N_9009,N_2518,N_210);
xor U9010 (N_9010,N_205,N_2466);
nand U9011 (N_9011,N_5730,N_5844);
nand U9012 (N_9012,N_1380,N_5974);
nand U9013 (N_9013,N_3672,N_1848);
or U9014 (N_9014,N_3547,N_925);
xor U9015 (N_9015,N_1622,N_3484);
nor U9016 (N_9016,N_851,N_659);
or U9017 (N_9017,N_1787,N_882);
nor U9018 (N_9018,N_2614,N_616);
and U9019 (N_9019,N_5129,N_872);
nor U9020 (N_9020,N_2283,N_5989);
or U9021 (N_9021,N_4196,N_853);
nand U9022 (N_9022,N_4623,N_4492);
xor U9023 (N_9023,N_4019,N_802);
nand U9024 (N_9024,N_3996,N_2230);
xor U9025 (N_9025,N_4366,N_853);
or U9026 (N_9026,N_341,N_4299);
nor U9027 (N_9027,N_4216,N_1562);
and U9028 (N_9028,N_2331,N_936);
or U9029 (N_9029,N_3900,N_1361);
nand U9030 (N_9030,N_5960,N_3961);
nor U9031 (N_9031,N_875,N_118);
nor U9032 (N_9032,N_1392,N_2726);
and U9033 (N_9033,N_5421,N_4315);
xnor U9034 (N_9034,N_1388,N_3148);
or U9035 (N_9035,N_3156,N_3091);
or U9036 (N_9036,N_3986,N_5469);
or U9037 (N_9037,N_2961,N_5428);
nand U9038 (N_9038,N_2510,N_562);
nor U9039 (N_9039,N_3406,N_4785);
nor U9040 (N_9040,N_2935,N_3761);
or U9041 (N_9041,N_1971,N_1551);
and U9042 (N_9042,N_707,N_4999);
or U9043 (N_9043,N_4993,N_5891);
nand U9044 (N_9044,N_5029,N_2638);
nor U9045 (N_9045,N_3038,N_335);
nand U9046 (N_9046,N_4632,N_5314);
and U9047 (N_9047,N_779,N_1454);
or U9048 (N_9048,N_2906,N_2118);
or U9049 (N_9049,N_5100,N_1316);
nor U9050 (N_9050,N_5897,N_2768);
nand U9051 (N_9051,N_4436,N_4245);
nor U9052 (N_9052,N_681,N_116);
xnor U9053 (N_9053,N_1920,N_3985);
nor U9054 (N_9054,N_4129,N_4932);
xor U9055 (N_9055,N_1668,N_692);
and U9056 (N_9056,N_998,N_3147);
or U9057 (N_9057,N_4924,N_4590);
and U9058 (N_9058,N_1031,N_793);
or U9059 (N_9059,N_1458,N_444);
nor U9060 (N_9060,N_4611,N_2916);
nor U9061 (N_9061,N_4804,N_2274);
nand U9062 (N_9062,N_2354,N_930);
nand U9063 (N_9063,N_1172,N_258);
nor U9064 (N_9064,N_3438,N_4058);
or U9065 (N_9065,N_569,N_1729);
or U9066 (N_9066,N_3045,N_2392);
and U9067 (N_9067,N_5563,N_706);
nand U9068 (N_9068,N_2355,N_2939);
nand U9069 (N_9069,N_3166,N_350);
or U9070 (N_9070,N_2772,N_1044);
nor U9071 (N_9071,N_3579,N_1731);
nand U9072 (N_9072,N_267,N_4962);
xor U9073 (N_9073,N_139,N_2711);
nand U9074 (N_9074,N_3060,N_1322);
or U9075 (N_9075,N_3320,N_5945);
or U9076 (N_9076,N_1724,N_3934);
nor U9077 (N_9077,N_2444,N_5771);
or U9078 (N_9078,N_243,N_4015);
xor U9079 (N_9079,N_3981,N_2491);
or U9080 (N_9080,N_3764,N_138);
or U9081 (N_9081,N_2555,N_5706);
or U9082 (N_9082,N_5761,N_3053);
and U9083 (N_9083,N_1760,N_1641);
or U9084 (N_9084,N_836,N_5854);
nand U9085 (N_9085,N_2545,N_4492);
nor U9086 (N_9086,N_5385,N_2337);
xnor U9087 (N_9087,N_1183,N_2984);
nand U9088 (N_9088,N_2404,N_3071);
xor U9089 (N_9089,N_3014,N_3033);
nor U9090 (N_9090,N_381,N_2976);
nor U9091 (N_9091,N_550,N_5384);
nor U9092 (N_9092,N_3756,N_2651);
or U9093 (N_9093,N_2285,N_1241);
xor U9094 (N_9094,N_2261,N_1624);
nand U9095 (N_9095,N_586,N_1654);
nand U9096 (N_9096,N_4722,N_3001);
or U9097 (N_9097,N_5425,N_5868);
nand U9098 (N_9098,N_4928,N_3399);
nand U9099 (N_9099,N_4059,N_5962);
xnor U9100 (N_9100,N_3812,N_2970);
or U9101 (N_9101,N_4718,N_5104);
nand U9102 (N_9102,N_675,N_716);
and U9103 (N_9103,N_793,N_15);
xor U9104 (N_9104,N_3944,N_194);
and U9105 (N_9105,N_3989,N_5378);
xor U9106 (N_9106,N_2984,N_1451);
nand U9107 (N_9107,N_2618,N_1627);
xor U9108 (N_9108,N_3251,N_4493);
nor U9109 (N_9109,N_2986,N_5927);
nor U9110 (N_9110,N_4260,N_2189);
nand U9111 (N_9111,N_5797,N_4771);
nand U9112 (N_9112,N_579,N_1985);
nor U9113 (N_9113,N_4413,N_5719);
and U9114 (N_9114,N_5051,N_292);
xor U9115 (N_9115,N_1887,N_5708);
xor U9116 (N_9116,N_814,N_2127);
nor U9117 (N_9117,N_936,N_3085);
or U9118 (N_9118,N_963,N_764);
nand U9119 (N_9119,N_1564,N_706);
nor U9120 (N_9120,N_4467,N_3918);
and U9121 (N_9121,N_1855,N_4588);
nor U9122 (N_9122,N_4505,N_2512);
xor U9123 (N_9123,N_2795,N_1650);
nand U9124 (N_9124,N_3710,N_1850);
nand U9125 (N_9125,N_2279,N_5857);
xor U9126 (N_9126,N_4423,N_3560);
xnor U9127 (N_9127,N_112,N_1254);
and U9128 (N_9128,N_4132,N_690);
or U9129 (N_9129,N_912,N_1944);
and U9130 (N_9130,N_130,N_4977);
or U9131 (N_9131,N_4767,N_4120);
nand U9132 (N_9132,N_5164,N_5473);
nand U9133 (N_9133,N_4033,N_2193);
xnor U9134 (N_9134,N_5328,N_1695);
and U9135 (N_9135,N_109,N_51);
or U9136 (N_9136,N_1301,N_3022);
xnor U9137 (N_9137,N_4360,N_5366);
and U9138 (N_9138,N_5570,N_5785);
nor U9139 (N_9139,N_2670,N_2904);
or U9140 (N_9140,N_3189,N_716);
or U9141 (N_9141,N_523,N_5477);
and U9142 (N_9142,N_390,N_239);
xor U9143 (N_9143,N_1433,N_1372);
xor U9144 (N_9144,N_2020,N_5679);
xnor U9145 (N_9145,N_2611,N_4590);
nand U9146 (N_9146,N_5174,N_4142);
or U9147 (N_9147,N_2561,N_1177);
and U9148 (N_9148,N_4466,N_1353);
nor U9149 (N_9149,N_2380,N_2427);
xnor U9150 (N_9150,N_2895,N_285);
nor U9151 (N_9151,N_998,N_1682);
nor U9152 (N_9152,N_5659,N_2981);
nand U9153 (N_9153,N_5351,N_1732);
nand U9154 (N_9154,N_2798,N_3085);
or U9155 (N_9155,N_338,N_4947);
nand U9156 (N_9156,N_2984,N_204);
nor U9157 (N_9157,N_3604,N_3474);
xnor U9158 (N_9158,N_4084,N_4031);
or U9159 (N_9159,N_7,N_870);
nor U9160 (N_9160,N_3857,N_4634);
nor U9161 (N_9161,N_4894,N_3397);
or U9162 (N_9162,N_585,N_442);
nor U9163 (N_9163,N_4707,N_2536);
or U9164 (N_9164,N_4919,N_41);
or U9165 (N_9165,N_655,N_3077);
or U9166 (N_9166,N_1273,N_203);
and U9167 (N_9167,N_3663,N_384);
and U9168 (N_9168,N_4749,N_5274);
xor U9169 (N_9169,N_455,N_2262);
nor U9170 (N_9170,N_3035,N_3990);
and U9171 (N_9171,N_2759,N_2764);
or U9172 (N_9172,N_1831,N_1403);
and U9173 (N_9173,N_4915,N_3545);
or U9174 (N_9174,N_2444,N_1405);
xor U9175 (N_9175,N_2230,N_5794);
nor U9176 (N_9176,N_4502,N_3492);
and U9177 (N_9177,N_5329,N_3829);
nor U9178 (N_9178,N_4644,N_5170);
or U9179 (N_9179,N_491,N_765);
and U9180 (N_9180,N_4681,N_4229);
nand U9181 (N_9181,N_5368,N_3387);
nor U9182 (N_9182,N_4775,N_352);
or U9183 (N_9183,N_4019,N_874);
nor U9184 (N_9184,N_4222,N_3372);
nor U9185 (N_9185,N_4732,N_409);
and U9186 (N_9186,N_734,N_963);
nor U9187 (N_9187,N_1751,N_5788);
nand U9188 (N_9188,N_5648,N_3595);
nand U9189 (N_9189,N_5947,N_4305);
xor U9190 (N_9190,N_2578,N_1727);
nand U9191 (N_9191,N_2957,N_1676);
nor U9192 (N_9192,N_3203,N_1118);
nor U9193 (N_9193,N_5440,N_1347);
nor U9194 (N_9194,N_1276,N_4082);
nor U9195 (N_9195,N_2219,N_2121);
and U9196 (N_9196,N_39,N_4553);
nand U9197 (N_9197,N_5419,N_2178);
or U9198 (N_9198,N_4021,N_4265);
or U9199 (N_9199,N_4573,N_5849);
nand U9200 (N_9200,N_594,N_1743);
or U9201 (N_9201,N_5810,N_5385);
nor U9202 (N_9202,N_4224,N_114);
or U9203 (N_9203,N_5348,N_2108);
xnor U9204 (N_9204,N_213,N_1188);
or U9205 (N_9205,N_2714,N_2507);
nor U9206 (N_9206,N_3161,N_3466);
and U9207 (N_9207,N_5514,N_5366);
xnor U9208 (N_9208,N_1459,N_399);
or U9209 (N_9209,N_4398,N_4489);
xnor U9210 (N_9210,N_3137,N_408);
or U9211 (N_9211,N_1150,N_5477);
nand U9212 (N_9212,N_3122,N_5684);
nand U9213 (N_9213,N_3336,N_1227);
xnor U9214 (N_9214,N_2375,N_1645);
and U9215 (N_9215,N_5898,N_4647);
or U9216 (N_9216,N_3950,N_2190);
and U9217 (N_9217,N_5102,N_5204);
xnor U9218 (N_9218,N_4715,N_3883);
xor U9219 (N_9219,N_222,N_3590);
nor U9220 (N_9220,N_3910,N_3792);
xor U9221 (N_9221,N_4862,N_2771);
xnor U9222 (N_9222,N_1468,N_2352);
or U9223 (N_9223,N_384,N_3986);
nor U9224 (N_9224,N_2771,N_5339);
nand U9225 (N_9225,N_5771,N_2814);
nor U9226 (N_9226,N_584,N_3432);
xor U9227 (N_9227,N_2046,N_4432);
and U9228 (N_9228,N_5882,N_1910);
or U9229 (N_9229,N_4550,N_4021);
nor U9230 (N_9230,N_3663,N_4794);
nor U9231 (N_9231,N_3004,N_5202);
xor U9232 (N_9232,N_3810,N_1742);
xnor U9233 (N_9233,N_158,N_840);
and U9234 (N_9234,N_3431,N_5814);
and U9235 (N_9235,N_5702,N_5069);
and U9236 (N_9236,N_2951,N_2763);
nor U9237 (N_9237,N_644,N_1568);
nor U9238 (N_9238,N_891,N_3322);
nand U9239 (N_9239,N_2825,N_4041);
and U9240 (N_9240,N_730,N_4271);
xor U9241 (N_9241,N_1361,N_5115);
xnor U9242 (N_9242,N_3632,N_756);
nor U9243 (N_9243,N_3300,N_4280);
and U9244 (N_9244,N_5479,N_3505);
and U9245 (N_9245,N_455,N_1378);
and U9246 (N_9246,N_3516,N_4639);
xor U9247 (N_9247,N_1597,N_2935);
xnor U9248 (N_9248,N_3873,N_2842);
and U9249 (N_9249,N_1253,N_711);
xor U9250 (N_9250,N_5690,N_1538);
nand U9251 (N_9251,N_844,N_3803);
nand U9252 (N_9252,N_4485,N_115);
nand U9253 (N_9253,N_5103,N_5241);
and U9254 (N_9254,N_2088,N_3543);
xor U9255 (N_9255,N_5755,N_3890);
nand U9256 (N_9256,N_1374,N_3801);
or U9257 (N_9257,N_5768,N_4348);
nand U9258 (N_9258,N_4980,N_4078);
nor U9259 (N_9259,N_4486,N_2188);
and U9260 (N_9260,N_1484,N_1233);
or U9261 (N_9261,N_3625,N_4157);
nor U9262 (N_9262,N_3029,N_463);
nand U9263 (N_9263,N_5879,N_2967);
or U9264 (N_9264,N_5539,N_225);
or U9265 (N_9265,N_2933,N_1750);
and U9266 (N_9266,N_5756,N_3309);
xor U9267 (N_9267,N_3972,N_2783);
nor U9268 (N_9268,N_1473,N_2241);
nand U9269 (N_9269,N_4790,N_875);
nand U9270 (N_9270,N_3299,N_5738);
or U9271 (N_9271,N_293,N_5952);
and U9272 (N_9272,N_2586,N_1940);
nand U9273 (N_9273,N_5965,N_5249);
and U9274 (N_9274,N_316,N_605);
and U9275 (N_9275,N_1904,N_870);
or U9276 (N_9276,N_4398,N_1469);
nor U9277 (N_9277,N_968,N_4710);
xor U9278 (N_9278,N_5720,N_1341);
and U9279 (N_9279,N_1792,N_4022);
or U9280 (N_9280,N_5308,N_1071);
and U9281 (N_9281,N_1795,N_1788);
xnor U9282 (N_9282,N_4892,N_3394);
nand U9283 (N_9283,N_1912,N_4277);
or U9284 (N_9284,N_2842,N_3335);
and U9285 (N_9285,N_1714,N_1943);
and U9286 (N_9286,N_1952,N_206);
and U9287 (N_9287,N_4398,N_5912);
and U9288 (N_9288,N_5153,N_1940);
or U9289 (N_9289,N_2765,N_5262);
or U9290 (N_9290,N_3240,N_606);
or U9291 (N_9291,N_1936,N_2463);
nand U9292 (N_9292,N_2278,N_4833);
nor U9293 (N_9293,N_371,N_299);
nor U9294 (N_9294,N_4699,N_1271);
nor U9295 (N_9295,N_4134,N_4092);
xnor U9296 (N_9296,N_2283,N_5528);
and U9297 (N_9297,N_4805,N_3319);
nor U9298 (N_9298,N_4449,N_4090);
and U9299 (N_9299,N_1537,N_2675);
and U9300 (N_9300,N_5359,N_4206);
or U9301 (N_9301,N_3248,N_3969);
nand U9302 (N_9302,N_3133,N_1886);
xnor U9303 (N_9303,N_3180,N_3627);
and U9304 (N_9304,N_589,N_4053);
or U9305 (N_9305,N_4188,N_913);
and U9306 (N_9306,N_4639,N_5575);
nand U9307 (N_9307,N_4826,N_4982);
nand U9308 (N_9308,N_1804,N_1246);
nand U9309 (N_9309,N_4074,N_96);
or U9310 (N_9310,N_4795,N_4765);
nor U9311 (N_9311,N_690,N_1394);
xnor U9312 (N_9312,N_3855,N_4277);
and U9313 (N_9313,N_310,N_838);
or U9314 (N_9314,N_1160,N_1785);
and U9315 (N_9315,N_4729,N_4849);
or U9316 (N_9316,N_5467,N_2971);
nor U9317 (N_9317,N_2863,N_617);
nand U9318 (N_9318,N_1325,N_341);
or U9319 (N_9319,N_1990,N_5432);
nand U9320 (N_9320,N_5020,N_2500);
nor U9321 (N_9321,N_5235,N_5709);
xor U9322 (N_9322,N_366,N_502);
nor U9323 (N_9323,N_1420,N_170);
and U9324 (N_9324,N_596,N_5141);
nor U9325 (N_9325,N_3008,N_3843);
or U9326 (N_9326,N_5399,N_1625);
xnor U9327 (N_9327,N_4412,N_5349);
and U9328 (N_9328,N_3480,N_5063);
nand U9329 (N_9329,N_3670,N_4969);
or U9330 (N_9330,N_3204,N_123);
xor U9331 (N_9331,N_539,N_5328);
nand U9332 (N_9332,N_2990,N_5030);
and U9333 (N_9333,N_5053,N_2658);
nand U9334 (N_9334,N_2753,N_243);
nand U9335 (N_9335,N_5127,N_737);
and U9336 (N_9336,N_2812,N_3704);
nand U9337 (N_9337,N_3148,N_48);
nand U9338 (N_9338,N_2630,N_392);
or U9339 (N_9339,N_413,N_5248);
and U9340 (N_9340,N_2556,N_2428);
nor U9341 (N_9341,N_1259,N_5990);
nand U9342 (N_9342,N_2594,N_5029);
nand U9343 (N_9343,N_3992,N_3498);
nand U9344 (N_9344,N_2051,N_3992);
nor U9345 (N_9345,N_474,N_839);
or U9346 (N_9346,N_1693,N_3024);
xnor U9347 (N_9347,N_1686,N_715);
and U9348 (N_9348,N_2907,N_2458);
and U9349 (N_9349,N_1901,N_3984);
xor U9350 (N_9350,N_1934,N_1950);
xor U9351 (N_9351,N_5606,N_659);
xor U9352 (N_9352,N_3890,N_3014);
and U9353 (N_9353,N_3428,N_4288);
xor U9354 (N_9354,N_5162,N_3652);
nand U9355 (N_9355,N_5030,N_4871);
and U9356 (N_9356,N_1519,N_4731);
or U9357 (N_9357,N_3726,N_4772);
xnor U9358 (N_9358,N_2879,N_5165);
xor U9359 (N_9359,N_2871,N_4480);
nor U9360 (N_9360,N_1753,N_2629);
nor U9361 (N_9361,N_3829,N_169);
nor U9362 (N_9362,N_5432,N_5308);
nand U9363 (N_9363,N_5605,N_856);
nand U9364 (N_9364,N_1398,N_144);
nand U9365 (N_9365,N_4105,N_2210);
xnor U9366 (N_9366,N_4728,N_4485);
or U9367 (N_9367,N_5223,N_4757);
and U9368 (N_9368,N_1802,N_3998);
nor U9369 (N_9369,N_4121,N_1710);
or U9370 (N_9370,N_3223,N_542);
nand U9371 (N_9371,N_4464,N_5203);
xor U9372 (N_9372,N_2604,N_2404);
and U9373 (N_9373,N_5196,N_72);
or U9374 (N_9374,N_1971,N_2283);
nor U9375 (N_9375,N_267,N_5370);
or U9376 (N_9376,N_259,N_4745);
nor U9377 (N_9377,N_4777,N_3582);
nand U9378 (N_9378,N_4158,N_590);
nand U9379 (N_9379,N_814,N_4715);
nand U9380 (N_9380,N_5228,N_1410);
xnor U9381 (N_9381,N_3442,N_2447);
and U9382 (N_9382,N_3563,N_3805);
nand U9383 (N_9383,N_5412,N_916);
nand U9384 (N_9384,N_4976,N_4623);
nand U9385 (N_9385,N_2092,N_3669);
xor U9386 (N_9386,N_1858,N_494);
xnor U9387 (N_9387,N_200,N_932);
or U9388 (N_9388,N_3742,N_2971);
nand U9389 (N_9389,N_4105,N_2874);
and U9390 (N_9390,N_1861,N_2923);
or U9391 (N_9391,N_932,N_2058);
nand U9392 (N_9392,N_1412,N_5855);
and U9393 (N_9393,N_1289,N_5033);
xnor U9394 (N_9394,N_2363,N_1906);
xnor U9395 (N_9395,N_998,N_4027);
nand U9396 (N_9396,N_4752,N_4469);
and U9397 (N_9397,N_5319,N_4810);
nand U9398 (N_9398,N_1447,N_128);
xor U9399 (N_9399,N_1552,N_331);
and U9400 (N_9400,N_832,N_2858);
xnor U9401 (N_9401,N_719,N_2953);
or U9402 (N_9402,N_4040,N_2785);
nor U9403 (N_9403,N_3581,N_4856);
nand U9404 (N_9404,N_4861,N_2382);
xnor U9405 (N_9405,N_1349,N_2984);
and U9406 (N_9406,N_3334,N_4663);
and U9407 (N_9407,N_2389,N_1130);
and U9408 (N_9408,N_386,N_633);
and U9409 (N_9409,N_2197,N_5431);
xor U9410 (N_9410,N_1532,N_1129);
nor U9411 (N_9411,N_2769,N_1371);
or U9412 (N_9412,N_4893,N_2837);
and U9413 (N_9413,N_1770,N_3194);
nand U9414 (N_9414,N_3355,N_2585);
or U9415 (N_9415,N_3436,N_3693);
or U9416 (N_9416,N_3549,N_3539);
xnor U9417 (N_9417,N_3314,N_2492);
xor U9418 (N_9418,N_4564,N_5895);
nor U9419 (N_9419,N_5515,N_5705);
nor U9420 (N_9420,N_4231,N_4119);
nand U9421 (N_9421,N_1868,N_1235);
and U9422 (N_9422,N_5389,N_5412);
nand U9423 (N_9423,N_1329,N_5446);
and U9424 (N_9424,N_4457,N_3970);
or U9425 (N_9425,N_391,N_1509);
or U9426 (N_9426,N_674,N_5811);
or U9427 (N_9427,N_2251,N_4701);
xor U9428 (N_9428,N_2933,N_390);
xnor U9429 (N_9429,N_3552,N_1667);
and U9430 (N_9430,N_3248,N_5578);
nor U9431 (N_9431,N_3934,N_3673);
nor U9432 (N_9432,N_4922,N_232);
and U9433 (N_9433,N_5910,N_62);
and U9434 (N_9434,N_3004,N_3398);
nand U9435 (N_9435,N_1021,N_3924);
nor U9436 (N_9436,N_1584,N_250);
or U9437 (N_9437,N_347,N_1143);
or U9438 (N_9438,N_1230,N_5846);
nand U9439 (N_9439,N_435,N_3052);
xor U9440 (N_9440,N_791,N_1910);
xnor U9441 (N_9441,N_2511,N_4554);
nand U9442 (N_9442,N_5484,N_5562);
nor U9443 (N_9443,N_3680,N_2840);
or U9444 (N_9444,N_4750,N_4291);
nand U9445 (N_9445,N_1886,N_1911);
nand U9446 (N_9446,N_1425,N_2211);
and U9447 (N_9447,N_3497,N_4783);
xor U9448 (N_9448,N_2997,N_693);
or U9449 (N_9449,N_4527,N_2902);
or U9450 (N_9450,N_42,N_2497);
and U9451 (N_9451,N_5350,N_1535);
or U9452 (N_9452,N_4814,N_2155);
and U9453 (N_9453,N_3581,N_4584);
xor U9454 (N_9454,N_5148,N_229);
or U9455 (N_9455,N_3147,N_5222);
nand U9456 (N_9456,N_4164,N_451);
nand U9457 (N_9457,N_5546,N_2625);
and U9458 (N_9458,N_5564,N_3907);
and U9459 (N_9459,N_1328,N_4871);
and U9460 (N_9460,N_2938,N_4317);
and U9461 (N_9461,N_499,N_5816);
and U9462 (N_9462,N_1564,N_595);
xnor U9463 (N_9463,N_5099,N_1144);
nor U9464 (N_9464,N_5029,N_3007);
and U9465 (N_9465,N_1283,N_1937);
xor U9466 (N_9466,N_2367,N_1449);
or U9467 (N_9467,N_3199,N_3812);
nor U9468 (N_9468,N_2870,N_832);
nor U9469 (N_9469,N_4458,N_3521);
nor U9470 (N_9470,N_4638,N_1316);
xnor U9471 (N_9471,N_1055,N_5648);
nand U9472 (N_9472,N_1451,N_2665);
nor U9473 (N_9473,N_637,N_5897);
xor U9474 (N_9474,N_434,N_3041);
xor U9475 (N_9475,N_958,N_5467);
or U9476 (N_9476,N_3312,N_709);
and U9477 (N_9477,N_2374,N_1569);
xnor U9478 (N_9478,N_5299,N_1330);
nor U9479 (N_9479,N_5058,N_169);
and U9480 (N_9480,N_2170,N_5984);
xor U9481 (N_9481,N_3239,N_4968);
or U9482 (N_9482,N_5927,N_178);
and U9483 (N_9483,N_453,N_4968);
nand U9484 (N_9484,N_5105,N_2446);
and U9485 (N_9485,N_3606,N_817);
nand U9486 (N_9486,N_3440,N_3076);
and U9487 (N_9487,N_2142,N_5887);
nand U9488 (N_9488,N_3778,N_2461);
xor U9489 (N_9489,N_594,N_2280);
and U9490 (N_9490,N_4773,N_1479);
nor U9491 (N_9491,N_4769,N_2428);
nand U9492 (N_9492,N_2958,N_578);
xnor U9493 (N_9493,N_1842,N_402);
nor U9494 (N_9494,N_4320,N_4508);
or U9495 (N_9495,N_1726,N_4480);
xnor U9496 (N_9496,N_4389,N_3802);
and U9497 (N_9497,N_3600,N_1687);
or U9498 (N_9498,N_1078,N_3150);
xnor U9499 (N_9499,N_2818,N_3620);
and U9500 (N_9500,N_396,N_5117);
nor U9501 (N_9501,N_4756,N_1765);
nor U9502 (N_9502,N_208,N_5121);
and U9503 (N_9503,N_4556,N_108);
nand U9504 (N_9504,N_1008,N_1654);
and U9505 (N_9505,N_5276,N_790);
or U9506 (N_9506,N_3751,N_5176);
nand U9507 (N_9507,N_723,N_1640);
and U9508 (N_9508,N_3191,N_125);
or U9509 (N_9509,N_3180,N_3337);
nand U9510 (N_9510,N_3491,N_2790);
or U9511 (N_9511,N_2309,N_2094);
or U9512 (N_9512,N_1254,N_5868);
xnor U9513 (N_9513,N_3568,N_2699);
nor U9514 (N_9514,N_3449,N_1032);
nor U9515 (N_9515,N_2528,N_3874);
and U9516 (N_9516,N_2963,N_1773);
xor U9517 (N_9517,N_3050,N_1830);
or U9518 (N_9518,N_3837,N_3282);
nor U9519 (N_9519,N_3285,N_4423);
and U9520 (N_9520,N_2815,N_1717);
nor U9521 (N_9521,N_1170,N_903);
xnor U9522 (N_9522,N_304,N_5035);
nand U9523 (N_9523,N_3552,N_3843);
xnor U9524 (N_9524,N_1606,N_4522);
xor U9525 (N_9525,N_1924,N_2813);
and U9526 (N_9526,N_5397,N_3124);
nand U9527 (N_9527,N_3598,N_5372);
nor U9528 (N_9528,N_2776,N_907);
nand U9529 (N_9529,N_5607,N_1428);
nand U9530 (N_9530,N_1827,N_3130);
xnor U9531 (N_9531,N_3180,N_2101);
and U9532 (N_9532,N_921,N_197);
or U9533 (N_9533,N_222,N_5265);
nor U9534 (N_9534,N_3946,N_1787);
nand U9535 (N_9535,N_312,N_1173);
nor U9536 (N_9536,N_1466,N_2001);
nor U9537 (N_9537,N_4461,N_3980);
nand U9538 (N_9538,N_1626,N_1262);
nand U9539 (N_9539,N_2547,N_2419);
nand U9540 (N_9540,N_2748,N_944);
xnor U9541 (N_9541,N_5728,N_5044);
and U9542 (N_9542,N_4006,N_3579);
nor U9543 (N_9543,N_5864,N_3893);
or U9544 (N_9544,N_4664,N_1947);
nor U9545 (N_9545,N_5626,N_59);
nand U9546 (N_9546,N_4283,N_1365);
nand U9547 (N_9547,N_727,N_5122);
nand U9548 (N_9548,N_4723,N_2303);
nor U9549 (N_9549,N_848,N_2575);
nand U9550 (N_9550,N_709,N_2613);
xor U9551 (N_9551,N_2818,N_2236);
nand U9552 (N_9552,N_1200,N_3539);
or U9553 (N_9553,N_5060,N_501);
xnor U9554 (N_9554,N_3780,N_1334);
or U9555 (N_9555,N_1170,N_229);
or U9556 (N_9556,N_5339,N_4189);
nor U9557 (N_9557,N_2271,N_5093);
nor U9558 (N_9558,N_897,N_1346);
xnor U9559 (N_9559,N_4952,N_2512);
and U9560 (N_9560,N_3812,N_2545);
nor U9561 (N_9561,N_3598,N_2869);
or U9562 (N_9562,N_3061,N_4143);
or U9563 (N_9563,N_1266,N_65);
or U9564 (N_9564,N_4870,N_4331);
nand U9565 (N_9565,N_3849,N_330);
or U9566 (N_9566,N_933,N_347);
or U9567 (N_9567,N_1214,N_186);
nor U9568 (N_9568,N_1958,N_3712);
xor U9569 (N_9569,N_1091,N_3729);
or U9570 (N_9570,N_1227,N_905);
and U9571 (N_9571,N_3812,N_4838);
xor U9572 (N_9572,N_4106,N_1637);
nor U9573 (N_9573,N_615,N_4878);
or U9574 (N_9574,N_4767,N_1668);
xor U9575 (N_9575,N_5186,N_3901);
nor U9576 (N_9576,N_186,N_1405);
nand U9577 (N_9577,N_5926,N_2375);
nand U9578 (N_9578,N_5406,N_5596);
xnor U9579 (N_9579,N_2779,N_838);
or U9580 (N_9580,N_4666,N_634);
or U9581 (N_9581,N_5089,N_4151);
xnor U9582 (N_9582,N_5867,N_3583);
nor U9583 (N_9583,N_1569,N_4907);
xnor U9584 (N_9584,N_4255,N_760);
nand U9585 (N_9585,N_2704,N_5177);
or U9586 (N_9586,N_3414,N_5422);
nand U9587 (N_9587,N_2975,N_3245);
or U9588 (N_9588,N_3395,N_2159);
nor U9589 (N_9589,N_5411,N_2677);
and U9590 (N_9590,N_4485,N_4070);
nor U9591 (N_9591,N_3933,N_3370);
xor U9592 (N_9592,N_5566,N_3752);
or U9593 (N_9593,N_488,N_4044);
nand U9594 (N_9594,N_975,N_4135);
nand U9595 (N_9595,N_3574,N_503);
nand U9596 (N_9596,N_2255,N_810);
nand U9597 (N_9597,N_5343,N_2881);
xor U9598 (N_9598,N_3375,N_1049);
nor U9599 (N_9599,N_2860,N_5803);
nand U9600 (N_9600,N_3861,N_1905);
or U9601 (N_9601,N_891,N_520);
nand U9602 (N_9602,N_2111,N_2301);
nand U9603 (N_9603,N_1449,N_4796);
or U9604 (N_9604,N_4838,N_4534);
nand U9605 (N_9605,N_258,N_3959);
nor U9606 (N_9606,N_4653,N_1060);
nor U9607 (N_9607,N_2370,N_932);
and U9608 (N_9608,N_4682,N_28);
nor U9609 (N_9609,N_3132,N_735);
and U9610 (N_9610,N_376,N_3500);
nand U9611 (N_9611,N_2977,N_908);
xor U9612 (N_9612,N_855,N_466);
nor U9613 (N_9613,N_3495,N_4875);
nor U9614 (N_9614,N_1578,N_2090);
and U9615 (N_9615,N_5768,N_4393);
nand U9616 (N_9616,N_107,N_1810);
nand U9617 (N_9617,N_2151,N_4470);
nand U9618 (N_9618,N_4077,N_959);
and U9619 (N_9619,N_5698,N_2297);
or U9620 (N_9620,N_5454,N_2714);
or U9621 (N_9621,N_5795,N_4039);
nor U9622 (N_9622,N_5355,N_3054);
nor U9623 (N_9623,N_5167,N_3223);
nor U9624 (N_9624,N_1487,N_3957);
or U9625 (N_9625,N_5596,N_2586);
and U9626 (N_9626,N_3179,N_5293);
nor U9627 (N_9627,N_2037,N_4137);
nor U9628 (N_9628,N_3000,N_109);
nor U9629 (N_9629,N_5081,N_2027);
and U9630 (N_9630,N_3218,N_3075);
or U9631 (N_9631,N_4251,N_3623);
nor U9632 (N_9632,N_2760,N_1194);
nor U9633 (N_9633,N_4386,N_5165);
nand U9634 (N_9634,N_80,N_2376);
or U9635 (N_9635,N_2548,N_2545);
or U9636 (N_9636,N_4524,N_4444);
nor U9637 (N_9637,N_5417,N_4846);
and U9638 (N_9638,N_4855,N_4275);
or U9639 (N_9639,N_5277,N_688);
and U9640 (N_9640,N_5230,N_2514);
nor U9641 (N_9641,N_1446,N_2478);
and U9642 (N_9642,N_117,N_5870);
nor U9643 (N_9643,N_1854,N_3345);
or U9644 (N_9644,N_392,N_342);
or U9645 (N_9645,N_4938,N_5209);
xor U9646 (N_9646,N_842,N_209);
and U9647 (N_9647,N_5770,N_2412);
xor U9648 (N_9648,N_5042,N_5290);
nor U9649 (N_9649,N_1146,N_2801);
xor U9650 (N_9650,N_4593,N_4717);
and U9651 (N_9651,N_459,N_150);
and U9652 (N_9652,N_984,N_2880);
and U9653 (N_9653,N_149,N_218);
or U9654 (N_9654,N_5710,N_3965);
and U9655 (N_9655,N_5456,N_4275);
xor U9656 (N_9656,N_2589,N_5024);
nand U9657 (N_9657,N_2274,N_4917);
nor U9658 (N_9658,N_2562,N_4936);
nor U9659 (N_9659,N_1206,N_1889);
xnor U9660 (N_9660,N_1770,N_3912);
and U9661 (N_9661,N_1305,N_2289);
xor U9662 (N_9662,N_1647,N_5901);
xor U9663 (N_9663,N_5538,N_2046);
or U9664 (N_9664,N_1888,N_711);
and U9665 (N_9665,N_1450,N_5762);
and U9666 (N_9666,N_3841,N_4353);
nor U9667 (N_9667,N_3446,N_1665);
nor U9668 (N_9668,N_2945,N_5207);
nor U9669 (N_9669,N_1441,N_4790);
xnor U9670 (N_9670,N_496,N_5650);
nand U9671 (N_9671,N_489,N_4243);
nand U9672 (N_9672,N_5803,N_2819);
and U9673 (N_9673,N_933,N_1084);
nor U9674 (N_9674,N_3548,N_4010);
or U9675 (N_9675,N_5665,N_2988);
or U9676 (N_9676,N_3561,N_4222);
or U9677 (N_9677,N_1156,N_4859);
or U9678 (N_9678,N_1727,N_294);
and U9679 (N_9679,N_73,N_3800);
nor U9680 (N_9680,N_1079,N_1963);
xnor U9681 (N_9681,N_155,N_3232);
nor U9682 (N_9682,N_2337,N_2830);
or U9683 (N_9683,N_4207,N_4191);
or U9684 (N_9684,N_1599,N_1658);
nor U9685 (N_9685,N_5954,N_2521);
nor U9686 (N_9686,N_2321,N_697);
nand U9687 (N_9687,N_1667,N_1390);
or U9688 (N_9688,N_1319,N_3986);
nor U9689 (N_9689,N_964,N_3472);
and U9690 (N_9690,N_173,N_5380);
xnor U9691 (N_9691,N_3578,N_1146);
nand U9692 (N_9692,N_5271,N_4917);
xnor U9693 (N_9693,N_2988,N_3266);
and U9694 (N_9694,N_433,N_1336);
nand U9695 (N_9695,N_2773,N_366);
nand U9696 (N_9696,N_1551,N_5541);
and U9697 (N_9697,N_4549,N_4694);
or U9698 (N_9698,N_2541,N_184);
nand U9699 (N_9699,N_3900,N_3179);
nor U9700 (N_9700,N_1092,N_3839);
or U9701 (N_9701,N_3996,N_3054);
xnor U9702 (N_9702,N_1784,N_558);
and U9703 (N_9703,N_3741,N_2151);
nand U9704 (N_9704,N_1986,N_402);
or U9705 (N_9705,N_2739,N_152);
and U9706 (N_9706,N_4043,N_668);
xnor U9707 (N_9707,N_1853,N_4197);
xnor U9708 (N_9708,N_99,N_3421);
and U9709 (N_9709,N_1602,N_3990);
nor U9710 (N_9710,N_5553,N_1507);
and U9711 (N_9711,N_3741,N_2666);
nand U9712 (N_9712,N_2972,N_4812);
or U9713 (N_9713,N_1568,N_4350);
nand U9714 (N_9714,N_1400,N_3742);
xnor U9715 (N_9715,N_3008,N_5824);
nand U9716 (N_9716,N_4423,N_9);
and U9717 (N_9717,N_836,N_826);
and U9718 (N_9718,N_2606,N_5041);
nand U9719 (N_9719,N_2867,N_3189);
and U9720 (N_9720,N_916,N_4653);
nor U9721 (N_9721,N_5860,N_828);
nor U9722 (N_9722,N_29,N_225);
xnor U9723 (N_9723,N_2993,N_1533);
or U9724 (N_9724,N_1404,N_4111);
xnor U9725 (N_9725,N_3498,N_4452);
nor U9726 (N_9726,N_3681,N_675);
or U9727 (N_9727,N_2958,N_4233);
and U9728 (N_9728,N_4063,N_1867);
nand U9729 (N_9729,N_408,N_3829);
xor U9730 (N_9730,N_5128,N_263);
and U9731 (N_9731,N_3270,N_5631);
nor U9732 (N_9732,N_230,N_1313);
nand U9733 (N_9733,N_3261,N_2535);
nand U9734 (N_9734,N_1,N_944);
xnor U9735 (N_9735,N_2770,N_1684);
nand U9736 (N_9736,N_1669,N_3773);
nand U9737 (N_9737,N_3012,N_4351);
and U9738 (N_9738,N_969,N_5451);
nor U9739 (N_9739,N_652,N_117);
or U9740 (N_9740,N_4569,N_2641);
nor U9741 (N_9741,N_5213,N_4389);
xnor U9742 (N_9742,N_4167,N_4840);
and U9743 (N_9743,N_504,N_1810);
nand U9744 (N_9744,N_848,N_2769);
nand U9745 (N_9745,N_2370,N_2154);
and U9746 (N_9746,N_303,N_3720);
xor U9747 (N_9747,N_583,N_4092);
nand U9748 (N_9748,N_1424,N_2195);
or U9749 (N_9749,N_5116,N_5742);
xnor U9750 (N_9750,N_3250,N_2973);
nand U9751 (N_9751,N_5877,N_791);
nand U9752 (N_9752,N_5899,N_2619);
or U9753 (N_9753,N_885,N_953);
or U9754 (N_9754,N_70,N_5237);
or U9755 (N_9755,N_2567,N_4274);
nand U9756 (N_9756,N_1946,N_266);
and U9757 (N_9757,N_570,N_4273);
xnor U9758 (N_9758,N_1167,N_5876);
nor U9759 (N_9759,N_4648,N_3159);
xor U9760 (N_9760,N_4764,N_3872);
nor U9761 (N_9761,N_5332,N_3967);
nor U9762 (N_9762,N_2712,N_801);
nand U9763 (N_9763,N_2856,N_5165);
nand U9764 (N_9764,N_4531,N_4608);
nor U9765 (N_9765,N_5113,N_4706);
or U9766 (N_9766,N_2288,N_3029);
nor U9767 (N_9767,N_632,N_4114);
and U9768 (N_9768,N_5213,N_5732);
xnor U9769 (N_9769,N_671,N_1983);
nand U9770 (N_9770,N_5772,N_1359);
or U9771 (N_9771,N_3845,N_4886);
and U9772 (N_9772,N_5817,N_456);
nor U9773 (N_9773,N_2552,N_3441);
or U9774 (N_9774,N_1322,N_2441);
xor U9775 (N_9775,N_1623,N_3816);
nand U9776 (N_9776,N_1011,N_4189);
nor U9777 (N_9777,N_5117,N_5842);
nor U9778 (N_9778,N_3479,N_942);
and U9779 (N_9779,N_55,N_5593);
and U9780 (N_9780,N_4251,N_545);
nor U9781 (N_9781,N_2958,N_2400);
or U9782 (N_9782,N_4938,N_1113);
or U9783 (N_9783,N_900,N_1893);
or U9784 (N_9784,N_1088,N_4172);
nand U9785 (N_9785,N_5293,N_3856);
nand U9786 (N_9786,N_318,N_2617);
or U9787 (N_9787,N_2863,N_2002);
xnor U9788 (N_9788,N_4824,N_2146);
and U9789 (N_9789,N_5075,N_1746);
nor U9790 (N_9790,N_1693,N_2421);
and U9791 (N_9791,N_2121,N_2383);
xor U9792 (N_9792,N_3279,N_3327);
nand U9793 (N_9793,N_1231,N_496);
xor U9794 (N_9794,N_3265,N_906);
xnor U9795 (N_9795,N_1486,N_5257);
nor U9796 (N_9796,N_1801,N_3710);
xor U9797 (N_9797,N_4142,N_772);
xor U9798 (N_9798,N_5558,N_3372);
nand U9799 (N_9799,N_3851,N_3713);
xor U9800 (N_9800,N_4621,N_5377);
nor U9801 (N_9801,N_1623,N_5402);
and U9802 (N_9802,N_152,N_1013);
nor U9803 (N_9803,N_4591,N_4003);
and U9804 (N_9804,N_3708,N_1324);
nand U9805 (N_9805,N_3652,N_4221);
xor U9806 (N_9806,N_3705,N_3434);
and U9807 (N_9807,N_3541,N_5340);
xnor U9808 (N_9808,N_4293,N_2643);
nand U9809 (N_9809,N_288,N_2627);
or U9810 (N_9810,N_3523,N_5427);
nand U9811 (N_9811,N_2659,N_632);
or U9812 (N_9812,N_2708,N_205);
nor U9813 (N_9813,N_3870,N_1530);
nor U9814 (N_9814,N_4839,N_2646);
or U9815 (N_9815,N_3861,N_887);
or U9816 (N_9816,N_2385,N_66);
nor U9817 (N_9817,N_4418,N_306);
nor U9818 (N_9818,N_5658,N_2456);
xnor U9819 (N_9819,N_842,N_4855);
xor U9820 (N_9820,N_3515,N_2015);
nor U9821 (N_9821,N_2337,N_664);
or U9822 (N_9822,N_1633,N_5254);
nand U9823 (N_9823,N_4623,N_1519);
or U9824 (N_9824,N_4246,N_2251);
nor U9825 (N_9825,N_5913,N_2014);
nand U9826 (N_9826,N_2578,N_3322);
and U9827 (N_9827,N_827,N_2041);
nor U9828 (N_9828,N_5329,N_5535);
nand U9829 (N_9829,N_2915,N_5318);
or U9830 (N_9830,N_2396,N_5350);
xor U9831 (N_9831,N_142,N_2972);
or U9832 (N_9832,N_3617,N_3244);
nand U9833 (N_9833,N_79,N_2741);
nand U9834 (N_9834,N_5599,N_394);
xnor U9835 (N_9835,N_4171,N_3929);
or U9836 (N_9836,N_3172,N_514);
or U9837 (N_9837,N_1417,N_4270);
xnor U9838 (N_9838,N_2318,N_5561);
nand U9839 (N_9839,N_2216,N_3485);
xnor U9840 (N_9840,N_2464,N_2890);
or U9841 (N_9841,N_270,N_5901);
or U9842 (N_9842,N_5866,N_4778);
nor U9843 (N_9843,N_2435,N_3871);
and U9844 (N_9844,N_4319,N_1553);
nor U9845 (N_9845,N_4137,N_2484);
nand U9846 (N_9846,N_351,N_3622);
nor U9847 (N_9847,N_2867,N_130);
xor U9848 (N_9848,N_171,N_3960);
nand U9849 (N_9849,N_388,N_5720);
nand U9850 (N_9850,N_2764,N_3420);
or U9851 (N_9851,N_1284,N_825);
xnor U9852 (N_9852,N_4613,N_2100);
nand U9853 (N_9853,N_137,N_2417);
and U9854 (N_9854,N_1322,N_1416);
nand U9855 (N_9855,N_1426,N_5907);
xor U9856 (N_9856,N_4909,N_4386);
xnor U9857 (N_9857,N_2315,N_623);
nand U9858 (N_9858,N_5761,N_5672);
and U9859 (N_9859,N_2702,N_4469);
nor U9860 (N_9860,N_4025,N_5515);
nor U9861 (N_9861,N_787,N_3337);
or U9862 (N_9862,N_5117,N_5823);
nor U9863 (N_9863,N_1836,N_4620);
xor U9864 (N_9864,N_5680,N_5210);
nand U9865 (N_9865,N_2606,N_2171);
nand U9866 (N_9866,N_1130,N_4976);
nand U9867 (N_9867,N_2380,N_2449);
xor U9868 (N_9868,N_883,N_3318);
xor U9869 (N_9869,N_1464,N_5647);
xor U9870 (N_9870,N_4412,N_5449);
or U9871 (N_9871,N_805,N_4686);
nand U9872 (N_9872,N_215,N_5555);
and U9873 (N_9873,N_1471,N_5561);
xor U9874 (N_9874,N_1441,N_3352);
xnor U9875 (N_9875,N_2779,N_1912);
and U9876 (N_9876,N_2886,N_125);
nand U9877 (N_9877,N_2488,N_1243);
or U9878 (N_9878,N_4020,N_983);
nand U9879 (N_9879,N_3955,N_3700);
or U9880 (N_9880,N_4789,N_1055);
nand U9881 (N_9881,N_2579,N_5696);
or U9882 (N_9882,N_5323,N_2256);
xnor U9883 (N_9883,N_500,N_8);
xor U9884 (N_9884,N_4616,N_4100);
xnor U9885 (N_9885,N_4104,N_3957);
nand U9886 (N_9886,N_4938,N_2638);
xor U9887 (N_9887,N_1795,N_3069);
nand U9888 (N_9888,N_5216,N_4144);
or U9889 (N_9889,N_3012,N_3963);
xor U9890 (N_9890,N_1939,N_1602);
or U9891 (N_9891,N_4353,N_5991);
xor U9892 (N_9892,N_3209,N_5751);
or U9893 (N_9893,N_3155,N_848);
xor U9894 (N_9894,N_1042,N_1640);
or U9895 (N_9895,N_2533,N_1088);
xor U9896 (N_9896,N_2696,N_603);
xnor U9897 (N_9897,N_4628,N_4957);
nand U9898 (N_9898,N_5383,N_2019);
nor U9899 (N_9899,N_2855,N_227);
nor U9900 (N_9900,N_4261,N_5042);
xnor U9901 (N_9901,N_1626,N_2633);
nor U9902 (N_9902,N_2493,N_2697);
nor U9903 (N_9903,N_1438,N_214);
and U9904 (N_9904,N_1765,N_2069);
and U9905 (N_9905,N_4170,N_1810);
xnor U9906 (N_9906,N_4383,N_838);
xnor U9907 (N_9907,N_4151,N_3022);
and U9908 (N_9908,N_5319,N_2901);
xor U9909 (N_9909,N_1503,N_4512);
or U9910 (N_9910,N_3923,N_2875);
and U9911 (N_9911,N_1202,N_1608);
xor U9912 (N_9912,N_78,N_3675);
or U9913 (N_9913,N_4499,N_2173);
or U9914 (N_9914,N_3877,N_2638);
or U9915 (N_9915,N_3399,N_5272);
nor U9916 (N_9916,N_3830,N_4164);
xor U9917 (N_9917,N_4035,N_1901);
nand U9918 (N_9918,N_2533,N_1625);
nor U9919 (N_9919,N_5709,N_2307);
nor U9920 (N_9920,N_3716,N_3776);
and U9921 (N_9921,N_4796,N_3211);
and U9922 (N_9922,N_1112,N_1371);
nand U9923 (N_9923,N_3231,N_224);
nand U9924 (N_9924,N_5050,N_2286);
xor U9925 (N_9925,N_2766,N_4600);
or U9926 (N_9926,N_3504,N_3529);
or U9927 (N_9927,N_2313,N_1118);
and U9928 (N_9928,N_3395,N_3055);
xor U9929 (N_9929,N_4466,N_2254);
or U9930 (N_9930,N_2291,N_292);
and U9931 (N_9931,N_2578,N_1489);
and U9932 (N_9932,N_4578,N_4491);
nor U9933 (N_9933,N_321,N_3359);
xnor U9934 (N_9934,N_1763,N_4442);
xnor U9935 (N_9935,N_4939,N_2477);
nand U9936 (N_9936,N_2437,N_3465);
nand U9937 (N_9937,N_3289,N_1722);
nor U9938 (N_9938,N_3273,N_5833);
nand U9939 (N_9939,N_2117,N_1758);
nor U9940 (N_9940,N_4849,N_3643);
xnor U9941 (N_9941,N_2436,N_4889);
nor U9942 (N_9942,N_5354,N_792);
and U9943 (N_9943,N_271,N_4827);
or U9944 (N_9944,N_5756,N_3130);
and U9945 (N_9945,N_87,N_1335);
and U9946 (N_9946,N_2295,N_543);
or U9947 (N_9947,N_144,N_2856);
or U9948 (N_9948,N_52,N_962);
and U9949 (N_9949,N_3820,N_5727);
nor U9950 (N_9950,N_1529,N_597);
or U9951 (N_9951,N_4930,N_2019);
nand U9952 (N_9952,N_1489,N_1620);
nand U9953 (N_9953,N_3939,N_2342);
or U9954 (N_9954,N_5797,N_1270);
xnor U9955 (N_9955,N_5796,N_3830);
xnor U9956 (N_9956,N_5524,N_1131);
nor U9957 (N_9957,N_2082,N_4585);
or U9958 (N_9958,N_395,N_1250);
and U9959 (N_9959,N_3999,N_4222);
or U9960 (N_9960,N_4944,N_2715);
nor U9961 (N_9961,N_3641,N_394);
and U9962 (N_9962,N_4673,N_3125);
xor U9963 (N_9963,N_5819,N_4080);
or U9964 (N_9964,N_489,N_1819);
and U9965 (N_9965,N_1601,N_1866);
and U9966 (N_9966,N_4292,N_423);
xnor U9967 (N_9967,N_3096,N_2990);
or U9968 (N_9968,N_4503,N_1237);
or U9969 (N_9969,N_4512,N_5652);
nand U9970 (N_9970,N_3831,N_282);
or U9971 (N_9971,N_3942,N_3985);
and U9972 (N_9972,N_2106,N_4644);
or U9973 (N_9973,N_2767,N_1213);
nor U9974 (N_9974,N_5381,N_4073);
or U9975 (N_9975,N_2060,N_1297);
and U9976 (N_9976,N_3985,N_2471);
or U9977 (N_9977,N_1216,N_3041);
nand U9978 (N_9978,N_2962,N_4165);
and U9979 (N_9979,N_5910,N_740);
and U9980 (N_9980,N_2311,N_4439);
nor U9981 (N_9981,N_2049,N_4254);
xnor U9982 (N_9982,N_4338,N_2193);
nand U9983 (N_9983,N_4726,N_2322);
xor U9984 (N_9984,N_4713,N_3805);
or U9985 (N_9985,N_2760,N_3213);
and U9986 (N_9986,N_3868,N_1628);
xor U9987 (N_9987,N_3449,N_5190);
and U9988 (N_9988,N_621,N_2724);
nor U9989 (N_9989,N_72,N_4659);
or U9990 (N_9990,N_143,N_3390);
nor U9991 (N_9991,N_1996,N_3924);
xor U9992 (N_9992,N_54,N_5446);
xnor U9993 (N_9993,N_1624,N_3048);
or U9994 (N_9994,N_5901,N_5228);
nand U9995 (N_9995,N_5731,N_2156);
nand U9996 (N_9996,N_1600,N_821);
nor U9997 (N_9997,N_3850,N_741);
xnor U9998 (N_9998,N_296,N_797);
xnor U9999 (N_9999,N_2302,N_2657);
and U10000 (N_10000,N_778,N_1066);
nand U10001 (N_10001,N_1647,N_2731);
nor U10002 (N_10002,N_5689,N_4117);
nor U10003 (N_10003,N_1158,N_4732);
xor U10004 (N_10004,N_755,N_4905);
nor U10005 (N_10005,N_2270,N_2083);
or U10006 (N_10006,N_2050,N_1426);
nand U10007 (N_10007,N_4789,N_1301);
nand U10008 (N_10008,N_4083,N_1915);
and U10009 (N_10009,N_108,N_133);
and U10010 (N_10010,N_4594,N_3827);
and U10011 (N_10011,N_3430,N_5482);
and U10012 (N_10012,N_5435,N_63);
nor U10013 (N_10013,N_1972,N_1101);
nand U10014 (N_10014,N_5929,N_5892);
and U10015 (N_10015,N_3955,N_196);
nor U10016 (N_10016,N_1354,N_2701);
or U10017 (N_10017,N_5797,N_5103);
and U10018 (N_10018,N_4102,N_4851);
and U10019 (N_10019,N_3332,N_5515);
nand U10020 (N_10020,N_5486,N_5094);
or U10021 (N_10021,N_583,N_5841);
xor U10022 (N_10022,N_3133,N_125);
nand U10023 (N_10023,N_3152,N_3431);
nor U10024 (N_10024,N_907,N_2960);
nand U10025 (N_10025,N_1999,N_440);
nand U10026 (N_10026,N_938,N_2500);
or U10027 (N_10027,N_1563,N_129);
and U10028 (N_10028,N_2963,N_5671);
and U10029 (N_10029,N_1859,N_56);
and U10030 (N_10030,N_2556,N_1267);
and U10031 (N_10031,N_5974,N_3669);
or U10032 (N_10032,N_5604,N_4295);
xor U10033 (N_10033,N_19,N_286);
nand U10034 (N_10034,N_1297,N_1334);
nand U10035 (N_10035,N_2356,N_4271);
and U10036 (N_10036,N_5389,N_5693);
nor U10037 (N_10037,N_2709,N_3352);
or U10038 (N_10038,N_3689,N_3924);
xor U10039 (N_10039,N_1554,N_1398);
nor U10040 (N_10040,N_674,N_1375);
xnor U10041 (N_10041,N_5200,N_4007);
or U10042 (N_10042,N_5288,N_2716);
or U10043 (N_10043,N_3058,N_5368);
nor U10044 (N_10044,N_5846,N_4420);
nor U10045 (N_10045,N_3932,N_4889);
xor U10046 (N_10046,N_1655,N_274);
nor U10047 (N_10047,N_1505,N_2054);
and U10048 (N_10048,N_5087,N_5268);
nor U10049 (N_10049,N_266,N_2908);
nand U10050 (N_10050,N_545,N_4668);
or U10051 (N_10051,N_525,N_1208);
or U10052 (N_10052,N_1410,N_4845);
or U10053 (N_10053,N_5312,N_1291);
and U10054 (N_10054,N_1246,N_806);
and U10055 (N_10055,N_5410,N_133);
and U10056 (N_10056,N_2273,N_4031);
nor U10057 (N_10057,N_3585,N_4360);
or U10058 (N_10058,N_4217,N_3091);
nor U10059 (N_10059,N_1299,N_2155);
nor U10060 (N_10060,N_3525,N_4140);
xnor U10061 (N_10061,N_2506,N_4345);
nand U10062 (N_10062,N_1266,N_1968);
nand U10063 (N_10063,N_1754,N_5745);
nand U10064 (N_10064,N_2921,N_4455);
and U10065 (N_10065,N_1149,N_2856);
or U10066 (N_10066,N_2114,N_4607);
and U10067 (N_10067,N_3508,N_2134);
xnor U10068 (N_10068,N_3008,N_3527);
nor U10069 (N_10069,N_4989,N_5415);
nor U10070 (N_10070,N_1556,N_5367);
and U10071 (N_10071,N_2088,N_2996);
or U10072 (N_10072,N_5398,N_2972);
xnor U10073 (N_10073,N_280,N_2697);
nor U10074 (N_10074,N_828,N_4623);
xor U10075 (N_10075,N_5939,N_2824);
and U10076 (N_10076,N_3251,N_5396);
nand U10077 (N_10077,N_5179,N_2847);
xor U10078 (N_10078,N_1445,N_1571);
nor U10079 (N_10079,N_4059,N_255);
xnor U10080 (N_10080,N_2628,N_3595);
nor U10081 (N_10081,N_722,N_4853);
xnor U10082 (N_10082,N_4991,N_3911);
nor U10083 (N_10083,N_1267,N_1481);
xor U10084 (N_10084,N_3183,N_3625);
nor U10085 (N_10085,N_994,N_1501);
and U10086 (N_10086,N_2232,N_2188);
and U10087 (N_10087,N_5682,N_1661);
or U10088 (N_10088,N_2243,N_1380);
xor U10089 (N_10089,N_5977,N_157);
nand U10090 (N_10090,N_4219,N_245);
nor U10091 (N_10091,N_2606,N_4583);
and U10092 (N_10092,N_391,N_3463);
nand U10093 (N_10093,N_867,N_1381);
nand U10094 (N_10094,N_72,N_5416);
xor U10095 (N_10095,N_2688,N_3447);
nor U10096 (N_10096,N_5237,N_610);
xor U10097 (N_10097,N_3574,N_5045);
or U10098 (N_10098,N_1797,N_4298);
or U10099 (N_10099,N_801,N_3460);
and U10100 (N_10100,N_5894,N_34);
nand U10101 (N_10101,N_5695,N_4093);
nor U10102 (N_10102,N_4621,N_1295);
nand U10103 (N_10103,N_5686,N_3076);
or U10104 (N_10104,N_3383,N_3260);
and U10105 (N_10105,N_2196,N_1237);
and U10106 (N_10106,N_218,N_1216);
nor U10107 (N_10107,N_3653,N_4532);
nor U10108 (N_10108,N_1198,N_4705);
nand U10109 (N_10109,N_3512,N_3204);
nor U10110 (N_10110,N_1533,N_3624);
and U10111 (N_10111,N_5359,N_5036);
nand U10112 (N_10112,N_5090,N_1025);
xor U10113 (N_10113,N_1462,N_2073);
nor U10114 (N_10114,N_3334,N_5744);
xnor U10115 (N_10115,N_1739,N_2550);
and U10116 (N_10116,N_1732,N_5251);
nor U10117 (N_10117,N_4589,N_4044);
xor U10118 (N_10118,N_5048,N_4548);
nor U10119 (N_10119,N_320,N_5163);
and U10120 (N_10120,N_5845,N_4365);
and U10121 (N_10121,N_5074,N_2249);
nor U10122 (N_10122,N_5833,N_19);
nor U10123 (N_10123,N_1570,N_1322);
xor U10124 (N_10124,N_4120,N_4090);
or U10125 (N_10125,N_5333,N_3355);
or U10126 (N_10126,N_2202,N_2335);
and U10127 (N_10127,N_5761,N_1751);
or U10128 (N_10128,N_2406,N_4977);
nor U10129 (N_10129,N_912,N_2077);
and U10130 (N_10130,N_3031,N_3375);
nor U10131 (N_10131,N_3515,N_1841);
nand U10132 (N_10132,N_1961,N_3631);
and U10133 (N_10133,N_5914,N_3371);
and U10134 (N_10134,N_5168,N_3484);
and U10135 (N_10135,N_779,N_5555);
xor U10136 (N_10136,N_2969,N_1715);
or U10137 (N_10137,N_4562,N_792);
nor U10138 (N_10138,N_4569,N_1804);
and U10139 (N_10139,N_5110,N_915);
nor U10140 (N_10140,N_2694,N_280);
nor U10141 (N_10141,N_5265,N_5411);
nand U10142 (N_10142,N_1065,N_2256);
or U10143 (N_10143,N_4919,N_2847);
xor U10144 (N_10144,N_1995,N_5666);
or U10145 (N_10145,N_288,N_928);
nand U10146 (N_10146,N_5134,N_3788);
or U10147 (N_10147,N_545,N_5516);
nor U10148 (N_10148,N_5799,N_727);
and U10149 (N_10149,N_5791,N_2624);
xnor U10150 (N_10150,N_190,N_5715);
nand U10151 (N_10151,N_3045,N_3921);
xnor U10152 (N_10152,N_1758,N_4998);
and U10153 (N_10153,N_5753,N_5081);
or U10154 (N_10154,N_2879,N_377);
nand U10155 (N_10155,N_180,N_839);
nor U10156 (N_10156,N_4775,N_5437);
or U10157 (N_10157,N_758,N_4283);
nor U10158 (N_10158,N_4101,N_3714);
and U10159 (N_10159,N_2378,N_803);
and U10160 (N_10160,N_3023,N_3176);
xor U10161 (N_10161,N_5797,N_2683);
and U10162 (N_10162,N_4074,N_2471);
nor U10163 (N_10163,N_2470,N_1740);
xor U10164 (N_10164,N_5136,N_1645);
nor U10165 (N_10165,N_5159,N_4379);
or U10166 (N_10166,N_5563,N_4743);
nand U10167 (N_10167,N_4789,N_2332);
xnor U10168 (N_10168,N_5187,N_1196);
xor U10169 (N_10169,N_376,N_4514);
nand U10170 (N_10170,N_885,N_4520);
or U10171 (N_10171,N_1358,N_5543);
nand U10172 (N_10172,N_958,N_1600);
or U10173 (N_10173,N_5745,N_3050);
and U10174 (N_10174,N_4953,N_1708);
xor U10175 (N_10175,N_2950,N_1529);
xor U10176 (N_10176,N_764,N_3289);
and U10177 (N_10177,N_2909,N_4191);
or U10178 (N_10178,N_3919,N_4467);
and U10179 (N_10179,N_3443,N_4334);
or U10180 (N_10180,N_974,N_2054);
xor U10181 (N_10181,N_2119,N_3107);
xor U10182 (N_10182,N_3651,N_102);
nand U10183 (N_10183,N_461,N_4767);
nand U10184 (N_10184,N_3236,N_870);
nor U10185 (N_10185,N_5687,N_2028);
or U10186 (N_10186,N_5979,N_5283);
or U10187 (N_10187,N_550,N_1730);
nor U10188 (N_10188,N_4018,N_662);
or U10189 (N_10189,N_1138,N_641);
nand U10190 (N_10190,N_5362,N_4577);
nand U10191 (N_10191,N_766,N_2781);
or U10192 (N_10192,N_1910,N_1070);
nor U10193 (N_10193,N_415,N_664);
nand U10194 (N_10194,N_4633,N_4309);
nor U10195 (N_10195,N_2805,N_2756);
nor U10196 (N_10196,N_5070,N_1223);
or U10197 (N_10197,N_2234,N_5869);
nor U10198 (N_10198,N_4301,N_5731);
nor U10199 (N_10199,N_1814,N_1575);
nand U10200 (N_10200,N_3695,N_2588);
or U10201 (N_10201,N_24,N_1420);
xor U10202 (N_10202,N_3179,N_3488);
nand U10203 (N_10203,N_2435,N_385);
xor U10204 (N_10204,N_4670,N_965);
xor U10205 (N_10205,N_1018,N_5664);
or U10206 (N_10206,N_5231,N_5219);
xor U10207 (N_10207,N_5881,N_254);
nand U10208 (N_10208,N_5613,N_1404);
or U10209 (N_10209,N_3721,N_3692);
and U10210 (N_10210,N_89,N_5450);
and U10211 (N_10211,N_1860,N_2398);
and U10212 (N_10212,N_2579,N_3175);
nand U10213 (N_10213,N_4332,N_2352);
or U10214 (N_10214,N_268,N_976);
nand U10215 (N_10215,N_101,N_1178);
and U10216 (N_10216,N_4539,N_2002);
nand U10217 (N_10217,N_1307,N_511);
nor U10218 (N_10218,N_1615,N_3713);
or U10219 (N_10219,N_662,N_884);
xnor U10220 (N_10220,N_4761,N_4435);
nor U10221 (N_10221,N_901,N_5292);
nor U10222 (N_10222,N_2479,N_2717);
nand U10223 (N_10223,N_1724,N_3278);
nand U10224 (N_10224,N_5108,N_2044);
or U10225 (N_10225,N_2633,N_927);
xor U10226 (N_10226,N_888,N_3573);
and U10227 (N_10227,N_3457,N_3227);
nand U10228 (N_10228,N_754,N_5038);
and U10229 (N_10229,N_2725,N_1683);
nand U10230 (N_10230,N_300,N_3913);
or U10231 (N_10231,N_4859,N_5068);
xnor U10232 (N_10232,N_5040,N_2267);
and U10233 (N_10233,N_1600,N_3999);
nor U10234 (N_10234,N_3888,N_1919);
nor U10235 (N_10235,N_2681,N_819);
xnor U10236 (N_10236,N_2508,N_4273);
or U10237 (N_10237,N_1565,N_4329);
or U10238 (N_10238,N_4607,N_5630);
and U10239 (N_10239,N_2099,N_4070);
xor U10240 (N_10240,N_2193,N_2975);
nor U10241 (N_10241,N_2812,N_1339);
or U10242 (N_10242,N_1761,N_5024);
and U10243 (N_10243,N_1517,N_1840);
nor U10244 (N_10244,N_3941,N_5089);
nor U10245 (N_10245,N_955,N_3020);
xor U10246 (N_10246,N_2822,N_434);
nor U10247 (N_10247,N_1503,N_1773);
nand U10248 (N_10248,N_2095,N_941);
or U10249 (N_10249,N_3211,N_4324);
nand U10250 (N_10250,N_5234,N_2862);
nor U10251 (N_10251,N_3627,N_1118);
nand U10252 (N_10252,N_3937,N_5915);
nand U10253 (N_10253,N_3725,N_1310);
xnor U10254 (N_10254,N_3140,N_4719);
xor U10255 (N_10255,N_4439,N_491);
nand U10256 (N_10256,N_4422,N_436);
or U10257 (N_10257,N_4363,N_4698);
xnor U10258 (N_10258,N_3890,N_3656);
or U10259 (N_10259,N_4341,N_1830);
and U10260 (N_10260,N_2908,N_341);
or U10261 (N_10261,N_5241,N_5215);
nand U10262 (N_10262,N_5307,N_2491);
or U10263 (N_10263,N_4418,N_1888);
xnor U10264 (N_10264,N_1529,N_2587);
xnor U10265 (N_10265,N_2968,N_3652);
and U10266 (N_10266,N_3630,N_881);
or U10267 (N_10267,N_4479,N_53);
nand U10268 (N_10268,N_2105,N_1838);
nand U10269 (N_10269,N_5391,N_5387);
nand U10270 (N_10270,N_4766,N_2595);
nor U10271 (N_10271,N_3771,N_3329);
or U10272 (N_10272,N_3782,N_215);
xor U10273 (N_10273,N_157,N_2176);
or U10274 (N_10274,N_4496,N_5965);
or U10275 (N_10275,N_2742,N_459);
nand U10276 (N_10276,N_2984,N_1705);
xnor U10277 (N_10277,N_2196,N_5310);
nor U10278 (N_10278,N_617,N_3184);
or U10279 (N_10279,N_1908,N_1720);
nand U10280 (N_10280,N_4861,N_512);
nor U10281 (N_10281,N_719,N_109);
and U10282 (N_10282,N_421,N_2315);
nand U10283 (N_10283,N_4444,N_5160);
xnor U10284 (N_10284,N_2074,N_881);
xor U10285 (N_10285,N_4530,N_5188);
or U10286 (N_10286,N_1058,N_4325);
or U10287 (N_10287,N_2186,N_5583);
or U10288 (N_10288,N_2694,N_5932);
nor U10289 (N_10289,N_2128,N_2109);
xor U10290 (N_10290,N_4655,N_79);
and U10291 (N_10291,N_1783,N_4253);
nor U10292 (N_10292,N_3794,N_3893);
nand U10293 (N_10293,N_2664,N_5150);
and U10294 (N_10294,N_4915,N_5191);
and U10295 (N_10295,N_4698,N_335);
or U10296 (N_10296,N_3987,N_1800);
nand U10297 (N_10297,N_1096,N_3396);
xor U10298 (N_10298,N_2489,N_2412);
nor U10299 (N_10299,N_1189,N_634);
and U10300 (N_10300,N_655,N_1457);
and U10301 (N_10301,N_1736,N_132);
nor U10302 (N_10302,N_1745,N_2266);
nand U10303 (N_10303,N_1549,N_4993);
nand U10304 (N_10304,N_3750,N_817);
or U10305 (N_10305,N_3669,N_1419);
xor U10306 (N_10306,N_2309,N_3423);
and U10307 (N_10307,N_2404,N_4485);
or U10308 (N_10308,N_2729,N_4206);
and U10309 (N_10309,N_5368,N_2147);
nand U10310 (N_10310,N_4198,N_3558);
nor U10311 (N_10311,N_3717,N_2355);
and U10312 (N_10312,N_436,N_4692);
xor U10313 (N_10313,N_5125,N_248);
or U10314 (N_10314,N_1483,N_3528);
or U10315 (N_10315,N_4399,N_3769);
xnor U10316 (N_10316,N_5903,N_4594);
or U10317 (N_10317,N_1889,N_3310);
xnor U10318 (N_10318,N_5858,N_1880);
nand U10319 (N_10319,N_1307,N_2559);
or U10320 (N_10320,N_4,N_3782);
and U10321 (N_10321,N_901,N_211);
and U10322 (N_10322,N_647,N_32);
xor U10323 (N_10323,N_5084,N_3229);
or U10324 (N_10324,N_2187,N_3006);
nor U10325 (N_10325,N_4565,N_282);
xor U10326 (N_10326,N_3772,N_5415);
and U10327 (N_10327,N_3838,N_539);
xor U10328 (N_10328,N_2266,N_2995);
xor U10329 (N_10329,N_1109,N_3194);
nor U10330 (N_10330,N_1886,N_5115);
xor U10331 (N_10331,N_5360,N_3276);
nor U10332 (N_10332,N_3175,N_1623);
or U10333 (N_10333,N_2957,N_2021);
nand U10334 (N_10334,N_4095,N_325);
and U10335 (N_10335,N_3377,N_3110);
or U10336 (N_10336,N_5275,N_3515);
xor U10337 (N_10337,N_3095,N_1875);
xnor U10338 (N_10338,N_3473,N_2361);
nand U10339 (N_10339,N_5457,N_500);
nor U10340 (N_10340,N_1396,N_775);
nor U10341 (N_10341,N_4340,N_5359);
or U10342 (N_10342,N_1180,N_3692);
or U10343 (N_10343,N_1274,N_153);
nand U10344 (N_10344,N_3650,N_3857);
nor U10345 (N_10345,N_430,N_5641);
nor U10346 (N_10346,N_5034,N_2438);
nor U10347 (N_10347,N_821,N_5904);
xor U10348 (N_10348,N_1665,N_5733);
nor U10349 (N_10349,N_1664,N_621);
or U10350 (N_10350,N_5745,N_24);
or U10351 (N_10351,N_1202,N_5209);
nand U10352 (N_10352,N_5817,N_5511);
and U10353 (N_10353,N_396,N_4016);
xor U10354 (N_10354,N_1886,N_5453);
xor U10355 (N_10355,N_4216,N_3514);
or U10356 (N_10356,N_4781,N_4462);
or U10357 (N_10357,N_5515,N_1);
nand U10358 (N_10358,N_5968,N_4174);
nor U10359 (N_10359,N_1264,N_2448);
nand U10360 (N_10360,N_1040,N_5161);
nor U10361 (N_10361,N_2982,N_1930);
and U10362 (N_10362,N_4659,N_4382);
nor U10363 (N_10363,N_332,N_1522);
nor U10364 (N_10364,N_5700,N_2862);
and U10365 (N_10365,N_562,N_1814);
and U10366 (N_10366,N_235,N_4774);
nand U10367 (N_10367,N_1560,N_2996);
nor U10368 (N_10368,N_1325,N_825);
xnor U10369 (N_10369,N_4890,N_1959);
xnor U10370 (N_10370,N_549,N_3812);
and U10371 (N_10371,N_2157,N_1395);
nand U10372 (N_10372,N_304,N_5920);
nand U10373 (N_10373,N_1740,N_4769);
nor U10374 (N_10374,N_2608,N_2923);
nand U10375 (N_10375,N_1502,N_3102);
and U10376 (N_10376,N_1904,N_233);
nand U10377 (N_10377,N_235,N_1700);
nor U10378 (N_10378,N_4596,N_4061);
xor U10379 (N_10379,N_3156,N_5604);
or U10380 (N_10380,N_1637,N_4679);
or U10381 (N_10381,N_1653,N_5558);
nor U10382 (N_10382,N_91,N_1212);
and U10383 (N_10383,N_794,N_4861);
nor U10384 (N_10384,N_1376,N_1675);
and U10385 (N_10385,N_3113,N_5003);
or U10386 (N_10386,N_3075,N_3336);
and U10387 (N_10387,N_3924,N_5112);
nand U10388 (N_10388,N_831,N_4150);
nand U10389 (N_10389,N_5790,N_3310);
xor U10390 (N_10390,N_92,N_3036);
or U10391 (N_10391,N_1855,N_2668);
nand U10392 (N_10392,N_870,N_4191);
or U10393 (N_10393,N_2881,N_5595);
nor U10394 (N_10394,N_1374,N_3593);
and U10395 (N_10395,N_957,N_3676);
xor U10396 (N_10396,N_3537,N_609);
nor U10397 (N_10397,N_5340,N_2552);
and U10398 (N_10398,N_487,N_2872);
xnor U10399 (N_10399,N_2406,N_5865);
xnor U10400 (N_10400,N_5783,N_4514);
and U10401 (N_10401,N_1086,N_4270);
and U10402 (N_10402,N_5680,N_260);
or U10403 (N_10403,N_4358,N_3866);
xor U10404 (N_10404,N_4564,N_5352);
nand U10405 (N_10405,N_5161,N_1368);
or U10406 (N_10406,N_9,N_2216);
or U10407 (N_10407,N_1634,N_5457);
nor U10408 (N_10408,N_1669,N_2009);
nand U10409 (N_10409,N_851,N_3969);
nand U10410 (N_10410,N_4670,N_2252);
nor U10411 (N_10411,N_460,N_5980);
or U10412 (N_10412,N_2923,N_2634);
xor U10413 (N_10413,N_3477,N_351);
nor U10414 (N_10414,N_1381,N_1012);
or U10415 (N_10415,N_5694,N_1580);
and U10416 (N_10416,N_1363,N_4617);
nor U10417 (N_10417,N_4002,N_372);
nand U10418 (N_10418,N_741,N_4284);
and U10419 (N_10419,N_744,N_2827);
xnor U10420 (N_10420,N_2251,N_2186);
and U10421 (N_10421,N_3823,N_2109);
xor U10422 (N_10422,N_3298,N_5828);
nor U10423 (N_10423,N_2250,N_855);
or U10424 (N_10424,N_3260,N_219);
or U10425 (N_10425,N_5366,N_4331);
and U10426 (N_10426,N_5909,N_114);
or U10427 (N_10427,N_2041,N_5810);
nor U10428 (N_10428,N_5667,N_3862);
xor U10429 (N_10429,N_413,N_1529);
xnor U10430 (N_10430,N_548,N_2557);
nor U10431 (N_10431,N_1416,N_4585);
nor U10432 (N_10432,N_2862,N_4975);
or U10433 (N_10433,N_4821,N_2026);
nand U10434 (N_10434,N_753,N_2163);
and U10435 (N_10435,N_2336,N_5542);
xnor U10436 (N_10436,N_5953,N_1126);
xor U10437 (N_10437,N_285,N_2107);
and U10438 (N_10438,N_3786,N_3876);
and U10439 (N_10439,N_3609,N_5313);
nand U10440 (N_10440,N_652,N_752);
nor U10441 (N_10441,N_3106,N_5081);
xnor U10442 (N_10442,N_1217,N_4189);
xor U10443 (N_10443,N_5532,N_1408);
or U10444 (N_10444,N_514,N_5390);
or U10445 (N_10445,N_5344,N_5987);
or U10446 (N_10446,N_298,N_5221);
or U10447 (N_10447,N_809,N_3747);
xor U10448 (N_10448,N_3940,N_3476);
or U10449 (N_10449,N_3899,N_4781);
xnor U10450 (N_10450,N_5077,N_1051);
and U10451 (N_10451,N_717,N_662);
or U10452 (N_10452,N_523,N_1994);
nand U10453 (N_10453,N_5940,N_3447);
nand U10454 (N_10454,N_1578,N_2762);
or U10455 (N_10455,N_5010,N_118);
or U10456 (N_10456,N_398,N_1561);
and U10457 (N_10457,N_3700,N_3239);
nand U10458 (N_10458,N_4630,N_816);
and U10459 (N_10459,N_4958,N_5305);
and U10460 (N_10460,N_4125,N_1396);
nor U10461 (N_10461,N_2863,N_3818);
and U10462 (N_10462,N_5887,N_5556);
nor U10463 (N_10463,N_4443,N_4411);
nor U10464 (N_10464,N_3058,N_2692);
nor U10465 (N_10465,N_4262,N_5093);
or U10466 (N_10466,N_1029,N_165);
and U10467 (N_10467,N_1294,N_1235);
xnor U10468 (N_10468,N_2197,N_5591);
xor U10469 (N_10469,N_4660,N_1257);
nand U10470 (N_10470,N_571,N_3976);
xor U10471 (N_10471,N_3385,N_2571);
xnor U10472 (N_10472,N_4709,N_884);
xor U10473 (N_10473,N_183,N_4539);
or U10474 (N_10474,N_3054,N_3917);
and U10475 (N_10475,N_2064,N_3803);
or U10476 (N_10476,N_342,N_3184);
or U10477 (N_10477,N_2629,N_1483);
and U10478 (N_10478,N_2464,N_4755);
xor U10479 (N_10479,N_4259,N_706);
or U10480 (N_10480,N_1202,N_5472);
and U10481 (N_10481,N_800,N_2501);
xnor U10482 (N_10482,N_2928,N_4740);
xor U10483 (N_10483,N_3342,N_3021);
and U10484 (N_10484,N_5414,N_19);
and U10485 (N_10485,N_4605,N_5587);
nor U10486 (N_10486,N_2711,N_809);
nor U10487 (N_10487,N_1690,N_1766);
or U10488 (N_10488,N_2468,N_690);
nor U10489 (N_10489,N_1998,N_1683);
and U10490 (N_10490,N_4480,N_47);
nor U10491 (N_10491,N_3857,N_5577);
and U10492 (N_10492,N_5072,N_711);
or U10493 (N_10493,N_2775,N_3755);
nand U10494 (N_10494,N_3811,N_2183);
and U10495 (N_10495,N_4410,N_5229);
xor U10496 (N_10496,N_2771,N_2976);
nand U10497 (N_10497,N_5519,N_3696);
or U10498 (N_10498,N_3019,N_5358);
and U10499 (N_10499,N_2726,N_2550);
or U10500 (N_10500,N_2002,N_1516);
nor U10501 (N_10501,N_4702,N_980);
xor U10502 (N_10502,N_3670,N_2875);
or U10503 (N_10503,N_813,N_5497);
xnor U10504 (N_10504,N_5789,N_976);
or U10505 (N_10505,N_51,N_5129);
and U10506 (N_10506,N_93,N_5312);
nor U10507 (N_10507,N_3214,N_252);
nand U10508 (N_10508,N_2684,N_5806);
and U10509 (N_10509,N_25,N_2650);
nor U10510 (N_10510,N_3586,N_471);
xnor U10511 (N_10511,N_3387,N_4044);
nor U10512 (N_10512,N_1656,N_1009);
and U10513 (N_10513,N_3896,N_2449);
and U10514 (N_10514,N_3551,N_5163);
xor U10515 (N_10515,N_1659,N_3185);
xor U10516 (N_10516,N_1114,N_975);
and U10517 (N_10517,N_4883,N_3641);
nand U10518 (N_10518,N_1780,N_4343);
xor U10519 (N_10519,N_1541,N_4818);
xor U10520 (N_10520,N_899,N_4061);
or U10521 (N_10521,N_3886,N_146);
nand U10522 (N_10522,N_1524,N_5539);
xor U10523 (N_10523,N_3525,N_2266);
nand U10524 (N_10524,N_4301,N_5211);
xor U10525 (N_10525,N_3465,N_3611);
xor U10526 (N_10526,N_5661,N_2533);
xnor U10527 (N_10527,N_1171,N_2848);
nand U10528 (N_10528,N_57,N_668);
or U10529 (N_10529,N_4756,N_4351);
nor U10530 (N_10530,N_2272,N_4293);
nor U10531 (N_10531,N_2548,N_5231);
xnor U10532 (N_10532,N_5489,N_3619);
nor U10533 (N_10533,N_1975,N_622);
nor U10534 (N_10534,N_5169,N_1194);
or U10535 (N_10535,N_5021,N_4493);
nand U10536 (N_10536,N_559,N_2845);
or U10537 (N_10537,N_4762,N_4076);
and U10538 (N_10538,N_4943,N_315);
or U10539 (N_10539,N_3080,N_4780);
and U10540 (N_10540,N_5612,N_2915);
nand U10541 (N_10541,N_1009,N_722);
or U10542 (N_10542,N_5298,N_2021);
or U10543 (N_10543,N_4303,N_5283);
xnor U10544 (N_10544,N_1916,N_3543);
and U10545 (N_10545,N_3442,N_4242);
or U10546 (N_10546,N_3497,N_4870);
nor U10547 (N_10547,N_4582,N_2929);
nand U10548 (N_10548,N_3767,N_4442);
or U10549 (N_10549,N_4772,N_331);
xor U10550 (N_10550,N_3828,N_3730);
nor U10551 (N_10551,N_1724,N_1351);
nor U10552 (N_10552,N_3674,N_2328);
nor U10553 (N_10553,N_1683,N_5677);
xnor U10554 (N_10554,N_2392,N_4837);
xnor U10555 (N_10555,N_1068,N_2019);
or U10556 (N_10556,N_3975,N_4999);
or U10557 (N_10557,N_3545,N_1046);
xor U10558 (N_10558,N_3355,N_3047);
xor U10559 (N_10559,N_1729,N_3914);
or U10560 (N_10560,N_5259,N_2711);
nand U10561 (N_10561,N_5621,N_2390);
nand U10562 (N_10562,N_3138,N_5780);
nand U10563 (N_10563,N_4396,N_1953);
nor U10564 (N_10564,N_3005,N_2042);
or U10565 (N_10565,N_1634,N_473);
and U10566 (N_10566,N_3700,N_4589);
or U10567 (N_10567,N_172,N_667);
and U10568 (N_10568,N_3397,N_5472);
xor U10569 (N_10569,N_5453,N_5736);
xor U10570 (N_10570,N_184,N_1990);
xor U10571 (N_10571,N_5188,N_1499);
nor U10572 (N_10572,N_2627,N_4880);
nand U10573 (N_10573,N_401,N_2345);
and U10574 (N_10574,N_2507,N_3503);
and U10575 (N_10575,N_3717,N_3016);
xor U10576 (N_10576,N_1056,N_4911);
nor U10577 (N_10577,N_3662,N_3294);
nand U10578 (N_10578,N_3944,N_3846);
or U10579 (N_10579,N_5010,N_1816);
nand U10580 (N_10580,N_3693,N_3449);
xor U10581 (N_10581,N_127,N_5097);
and U10582 (N_10582,N_3858,N_4452);
or U10583 (N_10583,N_5806,N_764);
nor U10584 (N_10584,N_2124,N_4512);
nand U10585 (N_10585,N_5245,N_3359);
and U10586 (N_10586,N_1048,N_4961);
and U10587 (N_10587,N_1862,N_4697);
nor U10588 (N_10588,N_43,N_218);
nor U10589 (N_10589,N_1972,N_4710);
nor U10590 (N_10590,N_349,N_815);
and U10591 (N_10591,N_1755,N_3907);
or U10592 (N_10592,N_2734,N_132);
or U10593 (N_10593,N_3086,N_5357);
or U10594 (N_10594,N_3751,N_239);
nor U10595 (N_10595,N_3134,N_5984);
or U10596 (N_10596,N_1610,N_1904);
nor U10597 (N_10597,N_4011,N_4951);
and U10598 (N_10598,N_4684,N_4012);
or U10599 (N_10599,N_3401,N_596);
xor U10600 (N_10600,N_94,N_2291);
nand U10601 (N_10601,N_5784,N_3139);
xnor U10602 (N_10602,N_5936,N_5644);
xor U10603 (N_10603,N_1697,N_5277);
or U10604 (N_10604,N_3155,N_4442);
nand U10605 (N_10605,N_3371,N_5809);
and U10606 (N_10606,N_1960,N_1200);
xor U10607 (N_10607,N_379,N_80);
xnor U10608 (N_10608,N_2705,N_3042);
and U10609 (N_10609,N_4772,N_3016);
or U10610 (N_10610,N_1232,N_378);
or U10611 (N_10611,N_2390,N_75);
or U10612 (N_10612,N_702,N_2691);
and U10613 (N_10613,N_2089,N_4337);
nand U10614 (N_10614,N_3169,N_4086);
and U10615 (N_10615,N_944,N_365);
xnor U10616 (N_10616,N_5149,N_496);
or U10617 (N_10617,N_137,N_2131);
xnor U10618 (N_10618,N_3269,N_3364);
or U10619 (N_10619,N_366,N_941);
nor U10620 (N_10620,N_3903,N_902);
nand U10621 (N_10621,N_262,N_3886);
xor U10622 (N_10622,N_2712,N_5555);
nand U10623 (N_10623,N_4732,N_5762);
and U10624 (N_10624,N_3269,N_5595);
and U10625 (N_10625,N_904,N_881);
xor U10626 (N_10626,N_4418,N_5700);
and U10627 (N_10627,N_1422,N_5542);
xor U10628 (N_10628,N_1366,N_1389);
nor U10629 (N_10629,N_3222,N_4886);
or U10630 (N_10630,N_4294,N_175);
nand U10631 (N_10631,N_5376,N_2275);
or U10632 (N_10632,N_4177,N_5119);
and U10633 (N_10633,N_316,N_4921);
nand U10634 (N_10634,N_146,N_5224);
xor U10635 (N_10635,N_2445,N_5013);
nor U10636 (N_10636,N_3152,N_2085);
or U10637 (N_10637,N_4725,N_4372);
nor U10638 (N_10638,N_2513,N_604);
and U10639 (N_10639,N_4256,N_4015);
xnor U10640 (N_10640,N_62,N_380);
or U10641 (N_10641,N_411,N_5980);
and U10642 (N_10642,N_4828,N_2330);
or U10643 (N_10643,N_5213,N_740);
or U10644 (N_10644,N_2499,N_2836);
nand U10645 (N_10645,N_5483,N_1245);
nand U10646 (N_10646,N_4580,N_4847);
xnor U10647 (N_10647,N_1412,N_4848);
or U10648 (N_10648,N_4514,N_2032);
xor U10649 (N_10649,N_4741,N_1838);
or U10650 (N_10650,N_5284,N_2728);
nor U10651 (N_10651,N_1909,N_2602);
xnor U10652 (N_10652,N_8,N_5683);
nor U10653 (N_10653,N_4355,N_5133);
xor U10654 (N_10654,N_5345,N_2499);
nor U10655 (N_10655,N_2227,N_703);
and U10656 (N_10656,N_5046,N_1291);
or U10657 (N_10657,N_247,N_2802);
nand U10658 (N_10658,N_1475,N_3262);
nor U10659 (N_10659,N_2861,N_1630);
nor U10660 (N_10660,N_3642,N_3077);
nand U10661 (N_10661,N_5380,N_998);
xor U10662 (N_10662,N_4567,N_3056);
nand U10663 (N_10663,N_47,N_4988);
xnor U10664 (N_10664,N_463,N_3381);
or U10665 (N_10665,N_1521,N_2864);
nor U10666 (N_10666,N_5188,N_1942);
nor U10667 (N_10667,N_115,N_4871);
nand U10668 (N_10668,N_1357,N_471);
or U10669 (N_10669,N_5673,N_1012);
nand U10670 (N_10670,N_3128,N_3645);
xnor U10671 (N_10671,N_4108,N_3602);
or U10672 (N_10672,N_298,N_4387);
or U10673 (N_10673,N_1979,N_3257);
and U10674 (N_10674,N_4992,N_4943);
nor U10675 (N_10675,N_4612,N_2774);
nor U10676 (N_10676,N_5227,N_2690);
and U10677 (N_10677,N_5785,N_4630);
or U10678 (N_10678,N_2426,N_3580);
and U10679 (N_10679,N_4782,N_375);
or U10680 (N_10680,N_417,N_4170);
or U10681 (N_10681,N_4709,N_3889);
and U10682 (N_10682,N_2039,N_3301);
nand U10683 (N_10683,N_842,N_5127);
and U10684 (N_10684,N_2822,N_3991);
or U10685 (N_10685,N_4571,N_3693);
xnor U10686 (N_10686,N_3984,N_3472);
and U10687 (N_10687,N_663,N_4423);
nor U10688 (N_10688,N_1828,N_5183);
xor U10689 (N_10689,N_5525,N_2317);
and U10690 (N_10690,N_5995,N_3232);
nand U10691 (N_10691,N_2227,N_4979);
or U10692 (N_10692,N_569,N_771);
or U10693 (N_10693,N_1687,N_3059);
and U10694 (N_10694,N_5661,N_3046);
or U10695 (N_10695,N_1823,N_4167);
and U10696 (N_10696,N_1896,N_129);
nand U10697 (N_10697,N_5028,N_1901);
nor U10698 (N_10698,N_4573,N_5826);
nor U10699 (N_10699,N_153,N_5644);
nand U10700 (N_10700,N_86,N_3317);
xnor U10701 (N_10701,N_2327,N_5044);
nand U10702 (N_10702,N_549,N_5884);
and U10703 (N_10703,N_748,N_582);
xnor U10704 (N_10704,N_140,N_5111);
and U10705 (N_10705,N_3742,N_1676);
nor U10706 (N_10706,N_3941,N_3043);
and U10707 (N_10707,N_5365,N_4854);
or U10708 (N_10708,N_5964,N_5205);
or U10709 (N_10709,N_1380,N_2762);
xor U10710 (N_10710,N_1450,N_401);
and U10711 (N_10711,N_87,N_2500);
nor U10712 (N_10712,N_1070,N_3388);
nand U10713 (N_10713,N_816,N_5904);
nand U10714 (N_10714,N_1143,N_2283);
or U10715 (N_10715,N_5114,N_3671);
nand U10716 (N_10716,N_4827,N_3484);
nand U10717 (N_10717,N_3113,N_5271);
or U10718 (N_10718,N_3804,N_1762);
xnor U10719 (N_10719,N_3617,N_210);
xor U10720 (N_10720,N_4240,N_926);
xnor U10721 (N_10721,N_3484,N_2611);
xnor U10722 (N_10722,N_2114,N_5073);
nand U10723 (N_10723,N_1367,N_1266);
xnor U10724 (N_10724,N_2153,N_4439);
or U10725 (N_10725,N_1072,N_3508);
xor U10726 (N_10726,N_5963,N_2882);
or U10727 (N_10727,N_4842,N_4788);
nor U10728 (N_10728,N_4671,N_5704);
nor U10729 (N_10729,N_3546,N_3767);
and U10730 (N_10730,N_1391,N_4624);
or U10731 (N_10731,N_1563,N_515);
xnor U10732 (N_10732,N_813,N_1603);
and U10733 (N_10733,N_3508,N_2082);
or U10734 (N_10734,N_1082,N_2132);
or U10735 (N_10735,N_4631,N_2672);
nor U10736 (N_10736,N_4761,N_5894);
xor U10737 (N_10737,N_5350,N_2268);
or U10738 (N_10738,N_1693,N_1147);
and U10739 (N_10739,N_47,N_4446);
and U10740 (N_10740,N_1085,N_2244);
xnor U10741 (N_10741,N_4768,N_3513);
or U10742 (N_10742,N_470,N_4200);
nand U10743 (N_10743,N_707,N_5905);
xnor U10744 (N_10744,N_1430,N_2121);
or U10745 (N_10745,N_1502,N_1435);
nor U10746 (N_10746,N_1990,N_5811);
nor U10747 (N_10747,N_1568,N_1886);
nand U10748 (N_10748,N_203,N_324);
and U10749 (N_10749,N_4283,N_3512);
nor U10750 (N_10750,N_932,N_1818);
nor U10751 (N_10751,N_1685,N_5048);
and U10752 (N_10752,N_1550,N_4892);
or U10753 (N_10753,N_5347,N_5915);
nand U10754 (N_10754,N_4577,N_5855);
xor U10755 (N_10755,N_1503,N_265);
and U10756 (N_10756,N_1381,N_1266);
or U10757 (N_10757,N_1799,N_686);
or U10758 (N_10758,N_3110,N_2840);
xnor U10759 (N_10759,N_291,N_1787);
and U10760 (N_10760,N_2863,N_4325);
and U10761 (N_10761,N_4988,N_3961);
xnor U10762 (N_10762,N_2059,N_1189);
and U10763 (N_10763,N_3836,N_4342);
nor U10764 (N_10764,N_248,N_3576);
nand U10765 (N_10765,N_4725,N_4822);
nor U10766 (N_10766,N_5054,N_1160);
xnor U10767 (N_10767,N_290,N_5566);
or U10768 (N_10768,N_3406,N_784);
nor U10769 (N_10769,N_4858,N_5597);
and U10770 (N_10770,N_5663,N_1270);
or U10771 (N_10771,N_3864,N_4728);
nand U10772 (N_10772,N_5331,N_1465);
or U10773 (N_10773,N_4047,N_2588);
nor U10774 (N_10774,N_5494,N_1816);
or U10775 (N_10775,N_4273,N_3630);
xnor U10776 (N_10776,N_4380,N_1306);
and U10777 (N_10777,N_2947,N_5043);
and U10778 (N_10778,N_4065,N_4064);
or U10779 (N_10779,N_4214,N_1558);
or U10780 (N_10780,N_4178,N_5511);
and U10781 (N_10781,N_5659,N_3148);
and U10782 (N_10782,N_2042,N_1209);
xor U10783 (N_10783,N_1301,N_2443);
nor U10784 (N_10784,N_2040,N_2327);
and U10785 (N_10785,N_1986,N_1940);
or U10786 (N_10786,N_448,N_625);
nand U10787 (N_10787,N_4316,N_634);
and U10788 (N_10788,N_981,N_2124);
nand U10789 (N_10789,N_3297,N_765);
nand U10790 (N_10790,N_2642,N_5270);
and U10791 (N_10791,N_4980,N_5198);
nand U10792 (N_10792,N_3951,N_534);
or U10793 (N_10793,N_4147,N_4049);
nand U10794 (N_10794,N_784,N_788);
or U10795 (N_10795,N_4514,N_1852);
xnor U10796 (N_10796,N_1137,N_834);
nand U10797 (N_10797,N_2550,N_3288);
or U10798 (N_10798,N_970,N_625);
or U10799 (N_10799,N_1899,N_1263);
or U10800 (N_10800,N_303,N_5325);
nor U10801 (N_10801,N_5043,N_2824);
and U10802 (N_10802,N_5026,N_2383);
and U10803 (N_10803,N_4967,N_424);
or U10804 (N_10804,N_4223,N_771);
nor U10805 (N_10805,N_1027,N_3917);
nand U10806 (N_10806,N_118,N_618);
nand U10807 (N_10807,N_5081,N_1526);
and U10808 (N_10808,N_3035,N_2089);
nor U10809 (N_10809,N_1495,N_2690);
or U10810 (N_10810,N_5511,N_3080);
or U10811 (N_10811,N_2039,N_5932);
or U10812 (N_10812,N_2820,N_2766);
nor U10813 (N_10813,N_832,N_2933);
nand U10814 (N_10814,N_3789,N_5763);
or U10815 (N_10815,N_4762,N_636);
nand U10816 (N_10816,N_1224,N_1273);
xnor U10817 (N_10817,N_1647,N_1271);
or U10818 (N_10818,N_4365,N_5156);
nand U10819 (N_10819,N_5831,N_2794);
and U10820 (N_10820,N_2938,N_4291);
and U10821 (N_10821,N_4168,N_5335);
and U10822 (N_10822,N_2605,N_3996);
or U10823 (N_10823,N_984,N_784);
nand U10824 (N_10824,N_4537,N_1621);
nor U10825 (N_10825,N_503,N_5742);
nand U10826 (N_10826,N_349,N_915);
and U10827 (N_10827,N_5180,N_5856);
nor U10828 (N_10828,N_1386,N_210);
or U10829 (N_10829,N_3792,N_1446);
nand U10830 (N_10830,N_2107,N_2709);
and U10831 (N_10831,N_1830,N_5176);
nand U10832 (N_10832,N_2026,N_436);
nand U10833 (N_10833,N_1323,N_398);
nand U10834 (N_10834,N_4439,N_3035);
xnor U10835 (N_10835,N_1298,N_4708);
and U10836 (N_10836,N_185,N_5734);
nor U10837 (N_10837,N_1865,N_183);
xnor U10838 (N_10838,N_5359,N_4387);
nand U10839 (N_10839,N_1347,N_5064);
nand U10840 (N_10840,N_5660,N_3581);
or U10841 (N_10841,N_3017,N_875);
nor U10842 (N_10842,N_5575,N_4817);
nand U10843 (N_10843,N_3917,N_923);
and U10844 (N_10844,N_1040,N_3642);
and U10845 (N_10845,N_4111,N_2258);
xor U10846 (N_10846,N_4300,N_2177);
xnor U10847 (N_10847,N_4424,N_1933);
nor U10848 (N_10848,N_471,N_5235);
and U10849 (N_10849,N_4421,N_3990);
xnor U10850 (N_10850,N_5920,N_167);
nand U10851 (N_10851,N_4375,N_3306);
nor U10852 (N_10852,N_2955,N_468);
or U10853 (N_10853,N_4551,N_2452);
xor U10854 (N_10854,N_4699,N_3895);
nor U10855 (N_10855,N_5050,N_2034);
nand U10856 (N_10856,N_1491,N_3759);
nor U10857 (N_10857,N_3122,N_3541);
xor U10858 (N_10858,N_1762,N_5610);
or U10859 (N_10859,N_863,N_2959);
and U10860 (N_10860,N_4038,N_5450);
and U10861 (N_10861,N_3643,N_3936);
nor U10862 (N_10862,N_2513,N_1760);
xor U10863 (N_10863,N_3527,N_4701);
nor U10864 (N_10864,N_5053,N_1504);
xnor U10865 (N_10865,N_518,N_3610);
nor U10866 (N_10866,N_2298,N_1430);
and U10867 (N_10867,N_660,N_1899);
xor U10868 (N_10868,N_1573,N_1286);
nor U10869 (N_10869,N_3448,N_4367);
and U10870 (N_10870,N_472,N_348);
and U10871 (N_10871,N_323,N_5897);
nor U10872 (N_10872,N_5861,N_2953);
or U10873 (N_10873,N_3705,N_3783);
xor U10874 (N_10874,N_1735,N_891);
or U10875 (N_10875,N_3904,N_2391);
and U10876 (N_10876,N_240,N_2814);
xnor U10877 (N_10877,N_5178,N_414);
nor U10878 (N_10878,N_2797,N_4519);
and U10879 (N_10879,N_2499,N_567);
and U10880 (N_10880,N_4651,N_3079);
or U10881 (N_10881,N_2143,N_2865);
nand U10882 (N_10882,N_5910,N_1111);
nor U10883 (N_10883,N_1839,N_2464);
or U10884 (N_10884,N_5127,N_2670);
or U10885 (N_10885,N_1292,N_3015);
nand U10886 (N_10886,N_5236,N_4503);
nor U10887 (N_10887,N_3216,N_281);
and U10888 (N_10888,N_2377,N_4209);
or U10889 (N_10889,N_3226,N_1833);
or U10890 (N_10890,N_5835,N_4123);
nor U10891 (N_10891,N_4282,N_3504);
nor U10892 (N_10892,N_2822,N_3982);
or U10893 (N_10893,N_4403,N_558);
or U10894 (N_10894,N_176,N_4939);
xnor U10895 (N_10895,N_2164,N_946);
nor U10896 (N_10896,N_1720,N_3253);
xnor U10897 (N_10897,N_5717,N_781);
nand U10898 (N_10898,N_665,N_989);
or U10899 (N_10899,N_3129,N_4914);
nand U10900 (N_10900,N_2965,N_2715);
xnor U10901 (N_10901,N_5424,N_64);
nor U10902 (N_10902,N_4571,N_1733);
nor U10903 (N_10903,N_3322,N_3834);
nand U10904 (N_10904,N_2149,N_5284);
nand U10905 (N_10905,N_369,N_3528);
or U10906 (N_10906,N_4007,N_3128);
nor U10907 (N_10907,N_3611,N_259);
nor U10908 (N_10908,N_971,N_2890);
and U10909 (N_10909,N_597,N_2067);
and U10910 (N_10910,N_660,N_1911);
nor U10911 (N_10911,N_5570,N_2540);
xnor U10912 (N_10912,N_720,N_2880);
nand U10913 (N_10913,N_4679,N_382);
nand U10914 (N_10914,N_3881,N_2784);
nand U10915 (N_10915,N_2459,N_1058);
nand U10916 (N_10916,N_4025,N_2761);
xnor U10917 (N_10917,N_2698,N_5189);
and U10918 (N_10918,N_3621,N_4841);
nor U10919 (N_10919,N_2793,N_5590);
and U10920 (N_10920,N_2298,N_2728);
and U10921 (N_10921,N_503,N_343);
nand U10922 (N_10922,N_4351,N_1916);
xor U10923 (N_10923,N_1917,N_3415);
and U10924 (N_10924,N_5309,N_422);
or U10925 (N_10925,N_2493,N_2231);
nand U10926 (N_10926,N_84,N_5241);
xnor U10927 (N_10927,N_1920,N_5280);
or U10928 (N_10928,N_3189,N_504);
and U10929 (N_10929,N_4339,N_1532);
or U10930 (N_10930,N_386,N_3974);
nor U10931 (N_10931,N_280,N_5914);
and U10932 (N_10932,N_110,N_1125);
xor U10933 (N_10933,N_5268,N_4813);
nor U10934 (N_10934,N_4762,N_2275);
nor U10935 (N_10935,N_1480,N_4580);
and U10936 (N_10936,N_3544,N_2275);
nor U10937 (N_10937,N_2376,N_1862);
nand U10938 (N_10938,N_3843,N_194);
nor U10939 (N_10939,N_5529,N_805);
or U10940 (N_10940,N_1644,N_240);
or U10941 (N_10941,N_133,N_1258);
nand U10942 (N_10942,N_3227,N_5126);
and U10943 (N_10943,N_4592,N_44);
or U10944 (N_10944,N_3904,N_4041);
or U10945 (N_10945,N_5803,N_1096);
xor U10946 (N_10946,N_1384,N_7);
xnor U10947 (N_10947,N_453,N_1648);
and U10948 (N_10948,N_5108,N_1524);
nand U10949 (N_10949,N_3100,N_3726);
and U10950 (N_10950,N_4278,N_1752);
nand U10951 (N_10951,N_436,N_5022);
or U10952 (N_10952,N_4139,N_5988);
or U10953 (N_10953,N_110,N_408);
nand U10954 (N_10954,N_3412,N_3409);
or U10955 (N_10955,N_4356,N_2170);
xor U10956 (N_10956,N_759,N_5396);
xor U10957 (N_10957,N_2731,N_1397);
nor U10958 (N_10958,N_1551,N_4943);
or U10959 (N_10959,N_5221,N_4849);
or U10960 (N_10960,N_1020,N_1516);
xnor U10961 (N_10961,N_5936,N_1659);
nor U10962 (N_10962,N_4426,N_5251);
xor U10963 (N_10963,N_1839,N_527);
nor U10964 (N_10964,N_4236,N_5169);
nor U10965 (N_10965,N_4989,N_2333);
or U10966 (N_10966,N_1284,N_4493);
and U10967 (N_10967,N_5774,N_5227);
nand U10968 (N_10968,N_2379,N_4026);
nor U10969 (N_10969,N_1935,N_3129);
and U10970 (N_10970,N_2091,N_4129);
xnor U10971 (N_10971,N_1457,N_5607);
xor U10972 (N_10972,N_2440,N_5841);
or U10973 (N_10973,N_44,N_3873);
xnor U10974 (N_10974,N_3408,N_1576);
xnor U10975 (N_10975,N_2198,N_4263);
and U10976 (N_10976,N_159,N_5347);
nor U10977 (N_10977,N_1869,N_1082);
nand U10978 (N_10978,N_954,N_4421);
xor U10979 (N_10979,N_3153,N_4236);
nand U10980 (N_10980,N_2103,N_1033);
and U10981 (N_10981,N_2853,N_593);
nor U10982 (N_10982,N_3987,N_8);
or U10983 (N_10983,N_3089,N_5229);
nand U10984 (N_10984,N_5067,N_5193);
xnor U10985 (N_10985,N_260,N_3696);
and U10986 (N_10986,N_5069,N_489);
and U10987 (N_10987,N_2100,N_2012);
or U10988 (N_10988,N_4846,N_4171);
nand U10989 (N_10989,N_1263,N_1550);
or U10990 (N_10990,N_5884,N_1288);
xnor U10991 (N_10991,N_1263,N_5004);
and U10992 (N_10992,N_3729,N_3174);
nor U10993 (N_10993,N_1752,N_5189);
xnor U10994 (N_10994,N_5311,N_5401);
and U10995 (N_10995,N_278,N_2243);
and U10996 (N_10996,N_2232,N_5419);
nor U10997 (N_10997,N_1483,N_5418);
and U10998 (N_10998,N_5299,N_2417);
xnor U10999 (N_10999,N_3720,N_4486);
nand U11000 (N_11000,N_1246,N_4333);
nand U11001 (N_11001,N_135,N_5999);
or U11002 (N_11002,N_1127,N_4258);
nor U11003 (N_11003,N_5766,N_97);
and U11004 (N_11004,N_4252,N_1325);
nor U11005 (N_11005,N_5096,N_1803);
nor U11006 (N_11006,N_377,N_1964);
nor U11007 (N_11007,N_800,N_1719);
xor U11008 (N_11008,N_1388,N_73);
or U11009 (N_11009,N_271,N_3293);
xor U11010 (N_11010,N_3848,N_205);
and U11011 (N_11011,N_3132,N_146);
xor U11012 (N_11012,N_1795,N_766);
and U11013 (N_11013,N_539,N_511);
and U11014 (N_11014,N_3351,N_3944);
and U11015 (N_11015,N_5528,N_1314);
nand U11016 (N_11016,N_4378,N_3060);
and U11017 (N_11017,N_2520,N_1743);
and U11018 (N_11018,N_4927,N_4519);
nand U11019 (N_11019,N_249,N_2796);
or U11020 (N_11020,N_3709,N_1851);
or U11021 (N_11021,N_3850,N_5174);
or U11022 (N_11022,N_995,N_3790);
nor U11023 (N_11023,N_3229,N_5011);
and U11024 (N_11024,N_2350,N_3262);
or U11025 (N_11025,N_2958,N_1370);
and U11026 (N_11026,N_3737,N_2359);
xor U11027 (N_11027,N_5021,N_2012);
xor U11028 (N_11028,N_3782,N_3441);
and U11029 (N_11029,N_5004,N_4142);
and U11030 (N_11030,N_665,N_3076);
nand U11031 (N_11031,N_3482,N_5358);
xor U11032 (N_11032,N_5909,N_4520);
nand U11033 (N_11033,N_2783,N_545);
nand U11034 (N_11034,N_1839,N_1400);
nand U11035 (N_11035,N_56,N_61);
xor U11036 (N_11036,N_5803,N_5936);
xnor U11037 (N_11037,N_5752,N_982);
nor U11038 (N_11038,N_5611,N_1191);
and U11039 (N_11039,N_1413,N_741);
nor U11040 (N_11040,N_3275,N_5424);
nand U11041 (N_11041,N_3208,N_541);
xnor U11042 (N_11042,N_4080,N_3332);
or U11043 (N_11043,N_3276,N_1626);
or U11044 (N_11044,N_5500,N_4296);
xnor U11045 (N_11045,N_23,N_2621);
nand U11046 (N_11046,N_528,N_3708);
xnor U11047 (N_11047,N_430,N_3161);
and U11048 (N_11048,N_4747,N_981);
or U11049 (N_11049,N_3255,N_971);
and U11050 (N_11050,N_815,N_1189);
nand U11051 (N_11051,N_1433,N_5952);
nand U11052 (N_11052,N_4009,N_4700);
xnor U11053 (N_11053,N_150,N_2155);
xnor U11054 (N_11054,N_2071,N_5020);
nand U11055 (N_11055,N_764,N_769);
nor U11056 (N_11056,N_3115,N_72);
nor U11057 (N_11057,N_1147,N_180);
nand U11058 (N_11058,N_4119,N_5897);
or U11059 (N_11059,N_2830,N_1658);
xnor U11060 (N_11060,N_435,N_420);
xor U11061 (N_11061,N_5318,N_1123);
xor U11062 (N_11062,N_5762,N_359);
or U11063 (N_11063,N_5041,N_5742);
nand U11064 (N_11064,N_4605,N_2321);
nand U11065 (N_11065,N_4924,N_4469);
nand U11066 (N_11066,N_506,N_4157);
xor U11067 (N_11067,N_3260,N_5154);
nor U11068 (N_11068,N_4555,N_3716);
nor U11069 (N_11069,N_3301,N_3425);
xnor U11070 (N_11070,N_5553,N_1016);
nor U11071 (N_11071,N_1611,N_3814);
and U11072 (N_11072,N_5642,N_4805);
nor U11073 (N_11073,N_1434,N_5676);
or U11074 (N_11074,N_2826,N_1827);
or U11075 (N_11075,N_1258,N_82);
or U11076 (N_11076,N_3976,N_5060);
or U11077 (N_11077,N_5844,N_1705);
nor U11078 (N_11078,N_5135,N_4326);
or U11079 (N_11079,N_2958,N_1224);
and U11080 (N_11080,N_3883,N_496);
or U11081 (N_11081,N_1192,N_4085);
nor U11082 (N_11082,N_4585,N_1632);
nor U11083 (N_11083,N_2391,N_3657);
and U11084 (N_11084,N_4994,N_3298);
nor U11085 (N_11085,N_3659,N_1440);
and U11086 (N_11086,N_4627,N_4428);
nor U11087 (N_11087,N_664,N_5680);
nand U11088 (N_11088,N_4190,N_2634);
and U11089 (N_11089,N_3731,N_471);
xnor U11090 (N_11090,N_5452,N_2919);
and U11091 (N_11091,N_5491,N_3145);
and U11092 (N_11092,N_2972,N_4039);
nor U11093 (N_11093,N_176,N_3360);
nor U11094 (N_11094,N_1726,N_5526);
nor U11095 (N_11095,N_5068,N_2074);
nor U11096 (N_11096,N_5820,N_2873);
nor U11097 (N_11097,N_2271,N_2855);
nor U11098 (N_11098,N_1526,N_3845);
xnor U11099 (N_11099,N_4467,N_5858);
and U11100 (N_11100,N_5621,N_5324);
nand U11101 (N_11101,N_408,N_295);
nor U11102 (N_11102,N_782,N_2583);
or U11103 (N_11103,N_862,N_834);
xor U11104 (N_11104,N_1457,N_2235);
nor U11105 (N_11105,N_1876,N_4293);
and U11106 (N_11106,N_62,N_1575);
and U11107 (N_11107,N_223,N_3721);
and U11108 (N_11108,N_4781,N_4832);
xnor U11109 (N_11109,N_4118,N_4028);
nor U11110 (N_11110,N_1364,N_5478);
and U11111 (N_11111,N_2834,N_102);
xor U11112 (N_11112,N_3916,N_2331);
xor U11113 (N_11113,N_805,N_2426);
nor U11114 (N_11114,N_3675,N_4210);
or U11115 (N_11115,N_3649,N_1515);
xnor U11116 (N_11116,N_4656,N_2014);
and U11117 (N_11117,N_4726,N_3527);
nor U11118 (N_11118,N_491,N_93);
xor U11119 (N_11119,N_94,N_1728);
nand U11120 (N_11120,N_2140,N_3063);
nand U11121 (N_11121,N_90,N_3872);
xnor U11122 (N_11122,N_4899,N_310);
xor U11123 (N_11123,N_5489,N_1709);
or U11124 (N_11124,N_4716,N_1432);
or U11125 (N_11125,N_2618,N_424);
and U11126 (N_11126,N_4614,N_5660);
nand U11127 (N_11127,N_4406,N_5242);
nand U11128 (N_11128,N_2886,N_2204);
nor U11129 (N_11129,N_2247,N_426);
nor U11130 (N_11130,N_3435,N_130);
and U11131 (N_11131,N_2550,N_5181);
nor U11132 (N_11132,N_4943,N_4524);
or U11133 (N_11133,N_1164,N_4547);
nand U11134 (N_11134,N_5600,N_3243);
xnor U11135 (N_11135,N_1703,N_1217);
and U11136 (N_11136,N_2638,N_3933);
and U11137 (N_11137,N_4334,N_2585);
xnor U11138 (N_11138,N_5182,N_3653);
nor U11139 (N_11139,N_1690,N_1944);
xor U11140 (N_11140,N_3785,N_1485);
or U11141 (N_11141,N_5995,N_2489);
nand U11142 (N_11142,N_5219,N_3203);
nand U11143 (N_11143,N_425,N_1755);
xnor U11144 (N_11144,N_5911,N_4919);
and U11145 (N_11145,N_5763,N_3142);
and U11146 (N_11146,N_2283,N_1382);
and U11147 (N_11147,N_3984,N_4659);
xor U11148 (N_11148,N_3692,N_1697);
xor U11149 (N_11149,N_790,N_5702);
nand U11150 (N_11150,N_4414,N_5489);
or U11151 (N_11151,N_4061,N_4920);
nand U11152 (N_11152,N_2771,N_4152);
and U11153 (N_11153,N_845,N_3104);
xor U11154 (N_11154,N_1883,N_245);
or U11155 (N_11155,N_5661,N_1545);
nand U11156 (N_11156,N_3421,N_5303);
nand U11157 (N_11157,N_5122,N_3110);
or U11158 (N_11158,N_1007,N_2467);
or U11159 (N_11159,N_5640,N_2786);
xnor U11160 (N_11160,N_5882,N_2883);
or U11161 (N_11161,N_1572,N_5558);
nand U11162 (N_11162,N_4063,N_3779);
xnor U11163 (N_11163,N_841,N_3902);
or U11164 (N_11164,N_5781,N_3752);
nand U11165 (N_11165,N_4735,N_710);
and U11166 (N_11166,N_4544,N_109);
nand U11167 (N_11167,N_1310,N_4243);
nor U11168 (N_11168,N_4609,N_2392);
nand U11169 (N_11169,N_55,N_4966);
and U11170 (N_11170,N_1547,N_1664);
nand U11171 (N_11171,N_2359,N_906);
or U11172 (N_11172,N_2289,N_5392);
xor U11173 (N_11173,N_4128,N_3768);
nor U11174 (N_11174,N_2513,N_2375);
or U11175 (N_11175,N_2977,N_2954);
xnor U11176 (N_11176,N_2135,N_191);
nand U11177 (N_11177,N_5315,N_3548);
xnor U11178 (N_11178,N_1223,N_3927);
and U11179 (N_11179,N_4882,N_5223);
nand U11180 (N_11180,N_1065,N_5698);
nor U11181 (N_11181,N_3869,N_1400);
nand U11182 (N_11182,N_1828,N_2374);
or U11183 (N_11183,N_2723,N_3296);
nor U11184 (N_11184,N_1512,N_2991);
and U11185 (N_11185,N_394,N_1720);
nor U11186 (N_11186,N_1803,N_5284);
xnor U11187 (N_11187,N_4056,N_823);
or U11188 (N_11188,N_3607,N_2608);
and U11189 (N_11189,N_413,N_3365);
or U11190 (N_11190,N_1538,N_4991);
nand U11191 (N_11191,N_1474,N_4971);
and U11192 (N_11192,N_3248,N_5642);
xor U11193 (N_11193,N_4702,N_2690);
and U11194 (N_11194,N_1222,N_3027);
or U11195 (N_11195,N_3608,N_2226);
or U11196 (N_11196,N_5734,N_3633);
or U11197 (N_11197,N_2647,N_444);
nor U11198 (N_11198,N_4325,N_5038);
nand U11199 (N_11199,N_2712,N_1926);
nand U11200 (N_11200,N_3837,N_1227);
xnor U11201 (N_11201,N_2626,N_1358);
or U11202 (N_11202,N_5816,N_3736);
nand U11203 (N_11203,N_534,N_1552);
nor U11204 (N_11204,N_3188,N_3658);
xor U11205 (N_11205,N_187,N_4984);
or U11206 (N_11206,N_2530,N_740);
xnor U11207 (N_11207,N_2022,N_4876);
xnor U11208 (N_11208,N_3426,N_3230);
and U11209 (N_11209,N_1557,N_4403);
xnor U11210 (N_11210,N_2229,N_5315);
nand U11211 (N_11211,N_5429,N_1656);
nand U11212 (N_11212,N_2170,N_5340);
nor U11213 (N_11213,N_2137,N_2408);
xnor U11214 (N_11214,N_2033,N_797);
nand U11215 (N_11215,N_3919,N_1459);
and U11216 (N_11216,N_5203,N_2530);
nand U11217 (N_11217,N_1720,N_1874);
nand U11218 (N_11218,N_4909,N_4180);
xnor U11219 (N_11219,N_3351,N_2151);
xor U11220 (N_11220,N_1245,N_4488);
xnor U11221 (N_11221,N_1717,N_1521);
nor U11222 (N_11222,N_3440,N_4674);
nor U11223 (N_11223,N_5652,N_2048);
xor U11224 (N_11224,N_4670,N_5325);
or U11225 (N_11225,N_2985,N_5600);
nor U11226 (N_11226,N_510,N_1863);
and U11227 (N_11227,N_5790,N_3831);
and U11228 (N_11228,N_246,N_5898);
and U11229 (N_11229,N_2011,N_1609);
and U11230 (N_11230,N_3799,N_4378);
xnor U11231 (N_11231,N_3452,N_1193);
nand U11232 (N_11232,N_1244,N_2346);
nor U11233 (N_11233,N_4915,N_2888);
xor U11234 (N_11234,N_5802,N_508);
xor U11235 (N_11235,N_3039,N_1953);
nor U11236 (N_11236,N_5826,N_2022);
or U11237 (N_11237,N_222,N_519);
xnor U11238 (N_11238,N_4348,N_1521);
xnor U11239 (N_11239,N_2386,N_5615);
nand U11240 (N_11240,N_1541,N_4308);
or U11241 (N_11241,N_1738,N_3758);
and U11242 (N_11242,N_4993,N_1624);
and U11243 (N_11243,N_4059,N_5822);
xnor U11244 (N_11244,N_5410,N_5890);
and U11245 (N_11245,N_327,N_2030);
or U11246 (N_11246,N_1560,N_2965);
and U11247 (N_11247,N_2019,N_1600);
nor U11248 (N_11248,N_4068,N_4325);
nand U11249 (N_11249,N_2539,N_4807);
xnor U11250 (N_11250,N_4755,N_4403);
xor U11251 (N_11251,N_751,N_3255);
nor U11252 (N_11252,N_4754,N_4312);
or U11253 (N_11253,N_3152,N_691);
xnor U11254 (N_11254,N_655,N_3755);
or U11255 (N_11255,N_5134,N_3934);
xnor U11256 (N_11256,N_1101,N_1565);
nor U11257 (N_11257,N_4939,N_1342);
and U11258 (N_11258,N_2350,N_152);
nor U11259 (N_11259,N_1163,N_5283);
or U11260 (N_11260,N_4268,N_3003);
or U11261 (N_11261,N_2356,N_926);
nand U11262 (N_11262,N_1689,N_4482);
or U11263 (N_11263,N_1750,N_3586);
or U11264 (N_11264,N_4810,N_4114);
xnor U11265 (N_11265,N_794,N_4029);
nand U11266 (N_11266,N_594,N_1590);
and U11267 (N_11267,N_1188,N_5996);
xnor U11268 (N_11268,N_69,N_1672);
nand U11269 (N_11269,N_4207,N_1390);
xnor U11270 (N_11270,N_748,N_5399);
and U11271 (N_11271,N_3237,N_5671);
or U11272 (N_11272,N_840,N_5947);
and U11273 (N_11273,N_1236,N_3747);
or U11274 (N_11274,N_225,N_4717);
xnor U11275 (N_11275,N_796,N_2226);
nand U11276 (N_11276,N_3874,N_3387);
xor U11277 (N_11277,N_4815,N_3916);
and U11278 (N_11278,N_4545,N_251);
and U11279 (N_11279,N_1328,N_2366);
nor U11280 (N_11280,N_4795,N_1725);
nor U11281 (N_11281,N_2779,N_5820);
or U11282 (N_11282,N_3336,N_2769);
nor U11283 (N_11283,N_4831,N_683);
or U11284 (N_11284,N_2418,N_2626);
nor U11285 (N_11285,N_385,N_5619);
xnor U11286 (N_11286,N_37,N_3617);
and U11287 (N_11287,N_5499,N_1396);
and U11288 (N_11288,N_4647,N_4891);
nand U11289 (N_11289,N_2962,N_1267);
or U11290 (N_11290,N_3074,N_1239);
xor U11291 (N_11291,N_4306,N_3022);
xnor U11292 (N_11292,N_1870,N_2884);
nor U11293 (N_11293,N_3296,N_590);
and U11294 (N_11294,N_5814,N_3712);
or U11295 (N_11295,N_2678,N_1029);
nor U11296 (N_11296,N_5013,N_1746);
and U11297 (N_11297,N_3887,N_4876);
nand U11298 (N_11298,N_4959,N_1303);
or U11299 (N_11299,N_1829,N_5220);
xor U11300 (N_11300,N_5802,N_284);
xor U11301 (N_11301,N_1208,N_4163);
nand U11302 (N_11302,N_1812,N_1448);
nor U11303 (N_11303,N_2591,N_1019);
xnor U11304 (N_11304,N_1189,N_3110);
nor U11305 (N_11305,N_2716,N_3683);
xor U11306 (N_11306,N_5263,N_1557);
nand U11307 (N_11307,N_3132,N_2958);
and U11308 (N_11308,N_2805,N_988);
or U11309 (N_11309,N_54,N_2073);
nand U11310 (N_11310,N_815,N_2447);
xor U11311 (N_11311,N_108,N_1752);
nor U11312 (N_11312,N_1097,N_2903);
or U11313 (N_11313,N_5471,N_4471);
or U11314 (N_11314,N_4305,N_5878);
nand U11315 (N_11315,N_611,N_5454);
or U11316 (N_11316,N_5562,N_3613);
nor U11317 (N_11317,N_2120,N_3045);
or U11318 (N_11318,N_4021,N_5914);
and U11319 (N_11319,N_5692,N_5517);
and U11320 (N_11320,N_578,N_443);
and U11321 (N_11321,N_1296,N_1248);
nand U11322 (N_11322,N_3446,N_1867);
xnor U11323 (N_11323,N_4859,N_2927);
or U11324 (N_11324,N_2499,N_3466);
nor U11325 (N_11325,N_1976,N_5684);
xnor U11326 (N_11326,N_2550,N_527);
xnor U11327 (N_11327,N_4598,N_5089);
nor U11328 (N_11328,N_2618,N_5439);
or U11329 (N_11329,N_5434,N_2802);
nor U11330 (N_11330,N_722,N_1170);
nor U11331 (N_11331,N_3284,N_4580);
nor U11332 (N_11332,N_3854,N_2712);
nand U11333 (N_11333,N_3033,N_1834);
xnor U11334 (N_11334,N_2025,N_5380);
nor U11335 (N_11335,N_1724,N_2980);
and U11336 (N_11336,N_3007,N_3153);
or U11337 (N_11337,N_583,N_52);
xnor U11338 (N_11338,N_1160,N_765);
nor U11339 (N_11339,N_1346,N_4720);
nor U11340 (N_11340,N_4516,N_3063);
xnor U11341 (N_11341,N_1990,N_2505);
nand U11342 (N_11342,N_3238,N_2454);
xnor U11343 (N_11343,N_2985,N_531);
or U11344 (N_11344,N_4824,N_4419);
or U11345 (N_11345,N_1705,N_4620);
nor U11346 (N_11346,N_2827,N_2765);
and U11347 (N_11347,N_472,N_3124);
nor U11348 (N_11348,N_2274,N_1103);
or U11349 (N_11349,N_150,N_3775);
and U11350 (N_11350,N_32,N_284);
nor U11351 (N_11351,N_3431,N_237);
and U11352 (N_11352,N_3485,N_3024);
and U11353 (N_11353,N_1568,N_194);
or U11354 (N_11354,N_3856,N_1899);
xor U11355 (N_11355,N_5997,N_679);
xnor U11356 (N_11356,N_5704,N_3794);
xor U11357 (N_11357,N_1080,N_5803);
xor U11358 (N_11358,N_3313,N_3189);
nand U11359 (N_11359,N_3327,N_4241);
nor U11360 (N_11360,N_2234,N_3585);
or U11361 (N_11361,N_3249,N_3275);
nor U11362 (N_11362,N_411,N_2676);
nand U11363 (N_11363,N_3634,N_2262);
nand U11364 (N_11364,N_3760,N_5072);
and U11365 (N_11365,N_4427,N_5380);
nand U11366 (N_11366,N_3080,N_1942);
nor U11367 (N_11367,N_4607,N_213);
or U11368 (N_11368,N_373,N_406);
xor U11369 (N_11369,N_3329,N_2087);
nand U11370 (N_11370,N_1891,N_2116);
or U11371 (N_11371,N_4135,N_5612);
or U11372 (N_11372,N_1012,N_2954);
nand U11373 (N_11373,N_5144,N_3280);
nand U11374 (N_11374,N_3348,N_342);
and U11375 (N_11375,N_1324,N_5710);
nor U11376 (N_11376,N_4315,N_3963);
and U11377 (N_11377,N_5338,N_1392);
and U11378 (N_11378,N_5170,N_3888);
nor U11379 (N_11379,N_2750,N_4330);
nand U11380 (N_11380,N_1407,N_3256);
or U11381 (N_11381,N_4223,N_3242);
and U11382 (N_11382,N_2530,N_4699);
nand U11383 (N_11383,N_472,N_169);
xnor U11384 (N_11384,N_5570,N_3518);
and U11385 (N_11385,N_1719,N_123);
or U11386 (N_11386,N_4991,N_4363);
xor U11387 (N_11387,N_1764,N_5904);
xnor U11388 (N_11388,N_5153,N_5411);
xnor U11389 (N_11389,N_3366,N_719);
xor U11390 (N_11390,N_4872,N_2197);
nand U11391 (N_11391,N_3103,N_5662);
nor U11392 (N_11392,N_2033,N_3023);
xor U11393 (N_11393,N_3275,N_4064);
xnor U11394 (N_11394,N_5141,N_4594);
nand U11395 (N_11395,N_5335,N_664);
xnor U11396 (N_11396,N_1085,N_5708);
xor U11397 (N_11397,N_62,N_3770);
and U11398 (N_11398,N_278,N_2782);
xor U11399 (N_11399,N_1047,N_2799);
nand U11400 (N_11400,N_1895,N_4312);
or U11401 (N_11401,N_4868,N_4712);
nor U11402 (N_11402,N_2821,N_3882);
xor U11403 (N_11403,N_1052,N_5809);
xnor U11404 (N_11404,N_3205,N_2293);
nand U11405 (N_11405,N_4938,N_2855);
or U11406 (N_11406,N_1175,N_249);
nor U11407 (N_11407,N_4336,N_2886);
nand U11408 (N_11408,N_1727,N_4471);
nand U11409 (N_11409,N_2134,N_5282);
nor U11410 (N_11410,N_3209,N_4369);
nor U11411 (N_11411,N_340,N_1512);
nand U11412 (N_11412,N_2541,N_48);
or U11413 (N_11413,N_2301,N_3645);
xnor U11414 (N_11414,N_2513,N_3148);
nand U11415 (N_11415,N_2427,N_5639);
and U11416 (N_11416,N_2166,N_4464);
nor U11417 (N_11417,N_5203,N_2251);
and U11418 (N_11418,N_2547,N_2512);
or U11419 (N_11419,N_1334,N_3061);
xnor U11420 (N_11420,N_2694,N_1319);
and U11421 (N_11421,N_4726,N_5257);
and U11422 (N_11422,N_2376,N_4422);
xnor U11423 (N_11423,N_2367,N_2689);
nand U11424 (N_11424,N_30,N_5490);
or U11425 (N_11425,N_5414,N_4390);
nor U11426 (N_11426,N_2997,N_792);
or U11427 (N_11427,N_2331,N_2732);
nor U11428 (N_11428,N_5286,N_1198);
or U11429 (N_11429,N_2574,N_4199);
nor U11430 (N_11430,N_3968,N_2615);
and U11431 (N_11431,N_733,N_5838);
nor U11432 (N_11432,N_2931,N_5090);
nand U11433 (N_11433,N_1045,N_5179);
nand U11434 (N_11434,N_4098,N_5222);
or U11435 (N_11435,N_2039,N_44);
and U11436 (N_11436,N_5459,N_3517);
nand U11437 (N_11437,N_3798,N_5679);
or U11438 (N_11438,N_1497,N_4484);
nor U11439 (N_11439,N_357,N_2061);
nand U11440 (N_11440,N_2488,N_4528);
or U11441 (N_11441,N_3999,N_1085);
and U11442 (N_11442,N_4397,N_1538);
xnor U11443 (N_11443,N_352,N_5790);
nor U11444 (N_11444,N_89,N_292);
nand U11445 (N_11445,N_2811,N_3212);
or U11446 (N_11446,N_5306,N_3834);
xnor U11447 (N_11447,N_1021,N_1037);
and U11448 (N_11448,N_4734,N_4064);
or U11449 (N_11449,N_280,N_639);
xor U11450 (N_11450,N_5041,N_1365);
xor U11451 (N_11451,N_2412,N_3941);
and U11452 (N_11452,N_2500,N_662);
and U11453 (N_11453,N_3012,N_4776);
nand U11454 (N_11454,N_1519,N_161);
nor U11455 (N_11455,N_4331,N_1213);
and U11456 (N_11456,N_5022,N_1402);
and U11457 (N_11457,N_4109,N_973);
xnor U11458 (N_11458,N_3222,N_3174);
xnor U11459 (N_11459,N_3101,N_943);
or U11460 (N_11460,N_1177,N_1648);
nand U11461 (N_11461,N_2286,N_2041);
nand U11462 (N_11462,N_4016,N_4554);
nand U11463 (N_11463,N_211,N_3671);
nor U11464 (N_11464,N_4490,N_4866);
nor U11465 (N_11465,N_5702,N_4797);
or U11466 (N_11466,N_2478,N_433);
or U11467 (N_11467,N_1857,N_33);
nor U11468 (N_11468,N_3756,N_2671);
nor U11469 (N_11469,N_3129,N_3220);
or U11470 (N_11470,N_5434,N_4321);
and U11471 (N_11471,N_3611,N_2966);
xnor U11472 (N_11472,N_4870,N_3254);
xor U11473 (N_11473,N_1028,N_4505);
nand U11474 (N_11474,N_4516,N_330);
or U11475 (N_11475,N_65,N_61);
xor U11476 (N_11476,N_407,N_1759);
nand U11477 (N_11477,N_2282,N_2428);
nand U11478 (N_11478,N_4214,N_611);
nand U11479 (N_11479,N_1825,N_4891);
and U11480 (N_11480,N_1817,N_403);
or U11481 (N_11481,N_5597,N_4302);
nand U11482 (N_11482,N_3377,N_2066);
and U11483 (N_11483,N_5324,N_258);
or U11484 (N_11484,N_1254,N_2565);
xnor U11485 (N_11485,N_2866,N_1525);
or U11486 (N_11486,N_634,N_5204);
xor U11487 (N_11487,N_406,N_1748);
nand U11488 (N_11488,N_3056,N_2197);
or U11489 (N_11489,N_3765,N_3468);
or U11490 (N_11490,N_3449,N_573);
and U11491 (N_11491,N_1069,N_3739);
nand U11492 (N_11492,N_5377,N_844);
or U11493 (N_11493,N_16,N_3758);
nand U11494 (N_11494,N_1077,N_2636);
or U11495 (N_11495,N_4177,N_1441);
nand U11496 (N_11496,N_2880,N_5201);
nor U11497 (N_11497,N_4766,N_3609);
or U11498 (N_11498,N_1933,N_407);
and U11499 (N_11499,N_1778,N_2107);
and U11500 (N_11500,N_5155,N_3112);
nor U11501 (N_11501,N_4211,N_2101);
xnor U11502 (N_11502,N_935,N_847);
and U11503 (N_11503,N_2666,N_223);
nor U11504 (N_11504,N_5777,N_5135);
nor U11505 (N_11505,N_3953,N_3694);
nor U11506 (N_11506,N_3824,N_4635);
xor U11507 (N_11507,N_1693,N_2281);
nand U11508 (N_11508,N_440,N_1312);
and U11509 (N_11509,N_756,N_5723);
nor U11510 (N_11510,N_411,N_3077);
xnor U11511 (N_11511,N_2491,N_4124);
and U11512 (N_11512,N_3851,N_188);
nand U11513 (N_11513,N_4319,N_2082);
xor U11514 (N_11514,N_2012,N_2208);
nor U11515 (N_11515,N_4442,N_4010);
and U11516 (N_11516,N_4413,N_4616);
or U11517 (N_11517,N_4717,N_2196);
xor U11518 (N_11518,N_2221,N_4031);
xnor U11519 (N_11519,N_164,N_2684);
nand U11520 (N_11520,N_1194,N_4162);
nor U11521 (N_11521,N_4902,N_445);
and U11522 (N_11522,N_1536,N_4444);
xnor U11523 (N_11523,N_841,N_4916);
nand U11524 (N_11524,N_1459,N_4363);
nand U11525 (N_11525,N_3386,N_1819);
or U11526 (N_11526,N_2082,N_4165);
and U11527 (N_11527,N_3195,N_2187);
nor U11528 (N_11528,N_1429,N_4537);
xnor U11529 (N_11529,N_3485,N_5797);
xor U11530 (N_11530,N_2962,N_5349);
nor U11531 (N_11531,N_2089,N_3495);
xnor U11532 (N_11532,N_1726,N_1250);
or U11533 (N_11533,N_1888,N_1334);
nor U11534 (N_11534,N_1344,N_713);
or U11535 (N_11535,N_2397,N_5970);
or U11536 (N_11536,N_4410,N_1372);
xnor U11537 (N_11537,N_681,N_3392);
nand U11538 (N_11538,N_2846,N_3798);
xnor U11539 (N_11539,N_3400,N_2909);
and U11540 (N_11540,N_1997,N_3733);
nor U11541 (N_11541,N_556,N_4233);
or U11542 (N_11542,N_677,N_4928);
and U11543 (N_11543,N_4438,N_877);
and U11544 (N_11544,N_5493,N_5340);
xnor U11545 (N_11545,N_1543,N_834);
nand U11546 (N_11546,N_1860,N_2256);
nand U11547 (N_11547,N_1878,N_1286);
nand U11548 (N_11548,N_1733,N_1167);
xnor U11549 (N_11549,N_5022,N_2881);
xnor U11550 (N_11550,N_5275,N_5380);
nor U11551 (N_11551,N_4832,N_1232);
nor U11552 (N_11552,N_5055,N_750);
nand U11553 (N_11553,N_4431,N_616);
xor U11554 (N_11554,N_1161,N_2146);
nor U11555 (N_11555,N_5002,N_3377);
nand U11556 (N_11556,N_2584,N_246);
nor U11557 (N_11557,N_5928,N_5561);
and U11558 (N_11558,N_2255,N_4348);
xnor U11559 (N_11559,N_2129,N_1776);
xor U11560 (N_11560,N_1131,N_1688);
and U11561 (N_11561,N_5092,N_5708);
nor U11562 (N_11562,N_4181,N_1608);
nand U11563 (N_11563,N_2732,N_3598);
nor U11564 (N_11564,N_5967,N_2723);
xor U11565 (N_11565,N_3322,N_3936);
and U11566 (N_11566,N_2592,N_2480);
xor U11567 (N_11567,N_891,N_3725);
or U11568 (N_11568,N_5298,N_3190);
nor U11569 (N_11569,N_2493,N_5080);
or U11570 (N_11570,N_1248,N_5572);
or U11571 (N_11571,N_2394,N_4117);
or U11572 (N_11572,N_3193,N_2146);
or U11573 (N_11573,N_4461,N_3679);
nand U11574 (N_11574,N_198,N_4529);
nand U11575 (N_11575,N_3613,N_678);
xnor U11576 (N_11576,N_3434,N_2952);
nand U11577 (N_11577,N_3997,N_3591);
and U11578 (N_11578,N_4052,N_4001);
xnor U11579 (N_11579,N_3957,N_5586);
xor U11580 (N_11580,N_4959,N_7);
or U11581 (N_11581,N_1741,N_5625);
nand U11582 (N_11582,N_519,N_2030);
nand U11583 (N_11583,N_1231,N_2610);
nand U11584 (N_11584,N_4954,N_5410);
xor U11585 (N_11585,N_3498,N_3468);
and U11586 (N_11586,N_4009,N_4235);
nor U11587 (N_11587,N_3782,N_1107);
nand U11588 (N_11588,N_2964,N_3198);
xor U11589 (N_11589,N_4018,N_3501);
nor U11590 (N_11590,N_160,N_4555);
nand U11591 (N_11591,N_3948,N_403);
nand U11592 (N_11592,N_618,N_3114);
xnor U11593 (N_11593,N_5379,N_1772);
and U11594 (N_11594,N_2539,N_192);
and U11595 (N_11595,N_5151,N_4417);
or U11596 (N_11596,N_729,N_5131);
xor U11597 (N_11597,N_1355,N_2900);
and U11598 (N_11598,N_3410,N_1295);
and U11599 (N_11599,N_1402,N_4045);
and U11600 (N_11600,N_1638,N_5030);
nand U11601 (N_11601,N_1886,N_5521);
and U11602 (N_11602,N_205,N_2668);
or U11603 (N_11603,N_2930,N_2055);
and U11604 (N_11604,N_3526,N_3089);
and U11605 (N_11605,N_5936,N_2678);
or U11606 (N_11606,N_3419,N_484);
nor U11607 (N_11607,N_1698,N_3681);
nand U11608 (N_11608,N_5461,N_1854);
nand U11609 (N_11609,N_2289,N_4461);
and U11610 (N_11610,N_1377,N_3875);
or U11611 (N_11611,N_586,N_3235);
or U11612 (N_11612,N_2071,N_4063);
xnor U11613 (N_11613,N_5574,N_4812);
and U11614 (N_11614,N_2492,N_2317);
nand U11615 (N_11615,N_3375,N_4907);
nor U11616 (N_11616,N_3489,N_796);
nand U11617 (N_11617,N_1279,N_3703);
xnor U11618 (N_11618,N_1579,N_833);
nand U11619 (N_11619,N_4318,N_2093);
xnor U11620 (N_11620,N_1342,N_5026);
or U11621 (N_11621,N_5608,N_4967);
and U11622 (N_11622,N_951,N_3446);
nor U11623 (N_11623,N_435,N_4611);
nor U11624 (N_11624,N_740,N_1618);
or U11625 (N_11625,N_773,N_3392);
nor U11626 (N_11626,N_2434,N_3360);
xor U11627 (N_11627,N_5425,N_2259);
or U11628 (N_11628,N_1068,N_5824);
and U11629 (N_11629,N_3274,N_3259);
xnor U11630 (N_11630,N_1854,N_5637);
xnor U11631 (N_11631,N_369,N_5304);
and U11632 (N_11632,N_2464,N_2460);
or U11633 (N_11633,N_3845,N_3403);
nor U11634 (N_11634,N_4666,N_2249);
and U11635 (N_11635,N_377,N_2090);
xor U11636 (N_11636,N_5470,N_5399);
nor U11637 (N_11637,N_3999,N_2320);
nand U11638 (N_11638,N_3263,N_1430);
or U11639 (N_11639,N_4553,N_1855);
xnor U11640 (N_11640,N_2282,N_5455);
or U11641 (N_11641,N_1392,N_4352);
nor U11642 (N_11642,N_3195,N_1315);
or U11643 (N_11643,N_5834,N_826);
and U11644 (N_11644,N_332,N_1391);
nor U11645 (N_11645,N_2757,N_115);
xnor U11646 (N_11646,N_5579,N_1657);
and U11647 (N_11647,N_3318,N_199);
and U11648 (N_11648,N_274,N_3097);
xnor U11649 (N_11649,N_1603,N_4824);
nor U11650 (N_11650,N_4072,N_546);
or U11651 (N_11651,N_4410,N_892);
xor U11652 (N_11652,N_3456,N_2642);
and U11653 (N_11653,N_3734,N_5694);
or U11654 (N_11654,N_282,N_61);
or U11655 (N_11655,N_4604,N_3898);
nand U11656 (N_11656,N_1790,N_2188);
nand U11657 (N_11657,N_2077,N_2146);
nand U11658 (N_11658,N_1736,N_4376);
xnor U11659 (N_11659,N_752,N_2980);
or U11660 (N_11660,N_5156,N_2858);
nand U11661 (N_11661,N_1553,N_5572);
and U11662 (N_11662,N_1393,N_3431);
nor U11663 (N_11663,N_4477,N_828);
nor U11664 (N_11664,N_5321,N_1086);
or U11665 (N_11665,N_4488,N_4721);
nor U11666 (N_11666,N_1899,N_5554);
or U11667 (N_11667,N_1043,N_3847);
and U11668 (N_11668,N_5661,N_2976);
or U11669 (N_11669,N_3152,N_2682);
nand U11670 (N_11670,N_2479,N_1001);
and U11671 (N_11671,N_5876,N_5021);
xnor U11672 (N_11672,N_212,N_14);
nand U11673 (N_11673,N_4161,N_3894);
or U11674 (N_11674,N_4062,N_1271);
xor U11675 (N_11675,N_1781,N_2270);
nand U11676 (N_11676,N_4114,N_5193);
nor U11677 (N_11677,N_844,N_3557);
nand U11678 (N_11678,N_2353,N_1129);
and U11679 (N_11679,N_4459,N_4487);
xnor U11680 (N_11680,N_3672,N_5648);
xor U11681 (N_11681,N_1411,N_2480);
or U11682 (N_11682,N_252,N_4231);
and U11683 (N_11683,N_5391,N_5682);
and U11684 (N_11684,N_1571,N_228);
nand U11685 (N_11685,N_4219,N_5598);
nor U11686 (N_11686,N_911,N_4864);
or U11687 (N_11687,N_920,N_1431);
nand U11688 (N_11688,N_3719,N_2940);
and U11689 (N_11689,N_2728,N_3440);
and U11690 (N_11690,N_4545,N_1291);
xor U11691 (N_11691,N_3060,N_1949);
or U11692 (N_11692,N_3278,N_581);
or U11693 (N_11693,N_1039,N_804);
or U11694 (N_11694,N_5208,N_4628);
or U11695 (N_11695,N_1326,N_5741);
nor U11696 (N_11696,N_1310,N_3324);
and U11697 (N_11697,N_5905,N_5011);
and U11698 (N_11698,N_3619,N_3800);
xor U11699 (N_11699,N_3446,N_350);
and U11700 (N_11700,N_1091,N_5334);
and U11701 (N_11701,N_3469,N_1972);
nand U11702 (N_11702,N_4095,N_2135);
and U11703 (N_11703,N_255,N_1590);
nand U11704 (N_11704,N_2985,N_3393);
or U11705 (N_11705,N_4172,N_2347);
nand U11706 (N_11706,N_3522,N_2607);
xor U11707 (N_11707,N_697,N_1412);
xnor U11708 (N_11708,N_2,N_86);
nand U11709 (N_11709,N_1723,N_5047);
and U11710 (N_11710,N_3776,N_2461);
nand U11711 (N_11711,N_3361,N_1608);
or U11712 (N_11712,N_4374,N_2001);
xnor U11713 (N_11713,N_806,N_4406);
xnor U11714 (N_11714,N_1956,N_2294);
or U11715 (N_11715,N_1217,N_1926);
xor U11716 (N_11716,N_3109,N_5753);
and U11717 (N_11717,N_5498,N_2471);
nand U11718 (N_11718,N_5461,N_4476);
nand U11719 (N_11719,N_2201,N_2669);
nand U11720 (N_11720,N_2909,N_922);
xnor U11721 (N_11721,N_880,N_3816);
or U11722 (N_11722,N_5453,N_735);
or U11723 (N_11723,N_2407,N_894);
and U11724 (N_11724,N_1778,N_1275);
or U11725 (N_11725,N_537,N_4475);
nor U11726 (N_11726,N_581,N_5584);
xnor U11727 (N_11727,N_5160,N_2324);
xor U11728 (N_11728,N_2221,N_1015);
and U11729 (N_11729,N_1024,N_5375);
xor U11730 (N_11730,N_3696,N_2800);
nor U11731 (N_11731,N_2038,N_4183);
xnor U11732 (N_11732,N_3412,N_3780);
or U11733 (N_11733,N_2347,N_4222);
and U11734 (N_11734,N_4907,N_117);
and U11735 (N_11735,N_135,N_1010);
and U11736 (N_11736,N_2735,N_5778);
nand U11737 (N_11737,N_3257,N_3597);
xor U11738 (N_11738,N_2049,N_719);
and U11739 (N_11739,N_3463,N_3532);
and U11740 (N_11740,N_3219,N_185);
or U11741 (N_11741,N_1593,N_5755);
or U11742 (N_11742,N_2397,N_5680);
xnor U11743 (N_11743,N_4416,N_1012);
nand U11744 (N_11744,N_115,N_2524);
and U11745 (N_11745,N_1660,N_1954);
nor U11746 (N_11746,N_5191,N_3051);
xnor U11747 (N_11747,N_3037,N_1859);
nor U11748 (N_11748,N_1310,N_803);
nand U11749 (N_11749,N_4390,N_4277);
nor U11750 (N_11750,N_3367,N_2464);
nand U11751 (N_11751,N_2606,N_253);
nor U11752 (N_11752,N_3328,N_2428);
nor U11753 (N_11753,N_4751,N_2473);
or U11754 (N_11754,N_5295,N_3421);
nor U11755 (N_11755,N_3609,N_3244);
and U11756 (N_11756,N_5182,N_5306);
nor U11757 (N_11757,N_4284,N_751);
nand U11758 (N_11758,N_3309,N_2443);
xor U11759 (N_11759,N_1789,N_3018);
and U11760 (N_11760,N_2774,N_3637);
or U11761 (N_11761,N_480,N_2615);
nor U11762 (N_11762,N_4712,N_1947);
nand U11763 (N_11763,N_2151,N_901);
nor U11764 (N_11764,N_253,N_2497);
xnor U11765 (N_11765,N_3202,N_4043);
xor U11766 (N_11766,N_4456,N_2694);
xnor U11767 (N_11767,N_301,N_5961);
or U11768 (N_11768,N_1551,N_68);
nor U11769 (N_11769,N_2628,N_4477);
xnor U11770 (N_11770,N_5325,N_2432);
xnor U11771 (N_11771,N_2901,N_2723);
nand U11772 (N_11772,N_37,N_4149);
nor U11773 (N_11773,N_4168,N_3510);
xor U11774 (N_11774,N_723,N_4809);
nand U11775 (N_11775,N_3638,N_4899);
nand U11776 (N_11776,N_2317,N_5724);
and U11777 (N_11777,N_3128,N_3442);
xor U11778 (N_11778,N_5946,N_1192);
and U11779 (N_11779,N_2350,N_1038);
nand U11780 (N_11780,N_4381,N_3473);
xnor U11781 (N_11781,N_384,N_2291);
and U11782 (N_11782,N_3727,N_5544);
nand U11783 (N_11783,N_4098,N_5939);
and U11784 (N_11784,N_876,N_5924);
and U11785 (N_11785,N_3433,N_1294);
xnor U11786 (N_11786,N_3304,N_4159);
or U11787 (N_11787,N_5919,N_3408);
or U11788 (N_11788,N_273,N_1745);
and U11789 (N_11789,N_1352,N_2228);
nand U11790 (N_11790,N_5981,N_4659);
and U11791 (N_11791,N_4338,N_4472);
and U11792 (N_11792,N_2449,N_5948);
nand U11793 (N_11793,N_4162,N_3419);
and U11794 (N_11794,N_5834,N_4828);
or U11795 (N_11795,N_4378,N_2240);
nand U11796 (N_11796,N_4426,N_1203);
or U11797 (N_11797,N_3069,N_771);
and U11798 (N_11798,N_2783,N_2501);
xnor U11799 (N_11799,N_442,N_1443);
nor U11800 (N_11800,N_1761,N_3232);
nor U11801 (N_11801,N_2092,N_5890);
nand U11802 (N_11802,N_2678,N_2630);
and U11803 (N_11803,N_5958,N_4098);
nor U11804 (N_11804,N_4391,N_3733);
xnor U11805 (N_11805,N_842,N_5154);
or U11806 (N_11806,N_4977,N_1545);
nand U11807 (N_11807,N_4430,N_5614);
xnor U11808 (N_11808,N_4735,N_1379);
nor U11809 (N_11809,N_4808,N_3634);
and U11810 (N_11810,N_3333,N_2572);
nor U11811 (N_11811,N_1001,N_4952);
nand U11812 (N_11812,N_5548,N_1380);
or U11813 (N_11813,N_1146,N_1051);
nand U11814 (N_11814,N_1943,N_2968);
nand U11815 (N_11815,N_5766,N_211);
nand U11816 (N_11816,N_2640,N_785);
and U11817 (N_11817,N_5653,N_2477);
nor U11818 (N_11818,N_4252,N_1863);
or U11819 (N_11819,N_4416,N_3159);
nand U11820 (N_11820,N_1388,N_3435);
nand U11821 (N_11821,N_5385,N_3922);
or U11822 (N_11822,N_1123,N_2646);
nor U11823 (N_11823,N_800,N_4087);
nor U11824 (N_11824,N_703,N_4899);
xor U11825 (N_11825,N_5515,N_1188);
xnor U11826 (N_11826,N_4320,N_55);
nor U11827 (N_11827,N_1387,N_906);
xnor U11828 (N_11828,N_505,N_4599);
nand U11829 (N_11829,N_4096,N_5722);
or U11830 (N_11830,N_4307,N_144);
and U11831 (N_11831,N_3229,N_2693);
or U11832 (N_11832,N_5166,N_4465);
nand U11833 (N_11833,N_2553,N_3695);
xor U11834 (N_11834,N_3031,N_253);
and U11835 (N_11835,N_2180,N_4262);
and U11836 (N_11836,N_1192,N_1808);
xnor U11837 (N_11837,N_4286,N_205);
and U11838 (N_11838,N_4424,N_3702);
xnor U11839 (N_11839,N_2651,N_3778);
and U11840 (N_11840,N_2419,N_822);
nor U11841 (N_11841,N_3215,N_4237);
or U11842 (N_11842,N_1912,N_3644);
or U11843 (N_11843,N_1807,N_4338);
nand U11844 (N_11844,N_5328,N_1681);
or U11845 (N_11845,N_5253,N_5618);
xnor U11846 (N_11846,N_5725,N_4619);
nand U11847 (N_11847,N_1610,N_5575);
nor U11848 (N_11848,N_4766,N_2311);
or U11849 (N_11849,N_2879,N_1233);
nor U11850 (N_11850,N_5528,N_2296);
or U11851 (N_11851,N_551,N_5523);
nor U11852 (N_11852,N_1318,N_1649);
nor U11853 (N_11853,N_4475,N_1960);
xnor U11854 (N_11854,N_1,N_4234);
or U11855 (N_11855,N_5477,N_5272);
and U11856 (N_11856,N_4447,N_1091);
or U11857 (N_11857,N_4565,N_2140);
and U11858 (N_11858,N_2770,N_3246);
xor U11859 (N_11859,N_1273,N_1959);
xnor U11860 (N_11860,N_241,N_981);
and U11861 (N_11861,N_4305,N_2866);
nand U11862 (N_11862,N_2261,N_5760);
or U11863 (N_11863,N_1354,N_3223);
xnor U11864 (N_11864,N_4152,N_1348);
nor U11865 (N_11865,N_5406,N_515);
nor U11866 (N_11866,N_5023,N_2433);
nor U11867 (N_11867,N_1073,N_4145);
nor U11868 (N_11868,N_1130,N_4175);
xor U11869 (N_11869,N_895,N_537);
xor U11870 (N_11870,N_2851,N_3879);
nand U11871 (N_11871,N_1645,N_3102);
and U11872 (N_11872,N_872,N_405);
nor U11873 (N_11873,N_3453,N_2496);
nor U11874 (N_11874,N_3699,N_3150);
or U11875 (N_11875,N_929,N_4004);
nor U11876 (N_11876,N_731,N_5560);
and U11877 (N_11877,N_5666,N_2117);
and U11878 (N_11878,N_234,N_4771);
nor U11879 (N_11879,N_2293,N_3329);
xor U11880 (N_11880,N_5862,N_4477);
xor U11881 (N_11881,N_5217,N_2120);
or U11882 (N_11882,N_3417,N_5689);
and U11883 (N_11883,N_3384,N_1270);
nand U11884 (N_11884,N_2435,N_370);
or U11885 (N_11885,N_3916,N_5336);
or U11886 (N_11886,N_5649,N_1891);
nand U11887 (N_11887,N_4177,N_3029);
nand U11888 (N_11888,N_913,N_4209);
nor U11889 (N_11889,N_1829,N_3142);
nor U11890 (N_11890,N_1796,N_1013);
nand U11891 (N_11891,N_1263,N_3539);
xnor U11892 (N_11892,N_2046,N_1036);
and U11893 (N_11893,N_835,N_1586);
nand U11894 (N_11894,N_518,N_287);
and U11895 (N_11895,N_4087,N_2833);
nand U11896 (N_11896,N_1473,N_38);
nor U11897 (N_11897,N_2975,N_3966);
and U11898 (N_11898,N_3885,N_421);
xnor U11899 (N_11899,N_4496,N_4659);
nand U11900 (N_11900,N_5622,N_3468);
and U11901 (N_11901,N_891,N_1297);
nand U11902 (N_11902,N_4890,N_2226);
and U11903 (N_11903,N_2367,N_1257);
xnor U11904 (N_11904,N_167,N_3950);
or U11905 (N_11905,N_425,N_5246);
and U11906 (N_11906,N_4806,N_2441);
nor U11907 (N_11907,N_113,N_5250);
xnor U11908 (N_11908,N_1294,N_476);
nand U11909 (N_11909,N_2735,N_2892);
nor U11910 (N_11910,N_855,N_4919);
and U11911 (N_11911,N_4702,N_4269);
or U11912 (N_11912,N_345,N_3987);
nand U11913 (N_11913,N_4625,N_637);
xor U11914 (N_11914,N_2760,N_1630);
nor U11915 (N_11915,N_5143,N_873);
or U11916 (N_11916,N_799,N_1924);
and U11917 (N_11917,N_3045,N_5876);
or U11918 (N_11918,N_4956,N_5819);
and U11919 (N_11919,N_1315,N_8);
nand U11920 (N_11920,N_4309,N_1062);
xor U11921 (N_11921,N_1210,N_5309);
xor U11922 (N_11922,N_373,N_3084);
nor U11923 (N_11923,N_3959,N_2308);
and U11924 (N_11924,N_3019,N_4758);
or U11925 (N_11925,N_4086,N_2310);
nand U11926 (N_11926,N_1015,N_5929);
nand U11927 (N_11927,N_3745,N_4030);
and U11928 (N_11928,N_537,N_2361);
or U11929 (N_11929,N_5410,N_236);
nand U11930 (N_11930,N_1791,N_2235);
xnor U11931 (N_11931,N_4390,N_4217);
or U11932 (N_11932,N_1077,N_2509);
xor U11933 (N_11933,N_4798,N_4255);
and U11934 (N_11934,N_1737,N_315);
or U11935 (N_11935,N_2186,N_3653);
nand U11936 (N_11936,N_367,N_4153);
or U11937 (N_11937,N_4666,N_2934);
nand U11938 (N_11938,N_307,N_146);
or U11939 (N_11939,N_5125,N_133);
nand U11940 (N_11940,N_2400,N_4734);
nor U11941 (N_11941,N_510,N_1826);
and U11942 (N_11942,N_3942,N_2968);
and U11943 (N_11943,N_1336,N_5682);
and U11944 (N_11944,N_2680,N_554);
or U11945 (N_11945,N_3728,N_2497);
nand U11946 (N_11946,N_1356,N_5931);
xnor U11947 (N_11947,N_4477,N_4591);
or U11948 (N_11948,N_3037,N_1513);
or U11949 (N_11949,N_3557,N_3540);
and U11950 (N_11950,N_1940,N_35);
nand U11951 (N_11951,N_3122,N_4529);
xor U11952 (N_11952,N_2507,N_5112);
nor U11953 (N_11953,N_5417,N_4229);
nand U11954 (N_11954,N_196,N_1481);
or U11955 (N_11955,N_4523,N_5056);
or U11956 (N_11956,N_3704,N_3617);
and U11957 (N_11957,N_4260,N_5707);
nor U11958 (N_11958,N_2235,N_366);
xnor U11959 (N_11959,N_3782,N_983);
and U11960 (N_11960,N_1660,N_2479);
or U11961 (N_11961,N_5730,N_5115);
or U11962 (N_11962,N_4943,N_1014);
nor U11963 (N_11963,N_2025,N_5381);
nor U11964 (N_11964,N_230,N_2712);
nand U11965 (N_11965,N_2397,N_3416);
or U11966 (N_11966,N_1623,N_1163);
nor U11967 (N_11967,N_282,N_5338);
or U11968 (N_11968,N_3578,N_2979);
and U11969 (N_11969,N_302,N_4156);
nand U11970 (N_11970,N_202,N_5657);
or U11971 (N_11971,N_4583,N_34);
and U11972 (N_11972,N_1833,N_2507);
and U11973 (N_11973,N_236,N_3928);
or U11974 (N_11974,N_1728,N_4066);
nor U11975 (N_11975,N_2504,N_5992);
or U11976 (N_11976,N_1465,N_2993);
nand U11977 (N_11977,N_1706,N_3006);
nand U11978 (N_11978,N_4742,N_2422);
nand U11979 (N_11979,N_4854,N_1713);
or U11980 (N_11980,N_964,N_5226);
nand U11981 (N_11981,N_1592,N_5829);
xnor U11982 (N_11982,N_5215,N_2420);
or U11983 (N_11983,N_4548,N_5797);
nor U11984 (N_11984,N_1163,N_1585);
nand U11985 (N_11985,N_1016,N_5500);
nor U11986 (N_11986,N_2816,N_4799);
and U11987 (N_11987,N_5388,N_2106);
or U11988 (N_11988,N_2471,N_2550);
nor U11989 (N_11989,N_3842,N_1279);
nand U11990 (N_11990,N_3007,N_1049);
or U11991 (N_11991,N_5490,N_2979);
nand U11992 (N_11992,N_4930,N_4592);
and U11993 (N_11993,N_2552,N_3406);
and U11994 (N_11994,N_3164,N_409);
and U11995 (N_11995,N_471,N_3990);
xnor U11996 (N_11996,N_1595,N_3098);
nor U11997 (N_11997,N_3342,N_4200);
and U11998 (N_11998,N_1640,N_798);
and U11999 (N_11999,N_1750,N_5079);
xnor U12000 (N_12000,N_11893,N_8346);
nand U12001 (N_12001,N_7929,N_8351);
xor U12002 (N_12002,N_9632,N_11186);
and U12003 (N_12003,N_11384,N_10010);
or U12004 (N_12004,N_9789,N_9749);
and U12005 (N_12005,N_9159,N_11951);
or U12006 (N_12006,N_10113,N_6448);
or U12007 (N_12007,N_9271,N_9331);
xor U12008 (N_12008,N_6818,N_10450);
nor U12009 (N_12009,N_10588,N_10348);
and U12010 (N_12010,N_11700,N_7321);
or U12011 (N_12011,N_11521,N_11329);
and U12012 (N_12012,N_6174,N_7198);
or U12013 (N_12013,N_6767,N_9160);
xnor U12014 (N_12014,N_7390,N_9548);
xnor U12015 (N_12015,N_9965,N_11537);
xnor U12016 (N_12016,N_6695,N_7746);
and U12017 (N_12017,N_9065,N_11415);
nand U12018 (N_12018,N_7446,N_7550);
xnor U12019 (N_12019,N_10827,N_8960);
or U12020 (N_12020,N_11802,N_11523);
or U12021 (N_12021,N_10448,N_9492);
xnor U12022 (N_12022,N_11484,N_7754);
nor U12023 (N_12023,N_10037,N_8686);
xor U12024 (N_12024,N_8427,N_11784);
nand U12025 (N_12025,N_11269,N_9772);
nand U12026 (N_12026,N_10093,N_9234);
nand U12027 (N_12027,N_9799,N_9531);
nor U12028 (N_12028,N_6846,N_6103);
xor U12029 (N_12029,N_10259,N_11930);
and U12030 (N_12030,N_9577,N_8554);
and U12031 (N_12031,N_9896,N_8943);
nor U12032 (N_12032,N_7978,N_7745);
nand U12033 (N_12033,N_8716,N_10521);
or U12034 (N_12034,N_10011,N_7666);
xor U12035 (N_12035,N_10822,N_11495);
xnor U12036 (N_12036,N_7069,N_11796);
nand U12037 (N_12037,N_9472,N_9400);
and U12038 (N_12038,N_9635,N_6155);
nand U12039 (N_12039,N_10422,N_7961);
and U12040 (N_12040,N_6526,N_11702);
and U12041 (N_12041,N_10159,N_7246);
xnor U12042 (N_12042,N_10245,N_6552);
nor U12043 (N_12043,N_10921,N_7574);
xnor U12044 (N_12044,N_6218,N_10028);
nand U12045 (N_12045,N_6693,N_8200);
or U12046 (N_12046,N_6874,N_10511);
or U12047 (N_12047,N_10547,N_7134);
nand U12048 (N_12048,N_7096,N_11313);
xnor U12049 (N_12049,N_11445,N_11088);
and U12050 (N_12050,N_11426,N_8851);
nand U12051 (N_12051,N_10533,N_6081);
or U12052 (N_12052,N_8080,N_7848);
or U12053 (N_12053,N_7311,N_10768);
xor U12054 (N_12054,N_11576,N_10691);
nor U12055 (N_12055,N_7020,N_10463);
and U12056 (N_12056,N_11076,N_7620);
and U12057 (N_12057,N_9422,N_7384);
nor U12058 (N_12058,N_9328,N_7739);
and U12059 (N_12059,N_11752,N_9007);
nor U12060 (N_12060,N_8421,N_6434);
and U12061 (N_12061,N_9384,N_9618);
and U12062 (N_12062,N_10960,N_7217);
nor U12063 (N_12063,N_7553,N_6264);
or U12064 (N_12064,N_6186,N_6293);
and U12065 (N_12065,N_9615,N_6203);
nor U12066 (N_12066,N_8688,N_10050);
nor U12067 (N_12067,N_9236,N_8495);
xnor U12068 (N_12068,N_7082,N_6176);
nor U12069 (N_12069,N_11090,N_7726);
nand U12070 (N_12070,N_9725,N_8771);
or U12071 (N_12071,N_8619,N_11962);
nand U12072 (N_12072,N_7907,N_10627);
and U12073 (N_12073,N_8362,N_7532);
nor U12074 (N_12074,N_10544,N_8590);
xor U12075 (N_12075,N_9147,N_6784);
nor U12076 (N_12076,N_8594,N_8720);
nor U12077 (N_12077,N_7445,N_9945);
and U12078 (N_12078,N_7706,N_11937);
or U12079 (N_12079,N_10571,N_11001);
xor U12080 (N_12080,N_8354,N_11114);
nor U12081 (N_12081,N_6928,N_11008);
and U12082 (N_12082,N_6499,N_7972);
and U12083 (N_12083,N_7994,N_11773);
and U12084 (N_12084,N_6074,N_9465);
or U12085 (N_12085,N_7953,N_9258);
nor U12086 (N_12086,N_6646,N_8700);
nor U12087 (N_12087,N_9515,N_6905);
nand U12088 (N_12088,N_6788,N_6051);
nor U12089 (N_12089,N_7061,N_11189);
nor U12090 (N_12090,N_11050,N_11619);
xor U12091 (N_12091,N_7495,N_11869);
nor U12092 (N_12092,N_9148,N_7452);
nand U12093 (N_12093,N_10392,N_10455);
and U12094 (N_12094,N_9326,N_6345);
nand U12095 (N_12095,N_8244,N_7383);
xor U12096 (N_12096,N_9360,N_7345);
nand U12097 (N_12097,N_8772,N_10800);
and U12098 (N_12098,N_9304,N_11212);
or U12099 (N_12099,N_6990,N_8683);
and U12100 (N_12100,N_10877,N_9891);
or U12101 (N_12101,N_9638,N_7851);
xnor U12102 (N_12102,N_8301,N_8132);
nand U12103 (N_12103,N_10437,N_11643);
and U12104 (N_12104,N_6407,N_9685);
nor U12105 (N_12105,N_7300,N_7733);
and U12106 (N_12106,N_9091,N_6167);
and U12107 (N_12107,N_10480,N_6613);
nor U12108 (N_12108,N_8168,N_11213);
or U12109 (N_12109,N_10531,N_10252);
nand U12110 (N_12110,N_7177,N_10192);
xor U12111 (N_12111,N_8250,N_9867);
nor U12112 (N_12112,N_8744,N_8062);
nand U12113 (N_12113,N_7215,N_6503);
and U12114 (N_12114,N_11738,N_9922);
and U12115 (N_12115,N_8931,N_9766);
xor U12116 (N_12116,N_11424,N_11874);
xnor U12117 (N_12117,N_6758,N_8253);
nor U12118 (N_12118,N_6305,N_6873);
or U12119 (N_12119,N_9103,N_8852);
xnor U12120 (N_12120,N_8779,N_10896);
nand U12121 (N_12121,N_8607,N_7108);
or U12122 (N_12122,N_11648,N_7595);
nand U12123 (N_12123,N_9626,N_9043);
nand U12124 (N_12124,N_9373,N_10497);
and U12125 (N_12125,N_7890,N_8860);
nand U12126 (N_12126,N_6493,N_8798);
or U12127 (N_12127,N_7527,N_7404);
nor U12128 (N_12128,N_10312,N_7172);
and U12129 (N_12129,N_8794,N_10714);
or U12130 (N_12130,N_6603,N_10805);
or U12131 (N_12131,N_10841,N_9461);
nand U12132 (N_12132,N_9120,N_9957);
nand U12133 (N_12133,N_7387,N_8949);
or U12134 (N_12134,N_6986,N_7074);
and U12135 (N_12135,N_8310,N_11462);
or U12136 (N_12136,N_11955,N_11672);
and U12137 (N_12137,N_9066,N_8923);
nand U12138 (N_12138,N_10417,N_7583);
nand U12139 (N_12139,N_9033,N_11585);
or U12140 (N_12140,N_9785,N_7167);
nand U12141 (N_12141,N_9778,N_7344);
and U12142 (N_12142,N_10145,N_8566);
or U12143 (N_12143,N_6795,N_6994);
or U12144 (N_12144,N_10638,N_8681);
nand U12145 (N_12145,N_11662,N_6590);
and U12146 (N_12146,N_10632,N_11499);
nor U12147 (N_12147,N_10982,N_9901);
or U12148 (N_12148,N_10570,N_6346);
or U12149 (N_12149,N_11265,N_10489);
nand U12150 (N_12150,N_10490,N_8486);
or U12151 (N_12151,N_11765,N_9455);
nor U12152 (N_12152,N_6424,N_9296);
or U12153 (N_12153,N_10598,N_7434);
nor U12154 (N_12154,N_11519,N_11933);
or U12155 (N_12155,N_7989,N_8854);
nand U12156 (N_12156,N_9002,N_10869);
nor U12157 (N_12157,N_7515,N_10469);
and U12158 (N_12158,N_9324,N_11063);
nand U12159 (N_12159,N_10386,N_9289);
or U12160 (N_12160,N_7719,N_11291);
or U12161 (N_12161,N_10368,N_8534);
nand U12162 (N_12162,N_6200,N_7682);
nand U12163 (N_12163,N_8615,N_9740);
nand U12164 (N_12164,N_8012,N_6184);
nand U12165 (N_12165,N_8034,N_6809);
nand U12166 (N_12166,N_7054,N_6625);
xnor U12167 (N_12167,N_9267,N_8109);
and U12168 (N_12168,N_10327,N_9252);
or U12169 (N_12169,N_7269,N_6249);
nor U12170 (N_12170,N_11200,N_11655);
xor U12171 (N_12171,N_6022,N_8199);
nor U12172 (N_12172,N_10398,N_8343);
and U12173 (N_12173,N_6391,N_7511);
or U12174 (N_12174,N_6090,N_8041);
nor U12175 (N_12175,N_7212,N_8747);
nand U12176 (N_12176,N_11525,N_8298);
xnor U12177 (N_12177,N_9314,N_7443);
nand U12178 (N_12178,N_9392,N_8542);
nand U12179 (N_12179,N_11650,N_7471);
nand U12180 (N_12180,N_6385,N_9829);
and U12181 (N_12181,N_7457,N_7674);
or U12182 (N_12182,N_7474,N_9856);
xor U12183 (N_12183,N_8647,N_8289);
xnor U12184 (N_12184,N_11046,N_8536);
or U12185 (N_12185,N_10336,N_10901);
nand U12186 (N_12186,N_6820,N_8039);
nor U12187 (N_12187,N_7147,N_8711);
nand U12188 (N_12188,N_6122,N_6220);
and U12189 (N_12189,N_7165,N_8485);
nor U12190 (N_12190,N_8529,N_6876);
or U12191 (N_12191,N_11664,N_8904);
nand U12192 (N_12192,N_10472,N_9087);
and U12193 (N_12193,N_9463,N_6779);
or U12194 (N_12194,N_11266,N_11281);
nand U12195 (N_12195,N_9182,N_8826);
xnor U12196 (N_12196,N_6671,N_11304);
and U12197 (N_12197,N_10996,N_8708);
nor U12198 (N_12198,N_10746,N_8699);
nor U12199 (N_12199,N_7905,N_10859);
nor U12200 (N_12200,N_11982,N_7483);
nor U12201 (N_12201,N_10622,N_7777);
or U12202 (N_12202,N_6047,N_7124);
xnor U12203 (N_12203,N_6395,N_10042);
or U12204 (N_12204,N_9102,N_8028);
and U12205 (N_12205,N_7053,N_7716);
or U12206 (N_12206,N_7886,N_9157);
xor U12207 (N_12207,N_11887,N_8629);
and U12208 (N_12208,N_6916,N_7829);
or U12209 (N_12209,N_11161,N_8078);
nand U12210 (N_12210,N_10594,N_8477);
nand U12211 (N_12211,N_8161,N_8879);
xnor U12212 (N_12212,N_10180,N_9379);
or U12213 (N_12213,N_8287,N_9519);
xor U12214 (N_12214,N_6707,N_11449);
or U12215 (N_12215,N_11051,N_8183);
or U12216 (N_12216,N_10387,N_8783);
and U12217 (N_12217,N_9984,N_7658);
xnor U12218 (N_12218,N_11774,N_6984);
and U12219 (N_12219,N_7185,N_10015);
and U12220 (N_12220,N_9990,N_7615);
xor U12221 (N_12221,N_8651,N_9715);
and U12222 (N_12222,N_9469,N_6933);
or U12223 (N_12223,N_6796,N_11928);
nor U12224 (N_12224,N_7704,N_11427);
nand U12225 (N_12225,N_6531,N_10017);
nor U12226 (N_12226,N_9387,N_10224);
and U12227 (N_12227,N_7220,N_11214);
and U12228 (N_12228,N_7736,N_8908);
nor U12229 (N_12229,N_10767,N_11311);
or U12230 (N_12230,N_9171,N_7143);
nor U12231 (N_12231,N_7647,N_7343);
and U12232 (N_12232,N_6230,N_8696);
and U12233 (N_12233,N_7591,N_6881);
nor U12234 (N_12234,N_10051,N_8321);
nand U12235 (N_12235,N_11419,N_9843);
nor U12236 (N_12236,N_9985,N_6117);
nor U12237 (N_12237,N_10944,N_8913);
or U12238 (N_12238,N_7419,N_8442);
nor U12239 (N_12239,N_7657,N_6977);
xnor U12240 (N_12240,N_11152,N_7226);
and U12241 (N_12241,N_10049,N_6692);
nor U12242 (N_12242,N_8945,N_9050);
nand U12243 (N_12243,N_8983,N_9627);
or U12244 (N_12244,N_8220,N_11828);
and U12245 (N_12245,N_9124,N_7087);
nor U12246 (N_12246,N_6569,N_11609);
nand U12247 (N_12247,N_11489,N_11179);
nand U12248 (N_12248,N_6572,N_10194);
xnor U12249 (N_12249,N_11149,N_7031);
xnor U12250 (N_12250,N_8416,N_7364);
or U12251 (N_12251,N_9098,N_6265);
or U12252 (N_12252,N_7326,N_11135);
or U12253 (N_12253,N_10620,N_6900);
nand U12254 (N_12254,N_8029,N_11731);
or U12255 (N_12255,N_8571,N_10485);
xnor U12256 (N_12256,N_6555,N_7222);
and U12257 (N_12257,N_8045,N_10585);
xor U12258 (N_12258,N_7911,N_10951);
nor U12259 (N_12259,N_9952,N_7329);
and U12260 (N_12260,N_9562,N_10692);
or U12261 (N_12261,N_8773,N_8329);
nand U12262 (N_12262,N_7386,N_8487);
nand U12263 (N_12263,N_10792,N_10769);
xnor U12264 (N_12264,N_8277,N_11383);
and U12265 (N_12265,N_9707,N_10060);
nor U12266 (N_12266,N_11627,N_7502);
nor U12267 (N_12267,N_10395,N_9445);
and U12268 (N_12268,N_10376,N_10477);
or U12269 (N_12269,N_8947,N_6702);
or U12270 (N_12270,N_6248,N_10181);
or U12271 (N_12271,N_9316,N_11283);
xor U12272 (N_12272,N_6479,N_7123);
and U12273 (N_12273,N_11742,N_10968);
nand U12274 (N_12274,N_6457,N_9733);
xnor U12275 (N_12275,N_10932,N_9557);
xor U12276 (N_12276,N_10677,N_11148);
xnor U12277 (N_12277,N_10458,N_7439);
xnor U12278 (N_12278,N_10952,N_9564);
and U12279 (N_12279,N_8728,N_7315);
xor U12280 (N_12280,N_9288,N_11931);
and U12281 (N_12281,N_7297,N_10554);
nand U12282 (N_12282,N_6120,N_11351);
nand U12283 (N_12283,N_10488,N_11478);
nor U12284 (N_12284,N_10992,N_9964);
and U12285 (N_12285,N_11490,N_8901);
xnor U12286 (N_12286,N_8965,N_6492);
nor U12287 (N_12287,N_9462,N_9729);
xor U12288 (N_12288,N_8054,N_6347);
nor U12289 (N_12289,N_6845,N_11726);
or U12290 (N_12290,N_9467,N_8400);
and U12291 (N_12291,N_11592,N_6880);
nor U12292 (N_12292,N_11373,N_11814);
nor U12293 (N_12293,N_6106,N_10154);
or U12294 (N_12294,N_11369,N_9628);
or U12295 (N_12295,N_10758,N_7763);
nor U12296 (N_12296,N_8439,N_6631);
xor U12297 (N_12297,N_7490,N_11207);
and U12298 (N_12298,N_6199,N_10158);
nand U12299 (N_12299,N_9759,N_6417);
or U12300 (N_12300,N_11267,N_10880);
nor U12301 (N_12301,N_11472,N_6611);
or U12302 (N_12302,N_10962,N_9958);
nand U12303 (N_12303,N_9568,N_6617);
and U12304 (N_12304,N_6144,N_6680);
and U12305 (N_12305,N_10197,N_9405);
or U12306 (N_12306,N_11990,N_6383);
xnor U12307 (N_12307,N_8251,N_11981);
xor U12308 (N_12308,N_10102,N_9027);
or U12309 (N_12309,N_6018,N_6823);
or U12310 (N_12310,N_10296,N_10725);
xor U12311 (N_12311,N_10334,N_9613);
nand U12312 (N_12312,N_9230,N_11792);
and U12313 (N_12313,N_6770,N_8660);
and U12314 (N_12314,N_11584,N_6790);
xnor U12315 (N_12315,N_7309,N_11751);
nand U12316 (N_12316,N_11728,N_7433);
and U12317 (N_12317,N_11959,N_6319);
nand U12318 (N_12318,N_11316,N_11971);
or U12319 (N_12319,N_9943,N_8503);
or U12320 (N_12320,N_9172,N_9695);
xnor U12321 (N_12321,N_7155,N_8909);
or U12322 (N_12322,N_8994,N_6780);
nand U12323 (N_12323,N_11037,N_6044);
xor U12324 (N_12324,N_8762,N_6768);
and U12325 (N_12325,N_8602,N_7348);
xnor U12326 (N_12326,N_9318,N_9202);
xor U12327 (N_12327,N_8995,N_9374);
and U12328 (N_12328,N_10326,N_10825);
nand U12329 (N_12329,N_10143,N_10575);
or U12330 (N_12330,N_9481,N_9475);
nor U12331 (N_12331,N_10937,N_10675);
nand U12332 (N_12332,N_6255,N_10111);
nand U12333 (N_12333,N_7880,N_11442);
nand U12334 (N_12334,N_6140,N_8271);
and U12335 (N_12335,N_11446,N_10335);
nand U12336 (N_12336,N_9454,N_10058);
nor U12337 (N_12337,N_10200,N_6012);
nor U12338 (N_12338,N_11704,N_6127);
and U12339 (N_12339,N_11301,N_6473);
xor U12340 (N_12340,N_9015,N_8415);
xor U12341 (N_12341,N_8673,N_11696);
and U12342 (N_12342,N_10985,N_6029);
xnor U12343 (N_12343,N_7157,N_10849);
nor U12344 (N_12344,N_8030,N_7129);
or U12345 (N_12345,N_10628,N_7568);
or U12346 (N_12346,N_8757,N_6892);
or U12347 (N_12347,N_9427,N_6419);
and U12348 (N_12348,N_11902,N_8560);
nor U12349 (N_12349,N_9041,N_9972);
and U12350 (N_12350,N_7001,N_6589);
nand U12351 (N_12351,N_6476,N_6399);
xnor U12352 (N_12352,N_8840,N_8134);
nor U12353 (N_12353,N_11646,N_7359);
nor U12354 (N_12354,N_9689,N_6490);
xnor U12355 (N_12355,N_11407,N_8023);
nor U12356 (N_12356,N_10950,N_6551);
or U12357 (N_12357,N_7018,N_9804);
and U12358 (N_12358,N_6883,N_6902);
xor U12359 (N_12359,N_6313,N_11762);
and U12360 (N_12360,N_9827,N_9709);
nand U12361 (N_12361,N_7097,N_6240);
and U12362 (N_12362,N_9931,N_9642);
xnor U12363 (N_12363,N_11935,N_11676);
nand U12364 (N_12364,N_10664,N_8974);
or U12365 (N_12365,N_9645,N_10439);
or U12366 (N_12366,N_6480,N_10148);
xor U12367 (N_12367,N_6954,N_10790);
xnor U12368 (N_12368,N_9538,N_6773);
or U12369 (N_12369,N_10161,N_11502);
and U12370 (N_12370,N_8411,N_10121);
nand U12371 (N_12371,N_7512,N_6947);
nand U12372 (N_12372,N_11323,N_11901);
xnor U12373 (N_12373,N_9660,N_11541);
nand U12374 (N_12374,N_10946,N_10212);
xor U12375 (N_12375,N_8482,N_7995);
and U12376 (N_12376,N_10381,N_9136);
or U12377 (N_12377,N_9806,N_11864);
nand U12378 (N_12378,N_8971,N_11177);
xnor U12379 (N_12379,N_6262,N_7128);
and U12380 (N_12380,N_6483,N_9247);
and U12381 (N_12381,N_10260,N_6534);
or U12382 (N_12382,N_8569,N_8734);
and U12383 (N_12383,N_6001,N_10023);
nand U12384 (N_12384,N_6581,N_7284);
and U12385 (N_12385,N_7681,N_7522);
and U12386 (N_12386,N_7667,N_11385);
nand U12387 (N_12387,N_9128,N_11785);
xor U12388 (N_12388,N_8025,N_10857);
nor U12389 (N_12389,N_7058,N_6224);
or U12390 (N_12390,N_9070,N_6194);
and U12391 (N_12391,N_7196,N_6955);
or U12392 (N_12392,N_11980,N_11171);
xor U12393 (N_12393,N_6981,N_10779);
nor U12394 (N_12394,N_10004,N_6958);
xnor U12395 (N_12395,N_11544,N_8430);
xor U12396 (N_12396,N_8144,N_9812);
nor U12397 (N_12397,N_8816,N_8441);
and U12398 (N_12398,N_9418,N_11813);
nor U12399 (N_12399,N_7887,N_6325);
nand U12400 (N_12400,N_6504,N_8280);
xor U12401 (N_12401,N_11559,N_10660);
nand U12402 (N_12402,N_8214,N_6340);
or U12403 (N_12403,N_7033,N_6036);
and U12404 (N_12404,N_10771,N_8261);
nor U12405 (N_12405,N_8058,N_7025);
nor U12406 (N_12406,N_7413,N_7088);
nand U12407 (N_12407,N_6757,N_7347);
nor U12408 (N_12408,N_10634,N_7021);
nand U12409 (N_12409,N_11191,N_11049);
nand U12410 (N_12410,N_11043,N_7267);
nor U12411 (N_12411,N_7341,N_9190);
or U12412 (N_12412,N_9039,N_7679);
or U12413 (N_12413,N_11367,N_8981);
nand U12414 (N_12414,N_6663,N_7545);
nor U12415 (N_12415,N_11963,N_11572);
nand U12416 (N_12416,N_6887,N_6939);
xor U12417 (N_12417,N_10105,N_8274);
nor U12418 (N_12418,N_7424,N_10802);
xnor U12419 (N_12419,N_10645,N_9540);
or U12420 (N_12420,N_8309,N_7559);
or U12421 (N_12421,N_11938,N_6243);
xor U12422 (N_12422,N_9902,N_11258);
xor U12423 (N_12423,N_9381,N_7144);
nand U12424 (N_12424,N_11914,N_6777);
or U12425 (N_12425,N_10796,N_10855);
or U12426 (N_12426,N_9169,N_8722);
nand U12427 (N_12427,N_7987,N_7254);
xor U12428 (N_12428,N_10282,N_7769);
and U12429 (N_12429,N_11477,N_7428);
and U12430 (N_12430,N_10164,N_7785);
nand U12431 (N_12431,N_9504,N_6918);
nand U12432 (N_12432,N_8238,N_8268);
nand U12433 (N_12433,N_6351,N_8992);
or U12434 (N_12434,N_8610,N_6341);
or U12435 (N_12435,N_6885,N_9727);
xor U12436 (N_12436,N_9770,N_11885);
nor U12437 (N_12437,N_7426,N_7039);
nor U12438 (N_12438,N_8157,N_7320);
nor U12439 (N_12439,N_10256,N_11459);
nor U12440 (N_12440,N_7305,N_11569);
and U12441 (N_12441,N_6400,N_8827);
nor U12442 (N_12442,N_8702,N_8778);
xnor U12443 (N_12443,N_11228,N_11336);
nand U12444 (N_12444,N_6643,N_6263);
nand U12445 (N_12445,N_9139,N_6466);
xor U12446 (N_12446,N_7011,N_11382);
or U12447 (N_12447,N_8622,N_10528);
nor U12448 (N_12448,N_7022,N_6063);
xor U12449 (N_12449,N_9197,N_8880);
nand U12450 (N_12450,N_8800,N_11747);
nor U12451 (N_12451,N_6437,N_7788);
xnor U12452 (N_12452,N_9842,N_9000);
nand U12453 (N_12453,N_10516,N_10742);
nor U12454 (N_12454,N_8422,N_7870);
nand U12455 (N_12455,N_8489,N_6201);
and U12456 (N_12456,N_9704,N_10043);
and U12457 (N_12457,N_10353,N_9385);
xor U12458 (N_12458,N_10703,N_10211);
xnor U12459 (N_12459,N_8326,N_10208);
xor U12460 (N_12460,N_10887,N_9257);
xnor U12461 (N_12461,N_10191,N_10330);
xor U12462 (N_12462,N_6566,N_7955);
nor U12463 (N_12463,N_7919,N_6497);
nor U12464 (N_12464,N_10089,N_7524);
xor U12465 (N_12465,N_8742,N_9130);
xnor U12466 (N_12466,N_9711,N_7377);
nor U12467 (N_12467,N_11601,N_11325);
or U12468 (N_12468,N_6307,N_6826);
xnor U12469 (N_12469,N_8850,N_9292);
nor U12470 (N_12470,N_7997,N_10739);
nand U12471 (N_12471,N_7556,N_6629);
nand U12472 (N_12472,N_7187,N_8339);
and U12473 (N_12473,N_10989,N_7332);
xor U12474 (N_12474,N_7047,N_10278);
nand U12475 (N_12475,N_6785,N_6026);
xor U12476 (N_12476,N_8942,N_9231);
or U12477 (N_12477,N_6915,N_9476);
xor U12478 (N_12478,N_9233,N_11353);
and U12479 (N_12479,N_6907,N_10393);
nor U12480 (N_12480,N_11512,N_6300);
nor U12481 (N_12481,N_6416,N_10341);
nand U12482 (N_12482,N_9250,N_10349);
xnor U12483 (N_12483,N_10510,N_11168);
nor U12484 (N_12484,N_6519,N_11247);
and U12485 (N_12485,N_8438,N_6728);
or U12486 (N_12486,N_6435,N_6914);
xnor U12487 (N_12487,N_8266,N_11469);
or U12488 (N_12488,N_10636,N_8922);
nand U12489 (N_12489,N_11438,N_8944);
xnor U12490 (N_12490,N_6851,N_6573);
or U12491 (N_12491,N_9555,N_9137);
xnor U12492 (N_12492,N_6684,N_7569);
or U12493 (N_12493,N_11067,N_7612);
xnor U12494 (N_12494,N_11540,N_11327);
or U12495 (N_12495,N_10569,N_9364);
or U12496 (N_12496,N_6438,N_7100);
and U12497 (N_12497,N_11516,N_6676);
xnor U12498 (N_12498,N_6987,N_10374);
nand U12499 (N_12499,N_9080,N_8026);
or U12500 (N_12500,N_11416,N_10574);
or U12501 (N_12501,N_9441,N_7441);
and U12502 (N_12502,N_6060,N_11899);
and U12503 (N_12503,N_8726,N_7091);
and U12504 (N_12504,N_11256,N_7504);
and U12505 (N_12505,N_11209,N_7694);
nand U12506 (N_12506,N_8769,N_7869);
and U12507 (N_12507,N_10274,N_11766);
xor U12508 (N_12508,N_7581,N_6276);
or U12509 (N_12509,N_10608,N_6428);
xor U12510 (N_12510,N_7360,N_11966);
or U12511 (N_12511,N_6087,N_11968);
xor U12512 (N_12512,N_11337,N_10233);
xor U12513 (N_12513,N_9513,N_10815);
and U12514 (N_12514,N_9822,N_10958);
or U12515 (N_12515,N_8832,N_8525);
xor U12516 (N_12516,N_6587,N_7582);
nand U12517 (N_12517,N_9828,N_8636);
xor U12518 (N_12518,N_8278,N_10945);
xnor U12519 (N_12519,N_8225,N_9313);
nand U12520 (N_12520,N_7683,N_11432);
and U12521 (N_12521,N_9432,N_10774);
and U12522 (N_12522,N_6477,N_8518);
and U12523 (N_12523,N_8970,N_7194);
xnor U12524 (N_12524,N_11651,N_7864);
nand U12525 (N_12525,N_9067,N_9413);
nand U12526 (N_12526,N_9760,N_6545);
and U12527 (N_12527,N_10166,N_6041);
nor U12528 (N_12528,N_7285,N_10502);
and U12529 (N_12529,N_9437,N_10423);
nand U12530 (N_12530,N_6983,N_6339);
or U12531 (N_12531,N_11437,N_11831);
or U12532 (N_12532,N_8883,N_8016);
and U12533 (N_12533,N_8703,N_11736);
nor U12534 (N_12534,N_6333,N_8476);
nor U12535 (N_12535,N_6456,N_9341);
xor U12536 (N_12536,N_8040,N_7850);
and U12537 (N_12537,N_6565,N_9068);
nor U12538 (N_12538,N_10008,N_9419);
xor U12539 (N_12539,N_6733,N_8657);
and U12540 (N_12540,N_7463,N_8745);
nor U12541 (N_12541,N_10276,N_7132);
and U12542 (N_12542,N_9520,N_10639);
and U12543 (N_12543,N_11823,N_10063);
and U12544 (N_12544,N_9126,N_8820);
or U12545 (N_12545,N_8048,N_6371);
nor U12546 (N_12546,N_7002,N_9951);
nor U12547 (N_12547,N_10306,N_8894);
nand U12548 (N_12548,N_6148,N_6521);
and U12549 (N_12549,N_10474,N_11724);
nor U12550 (N_12550,N_6487,N_6562);
and U12551 (N_12551,N_8363,N_8043);
nor U12552 (N_12552,N_6927,N_11716);
nand U12553 (N_12553,N_11176,N_8240);
nand U12554 (N_12554,N_8998,N_11666);
nand U12555 (N_12555,N_10680,N_10559);
nand U12556 (N_12556,N_9356,N_7575);
nor U12557 (N_12557,N_7375,N_9163);
and U12558 (N_12558,N_6205,N_10493);
nand U12559 (N_12559,N_11216,N_6679);
xor U12560 (N_12560,N_7110,N_6213);
and U12561 (N_12561,N_7227,N_9755);
or U12562 (N_12562,N_9639,N_7770);
or U12563 (N_12563,N_9925,N_8870);
xor U12564 (N_12564,N_11605,N_9741);
and U12565 (N_12565,N_7302,N_9503);
nor U12566 (N_12566,N_7611,N_9062);
nor U12567 (N_12567,N_9084,N_10515);
nand U12568 (N_12568,N_11547,N_8233);
xnor U12569 (N_12569,N_6336,N_7420);
or U12570 (N_12570,N_7561,N_9542);
xnor U12571 (N_12571,N_10238,N_10473);
nor U12572 (N_12572,N_10241,N_7092);
nand U12573 (N_12573,N_9010,N_8083);
nand U12574 (N_12574,N_6494,N_7884);
nand U12575 (N_12575,N_9763,N_7689);
xor U12576 (N_12576,N_6257,N_11169);
or U12577 (N_12577,N_11003,N_10272);
nor U12578 (N_12578,N_6086,N_9798);
nand U12579 (N_12579,N_9866,N_11272);
xnor U12580 (N_12580,N_11860,N_6268);
nand U12581 (N_12581,N_6168,N_10470);
xor U12582 (N_12582,N_9042,N_7624);
nand U12583 (N_12583,N_9487,N_9658);
and U12584 (N_12584,N_6953,N_11652);
nand U12585 (N_12585,N_9040,N_7478);
nor U12586 (N_12586,N_7178,N_8364);
nand U12587 (N_12587,N_11720,N_11947);
nor U12588 (N_12588,N_6868,N_11110);
xor U12589 (N_12589,N_7161,N_10593);
or U12590 (N_12590,N_7567,N_9366);
or U12591 (N_12591,N_8706,N_9991);
xnor U12592 (N_12592,N_9332,N_8650);
xor U12593 (N_12593,N_6838,N_7715);
or U12594 (N_12594,N_6059,N_8481);
or U12595 (N_12595,N_8406,N_7056);
or U12596 (N_12596,N_11404,N_10797);
or U12597 (N_12597,N_7295,N_9121);
xnor U12598 (N_12598,N_11299,N_7889);
xnor U12599 (N_12599,N_9048,N_10509);
xor U12600 (N_12600,N_6231,N_8155);
or U12601 (N_12601,N_11918,N_6301);
and U12602 (N_12602,N_8808,N_7718);
nand U12603 (N_12603,N_6675,N_7742);
nor U12604 (N_12604,N_11024,N_11172);
xor U12605 (N_12605,N_7705,N_10209);
or U12606 (N_12606,N_11264,N_11492);
nand U12607 (N_12607,N_10449,N_8924);
or U12608 (N_12608,N_10451,N_6714);
nor U12609 (N_12609,N_8383,N_11362);
and U12610 (N_12610,N_8260,N_9301);
and U12611 (N_12611,N_11941,N_7952);
nor U12612 (N_12612,N_11689,N_8230);
or U12613 (N_12613,N_11355,N_6260);
and U12614 (N_12614,N_11005,N_8325);
or U12615 (N_12615,N_9929,N_7835);
nand U12616 (N_12616,N_10438,N_6781);
or U12617 (N_12617,N_8836,N_8100);
xor U12618 (N_12618,N_10481,N_10602);
nor U12619 (N_12619,N_8279,N_8597);
xor U12620 (N_12620,N_6115,N_7328);
or U12621 (N_12621,N_11221,N_11894);
or U12622 (N_12622,N_6342,N_9485);
xnor U12623 (N_12623,N_10651,N_9948);
nand U12624 (N_12624,N_11888,N_8055);
or U12625 (N_12625,N_11713,N_11878);
nor U12626 (N_12626,N_11589,N_8929);
or U12627 (N_12627,N_7412,N_10751);
and U12628 (N_12628,N_6420,N_9594);
and U12629 (N_12629,N_9295,N_8234);
or U12630 (N_12630,N_6119,N_11805);
xor U12631 (N_12631,N_6185,N_8725);
or U12632 (N_12632,N_7875,N_9162);
or U12633 (N_12633,N_9009,N_10924);
and U12634 (N_12634,N_11238,N_7505);
nand U12635 (N_12635,N_11359,N_8739);
nor U12636 (N_12636,N_6475,N_8685);
and U12637 (N_12637,N_9092,N_9498);
or U12638 (N_12638,N_7073,N_9205);
xnor U12639 (N_12639,N_10504,N_11170);
and U12640 (N_12640,N_11006,N_11760);
xnor U12641 (N_12641,N_10844,N_9100);
nor U12642 (N_12642,N_8581,N_7517);
nor U12643 (N_12643,N_7914,N_6748);
xor U12644 (N_12644,N_7594,N_7099);
xnor U12645 (N_12645,N_9662,N_6661);
or U12646 (N_12646,N_9337,N_7818);
nor U12647 (N_12647,N_11983,N_10879);
nand U12648 (N_12648,N_6935,N_11346);
or U12649 (N_12649,N_8307,N_9056);
nand U12650 (N_12650,N_9335,N_9983);
nor U12651 (N_12651,N_8410,N_7450);
nand U12652 (N_12652,N_8561,N_8129);
and U12653 (N_12653,N_7749,N_7346);
or U12654 (N_12654,N_7482,N_7133);
xnor U12655 (N_12655,N_9410,N_6172);
nand U12656 (N_12656,N_9889,N_7758);
or U12657 (N_12657,N_9508,N_6865);
and U12658 (N_12658,N_10316,N_10722);
and U12659 (N_12659,N_6429,N_6567);
nor U12660 (N_12660,N_11420,N_6583);
nor U12661 (N_12661,N_11710,N_9107);
or U12662 (N_12662,N_8502,N_7263);
nand U12663 (N_12663,N_8967,N_10610);
and U12664 (N_12664,N_10567,N_11780);
nand U12665 (N_12665,N_7977,N_6304);
xor U12666 (N_12666,N_8246,N_9681);
nor U12667 (N_12667,N_9488,N_7041);
or U12668 (N_12668,N_9637,N_11686);
nand U12669 (N_12669,N_8858,N_10428);
nand U12670 (N_12670,N_9758,N_9864);
nor U12671 (N_12671,N_10357,N_11638);
and U12672 (N_12672,N_8512,N_9722);
or U12673 (N_12673,N_9908,N_6258);
and U12674 (N_12674,N_9320,N_10617);
xor U12675 (N_12675,N_8599,N_6793);
nor U12676 (N_12676,N_11620,N_8844);
or U12677 (N_12677,N_10794,N_6645);
xnor U12678 (N_12678,N_11026,N_10899);
nor U12679 (N_12679,N_6251,N_6649);
xor U12680 (N_12680,N_10972,N_8049);
and U12681 (N_12681,N_11987,N_10858);
nor U12682 (N_12682,N_7492,N_7391);
and U12683 (N_12683,N_10123,N_7633);
and U12684 (N_12684,N_9807,N_9584);
nand U12685 (N_12685,N_10196,N_10538);
and U12686 (N_12686,N_6852,N_6112);
and U12687 (N_12687,N_8452,N_6458);
nand U12688 (N_12688,N_8419,N_10970);
and U12689 (N_12689,N_9001,N_9726);
xor U12690 (N_12690,N_11457,N_10993);
nor U12691 (N_12691,N_6208,N_11368);
xor U12692 (N_12692,N_10782,N_9914);
xnor U12693 (N_12693,N_9428,N_11131);
nor U12694 (N_12694,N_6815,N_7960);
nand U12695 (N_12695,N_9813,N_10957);
and U12696 (N_12696,N_10686,N_8148);
nor U12697 (N_12697,N_7324,N_9757);
nand U12698 (N_12698,N_8991,N_7009);
or U12699 (N_12699,N_8450,N_9344);
or U12700 (N_12700,N_7060,N_7685);
or U12701 (N_12701,N_7537,N_6975);
or U12702 (N_12702,N_11077,N_9305);
or U12703 (N_12703,N_7158,N_8127);
or U12704 (N_12704,N_8138,N_6666);
xor U12705 (N_12705,N_6053,N_8815);
and U12706 (N_12706,N_10812,N_6615);
and U12707 (N_12707,N_7005,N_7398);
nor U12708 (N_12708,N_6306,N_8130);
nand U12709 (N_12709,N_11846,N_9705);
nor U12710 (N_12710,N_10582,N_9302);
and U12711 (N_12711,N_8455,N_11522);
xnor U12712 (N_12712,N_9949,N_9123);
nor U12713 (N_12713,N_9291,N_8903);
or U12714 (N_12714,N_11839,N_7101);
or U12715 (N_12715,N_11772,N_7230);
and U12716 (N_12716,N_8665,N_8131);
or U12717 (N_12717,N_6363,N_6966);
or U12718 (N_12718,N_11232,N_7755);
and U12719 (N_12719,N_10459,N_11555);
or U12720 (N_12720,N_6376,N_10391);
and U12721 (N_12721,N_10611,N_9650);
nor U12722 (N_12722,N_9815,N_11259);
nand U12723 (N_12723,N_11042,N_11009);
nor U12724 (N_12724,N_7065,N_6909);
nand U12725 (N_12725,N_8499,N_11872);
nand U12726 (N_12726,N_11236,N_11687);
or U12727 (N_12727,N_10359,N_10317);
nor U12728 (N_12728,N_10400,N_6093);
and U12729 (N_12729,N_11140,N_11701);
nor U12730 (N_12730,N_7860,N_7898);
or U12731 (N_12731,N_10213,N_9213);
xor U12732 (N_12732,N_8878,N_6183);
nand U12733 (N_12733,N_6031,N_8368);
and U12734 (N_12734,N_7616,N_10119);
nor U12735 (N_12735,N_7003,N_10440);
or U12736 (N_12736,N_9906,N_7514);
nand U12737 (N_12737,N_11215,N_11621);
nand U12738 (N_12738,N_10864,N_7675);
nand U12739 (N_12739,N_6422,N_11546);
nand U12740 (N_12740,N_11029,N_10258);
or U12741 (N_12741,N_8318,N_8831);
and U12742 (N_12742,N_7649,N_11119);
nand U12743 (N_12743,N_9468,N_9380);
or U12744 (N_12744,N_6223,N_7654);
xor U12745 (N_12745,N_9082,N_7477);
or U12746 (N_12746,N_10814,N_7549);
nor U12747 (N_12747,N_9053,N_6929);
or U12748 (N_12748,N_7396,N_7935);
and U12749 (N_12749,N_11849,N_11750);
nor U12750 (N_12750,N_10925,N_7406);
nor U12751 (N_12751,N_9992,N_6832);
nand U12752 (N_12752,N_11429,N_7281);
nand U12753 (N_12753,N_11142,N_8197);
nand U12754 (N_12754,N_7044,N_6067);
and U12755 (N_12755,N_7663,N_8504);
or U12756 (N_12756,N_9449,N_10707);
and U12757 (N_12757,N_8408,N_10009);
xnor U12758 (N_12758,N_10412,N_10752);
nor U12759 (N_12759,N_6329,N_7824);
or U12760 (N_12760,N_8491,N_11085);
and U12761 (N_12761,N_9342,N_10709);
nand U12762 (N_12762,N_7479,N_7125);
or U12763 (N_12763,N_7713,N_10484);
xor U12764 (N_12764,N_8194,N_9880);
nor U12765 (N_12765,N_8295,N_6241);
and U12766 (N_12766,N_7029,N_10476);
nand U12767 (N_12767,N_6065,N_10524);
nor U12768 (N_12768,N_11753,N_6831);
or U12769 (N_12769,N_8635,N_9456);
xor U12770 (N_12770,N_11518,N_10726);
or U12771 (N_12771,N_8592,N_9730);
nor U12772 (N_12772,N_11358,N_8388);
and U12773 (N_12773,N_9640,N_7476);
nand U12774 (N_12774,N_9553,N_10118);
xor U12775 (N_12775,N_11571,N_8258);
and U12776 (N_12776,N_9141,N_11334);
xor U12777 (N_12777,N_6125,N_9928);
or U12778 (N_12778,N_6735,N_10319);
or U12779 (N_12779,N_8079,N_8857);
nand U12780 (N_12780,N_9491,N_7965);
nand U12781 (N_12781,N_11333,N_11206);
nor U12782 (N_12782,N_6651,N_10843);
nand U12783 (N_12783,N_11059,N_7949);
nor U12784 (N_12784,N_10615,N_9281);
or U12785 (N_12785,N_6017,N_11809);
and U12786 (N_12786,N_9699,N_9754);
and U12787 (N_12787,N_6621,N_6791);
and U12788 (N_12788,N_10984,N_6343);
or U12789 (N_12789,N_6980,N_11661);
or U12790 (N_12790,N_11591,N_10715);
nor U12791 (N_12791,N_9083,N_7557);
xor U12792 (N_12792,N_11321,N_6352);
nand U12793 (N_12793,N_10541,N_9037);
and U12794 (N_12794,N_10409,N_11767);
nor U12795 (N_12795,N_11098,N_8074);
nor U12796 (N_12796,N_11629,N_6049);
nand U12797 (N_12797,N_6898,N_10991);
nor U12798 (N_12798,N_8937,N_10838);
and U12799 (N_12799,N_6664,N_7454);
nand U12800 (N_12800,N_10532,N_8113);
or U12801 (N_12801,N_10922,N_7225);
and U12802 (N_12802,N_9057,N_8603);
and U12803 (N_12803,N_9151,N_10998);
or U12804 (N_12804,N_10505,N_11797);
nor U12805 (N_12805,N_9717,N_11628);
nand U12806 (N_12806,N_8373,N_9576);
nand U12807 (N_12807,N_7282,N_8588);
nor U12808 (N_12808,N_9207,N_11260);
nor U12809 (N_12809,N_6324,N_6653);
or U12810 (N_12810,N_9706,N_8024);
nor U12811 (N_12811,N_11579,N_11277);
and U12812 (N_12812,N_6974,N_10090);
and U12813 (N_12813,N_11280,N_7798);
nor U12814 (N_12814,N_9024,N_10916);
nand U12815 (N_12815,N_11357,N_6925);
xor U12816 (N_12816,N_9712,N_11365);
nor U12817 (N_12817,N_8361,N_11147);
nor U12818 (N_12818,N_9459,N_11433);
nor U12819 (N_12819,N_6212,N_6379);
nor U12820 (N_12820,N_6516,N_8933);
xnor U12821 (N_12821,N_8584,N_10137);
or U12822 (N_12822,N_8395,N_7563);
xor U12823 (N_12823,N_10783,N_8950);
and U12824 (N_12824,N_11391,N_6149);
xor U12825 (N_12825,N_11428,N_7808);
or U12826 (N_12826,N_7757,N_8705);
nand U12827 (N_12827,N_7336,N_8104);
and U12828 (N_12828,N_7393,N_6222);
or U12829 (N_12829,N_7270,N_6056);
and U12830 (N_12830,N_10734,N_10215);
xor U12831 (N_12831,N_10227,N_11513);
nand U12832 (N_12832,N_6712,N_9809);
xor U12833 (N_12833,N_10067,N_6266);
or U12834 (N_12834,N_11958,N_6283);
xnor U12835 (N_12835,N_11536,N_10874);
xnor U12836 (N_12836,N_9319,N_6131);
nor U12837 (N_12837,N_8212,N_6170);
xor U12838 (N_12838,N_6330,N_7485);
xnor U12839 (N_12839,N_6628,N_7598);
nor U12840 (N_12840,N_7127,N_10555);
nor U12841 (N_12841,N_7560,N_6096);
nor U12842 (N_12842,N_6111,N_11994);
xnor U12843 (N_12843,N_6606,N_10262);
and U12844 (N_12844,N_6278,N_8243);
xnor U12845 (N_12845,N_11349,N_8035);
and U12846 (N_12846,N_7636,N_8907);
xnor U12847 (N_12847,N_6292,N_8172);
nor U12848 (N_12848,N_10337,N_6235);
xnor U12849 (N_12849,N_10913,N_11242);
and U12850 (N_12850,N_8010,N_6275);
or U12851 (N_12851,N_9732,N_10983);
and U12852 (N_12852,N_8353,N_9811);
or U12853 (N_12853,N_10601,N_9966);
and U12854 (N_12854,N_8159,N_7917);
and U12855 (N_12855,N_8227,N_7578);
nand U12856 (N_12856,N_8577,N_10304);
or U12857 (N_12857,N_8145,N_6190);
xor U12858 (N_12858,N_6518,N_6959);
or U12859 (N_12859,N_10198,N_10182);
xor U12860 (N_12860,N_8544,N_9816);
xor U12861 (N_12861,N_7138,N_10325);
or U12862 (N_12862,N_9887,N_10152);
nor U12863 (N_12863,N_11164,N_6375);
and U12864 (N_12864,N_6299,N_9031);
nand U12865 (N_12865,N_8578,N_6270);
xor U12866 (N_12866,N_10003,N_9836);
nand U12867 (N_12867,N_9430,N_10609);
nand U12868 (N_12868,N_8765,N_11845);
nand U12869 (N_12869,N_9178,N_11717);
nor U12870 (N_12870,N_6731,N_7334);
nor U12871 (N_12871,N_11339,N_6050);
nand U12872 (N_12872,N_6601,N_6390);
xnor U12873 (N_12873,N_9382,N_6028);
and U12874 (N_12874,N_7520,N_8861);
nor U12875 (N_12875,N_9634,N_9044);
or U12876 (N_12876,N_9668,N_7152);
nor U12877 (N_12877,N_11632,N_9738);
and U12878 (N_12878,N_9187,N_11685);
and U12879 (N_12879,N_7200,N_11294);
and U12880 (N_12880,N_6159,N_6698);
nor U12881 (N_12881,N_9489,N_10128);
xor U12882 (N_12882,N_9377,N_8235);
xnor U12883 (N_12883,N_7696,N_8714);
nor U12884 (N_12884,N_11203,N_6740);
and U12885 (N_12885,N_8724,N_9072);
nand U12886 (N_12886,N_8807,N_8801);
nor U12887 (N_12887,N_10550,N_8846);
or U12888 (N_12888,N_11910,N_10867);
nor U12889 (N_12889,N_8663,N_6048);
nand U12890 (N_12890,N_7858,N_6334);
and U12891 (N_12891,N_11759,N_10046);
or U12892 (N_12892,N_7523,N_8604);
or U12893 (N_12893,N_10919,N_10630);
and U12894 (N_12894,N_6046,N_7941);
xor U12895 (N_12895,N_7974,N_11583);
nand U12896 (N_12896,N_8695,N_7827);
and U12897 (N_12897,N_9993,N_11607);
or U12898 (N_12898,N_8374,N_7380);
and U12899 (N_12899,N_7822,N_9938);
nand U12900 (N_12900,N_6030,N_9277);
nand U12901 (N_12901,N_11798,N_7286);
nand U12902 (N_12902,N_6574,N_10522);
or U12903 (N_12903,N_8961,N_9184);
xnor U12904 (N_12904,N_7817,N_8862);
nand U12905 (N_12905,N_9773,N_11233);
xor U12906 (N_12906,N_8473,N_11298);
nand U12907 (N_12907,N_7868,N_10527);
nor U12908 (N_12908,N_7182,N_11827);
nand U12909 (N_12909,N_9633,N_11905);
and U12910 (N_12910,N_10905,N_10851);
and U12911 (N_12911,N_7076,N_10070);
and U12912 (N_12912,N_6948,N_9268);
or U12913 (N_12913,N_6441,N_7233);
nand U12914 (N_12914,N_7855,N_7756);
nand U12915 (N_12915,N_10418,N_8869);
nand U12916 (N_12916,N_9978,N_8871);
xor U12917 (N_12917,N_11338,N_9654);
or U12918 (N_12918,N_6286,N_8445);
nand U12919 (N_12919,N_9526,N_11379);
nand U12920 (N_12920,N_10906,N_9198);
nor U12921 (N_12921,N_11771,N_6840);
nand U12922 (N_12922,N_9857,N_7802);
or U12923 (N_12923,N_6920,N_6052);
and U12924 (N_12924,N_8292,N_9223);
or U12925 (N_12925,N_8989,N_11310);
xor U12926 (N_12926,N_9293,N_6411);
nand U12927 (N_12927,N_9312,N_10175);
or U12928 (N_12928,N_8791,N_10577);
or U12929 (N_12929,N_9980,N_8732);
or U12930 (N_12930,N_8864,N_10205);
or U12931 (N_12931,N_7629,N_8316);
or U12932 (N_12932,N_6696,N_11450);
nor U12933 (N_12933,N_6510,N_8885);
xor U12934 (N_12934,N_7388,N_6743);
nand U12935 (N_12935,N_11486,N_6844);
xnor U12936 (N_12936,N_8263,N_11204);
nor U12937 (N_12937,N_8672,N_9907);
and U12938 (N_12938,N_9837,N_9831);
xor U12939 (N_12939,N_6273,N_11830);
xnor U12940 (N_12940,N_7555,N_9671);
nor U12941 (N_12941,N_8664,N_11719);
nand U12942 (N_12942,N_6467,N_8746);
nand U12943 (N_12943,N_7498,N_7507);
or U12944 (N_12944,N_10087,N_8165);
or U12945 (N_12945,N_7776,N_6607);
xnor U12946 (N_12946,N_7692,N_11178);
or U12947 (N_12947,N_11697,N_7918);
nand U12948 (N_12948,N_8417,N_10587);
xor U12949 (N_12949,N_10889,N_11586);
nand U12950 (N_12950,N_8213,N_9915);
or U12951 (N_12951,N_8494,N_10795);
xnor U12952 (N_12952,N_7460,N_8656);
xnor U12953 (N_12953,N_8290,N_7862);
xnor U12954 (N_12954,N_6776,N_9886);
or U12955 (N_12955,N_8071,N_7080);
nor U12956 (N_12956,N_10120,N_10606);
nand U12957 (N_12957,N_10749,N_7888);
or U12958 (N_12958,N_9795,N_10687);
nor U12959 (N_12959,N_7867,N_11468);
or U12960 (N_12960,N_6226,N_11671);
and U12961 (N_12961,N_11342,N_6801);
and U12962 (N_12962,N_11366,N_7181);
and U12963 (N_12963,N_7416,N_11900);
xnor U12964 (N_12964,N_8193,N_9134);
nor U12965 (N_12965,N_6505,N_9117);
or U12966 (N_12966,N_10710,N_8461);
and U12967 (N_12967,N_8188,N_7026);
nor U12968 (N_12968,N_6114,N_10633);
and U12969 (N_12969,N_9129,N_6365);
nor U12970 (N_12970,N_11239,N_8267);
xnor U12971 (N_12971,N_10007,N_10190);
nor U12972 (N_12972,N_11996,N_8833);
nand U12973 (N_12973,N_9306,N_11616);
and U12974 (N_12974,N_7095,N_11945);
xnor U12975 (N_12975,N_11808,N_8399);
nor U12976 (N_12976,N_10596,N_6083);
xnor U12977 (N_12977,N_8242,N_8759);
and U12978 (N_12978,N_7707,N_6522);
and U12979 (N_12979,N_10953,N_9916);
or U12980 (N_12980,N_10234,N_7600);
and U12981 (N_12981,N_7572,N_7274);
nor U12982 (N_12982,N_6949,N_6866);
and U12983 (N_12983,N_8204,N_9086);
xnor U12984 (N_12984,N_7702,N_9186);
and U12985 (N_12985,N_6403,N_9739);
nor U12986 (N_12986,N_7301,N_6669);
or U12987 (N_12987,N_10225,N_10371);
or U12988 (N_12988,N_7673,N_10014);
xnor U12989 (N_12989,N_10607,N_8954);
nand U12990 (N_12990,N_9858,N_7878);
nand U12991 (N_12991,N_11393,N_9933);
xor U12992 (N_12992,N_7686,N_11986);
and U12993 (N_12993,N_10713,N_9713);
nand U12994 (N_12994,N_10548,N_7023);
xnor U12995 (N_12995,N_9099,N_9478);
or U12996 (N_12996,N_10730,N_7231);
and U12997 (N_12997,N_8679,N_7842);
and U12998 (N_12998,N_10117,N_11013);
xnor U12999 (N_12999,N_9018,N_11565);
and U13000 (N_13000,N_11777,N_7437);
nand U13001 (N_13001,N_7503,N_8533);
and U13002 (N_13002,N_7422,N_8493);
xnor U13003 (N_13003,N_9549,N_9909);
nor U13004 (N_13004,N_9403,N_9448);
xor U13005 (N_13005,N_9200,N_9884);
or U13006 (N_13006,N_6934,N_7954);
and U13007 (N_13007,N_11066,N_11826);
nor U13008 (N_13008,N_10127,N_10292);
nand U13009 (N_13009,N_8086,N_6066);
nand U13010 (N_13010,N_6177,N_11506);
and U13011 (N_13011,N_6233,N_11234);
nand U13012 (N_13012,N_6996,N_9323);
xnor U13013 (N_13013,N_9073,N_6703);
nor U13014 (N_13014,N_9585,N_11999);
xnor U13015 (N_13015,N_6173,N_11534);
nor U13016 (N_13016,N_9409,N_7846);
and U13017 (N_13017,N_11240,N_7731);
xnor U13018 (N_13018,N_9954,N_11028);
nor U13019 (N_13019,N_8184,N_11122);
nand U13020 (N_13020,N_8149,N_6322);
or U13021 (N_13021,N_8389,N_6717);
nand U13022 (N_13022,N_8187,N_9093);
or U13023 (N_13023,N_8830,N_6323);
nand U13024 (N_13024,N_8176,N_7712);
nand U13025 (N_13025,N_10529,N_7804);
nand U13026 (N_13026,N_11754,N_10321);
nor U13027 (N_13027,N_6105,N_10735);
nor U13028 (N_13028,N_8117,N_10055);
nor U13029 (N_13029,N_11295,N_8146);
or U13030 (N_13030,N_10096,N_9682);
nand U13031 (N_13031,N_9095,N_6027);
and U13032 (N_13032,N_11927,N_8474);
xor U13033 (N_13033,N_8682,N_6107);
nor U13034 (N_13034,N_8729,N_6806);
and U13035 (N_13035,N_6038,N_9808);
and U13036 (N_13036,N_6461,N_9180);
xnor U13037 (N_13037,N_10204,N_6225);
and U13038 (N_13038,N_10149,N_9723);
xor U13039 (N_13039,N_7209,N_11644);
or U13040 (N_13040,N_6962,N_7266);
or U13041 (N_13041,N_10435,N_7410);
nor U13042 (N_13042,N_8576,N_7109);
nand U13043 (N_13043,N_9667,N_7540);
and U13044 (N_13044,N_11904,N_10731);
or U13045 (N_13045,N_6406,N_11422);
or U13046 (N_13046,N_8414,N_7455);
xnor U13047 (N_13047,N_11392,N_8073);
nor U13048 (N_13048,N_7085,N_8150);
and U13049 (N_13049,N_9581,N_6151);
and U13050 (N_13050,N_6863,N_9114);
or U13051 (N_13051,N_7779,N_8114);
xor U13052 (N_13052,N_11817,N_6620);
xnor U13053 (N_13053,N_11739,N_7548);
nor U13054 (N_13054,N_10022,N_11011);
nand U13055 (N_13055,N_7362,N_7933);
or U13056 (N_13056,N_10289,N_6807);
and U13057 (N_13057,N_9017,N_9663);
and U13058 (N_13058,N_7149,N_6500);
nor U13059 (N_13059,N_7265,N_11284);
nor U13060 (N_13060,N_9219,N_7807);
nand U13061 (N_13061,N_7609,N_11603);
and U13062 (N_13062,N_9604,N_9870);
or U13063 (N_13063,N_11528,N_7996);
nand U13064 (N_13064,N_6618,N_8559);
and U13065 (N_13065,N_8721,N_10144);
nor U13066 (N_13066,N_6827,N_10343);
and U13067 (N_13067,N_7007,N_10773);
nor U13068 (N_13068,N_11825,N_11151);
nand U13069 (N_13069,N_9383,N_11144);
xnor U13070 (N_13070,N_10074,N_11483);
and U13071 (N_13071,N_9611,N_6910);
or U13072 (N_13072,N_11113,N_11723);
or U13073 (N_13073,N_10285,N_11146);
nor U13074 (N_13074,N_6132,N_7985);
nand U13075 (N_13075,N_9868,N_7944);
or U13076 (N_13076,N_10377,N_8210);
nor U13077 (N_13077,N_11309,N_9834);
or U13078 (N_13078,N_8674,N_7783);
nand U13079 (N_13079,N_9138,N_9244);
nand U13080 (N_13080,N_10865,N_7680);
nor U13081 (N_13081,N_11562,N_10246);
and U13082 (N_13082,N_7541,N_9389);
and U13083 (N_13083,N_11890,N_7899);
nand U13084 (N_13084,N_8394,N_10741);
nand U13085 (N_13085,N_8372,N_7603);
nand U13086 (N_13086,N_9161,N_6783);
xnor U13087 (N_13087,N_6529,N_10290);
and U13088 (N_13088,N_9175,N_6644);
nand U13089 (N_13089,N_10909,N_8550);
nor U13090 (N_13090,N_11094,N_8050);
nor U13091 (N_13091,N_8111,N_7203);
and U13092 (N_13092,N_6861,N_8222);
nand U13093 (N_13093,N_6685,N_11195);
nand U13094 (N_13094,N_11097,N_7519);
xor U13095 (N_13095,N_10270,N_6630);
nor U13096 (N_13096,N_10604,N_8690);
xor U13097 (N_13097,N_6792,N_9359);
xnor U13098 (N_13098,N_10112,N_7538);
xnor U13099 (N_13099,N_6538,N_8467);
nor U13100 (N_13100,N_9317,N_11225);
nand U13101 (N_13101,N_10410,N_8910);
or U13102 (N_13102,N_10279,N_6998);
or U13103 (N_13103,N_6775,N_6101);
or U13104 (N_13104,N_8381,N_8999);
or U13105 (N_13105,N_6080,N_11593);
and U13106 (N_13106,N_6951,N_9693);
or U13107 (N_13107,N_8107,N_6162);
nor U13108 (N_13108,N_10492,N_11222);
nor U13109 (N_13109,N_8110,N_10557);
and U13110 (N_13110,N_8262,N_6471);
xor U13111 (N_13111,N_8370,N_9877);
and U13112 (N_13112,N_10347,N_10110);
and U13113 (N_13113,N_8819,N_11224);
and U13114 (N_13114,N_8628,N_10382);
nand U13115 (N_13115,N_11278,N_10142);
nor U13116 (N_13116,N_8463,N_8311);
or U13117 (N_13117,N_8535,N_10269);
or U13118 (N_13118,N_11165,N_11897);
nor U13119 (N_13119,N_6576,N_10904);
or U13120 (N_13120,N_7812,N_10101);
nor U13121 (N_13121,N_10975,N_9629);
nand U13122 (N_13122,N_7750,N_9483);
xor U13123 (N_13123,N_7721,N_10394);
or U13124 (N_13124,N_6627,N_9211);
nand U13125 (N_13125,N_11253,N_7411);
nor U13126 (N_13126,N_6297,N_8095);
nor U13127 (N_13127,N_7319,N_10589);
nor U13128 (N_13128,N_11903,N_11476);
nor U13129 (N_13129,N_6410,N_7312);
nor U13130 (N_13130,N_10508,N_10020);
nand U13131 (N_13131,N_10267,N_8443);
or U13132 (N_13132,N_10853,N_8490);
or U13133 (N_13133,N_8751,N_7103);
nor U13134 (N_13134,N_7920,N_11725);
nor U13135 (N_13135,N_10433,N_11314);
and U13136 (N_13136,N_10545,N_9591);
xor U13137 (N_13137,N_11744,N_11102);
and U13138 (N_13138,N_8497,N_9076);
nand U13139 (N_13139,N_6536,N_8538);
and U13140 (N_13140,N_9622,N_10328);
nand U13141 (N_13141,N_9371,N_9484);
nor U13142 (N_13142,N_11488,N_9330);
nor U13143 (N_13143,N_9500,N_7677);
nor U13144 (N_13144,N_9910,N_9596);
nand U13145 (N_13145,N_8162,N_10446);
nor U13146 (N_13146,N_10732,N_6976);
xnor U13147 (N_13147,N_10176,N_10518);
xnor U13148 (N_13148,N_6752,N_9307);
or U13149 (N_13149,N_9521,N_11466);
nor U13150 (N_13150,N_10702,N_11331);
and U13151 (N_13151,N_7516,N_9346);
or U13152 (N_13152,N_8617,N_11399);
or U13153 (N_13153,N_6856,N_10781);
and U13154 (N_13154,N_6726,N_9570);
and U13155 (N_13155,N_10995,N_11068);
or U13156 (N_13156,N_11776,N_11444);
or U13157 (N_13157,N_7699,N_8170);
or U13158 (N_13158,N_7508,N_6389);
or U13159 (N_13159,N_6498,N_9424);
or U13160 (N_13160,N_9833,N_11482);
nand U13161 (N_13161,N_9619,N_11340);
and U13162 (N_13162,N_6710,N_6686);
nand U13163 (N_13163,N_8344,N_11293);
nor U13164 (N_13164,N_10654,N_8275);
xor U13165 (N_13165,N_10875,N_10600);
xnor U13166 (N_13166,N_11153,N_9803);
nor U13167 (N_13167,N_11678,N_7229);
or U13168 (N_13168,N_8479,N_11560);
nor U13169 (N_13169,N_7371,N_7027);
nand U13170 (N_13170,N_9417,N_8166);
or U13171 (N_13171,N_6291,N_9075);
xor U13172 (N_13172,N_7740,N_11756);
or U13173 (N_13173,N_10345,N_8624);
or U13174 (N_13174,N_11150,N_7385);
and U13175 (N_13175,N_8839,N_11118);
and U13176 (N_13176,N_10429,N_9414);
or U13177 (N_13177,N_11061,N_6751);
nor U13178 (N_13178,N_10221,N_6584);
xor U13179 (N_13179,N_8382,N_10332);
nor U13180 (N_13180,N_8036,N_6769);
and U13181 (N_13181,N_10737,N_11804);
nor U13182 (N_13182,N_9845,N_7893);
or U13183 (N_13183,N_6720,N_8293);
nor U13184 (N_13184,N_7487,N_8761);
nand U13185 (N_13185,N_9574,N_8713);
nor U13186 (N_13186,N_8552,N_7098);
or U13187 (N_13187,N_8076,N_10263);
nand U13188 (N_13188,N_10591,N_10835);
nand U13189 (N_13189,N_8313,N_11350);
nand U13190 (N_13190,N_10890,N_6517);
nor U13191 (N_13191,N_11714,N_10943);
xnor U13192 (N_13192,N_8282,N_10069);
or U13193 (N_13193,N_11498,N_10637);
nand U13194 (N_13194,N_11158,N_9372);
xnor U13195 (N_13195,N_6141,N_6088);
xnor U13196 (N_13196,N_10358,N_9665);
or U13197 (N_13197,N_10699,N_11086);
nand U13198 (N_13198,N_8179,N_8818);
and U13199 (N_13199,N_7847,N_10082);
xnor U13200 (N_13200,N_11871,N_11056);
xnor U13201 (N_13201,N_8886,N_10673);
xor U13202 (N_13202,N_11322,N_11185);
nor U13203 (N_13203,N_8669,N_7631);
nand U13204 (N_13204,N_11936,N_8051);
xnor U13205 (N_13205,N_6502,N_8670);
or U13206 (N_13206,N_8116,N_6009);
nor U13207 (N_13207,N_10248,N_7734);
nor U13208 (N_13208,N_11121,N_11733);
and U13209 (N_13209,N_6579,N_11287);
nand U13210 (N_13210,N_8567,N_8003);
nor U13211 (N_13211,N_9641,N_8557);
and U13212 (N_13212,N_6875,N_11669);
nor U13213 (N_13213,N_11014,N_8255);
xnor U13214 (N_13214,N_11436,N_9370);
nand U13215 (N_13215,N_9096,N_8101);
nand U13216 (N_13216,N_7456,N_7844);
and U13217 (N_13217,N_10635,N_10882);
nand U13218 (N_13218,N_10818,N_10536);
nor U13219 (N_13219,N_8564,N_7164);
xor U13220 (N_13220,N_7877,N_7175);
xnor U13221 (N_13221,N_7392,N_6259);
or U13222 (N_13222,N_10040,N_7232);
xor U13223 (N_13223,N_9865,N_10115);
nor U13224 (N_13224,N_8872,N_6588);
xor U13225 (N_13225,N_10757,N_7500);
or U13226 (N_13226,N_7641,N_7444);
or U13227 (N_13227,N_6890,N_11250);
or U13228 (N_13228,N_6969,N_6945);
and U13229 (N_13229,N_8568,N_6332);
nand U13230 (N_13230,N_6409,N_11289);
and U13231 (N_13231,N_7939,N_11497);
or U13232 (N_13232,N_9060,N_8952);
and U13233 (N_13233,N_6386,N_7442);
xor U13234 (N_13234,N_6202,N_9976);
and U13235 (N_13235,N_10621,N_9623);
nand U13236 (N_13236,N_11292,N_10969);
nand U13237 (N_13237,N_11412,N_6901);
xnor U13238 (N_13238,N_9844,N_7170);
nor U13239 (N_13239,N_7526,N_7407);
nor U13240 (N_13240,N_7934,N_6040);
nor U13241 (N_13241,N_10787,N_6816);
or U13242 (N_13242,N_11842,N_9702);
and U13243 (N_13243,N_6540,N_10685);
and U13244 (N_13244,N_11493,N_9367);
nor U13245 (N_13245,N_7481,N_10426);
and U13246 (N_13246,N_6656,N_6970);
or U13247 (N_13247,N_10819,N_7014);
nor U13248 (N_13248,N_7016,N_7671);
or U13249 (N_13249,N_6098,N_11815);
xnor U13250 (N_13250,N_10491,N_10644);
xnor U13251 (N_13251,N_7421,N_11976);
and U13252 (N_13252,N_9412,N_9474);
and U13253 (N_13253,N_10791,N_6394);
or U13254 (N_13254,N_11973,N_9444);
or U13255 (N_13255,N_10174,N_9919);
or U13256 (N_13256,N_7071,N_7130);
nand U13257 (N_13257,N_8884,N_10760);
or U13258 (N_13258,N_11262,N_9664);
nand U13259 (N_13259,N_11296,N_6772);
xnor U13260 (N_13260,N_6077,N_6554);
and U13261 (N_13261,N_7323,N_8873);
nand U13262 (N_13262,N_6298,N_6469);
nor U13263 (N_13263,N_11448,N_10566);
and U13264 (N_13264,N_11180,N_7801);
and U13265 (N_13265,N_6713,N_6182);
nor U13266 (N_13266,N_6602,N_10778);
nor U13267 (N_13267,N_8484,N_7695);
xor U13268 (N_13268,N_11892,N_7587);
xnor U13269 (N_13269,N_10748,N_6045);
xnor U13270 (N_13270,N_6828,N_6765);
nor U13271 (N_13271,N_10979,N_11455);
and U13272 (N_13272,N_7784,N_7259);
and U13273 (N_13273,N_10681,N_7764);
nand U13274 (N_13274,N_6160,N_8169);
nand U13275 (N_13275,N_8802,N_7833);
nor U13276 (N_13276,N_10199,N_7223);
nand U13277 (N_13277,N_10661,N_7257);
nor U13278 (N_13278,N_10716,N_6835);
nand U13279 (N_13279,N_9426,N_8874);
xnor U13280 (N_13280,N_6253,N_8456);
or U13281 (N_13281,N_6965,N_7975);
nand U13282 (N_13282,N_11520,N_11035);
xnor U13283 (N_13283,N_11730,N_8480);
nor U13284 (N_13284,N_7643,N_10743);
nor U13285 (N_13285,N_8335,N_8340);
and U13286 (N_13286,N_11732,N_6348);
xor U13287 (N_13287,N_6850,N_6217);
nor U13288 (N_13288,N_8124,N_7430);
xor U13289 (N_13289,N_8972,N_8097);
nand U13290 (N_13290,N_11162,N_11105);
xor U13291 (N_13291,N_9167,N_11137);
nand U13292 (N_13292,N_9792,N_8631);
nor U13293 (N_13293,N_11111,N_8047);
xor U13294 (N_13294,N_9824,N_9708);
nor U13295 (N_13295,N_10124,N_9263);
nor U13296 (N_13296,N_11977,N_9871);
xor U13297 (N_13297,N_6687,N_11675);
nor U13298 (N_13298,N_6359,N_11360);
and U13299 (N_13299,N_6511,N_10076);
nor U13300 (N_13300,N_11507,N_6864);
nand U13301 (N_13301,N_8283,N_9351);
nor U13302 (N_13302,N_7640,N_6810);
nand U13303 (N_13303,N_11768,N_10576);
nand U13304 (N_13304,N_11821,N_9590);
nand U13305 (N_13305,N_9022,N_8330);
nor U13306 (N_13306,N_6745,N_10980);
xnor U13307 (N_13307,N_8687,N_11156);
xor U13308 (N_13308,N_6559,N_11538);
and U13309 (N_13309,N_7882,N_7883);
nand U13310 (N_13310,N_10114,N_11288);
xor U13311 (N_13311,N_6023,N_6553);
nand U13312 (N_13312,N_6250,N_7094);
or U13313 (N_13313,N_11588,N_10669);
and U13314 (N_13314,N_11984,N_6514);
and U13315 (N_13315,N_10202,N_9408);
and U13316 (N_13316,N_9486,N_11853);
and U13317 (N_13317,N_9575,N_6113);
or U13318 (N_13318,N_10445,N_7121);
nand U13319 (N_13319,N_7744,N_7278);
nor U13320 (N_13320,N_8541,N_8459);
xnor U13321 (N_13321,N_11371,N_11972);
nor U13322 (N_13322,N_6372,N_7687);
nand U13323 (N_13323,N_9893,N_10912);
nand U13324 (N_13324,N_11684,N_11254);
nand U13325 (N_13325,N_10900,N_6123);
nand U13326 (N_13326,N_9714,N_9875);
and U13327 (N_13327,N_7059,N_10978);
nand U13328 (N_13328,N_8156,N_8891);
xor U13329 (N_13329,N_11956,N_7173);
or U13330 (N_13330,N_9518,N_11882);
and U13331 (N_13331,N_6153,N_9750);
and U13332 (N_13332,N_6381,N_11193);
xor U13333 (N_13333,N_8701,N_7357);
or U13334 (N_13334,N_6632,N_10029);
and U13335 (N_13335,N_8926,N_6271);
or U13336 (N_13336,N_11282,N_9535);
and U13337 (N_13337,N_10898,N_6594);
and U13338 (N_13338,N_7043,N_9132);
and U13339 (N_13339,N_10729,N_7771);
nand U13340 (N_13340,N_11080,N_10310);
xnor U13341 (N_13341,N_8464,N_6841);
and U13342 (N_13342,N_11957,N_11654);
xor U13343 (N_13343,N_7224,N_11581);
or U13344 (N_13344,N_9677,N_8272);
or U13345 (N_13345,N_7904,N_10280);
or U13346 (N_13346,N_9494,N_7064);
nand U13347 (N_13347,N_6732,N_6247);
nand U13348 (N_13348,N_6756,N_6146);
and U13349 (N_13349,N_11174,N_11942);
and U13350 (N_13350,N_6481,N_11387);
xnor U13351 (N_13351,N_7967,N_7183);
or U13352 (N_13352,N_10396,N_9192);
and U13353 (N_13353,N_8237,N_6812);
nor U13354 (N_13354,N_6862,N_7908);
nor U13355 (N_13355,N_9697,N_6054);
or U13356 (N_13356,N_8245,N_9218);
xor U13357 (N_13357,N_7063,N_10886);
or U13358 (N_13358,N_11641,N_6532);
or U13359 (N_13359,N_11530,N_9657);
and U13360 (N_13360,N_8600,N_10892);
or U13361 (N_13361,N_10551,N_6206);
nand U13362 (N_13362,N_7535,N_8601);
xor U13363 (N_13363,N_8446,N_8447);
or U13364 (N_13364,N_9109,N_9077);
or U13365 (N_13365,N_6640,N_9670);
and U13366 (N_13366,N_6744,N_8719);
xnor U13367 (N_13367,N_6913,N_7303);
nor U13368 (N_13368,N_6488,N_11939);
and U13369 (N_13369,N_6401,N_7317);
or U13370 (N_13370,N_11326,N_7314);
xnor U13371 (N_13371,N_9631,N_11092);
nor U13372 (N_13372,N_10682,N_9674);
or U13373 (N_13373,N_10471,N_9653);
or U13374 (N_13374,N_9310,N_9869);
nand U13375 (N_13375,N_9647,N_6578);
nor U13376 (N_13376,N_8334,N_6755);
nor U13377 (N_13377,N_8526,N_8466);
or U13378 (N_13378,N_8217,N_7565);
nor U13379 (N_13379,N_8359,N_6337);
nand U13380 (N_13380,N_11464,N_9977);
nor U13381 (N_13381,N_9859,N_9544);
and U13382 (N_13382,N_10612,N_8823);
xnor U13383 (N_13383,N_10848,N_10708);
nor U13384 (N_13384,N_8595,N_6563);
or U13385 (N_13385,N_8709,N_9675);
xor U13386 (N_13386,N_8105,N_6709);
or U13387 (N_13387,N_11577,N_9579);
and U13388 (N_13388,N_8692,N_9340);
nand U13389 (N_13389,N_8940,N_11210);
xor U13390 (N_13390,N_7150,N_9780);
or U13391 (N_13391,N_11649,N_6368);
xor U13392 (N_13392,N_7024,N_6287);
or U13393 (N_13393,N_7451,N_10728);
xor U13394 (N_13394,N_7268,N_10653);
xor U13395 (N_13395,N_7205,N_6229);
or U13396 (N_13396,N_10549,N_6109);
nand U13397 (N_13397,N_10366,N_11474);
nor U13398 (N_13398,N_11920,N_11188);
and U13399 (N_13399,N_7958,N_11319);
nor U13400 (N_13400,N_9225,N_11463);
and U13401 (N_13401,N_7438,N_9490);
nand U13402 (N_13402,N_11244,N_10308);
nand U13403 (N_13403,N_6811,N_6921);
nand U13404 (N_13404,N_9299,N_9602);
and U13405 (N_13405,N_11361,N_6294);
nand U13406 (N_13406,N_6895,N_7436);
or U13407 (N_13407,N_11545,N_10871);
nor U13408 (N_13408,N_8264,N_11612);
nand U13409 (N_13409,N_6234,N_9950);
nor U13410 (N_13410,N_8180,N_8753);
and U13411 (N_13411,N_7448,N_6636);
or U13412 (N_13412,N_7828,N_6530);
and U13413 (N_13413,N_8216,N_8562);
or U13414 (N_13414,N_6585,N_7693);
and U13415 (N_13415,N_10064,N_9930);
and U13416 (N_13416,N_11344,N_11630);
xnor U13417 (N_13417,N_6415,N_11452);
and U13418 (N_13418,N_11356,N_11073);
and U13419 (N_13419,N_11932,N_10915);
nor U13420 (N_13420,N_6557,N_9460);
nor U13421 (N_13421,N_6821,N_8379);
nor U13422 (N_13422,N_9115,N_6169);
or U13423 (N_13423,N_11192,N_11549);
or U13424 (N_13424,N_8092,N_11041);
nand U13425 (N_13425,N_9338,N_10185);
nand U13426 (N_13426,N_8434,N_10804);
and U13427 (N_13427,N_6737,N_8413);
nand U13428 (N_13428,N_10454,N_6227);
xnor U13429 (N_13429,N_11614,N_10501);
nor U13430 (N_13430,N_11551,N_8841);
nand U13431 (N_13431,N_9735,N_10151);
or U13432 (N_13432,N_6452,N_7554);
nand U13433 (N_13433,N_7529,N_6734);
xor U13434 (N_13434,N_9423,N_6356);
nand U13435 (N_13435,N_8804,N_9255);
and U13436 (N_13436,N_9420,N_11182);
nand U13437 (N_13437,N_8139,N_7078);
and U13438 (N_13438,N_6116,N_11912);
and U13439 (N_13439,N_7668,N_10286);
or U13440 (N_13440,N_7036,N_8764);
and U13441 (N_13441,N_9636,N_7249);
xnor U13442 (N_13442,N_6917,N_7363);
xnor U13443 (N_13443,N_7761,N_7590);
nor U13444 (N_13444,N_8623,N_11335);
xnor U13445 (N_13445,N_6971,N_10759);
or U13446 (N_13446,N_11624,N_10525);
and U13447 (N_13447,N_11196,N_7139);
and U13448 (N_13448,N_6197,N_10562);
xor U13449 (N_13449,N_10535,N_11898);
nand U13450 (N_13450,N_7042,N_6754);
nor U13451 (N_13451,N_10006,N_8515);
xor U13452 (N_13452,N_11794,N_11706);
xnor U13453 (N_13453,N_6451,N_10860);
and U13454 (N_13454,N_6393,N_7432);
or U13455 (N_13455,N_6535,N_11117);
xor U13456 (N_13456,N_9439,N_9955);
or U13457 (N_13457,N_8586,N_10342);
nand U13458 (N_13458,N_9852,N_11268);
nor U13459 (N_13459,N_7493,N_8465);
or U13460 (N_13460,N_10375,N_6736);
xnor U13461 (N_13461,N_11812,N_6187);
or U13462 (N_13462,N_7051,N_8570);
nand U13463 (N_13463,N_11352,N_7619);
or U13464 (N_13464,N_7497,N_10756);
nor U13465 (N_13465,N_8208,N_6648);
xnor U13466 (N_13466,N_6309,N_7045);
nand U13467 (N_13467,N_9536,N_11100);
or U13468 (N_13468,N_11602,N_6704);
and U13469 (N_13469,N_8758,N_9251);
nor U13470 (N_13470,N_11257,N_11467);
nor U13471 (N_13471,N_11417,N_7982);
or U13472 (N_13472,N_7630,N_7484);
nor U13473 (N_13473,N_11674,N_7936);
nand U13474 (N_13474,N_8835,N_7093);
and U13475 (N_13475,N_9365,N_6550);
or U13476 (N_13476,N_8075,N_10231);
nor U13477 (N_13477,N_9145,N_9701);
nand U13478 (N_13478,N_7250,N_10462);
or U13479 (N_13479,N_9587,N_6414);
nor U13480 (N_13480,N_7964,N_7366);
and U13481 (N_13481,N_10745,N_11533);
and U13482 (N_13482,N_10961,N_7401);
nand U13483 (N_13483,N_11642,N_10688);
or U13484 (N_13484,N_9315,N_9363);
or U13485 (N_13485,N_8357,N_8008);
and U13486 (N_13486,N_9514,N_11795);
nand U13487 (N_13487,N_9195,N_10331);
and U13488 (N_13488,N_7857,N_7179);
and U13489 (N_13489,N_6771,N_7909);
and U13490 (N_13490,N_11916,N_6936);
nand U13491 (N_13491,N_9648,N_11526);
nand U13492 (N_13492,N_9228,N_10863);
and U13493 (N_13493,N_10106,N_6072);
nand U13494 (N_13494,N_10744,N_7894);
nor U13495 (N_13495,N_7340,N_7355);
and U13496 (N_13496,N_10498,N_11363);
and U13497 (N_13497,N_10881,N_11208);
nor U13498 (N_13498,N_8171,N_9235);
xor U13499 (N_13499,N_10251,N_11307);
xnor U13500 (N_13500,N_10229,N_9201);
and U13501 (N_13501,N_7871,N_9630);
nand U13502 (N_13502,N_6382,N_10281);
and U13503 (N_13503,N_11940,N_6057);
or U13504 (N_13504,N_10590,N_11578);
xnor U13505 (N_13505,N_9112,N_9603);
xor U13506 (N_13506,N_11343,N_11950);
xnor U13507 (N_13507,N_10044,N_7678);
nand U13508 (N_13508,N_7653,N_9533);
and U13509 (N_13509,N_8175,N_8052);
nor U13510 (N_13510,N_7397,N_9606);
or U13511 (N_13511,N_6527,N_8824);
or U13512 (N_13512,N_11108,N_7913);
or U13513 (N_13513,N_6279,N_9088);
or U13514 (N_13514,N_6455,N_9406);
nand U13515 (N_13515,N_10964,N_6303);
and U13516 (N_13516,N_6564,N_6035);
nand U13517 (N_13517,N_10942,N_7032);
nand U13518 (N_13518,N_6591,N_7963);
nand U13519 (N_13519,N_11761,N_9473);
nor U13520 (N_13520,N_9556,N_9703);
and U13521 (N_13521,N_11354,N_10126);
xor U13522 (N_13522,N_11670,N_8384);
and U13523 (N_13523,N_8644,N_9404);
xor U13524 (N_13524,N_10136,N_10667);
and U13525 (N_13525,N_8027,N_6425);
and U13526 (N_13526,N_10268,N_8231);
nand U13527 (N_13527,N_9569,N_8735);
nor U13528 (N_13528,N_9256,N_8684);
nor U13529 (N_13529,N_9153,N_10856);
and U13530 (N_13530,N_8565,N_11866);
nor U13531 (N_13531,N_8973,N_8797);
xor U13532 (N_13532,N_11608,N_7140);
xnor U13533 (N_13533,N_8385,N_9656);
nand U13534 (N_13534,N_6654,N_7288);
and U13535 (N_13535,N_9860,N_9376);
nand U13536 (N_13536,N_9530,N_11007);
or U13537 (N_13537,N_8108,N_6246);
nor U13538 (N_13538,N_7562,N_11851);
nand U13539 (N_13539,N_8630,N_6373);
xor U13540 (N_13540,N_9333,N_9154);
nand U13541 (N_13541,N_11748,N_10362);
nor U13542 (N_13542,N_10036,N_10379);
or U13543 (N_13543,N_9511,N_7381);
or U13544 (N_13544,N_7322,N_11231);
nand U13545 (N_13545,N_10237,N_10668);
nand U13546 (N_13546,N_10206,N_6100);
nand U13547 (N_13547,N_9345,N_7767);
nand U13548 (N_13548,N_6853,N_6888);
nand U13549 (N_13549,N_7915,N_7820);
xnor U13550 (N_13550,N_9006,N_7195);
xor U13551 (N_13551,N_7258,N_11645);
or U13552 (N_13552,N_11755,N_6432);
nor U13553 (N_13553,N_11862,N_10456);
and U13554 (N_13554,N_10257,N_6993);
nand U13555 (N_13555,N_9779,N_11439);
xor U13556 (N_13556,N_7984,N_9823);
nand U13557 (N_13557,N_7937,N_8959);
and U13558 (N_13558,N_8119,N_6688);
nand U13559 (N_13559,N_7176,N_10291);
xnor U13560 (N_13560,N_8691,N_7365);
and U13561 (N_13561,N_11230,N_10419);
nor U13562 (N_13562,N_6762,N_10816);
or U13563 (N_13563,N_7114,N_7892);
nand U13564 (N_13564,N_6133,N_8938);
xnor U13565 (N_13565,N_9563,N_7280);
or U13566 (N_13566,N_7589,N_8887);
nor U13567 (N_13567,N_9507,N_7361);
nor U13568 (N_13568,N_11954,N_8160);
nand U13569 (N_13569,N_10299,N_8782);
nand U13570 (N_13570,N_11542,N_6320);
or U13571 (N_13571,N_10642,N_8185);
and U13572 (N_13572,N_11861,N_10986);
nor U13573 (N_13573,N_8866,N_7486);
nand U13574 (N_13574,N_8391,N_11881);
or U13575 (N_13575,N_7879,N_8033);
xnor U13576 (N_13576,N_10378,N_11604);
xor U13577 (N_13577,N_11160,N_7701);
and U13578 (N_13578,N_10784,N_6623);
and U13579 (N_13579,N_11511,N_6142);
xor U13580 (N_13580,N_10153,N_7813);
or U13581 (N_13581,N_8591,N_11995);
and U13582 (N_13582,N_9534,N_10671);
or U13583 (N_13583,N_6171,N_7521);
xor U13584 (N_13584,N_9122,N_9989);
or U13585 (N_13585,N_7610,N_11667);
and U13586 (N_13586,N_7192,N_7494);
or U13587 (N_13587,N_8519,N_7925);
nand U13588 (N_13588,N_6214,N_10831);
nand U13589 (N_13589,N_10261,N_7162);
or U13590 (N_13590,N_9232,N_6571);
or U13591 (N_13591,N_8678,N_9694);
or U13592 (N_13592,N_7825,N_6110);
nor U13593 (N_13593,N_8641,N_6604);
nor U13594 (N_13594,N_7938,N_11636);
nand U13595 (N_13595,N_9259,N_8556);
xnor U13596 (N_13596,N_10625,N_9595);
nor U13597 (N_13597,N_11377,N_10976);
xor U13598 (N_13598,N_11345,N_9286);
and U13599 (N_13599,N_10581,N_6043);
and U13600 (N_13600,N_8780,N_10583);
xor U13601 (N_13601,N_7551,N_6931);
nor U13602 (N_13602,N_11891,N_7528);
or U13603 (N_13603,N_7593,N_6697);
nor U13604 (N_13604,N_10941,N_11096);
xnor U13605 (N_13605,N_11286,N_10526);
xor U13606 (N_13606,N_7057,N_7106);
nand U13607 (N_13607,N_8587,N_7310);
nor U13608 (N_13608,N_11879,N_10077);
or U13609 (N_13609,N_7586,N_9546);
nor U13610 (N_13610,N_11721,N_10523);
or U13611 (N_13611,N_6548,N_11402);
nand U13612 (N_13612,N_7370,N_7019);
or U13613 (N_13613,N_7180,N_6633);
and U13614 (N_13614,N_10931,N_9616);
and U13615 (N_13615,N_10806,N_10230);
and U13616 (N_13616,N_9768,N_6833);
nor U13617 (N_13617,N_8378,N_10054);
xor U13618 (N_13618,N_9961,N_11514);
nor U13619 (N_13619,N_6508,N_10803);
or U13620 (N_13620,N_8360,N_10586);
or U13621 (N_13621,N_7342,N_9224);
nor U13622 (N_13622,N_11139,N_9883);
and U13623 (N_13623,N_6908,N_8977);
and U13624 (N_13624,N_8128,N_8731);
nand U13625 (N_13625,N_8605,N_8956);
or U13626 (N_13626,N_8147,N_10294);
nor U13627 (N_13627,N_9004,N_11375);
nand U13628 (N_13628,N_11913,N_6496);
nand U13629 (N_13629,N_9917,N_10579);
or U13630 (N_13630,N_8448,N_10736);
and U13631 (N_13631,N_8986,N_9097);
or U13632 (N_13632,N_7998,N_6501);
and U13633 (N_13633,N_7752,N_8031);
xor U13634 (N_13634,N_6037,N_10820);
or U13635 (N_13635,N_9185,N_11943);
nor U13636 (N_13636,N_6967,N_6597);
xnor U13637 (N_13637,N_9026,N_11159);
nand U13638 (N_13638,N_9988,N_9539);
nand U13639 (N_13639,N_7634,N_9140);
nor U13640 (N_13640,N_10503,N_7352);
or U13641 (N_13641,N_9796,N_10026);
or U13642 (N_13642,N_6277,N_11509);
or U13643 (N_13643,N_10467,N_10297);
or U13644 (N_13644,N_9396,N_10452);
and U13645 (N_13645,N_8232,N_10141);
or U13646 (N_13646,N_7188,N_9721);
nand U13647 (N_13647,N_7617,N_10947);
or U13648 (N_13648,N_9411,N_11458);
or U13649 (N_13649,N_7730,N_9222);
or U13650 (N_13650,N_6463,N_10830);
nor U13651 (N_13651,N_7973,N_9862);
nand U13652 (N_13652,N_10324,N_10130);
and U13653 (N_13653,N_8099,N_9825);
or U13654 (N_13654,N_9254,N_9661);
nand U13655 (N_13655,N_11615,N_8877);
nand U13656 (N_13656,N_7423,N_8697);
nor U13657 (N_13657,N_9156,N_11623);
nor U13658 (N_13658,N_8717,N_6964);
nand U13659 (N_13659,N_8500,N_7418);
nor U13660 (N_13660,N_7000,N_7349);
nor U13661 (N_13661,N_10372,N_8813);
nand U13662 (N_13662,N_6870,N_8710);
xnor U13663 (N_13663,N_7415,N_7368);
nand U13664 (N_13664,N_10674,N_8975);
xor U13665 (N_13665,N_8126,N_8927);
or U13666 (N_13666,N_7942,N_9378);
and U13667 (N_13667,N_8469,N_9032);
and U13668 (N_13668,N_8297,N_10461);
nand U13669 (N_13669,N_11447,N_7141);
nor U13670 (N_13670,N_7664,N_7959);
and U13671 (N_13671,N_6622,N_10072);
and U13672 (N_13672,N_11855,N_11779);
and U13673 (N_13673,N_6570,N_8625);
or U13674 (N_13674,N_8386,N_7506);
nand U13675 (N_13675,N_6963,N_7543);
nand U13676 (N_13676,N_6665,N_10013);
nor U13677 (N_13677,N_7606,N_9282);
nor U13678 (N_13678,N_7293,N_7644);
nor U13679 (N_13679,N_11790,N_6008);
nand U13680 (N_13680,N_11510,N_10303);
nand U13681 (N_13681,N_7737,N_8829);
xnor U13682 (N_13682,N_10926,N_8404);
or U13683 (N_13683,N_9036,N_9270);
nand U13684 (N_13684,N_11886,N_10999);
nor U13685 (N_13685,N_6699,N_8917);
nor U13686 (N_13686,N_6741,N_9769);
or U13687 (N_13687,N_7796,N_6638);
and U13688 (N_13688,N_6157,N_10032);
nor U13689 (N_13689,N_7795,N_10024);
or U13690 (N_13690,N_10095,N_6673);
and U13691 (N_13691,N_10271,N_11793);
and U13692 (N_13692,N_8348,N_7727);
or U13693 (N_13693,N_6430,N_11832);
nor U13694 (N_13694,N_7831,N_6025);
xor U13695 (N_13695,N_8530,N_8549);
nand U13696 (N_13696,N_10401,N_8522);
nor U13697 (N_13697,N_8203,N_8662);
and U13698 (N_13698,N_7408,N_6539);
xor U13699 (N_13699,N_10056,N_11734);
nor U13700 (N_13700,N_8257,N_7638);
and U13701 (N_13701,N_6439,N_11127);
xnor U13702 (N_13702,N_11659,N_7010);
nor U13703 (N_13703,N_9308,N_9482);
xor U13704 (N_13704,N_6211,N_9853);
or U13705 (N_13705,N_11485,N_7004);
or U13706 (N_13706,N_8616,N_6128);
nor U13707 (N_13707,N_8990,N_11741);
nand U13708 (N_13708,N_9436,N_10564);
nand U13709 (N_13709,N_6912,N_6766);
nor U13710 (N_13710,N_6193,N_10724);
xor U13711 (N_13711,N_8336,N_7981);
nand U13712 (N_13712,N_8795,N_8440);
nor U13713 (N_13713,N_6830,N_9620);
nand U13714 (N_13714,N_7916,N_11953);
and U13715 (N_13715,N_8308,N_8115);
xor U13716 (N_13716,N_9038,N_6032);
nor U13717 (N_13717,N_10019,N_7866);
and U13718 (N_13718,N_9583,N_9011);
xor U13719 (N_13719,N_7079,N_10071);
or U13720 (N_13720,N_8409,N_8774);
or U13721 (N_13721,N_10178,N_8653);
xnor U13722 (N_13722,N_9986,N_11020);
xnor U13723 (N_13723,N_10534,N_8627);
and U13724 (N_13724,N_10507,N_8205);
nor U13725 (N_13725,N_9720,N_8315);
nand U13726 (N_13726,N_11163,N_9401);
xnor U13727 (N_13727,N_6891,N_6992);
and U13728 (N_13728,N_8935,N_11529);
nor U13729 (N_13729,N_8294,N_9443);
and U13730 (N_13730,N_9903,N_10301);
nor U13731 (N_13731,N_11594,N_6370);
xnor U13732 (N_13732,N_8658,N_10066);
or U13733 (N_13733,N_7107,N_10764);
and U13734 (N_13734,N_9835,N_11775);
xor U13735 (N_13735,N_11396,N_11347);
nor U13736 (N_13736,N_10872,N_10415);
nor U13737 (N_13737,N_10852,N_6104);
nand U13738 (N_13738,N_8638,N_11863);
xor U13739 (N_13739,N_9495,N_10873);
and U13740 (N_13740,N_7331,N_6677);
xnor U13741 (N_13741,N_10385,N_11501);
or U13742 (N_13742,N_7276,N_6489);
or U13743 (N_13743,N_11040,N_10990);
xor U13744 (N_13744,N_10648,N_9350);
nand U13745 (N_13745,N_6764,N_10168);
nand U13746 (N_13746,N_9765,N_7193);
nand U13747 (N_13747,N_9266,N_10000);
or U13748 (N_13748,N_7189,N_9947);
nand U13749 (N_13749,N_7803,N_7542);
and U13750 (N_13750,N_6091,N_6078);
nor U13751 (N_13751,N_10876,N_11575);
or U13752 (N_13752,N_10264,N_10189);
xnor U13753 (N_13753,N_10479,N_9311);
or U13754 (N_13754,N_10813,N_7906);
nand U13755 (N_13755,N_9593,N_10384);
or U13756 (N_13756,N_8892,N_7873);
nand U13757 (N_13757,N_8668,N_6150);
nand U13758 (N_13758,N_11320,N_6946);
or U13759 (N_13759,N_8766,N_11926);
nor U13760 (N_13760,N_7153,N_9600);
and U13761 (N_13761,N_9146,N_11708);
nor U13762 (N_13762,N_11907,N_11763);
nand U13763 (N_13763,N_11084,N_8918);
xnor U13764 (N_13764,N_10432,N_8809);
xor U13765 (N_13765,N_10603,N_11653);
nand U13766 (N_13766,N_11202,N_9447);
or U13767 (N_13767,N_10513,N_6092);
nor U13768 (N_13768,N_7821,N_8528);
nand U13769 (N_13769,N_10618,N_11064);
nor U13770 (N_13770,N_8241,N_10239);
nor U13771 (N_13771,N_6164,N_11430);
and U13772 (N_13772,N_9655,N_9527);
or U13773 (N_13773,N_10539,N_10894);
xor U13774 (N_13774,N_8598,N_8042);
xnor U13775 (N_13775,N_11770,N_10109);
and U13776 (N_13776,N_7703,N_6290);
and U13777 (N_13777,N_6210,N_9607);
xnor U13778 (N_13778,N_9249,N_6817);
and U13779 (N_13779,N_8152,N_8531);
nand U13780 (N_13780,N_6446,N_10284);
nor U13781 (N_13781,N_9273,N_6129);
nand U13782 (N_13782,N_7700,N_7684);
and U13783 (N_13783,N_9690,N_11699);
and U13784 (N_13784,N_8355,N_11398);
nor U13785 (N_13785,N_7509,N_6296);
and U13786 (N_13786,N_9797,N_6749);
nor U13787 (N_13787,N_9684,N_10173);
nand U13788 (N_13788,N_8153,N_7782);
and U13789 (N_13789,N_8796,N_6725);
xor U13790 (N_13790,N_8163,N_6843);
xnor U13791 (N_13791,N_7275,N_7264);
and U13792 (N_13792,N_11199,N_6650);
xor U13793 (N_13793,N_9431,N_9505);
and U13794 (N_13794,N_7932,N_10165);
and U13795 (N_13795,N_9214,N_7720);
or U13796 (N_13796,N_9220,N_10573);
nand U13797 (N_13797,N_7546,N_6094);
or U13798 (N_13798,N_7279,N_10364);
and U13799 (N_13799,N_8226,N_11865);
nand U13800 (N_13800,N_9936,N_7075);
nand U13801 (N_13801,N_6387,N_8611);
nor U13802 (N_13802,N_10081,N_8951);
or U13803 (N_13803,N_10186,N_6943);
nor U13804 (N_13804,N_11695,N_8671);
xnor U13805 (N_13805,N_8661,N_6228);
and U13806 (N_13806,N_10923,N_8514);
xnor U13807 (N_13807,N_7351,N_11556);
or U13808 (N_13808,N_11081,N_9905);
xor U13809 (N_13809,N_9368,N_8121);
nand U13810 (N_13810,N_8642,N_9598);
nand U13811 (N_13811,N_10254,N_6378);
nor U13812 (N_13812,N_11568,N_11471);
nand U13813 (N_13813,N_8498,N_9752);
xnor U13814 (N_13814,N_8420,N_7431);
nor U13815 (N_13815,N_9934,N_10599);
nand U13816 (N_13816,N_9586,N_7273);
nand U13817 (N_13817,N_9502,N_10801);
or U13818 (N_13818,N_8799,N_9832);
nor U13819 (N_13819,N_7665,N_11992);
nand U13820 (N_13820,N_7052,N_8286);
nor U13821 (N_13821,N_11856,N_9719);
nor U13822 (N_13822,N_11012,N_6256);
or U13823 (N_13823,N_6899,N_7081);
xor U13824 (N_13824,N_9105,N_6474);
or U13825 (N_13825,N_9386,N_6624);
and U13826 (N_13826,N_8317,N_9580);
and U13827 (N_13827,N_6803,N_9895);
and U13828 (N_13828,N_6070,N_6860);
or U13829 (N_13829,N_6715,N_9506);
xnor U13830 (N_13830,N_10179,N_10038);
and U13831 (N_13831,N_6520,N_10810);
or U13832 (N_13832,N_7247,N_10823);
and U13833 (N_13833,N_6318,N_7168);
nand U13834 (N_13834,N_6165,N_11044);
xor U13835 (N_13835,N_7382,N_6659);
nand U13836 (N_13836,N_6612,N_6402);
or U13837 (N_13837,N_10754,N_8001);
nor U13838 (N_13838,N_9973,N_6136);
nor U13839 (N_13839,N_9496,N_7028);
or U13840 (N_13840,N_11038,N_11570);
nor U13841 (N_13841,N_8786,N_8405);
or U13842 (N_13842,N_11840,N_11524);
nand U13843 (N_13843,N_10824,N_7768);
nor U13844 (N_13844,N_7228,N_7394);
xor U13845 (N_13845,N_10738,N_9545);
xor U13846 (N_13846,N_7239,N_7772);
and U13847 (N_13847,N_7646,N_11248);
or U13848 (N_13848,N_6024,N_10133);
and U13849 (N_13849,N_7201,N_7790);
and U13850 (N_13850,N_7294,N_7531);
and U13851 (N_13851,N_9691,N_10496);
nand U13852 (N_13852,N_7766,N_9745);
or U13853 (N_13853,N_8655,N_6034);
and U13854 (N_13854,N_8236,N_7841);
and U13855 (N_13855,N_7449,N_11680);
nand U13856 (N_13856,N_9058,N_7966);
or U13857 (N_13857,N_8392,N_7489);
and U13858 (N_13858,N_9051,N_11031);
or U13859 (N_13859,N_6405,N_6135);
xor U13860 (N_13860,N_6641,N_6893);
xor U13861 (N_13861,N_10954,N_11071);
nand U13862 (N_13862,N_9177,N_11057);
nor U13863 (N_13863,N_7272,N_11567);
xor U13864 (N_13864,N_8069,N_6782);
or U13865 (N_13865,N_10981,N_7151);
and U13866 (N_13866,N_8002,N_9116);
xnor U13867 (N_13867,N_10298,N_7979);
nand U13868 (N_13868,N_11103,N_11251);
nand U13869 (N_13869,N_6938,N_11852);
nor U13870 (N_13870,N_6335,N_6145);
nand U13871 (N_13871,N_11548,N_6763);
or U13872 (N_13872,N_10828,N_9578);
nor U13873 (N_13873,N_11453,N_9204);
nor U13874 (N_13874,N_11124,N_6614);
xnor U13875 (N_13875,N_10514,N_7467);
xnor U13876 (N_13876,N_9840,N_8507);
or U13877 (N_13877,N_6506,N_9588);
xnor U13878 (N_13878,N_9049,N_8680);
nand U13879 (N_13879,N_7083,N_9280);
nor U13880 (N_13880,N_9601,N_9395);
nand U13881 (N_13881,N_8789,N_6819);
xor U13882 (N_13882,N_9152,N_10846);
and U13883 (N_13883,N_11010,N_6207);
nor U13884 (N_13884,N_10494,N_8436);
and U13885 (N_13885,N_8380,N_6055);
or U13886 (N_13886,N_10475,N_9275);
nor U13887 (N_13887,N_7872,N_7453);
and U13888 (N_13888,N_7805,N_9956);
nor U13889 (N_13889,N_8895,N_10059);
and U13890 (N_13890,N_8750,N_7159);
nand U13891 (N_13891,N_11816,N_11315);
and U13892 (N_13892,N_7969,N_6328);
and U13893 (N_13893,N_10903,N_10698);
or U13894 (N_13894,N_9854,N_9962);
xnor U13895 (N_13895,N_11220,N_6858);
xor U13896 (N_13896,N_7809,N_11964);
and U13897 (N_13897,N_6789,N_6919);
and U13898 (N_13898,N_8328,N_9890);
and U13899 (N_13899,N_6005,N_10365);
xor U13900 (N_13900,N_7896,N_7291);
or U13901 (N_13901,N_8196,N_9470);
xnor U13902 (N_13902,N_7789,N_9191);
xnor U13903 (N_13903,N_11921,N_8930);
xor U13904 (N_13904,N_10543,N_8639);
xnor U13905 (N_13905,N_6872,N_9686);
nor U13906 (N_13906,N_8323,N_8338);
or U13907 (N_13907,N_9967,N_7256);
nand U13908 (N_13908,N_10537,N_6000);
or U13909 (N_13909,N_10399,N_10928);
xnor U13910 (N_13910,N_8167,N_10163);
and U13911 (N_13911,N_11201,N_10218);
nand U13912 (N_13912,N_11917,N_10116);
nand U13913 (N_13913,N_9325,N_6392);
and U13914 (N_13914,N_11691,N_11494);
and U13915 (N_13915,N_10693,N_9818);
xnor U13916 (N_13916,N_10862,N_7240);
or U13917 (N_13917,N_10275,N_11227);
nor U13918 (N_13918,N_11709,N_7605);
nand U13919 (N_13919,N_6464,N_9283);
nor U13920 (N_13920,N_11961,N_9683);
and U13921 (N_13921,N_11116,N_11243);
or U13922 (N_13922,N_9287,N_8341);
nor U13923 (N_13923,N_8898,N_10157);
nand U13924 (N_13924,N_9438,N_6886);
xor U13925 (N_13925,N_8106,N_11069);
nand U13926 (N_13926,N_9260,N_11991);
and U13927 (N_13927,N_10584,N_9016);
and U13928 (N_13928,N_7759,N_10021);
nand U13929 (N_13929,N_6834,N_11235);
xnor U13930 (N_13930,N_10705,N_10546);
or U13931 (N_13931,N_6691,N_7628);
xnor U13932 (N_13932,N_10125,N_8755);
or U13933 (N_13933,N_10210,N_8849);
nand U13934 (N_13934,N_11737,N_6236);
nand U13935 (N_13935,N_7625,N_8704);
nand U13936 (N_13936,N_6462,N_7604);
nor U13937 (N_13937,N_6166,N_10799);
nor U13938 (N_13938,N_8982,N_9240);
xor U13939 (N_13939,N_10676,N_9775);
nand U13940 (N_13940,N_6126,N_10002);
and U13941 (N_13941,N_8889,N_7946);
nand U13942 (N_13942,N_11255,N_9959);
nor U13943 (N_13943,N_9736,N_11508);
or U13944 (N_13944,N_6326,N_10706);
or U13945 (N_13945,N_6204,N_6689);
or U13946 (N_13946,N_10414,N_8396);
nor U13947 (N_13947,N_10085,N_6423);
or U13948 (N_13948,N_6089,N_11060);
nor U13949 (N_13949,N_8174,N_8020);
nand U13950 (N_13950,N_7861,N_6738);
and U13951 (N_13951,N_9440,N_10777);
or U13952 (N_13952,N_9924,N_10315);
nor U13953 (N_13953,N_10005,N_11587);
xnor U13954 (N_13954,N_10413,N_9678);
or U13955 (N_13955,N_8178,N_10719);
nand U13956 (N_13956,N_11799,N_8367);
nand U13957 (N_13957,N_11715,N_6284);
nor U13958 (N_13958,N_11757,N_8066);
nor U13959 (N_13959,N_6188,N_9471);
nand U13960 (N_13960,N_10107,N_8006);
and U13961 (N_13961,N_8546,N_9358);
and U13962 (N_13962,N_11173,N_6616);
nand U13963 (N_13963,N_9528,N_11884);
xnor U13964 (N_13964,N_9996,N_11034);
xor U13965 (N_13965,N_8964,N_6678);
xor U13966 (N_13966,N_8254,N_7660);
nor U13967 (N_13967,N_8648,N_9104);
and U13968 (N_13968,N_10039,N_8645);
xor U13969 (N_13969,N_6753,N_7199);
or U13970 (N_13970,N_6427,N_7470);
nor U13971 (N_13971,N_11663,N_11440);
xor U13972 (N_13972,N_7836,N_10420);
nand U13973 (N_13973,N_11791,N_11275);
or U13974 (N_13974,N_7838,N_6237);
nor U13975 (N_13975,N_6192,N_11908);
nor U13976 (N_13976,N_9971,N_10727);
nand U13977 (N_13977,N_11952,N_9565);
nand U13978 (N_13978,N_9920,N_8863);
xnor U13979 (N_13979,N_7793,N_7046);
nor U13980 (N_13980,N_11019,N_11911);
nand U13981 (N_13981,N_8593,N_7308);
and U13982 (N_13982,N_7853,N_7488);
nand U13983 (N_13983,N_8659,N_7369);
nor U13984 (N_13984,N_10338,N_9264);
nor U13985 (N_13985,N_11053,N_7592);
nand U13986 (N_13986,N_6837,N_6021);
xnor U13987 (N_13987,N_7618,N_6711);
nor U13988 (N_13988,N_11364,N_9003);
or U13989 (N_13989,N_8928,N_9209);
nand U13990 (N_13990,N_7816,N_10977);
and U13991 (N_13991,N_6121,N_6960);
xor U13992 (N_13992,N_11557,N_9567);
nand U13993 (N_13993,N_11625,N_10084);
nor U13994 (N_13994,N_11749,N_11389);
xor U13995 (N_13995,N_8077,N_7160);
or U13996 (N_13996,N_8453,N_10318);
and U13997 (N_13997,N_7659,N_7627);
or U13998 (N_13998,N_11563,N_9347);
nand U13999 (N_13999,N_7435,N_9045);
xor U14000 (N_14000,N_7241,N_7013);
or U14001 (N_14001,N_11500,N_11126);
nand U14002 (N_14002,N_9210,N_9687);
nor U14003 (N_14003,N_7102,N_8792);
or U14004 (N_14004,N_10658,N_6353);
xnor U14005 (N_14005,N_8314,N_10352);
and U14006 (N_14006,N_10605,N_9329);
nor U14007 (N_14007,N_7968,N_8881);
and U14008 (N_14008,N_11303,N_11692);
or U14009 (N_14009,N_9125,N_7832);
or U14010 (N_14010,N_8433,N_8470);
nor U14011 (N_14011,N_9810,N_6349);
xor U14012 (N_14012,N_11431,N_6577);
xnor U14013 (N_14013,N_11136,N_7171);
nand U14014 (N_14014,N_11919,N_11318);
and U14015 (N_14015,N_6544,N_7986);
and U14016 (N_14016,N_9676,N_10443);
or U14017 (N_14017,N_9761,N_10506);
or U14018 (N_14018,N_10808,N_10253);
xnor U14019 (N_14019,N_11786,N_7206);
nand U14020 (N_14020,N_7791,N_7723);
nor U14021 (N_14021,N_9904,N_11237);
xnor U14022 (N_14022,N_11062,N_9849);
nor U14023 (N_14023,N_10956,N_11120);
or U14024 (N_14024,N_8919,N_10243);
or U14025 (N_14025,N_10696,N_8899);
nor U14026 (N_14026,N_7480,N_11843);
nand U14027 (N_14027,N_9554,N_11435);
and U14028 (N_14028,N_9221,N_11858);
or U14029 (N_14029,N_9911,N_8920);
and U14030 (N_14030,N_7856,N_11597);
nor U14031 (N_14031,N_7676,N_8019);
nand U14032 (N_14032,N_7926,N_11441);
nor U14033 (N_14033,N_8553,N_11401);
or U14034 (N_14034,N_6647,N_7496);
nand U14035 (N_14035,N_8513,N_7131);
and U14036 (N_14036,N_11574,N_11844);
xnor U14037 (N_14037,N_11829,N_7208);
and U14038 (N_14038,N_9348,N_9873);
nor U14039 (N_14039,N_6282,N_11564);
xor U14040 (N_14040,N_10367,N_7711);
nand U14041 (N_14041,N_8609,N_11613);
nand U14042 (N_14042,N_11443,N_7826);
and U14043 (N_14043,N_10920,N_8775);
nor U14044 (N_14044,N_8429,N_6003);
or U14045 (N_14045,N_11039,N_11870);
or U14046 (N_14046,N_6670,N_6956);
nor U14047 (N_14047,N_10460,N_10798);
nor U14048 (N_14048,N_7778,N_9425);
and U14049 (N_14049,N_7050,N_10678);
nor U14050 (N_14050,N_11658,N_7126);
nor U14051 (N_14051,N_6189,N_9030);
nand U14052 (N_14052,N_9774,N_9688);
nand U14053 (N_14053,N_10242,N_11101);
xor U14054 (N_14054,N_8532,N_9046);
or U14055 (N_14055,N_7774,N_7204);
xnor U14056 (N_14056,N_11141,N_8821);
nand U14057 (N_14057,N_10416,N_7910);
and U14058 (N_14058,N_10048,N_10908);
and U14059 (N_14059,N_6760,N_6582);
xnor U14060 (N_14060,N_7197,N_7950);
and U14061 (N_14061,N_7781,N_7709);
nor U14062 (N_14062,N_9743,N_6369);
xor U14063 (N_14063,N_7066,N_9817);
xnor U14064 (N_14064,N_8013,N_6805);
and U14065 (N_14065,N_9724,N_7146);
nor U14066 (N_14066,N_8202,N_9509);
xor U14067 (N_14067,N_7120,N_7637);
xnor U14068 (N_14068,N_11906,N_6968);
nor U14069 (N_14069,N_9981,N_10078);
xor U14070 (N_14070,N_10346,N_6957);
nand U14071 (N_14071,N_11091,N_8843);
and U14072 (N_14072,N_7117,N_10486);
or U14073 (N_14073,N_7113,N_9696);
nand U14074 (N_14074,N_10030,N_11552);
nand U14075 (N_14075,N_10623,N_11683);
and U14076 (N_14076,N_10427,N_11707);
nand U14077 (N_14077,N_8122,N_8547);
and U14078 (N_14078,N_6923,N_9529);
nand U14079 (N_14079,N_7491,N_6315);
nor U14080 (N_14080,N_10893,N_6926);
xor U14081 (N_14081,N_8897,N_11743);
or U14082 (N_14082,N_9742,N_6486);
xor U14083 (N_14083,N_7086,N_6426);
and U14084 (N_14084,N_7840,N_8377);
and U14085 (N_14085,N_9782,N_6721);
nand U14086 (N_14086,N_7599,N_8939);
nor U14087 (N_14087,N_9142,N_10817);
or U14088 (N_14088,N_6642,N_7414);
xor U14089 (N_14089,N_6447,N_7956);
nand U14090 (N_14090,N_9241,N_10027);
or U14091 (N_14091,N_8806,N_6595);
xor U14092 (N_14092,N_11970,N_6453);
xor U14093 (N_14093,N_8390,N_11965);
xor U14094 (N_14094,N_6787,N_11348);
nand U14095 (N_14095,N_11000,N_10104);
xnor U14096 (N_14096,N_9927,N_10351);
and U14097 (N_14097,N_9666,N_9617);
and U14098 (N_14098,N_11969,N_8102);
nor U14099 (N_14099,N_7632,N_10080);
or U14100 (N_14100,N_9532,N_8893);
and U14101 (N_14101,N_10099,N_9987);
nor U14102 (N_14102,N_10666,N_8256);
or U14103 (N_14103,N_8957,N_7337);
or U14104 (N_14104,N_9416,N_8158);
nor U14105 (N_14105,N_11004,N_6124);
and U14106 (N_14106,N_9861,N_10936);
and U14107 (N_14107,N_9659,N_8555);
and U14108 (N_14108,N_7459,N_9127);
or U14109 (N_14109,N_11181,N_6849);
nor U14110 (N_14110,N_7154,N_10226);
nor U14111 (N_14111,N_11198,N_9265);
or U14112 (N_14112,N_7577,N_6295);
nand U14113 (N_14113,N_9543,N_8620);
and U14114 (N_14114,N_10655,N_11561);
xor U14115 (N_14115,N_6722,N_10150);
xnor U14116 (N_14116,N_10939,N_9402);
xor U14117 (N_14117,N_10973,N_6450);
nand U14118 (N_14118,N_6058,N_10390);
nor U14119 (N_14119,N_7652,N_6973);
nand U14120 (N_14120,N_9776,N_10287);
nor U14121 (N_14121,N_11300,N_11590);
and U14122 (N_14122,N_7691,N_8322);
nor U14123 (N_14123,N_6180,N_6799);
nor U14124 (N_14124,N_9398,N_9269);
nand U14125 (N_14125,N_9710,N_10955);
xnor U14126 (N_14126,N_8312,N_9119);
xnor U14127 (N_14127,N_9014,N_11787);
nor U14128 (N_14128,N_8239,N_8848);
xnor U14129 (N_14129,N_7922,N_11505);
or U14130 (N_14130,N_8979,N_8098);
nor U14131 (N_14131,N_11211,N_7089);
and U14132 (N_14132,N_9433,N_8081);
xnor U14133 (N_14133,N_6465,N_11665);
or U14134 (N_14134,N_10052,N_10184);
and U14135 (N_14135,N_10177,N_11729);
nand U14136 (N_14136,N_10195,N_10354);
and U14137 (N_14137,N_9560,N_7608);
or U14138 (N_14138,N_8089,N_6547);
and U14139 (N_14139,N_9111,N_10659);
nand U14140 (N_14140,N_6972,N_6362);
or U14141 (N_14141,N_6839,N_8596);
nand U14142 (N_14142,N_10761,N_6181);
and U14143 (N_14143,N_9767,N_10829);
and U14144 (N_14144,N_8387,N_8822);
or U14145 (N_14145,N_11527,N_7622);
xnor U14146 (N_14146,N_9898,N_8084);
nand U14147 (N_14147,N_9644,N_7621);
xor U14148 (N_14148,N_8777,N_6558);
xnor U14149 (N_14149,N_9059,N_8046);
nor U14150 (N_14150,N_10733,N_7429);
xor U14151 (N_14151,N_11017,N_7513);
nand U14152 (N_14152,N_8768,N_9355);
and U14153 (N_14153,N_11883,N_9777);
nand U14154 (N_14154,N_10519,N_11388);
xor U14155 (N_14155,N_7748,N_8580);
or U14156 (N_14156,N_11599,N_11025);
nor U14157 (N_14157,N_6245,N_9918);
nand U14158 (N_14158,N_10809,N_9510);
nor U14159 (N_14159,N_7976,N_6198);
and U14160 (N_14160,N_7714,N_10811);
or U14161 (N_14161,N_11810,N_10697);
xnor U14162 (N_14162,N_8743,N_9499);
or U14163 (N_14163,N_6377,N_11877);
nand U14164 (N_14164,N_10885,N_6690);
nor U14165 (N_14165,N_9975,N_7544);
nand U14166 (N_14166,N_9176,N_8776);
xnor U14167 (N_14167,N_8867,N_9442);
and U14168 (N_14168,N_6997,N_7874);
nand U14169 (N_14169,N_8375,N_7017);
nand U14170 (N_14170,N_8859,N_10933);
nor U14171 (N_14171,N_6442,N_7070);
xor U14172 (N_14172,N_7316,N_6484);
nor U14173 (N_14173,N_10883,N_9624);
or U14174 (N_14174,N_8583,N_6596);
nand U14175 (N_14175,N_8643,N_11895);
xnor U14176 (N_14176,N_8067,N_11223);
xnor U14177 (N_14177,N_7601,N_8707);
and U14178 (N_14178,N_6871,N_7338);
and U14179 (N_14179,N_8969,N_11386);
nand U14180 (N_14180,N_6396,N_11205);
and U14181 (N_14181,N_6154,N_6672);
and U14182 (N_14182,N_7525,N_7725);
nor U14183 (N_14183,N_8488,N_9968);
nand U14184 (N_14184,N_6312,N_8838);
nand U14185 (N_14185,N_11848,N_9284);
and U14186 (N_14186,N_7900,N_8896);
xor U14187 (N_14187,N_6730,N_9786);
or U14188 (N_14188,N_6657,N_10663);
nand U14189 (N_14189,N_7277,N_9497);
nor U14190 (N_14190,N_7708,N_6436);
and U14191 (N_14191,N_9819,N_8511);
and U14192 (N_14192,N_6191,N_8606);
nor U14193 (N_14193,N_9285,N_9643);
nand U14194 (N_14194,N_8934,N_10441);
and U14195 (N_14195,N_7186,N_11027);
or U14196 (N_14196,N_7313,N_6195);
or U14197 (N_14197,N_10086,N_7464);
xnor U14198 (N_14198,N_9229,N_6495);
and U14199 (N_14199,N_10302,N_6431);
or U14200 (N_14200,N_10091,N_11617);
or U14201 (N_14201,N_11397,N_6985);
xnor U14202 (N_14202,N_10558,N_11048);
or U14203 (N_14203,N_7865,N_9599);
and U14204 (N_14204,N_11975,N_11290);
nand U14205 (N_14205,N_8273,N_11948);
nor U14206 (N_14206,N_8347,N_9731);
xor U14207 (N_14207,N_9547,N_8209);
nand U14208 (N_14208,N_8980,N_8103);
and U14209 (N_14209,N_6513,N_9764);
nand U14210 (N_14210,N_10273,N_9878);
nand U14211 (N_14211,N_7536,N_9734);
and U14212 (N_14212,N_9979,N_9748);
xor U14213 (N_14213,N_6942,N_10062);
and U14214 (N_14214,N_10363,N_6244);
nor U14215 (N_14215,N_6560,N_8192);
nand U14216 (N_14216,N_8790,N_7697);
and U14217 (N_14217,N_11967,N_7405);
xnor U14218 (N_14218,N_11184,N_8900);
or U14219 (N_14219,N_9493,N_11532);
xor U14220 (N_14220,N_6366,N_8223);
nand U14221 (N_14221,N_9294,N_7378);
or U14222 (N_14222,N_8471,N_11461);
nor U14223 (N_14223,N_11558,N_7327);
or U14224 (N_14224,N_8219,N_7090);
xor U14225 (N_14225,N_10293,N_8785);
nand U14226 (N_14226,N_7547,N_10487);
or U14227 (N_14227,N_9047,N_7260);
xor U14228 (N_14228,N_9399,N_7307);
and U14229 (N_14229,N_7330,N_7773);
xor U14230 (N_14230,N_9612,N_6842);
nor U14231 (N_14231,N_11712,N_6660);
xor U14232 (N_14232,N_10934,N_11106);
and U14233 (N_14233,N_10466,N_7468);
nand U14234 (N_14234,N_11998,N_7626);
and U14235 (N_14235,N_7409,N_7717);
or U14236 (N_14236,N_8537,N_10578);
nor U14237 (N_14237,N_8009,N_10997);
and U14238 (N_14238,N_7030,N_9940);
nand U14239 (N_14239,N_8206,N_10329);
and U14240 (N_14240,N_7136,N_10247);
nand U14241 (N_14241,N_6178,N_7335);
or U14242 (N_14242,N_9932,N_7466);
nand U14243 (N_14243,N_6242,N_6716);
nand U14244 (N_14244,N_11475,N_7242);
and U14245 (N_14245,N_9133,N_8120);
xnor U14246 (N_14246,N_11015,N_6358);
and U14247 (N_14247,N_10309,N_8812);
and U14248 (N_14248,N_8088,N_11868);
nor U14249 (N_14249,N_11800,N_8063);
or U14250 (N_14250,N_9435,N_6904);
xnor U14251 (N_14251,N_11690,N_10193);
and U14252 (N_14252,N_8763,N_7379);
nand U14253 (N_14253,N_9838,N_6847);
or U14254 (N_14254,N_6797,N_8803);
nand U14255 (N_14255,N_6961,N_6561);
or U14256 (N_14256,N_6541,N_10425);
and U14257 (N_14257,N_10160,N_10436);
and U14258 (N_14258,N_10959,N_11924);
xnor U14259 (N_14259,N_10847,N_10641);
nor U14260 (N_14260,N_6421,N_10837);
xor U14261 (N_14261,N_10793,N_10911);
or U14262 (N_14262,N_8091,N_11465);
xnor U14263 (N_14263,N_8248,N_11539);
or U14264 (N_14264,N_7670,N_11693);
and U14265 (N_14265,N_7252,N_9846);
xor U14266 (N_14266,N_7245,N_8288);
nor U14267 (N_14267,N_6020,N_9415);
nor U14268 (N_14268,N_8516,N_7244);
xnor U14269 (N_14269,N_10146,N_11867);
nor U14270 (N_14270,N_11656,N_10434);
and U14271 (N_14271,N_10464,N_9278);
and U14272 (N_14272,N_9800,N_8845);
and U14273 (N_14273,N_11032,N_8985);
xnor U14274 (N_14274,N_11946,N_8082);
nand U14275 (N_14275,N_11138,N_9212);
or U14276 (N_14276,N_10967,N_6930);
xor U14277 (N_14277,N_11074,N_8182);
nor U14278 (N_14278,N_7289,N_9391);
and U14279 (N_14279,N_9390,N_7135);
and U14280 (N_14280,N_6626,N_8868);
xnor U14281 (N_14281,N_6289,N_8936);
or U14282 (N_14282,N_8693,N_6002);
nor U14283 (N_14283,N_11640,N_8211);
xnor U14284 (N_14284,N_11543,N_6808);
or U14285 (N_14285,N_11949,N_11125);
and U14286 (N_14286,N_7792,N_8563);
xnor U14287 (N_14287,N_8302,N_6470);
xor U14288 (N_14288,N_8837,N_9397);
and U14289 (N_14289,N_11668,N_9814);
nor U14290 (N_14290,N_8675,N_6137);
or U14291 (N_14291,N_6896,N_8324);
xnor U14292 (N_14292,N_11595,N_8955);
and U14293 (N_14293,N_9144,N_9751);
xor U14294 (N_14294,N_7579,N_6302);
xnor U14295 (N_14295,N_11109,N_6802);
xnor U14296 (N_14296,N_9790,N_6655);
nand U14297 (N_14297,N_6079,N_10560);
or U14298 (N_14298,N_10701,N_6156);
xor U14299 (N_14299,N_6232,N_10670);
nor U14300 (N_14300,N_9937,N_11694);
nand U14301 (N_14301,N_7354,N_9651);
or U14302 (N_14302,N_9787,N_10499);
nor U14303 (N_14303,N_8143,N_10520);
xor U14304 (N_14304,N_10169,N_10307);
xor U14305 (N_14305,N_10866,N_10249);
nor U14306 (N_14306,N_10305,N_11023);
and U14307 (N_14307,N_6281,N_8191);
nand U14308 (N_14308,N_7499,N_8748);
or U14309 (N_14309,N_8509,N_6988);
nor U14310 (N_14310,N_9874,N_11130);
nand U14311 (N_14311,N_8572,N_8626);
nand U14312 (N_14312,N_6739,N_9446);
nor U14313 (N_14313,N_11155,N_11781);
nand U14314 (N_14314,N_6549,N_9960);
and U14315 (N_14315,N_10320,N_6889);
xor U14316 (N_14316,N_8963,N_6460);
nor U14317 (N_14317,N_11285,N_7318);
xnor U14318 (N_14318,N_10646,N_7895);
and U14319 (N_14319,N_9453,N_11194);
nor U14320 (N_14320,N_7372,N_8449);
nand U14321 (N_14321,N_11246,N_11414);
xor U14322 (N_14322,N_8698,N_10217);
or U14323 (N_14323,N_8649,N_9215);
and U14324 (N_14324,N_11582,N_9094);
nor U14325 (N_14325,N_10895,N_10404);
nand U14326 (N_14326,N_10103,N_6357);
and U14327 (N_14327,N_10355,N_9199);
xnor U14328 (N_14328,N_11197,N_10723);
or U14329 (N_14329,N_10910,N_8198);
or U14330 (N_14330,N_10083,N_7202);
nor U14331 (N_14331,N_10187,N_7947);
and U14332 (N_14332,N_10001,N_6239);
or U14333 (N_14333,N_6440,N_7607);
xnor U14334 (N_14334,N_7118,N_11611);
nand U14335 (N_14335,N_10162,N_11410);
xnor U14336 (N_14336,N_9900,N_9375);
and U14337 (N_14337,N_10250,N_8021);
nand U14338 (N_14338,N_11249,N_11854);
or U14339 (N_14339,N_10568,N_11660);
or U14340 (N_14340,N_9802,N_11079);
nand U14341 (N_14341,N_11727,N_8579);
xnor U14342 (N_14342,N_6533,N_8000);
and U14343 (N_14343,N_11622,N_7845);
nor U14344 (N_14344,N_9118,N_9847);
nand U14345 (N_14345,N_6897,N_11553);
and U14346 (N_14346,N_11002,N_9253);
nand U14347 (N_14347,N_8888,N_8094);
or U14348 (N_14348,N_7876,N_8296);
and U14349 (N_14349,N_8221,N_10183);
and U14350 (N_14350,N_7145,N_10897);
or U14351 (N_14351,N_9781,N_8435);
or U14352 (N_14352,N_8847,N_9841);
and U14353 (N_14353,N_6311,N_7333);
or U14354 (N_14354,N_10403,N_8582);
nor U14355 (N_14355,N_11682,N_9997);
xor U14356 (N_14356,N_7115,N_9609);
xnor U14357 (N_14357,N_7417,N_11411);
xnor U14358 (N_14358,N_8190,N_9450);
nor U14359 (N_14359,N_7854,N_11413);
or U14360 (N_14360,N_8754,N_9457);
nand U14361 (N_14361,N_8633,N_7325);
and U14362 (N_14362,N_9881,N_8154);
nand U14363 (N_14363,N_11703,N_6380);
nand U14364 (N_14364,N_10228,N_8173);
nor U14365 (N_14365,N_10938,N_8781);
and U14366 (N_14366,N_6652,N_9034);
xnor U14367 (N_14367,N_7729,N_6006);
or U14368 (N_14368,N_8793,N_11838);
xor U14369 (N_14369,N_11718,N_6989);
nand U14370 (N_14370,N_6515,N_11302);
xnor U14371 (N_14371,N_7661,N_8756);
xnor U14372 (N_14372,N_8345,N_9746);
or U14373 (N_14373,N_10561,N_11677);
nand U14374 (N_14374,N_8521,N_11487);
xnor U14375 (N_14375,N_11896,N_10629);
nand U14376 (N_14376,N_9407,N_6877);
nand U14377 (N_14377,N_8151,N_9393);
or U14378 (N_14378,N_7576,N_10988);
nor U14379 (N_14379,N_8093,N_11425);
nand U14380 (N_14380,N_6449,N_6525);
nand U14381 (N_14381,N_9052,N_8558);
nor U14382 (N_14382,N_9851,N_8437);
and U14383 (N_14383,N_6575,N_11769);
and U14384 (N_14384,N_8916,N_6404);
xor U14385 (N_14385,N_11187,N_11929);
or U14386 (N_14386,N_7049,N_8403);
and U14387 (N_14387,N_6658,N_8123);
xnor U14388 (N_14388,N_9941,N_10167);
or U14389 (N_14389,N_6903,N_6102);
nor U14390 (N_14390,N_10765,N_8142);
nor U14391 (N_14391,N_6011,N_6016);
nand U14392 (N_14392,N_10840,N_7034);
or U14393 (N_14393,N_6894,N_8614);
xnor U14394 (N_14394,N_10649,N_6010);
nand U14395 (N_14395,N_9680,N_7564);
or U14396 (N_14396,N_10389,N_10266);
xor U14397 (N_14397,N_11083,N_10444);
and U14398 (N_14398,N_10672,N_9206);
or U14399 (N_14399,N_11835,N_9939);
or U14400 (N_14400,N_6076,N_9718);
or U14401 (N_14401,N_6592,N_10740);
or U14402 (N_14402,N_6061,N_6433);
or U14403 (N_14403,N_8136,N_9309);
and U14404 (N_14404,N_11078,N_6634);
or U14405 (N_14405,N_7038,N_7237);
or U14406 (N_14406,N_9261,N_11824);
nand U14407 (N_14407,N_9525,N_9143);
or U14408 (N_14408,N_11218,N_10753);
nand U14409 (N_14409,N_8401,N_6482);
xnor U14410 (N_14410,N_11021,N_9019);
and U14411 (N_14411,N_10613,N_6729);
and U14412 (N_14412,N_7800,N_6138);
nor U14413 (N_14413,N_8053,N_9673);
nor U14414 (N_14414,N_11128,N_6163);
nor U14415 (N_14415,N_9336,N_10553);
or U14416 (N_14416,N_6143,N_9303);
nor U14417 (N_14417,N_7055,N_8064);
or U14418 (N_14418,N_10987,N_7373);
nor U14419 (N_14419,N_10597,N_9055);
or U14420 (N_14420,N_10542,N_7376);
and U14421 (N_14421,N_11596,N_10971);
xnor U14422 (N_14422,N_10563,N_10380);
nor U14423 (N_14423,N_10057,N_11271);
nand U14424 (N_14424,N_8925,N_6097);
and U14425 (N_14425,N_7292,N_10530);
or U14426 (N_14426,N_8065,N_8736);
nor U14427 (N_14427,N_6443,N_7819);
or U14428 (N_14428,N_9885,N_7891);
nand U14429 (N_14429,N_9517,N_9274);
or U14430 (N_14430,N_7962,N_6209);
nor U14431 (N_14431,N_11764,N_8458);
and U14432 (N_14432,N_9737,N_6355);
or U14433 (N_14433,N_7762,N_9054);
and U14434 (N_14434,N_6580,N_9173);
nand U14435 (N_14435,N_8057,N_10035);
nand U14436 (N_14436,N_7901,N_9394);
nor U14437 (N_14437,N_7837,N_8090);
or U14438 (N_14438,N_6338,N_6978);
nand U14439 (N_14439,N_8070,N_11481);
nand U14440 (N_14440,N_8011,N_11380);
xor U14441 (N_14441,N_6674,N_6134);
xor U14442 (N_14442,N_8135,N_11421);
nor U14443 (N_14443,N_6941,N_7306);
nor U14444 (N_14444,N_11637,N_10402);
nor U14445 (N_14445,N_11104,N_10842);
xnor U14446 (N_14446,N_10854,N_6361);
and U14447 (N_14447,N_8510,N_11045);
or U14448 (N_14448,N_10592,N_10918);
and U14449 (N_14449,N_10785,N_6869);
nor U14450 (N_14450,N_11889,N_8752);
and U14451 (N_14451,N_8817,N_11154);
and U14452 (N_14452,N_10631,N_11859);
xor U14453 (N_14453,N_6485,N_10556);
xnor U14454 (N_14454,N_7743,N_7584);
nor U14455 (N_14455,N_9974,N_6598);
nor U14456 (N_14456,N_7951,N_11219);
nand U14457 (N_14457,N_6999,N_6824);
xor U14458 (N_14458,N_7849,N_6940);
nor U14459 (N_14459,N_10870,N_6706);
and U14460 (N_14460,N_7539,N_6331);
nor U14461 (N_14461,N_9237,N_7596);
nor U14462 (N_14462,N_9349,N_8855);
or U14463 (N_14463,N_11681,N_7048);
nand U14464 (N_14464,N_9369,N_10147);
or U14465 (N_14465,N_10406,N_10836);
and U14466 (N_14466,N_10657,N_11454);
or U14467 (N_14467,N_10772,N_11979);
or U14468 (N_14468,N_9552,N_6759);
nand U14469 (N_14469,N_10832,N_9541);
xnor U14470 (N_14470,N_9698,N_7650);
nand U14471 (N_14471,N_6095,N_10861);
and U14472 (N_14472,N_7533,N_7261);
and U14473 (N_14473,N_10431,N_9894);
and U14474 (N_14474,N_6360,N_8005);
nand U14475 (N_14475,N_11788,N_6019);
xnor U14476 (N_14476,N_9243,N_8291);
and U14477 (N_14477,N_11711,N_9821);
nor U14478 (N_14478,N_6701,N_7722);
nand U14479 (N_14479,N_10826,N_10689);
xor U14480 (N_14480,N_9756,N_7304);
xnor U14481 (N_14481,N_6139,N_8906);
xor U14482 (N_14482,N_8551,N_10100);
xnor U14483 (N_14483,N_10430,N_10850);
or U14484 (N_14484,N_10626,N_9352);
nand U14485 (N_14485,N_11252,N_7207);
nor U14486 (N_14486,N_9321,N_11922);
nand U14487 (N_14487,N_10963,N_6906);
and U14488 (N_14488,N_7927,N_10232);
nor U14489 (N_14489,N_9610,N_9131);
xor U14490 (N_14490,N_11634,N_6609);
nor U14491 (N_14491,N_7881,N_6321);
nor U14492 (N_14492,N_7040,N_11072);
xor U14493 (N_14493,N_8118,N_9855);
or U14494 (N_14494,N_9744,N_10650);
or U14495 (N_14495,N_8738,N_6364);
nand U14496 (N_14496,N_6600,N_8718);
nor U14497 (N_14497,N_11381,N_7815);
and U14498 (N_14498,N_6682,N_11837);
xor U14499 (N_14499,N_9262,N_10012);
nand U14500 (N_14500,N_8140,N_10776);
nor U14501 (N_14501,N_8814,N_8962);
and U14502 (N_14502,N_10373,N_10033);
nand U14503 (N_14503,N_8749,N_9362);
nor U14504 (N_14504,N_9551,N_11145);
or U14505 (N_14505,N_11075,N_10041);
nor U14506 (N_14506,N_7530,N_11783);
or U14507 (N_14507,N_8358,N_9783);
nor U14508 (N_14508,N_10478,N_8520);
or U14509 (N_14509,N_9558,N_8229);
and U14510 (N_14510,N_11332,N_10940);
and U14511 (N_14511,N_11978,N_6398);
and U14512 (N_14512,N_9203,N_11107);
nand U14513 (N_14513,N_10094,N_10140);
and U14514 (N_14514,N_9793,N_8270);
nor U14515 (N_14515,N_11297,N_10222);
nand U14516 (N_14516,N_8407,N_9135);
nand U14517 (N_14517,N_8646,N_6354);
xor U14518 (N_14518,N_11934,N_11820);
or U14519 (N_14519,N_11847,N_6509);
or U14520 (N_14520,N_9999,N_8996);
xnor U14521 (N_14521,N_7945,N_10236);
or U14522 (N_14522,N_8402,N_9899);
xor U14523 (N_14523,N_11566,N_11554);
nor U14524 (N_14524,N_9090,N_7859);
nand U14525 (N_14525,N_8014,N_7930);
and U14526 (N_14526,N_8331,N_10134);
and U14527 (N_14527,N_10061,N_11517);
nor U14528 (N_14528,N_6221,N_7992);
nor U14529 (N_14529,N_6995,N_6528);
nor U14530 (N_14530,N_7067,N_9208);
and U14531 (N_14531,N_7287,N_8056);
xnor U14532 (N_14532,N_6761,N_8875);
nand U14533 (N_14533,N_6491,N_10339);
nor U14534 (N_14534,N_7645,N_6708);
nand U14535 (N_14535,N_7122,N_9170);
nand U14536 (N_14536,N_10333,N_8825);
nor U14537 (N_14537,N_10717,N_11409);
and U14538 (N_14538,N_10891,N_6272);
nand U14539 (N_14539,N_6344,N_6108);
and U14540 (N_14540,N_8247,N_9716);
xor U14541 (N_14541,N_9242,N_9078);
xor U14542 (N_14542,N_7597,N_10643);
nand U14543 (N_14543,N_9276,N_6408);
xor U14544 (N_14544,N_9953,N_6152);
xnor U14545 (N_14545,N_8371,N_10750);
and U14546 (N_14546,N_6397,N_6798);
and U14547 (N_14547,N_8087,N_6468);
nand U14548 (N_14548,N_7374,N_6317);
xnor U14549 (N_14549,N_11115,N_7570);
and U14550 (N_14550,N_7184,N_9608);
or U14551 (N_14551,N_6288,N_7238);
or U14552 (N_14552,N_10350,N_11944);
nand U14553 (N_14553,N_7970,N_10424);
or U14554 (N_14554,N_6013,N_9079);
or U14555 (N_14555,N_11496,N_8902);
and U14556 (N_14556,N_10300,N_6542);
xnor U14557 (N_14557,N_8304,N_10845);
nor U14558 (N_14558,N_6084,N_8215);
nand U14559 (N_14559,N_11134,N_10075);
and U14560 (N_14560,N_7806,N_6007);
nand U14561 (N_14561,N_8968,N_11989);
nand U14562 (N_14562,N_8523,N_8356);
nor U14563 (N_14563,N_10994,N_7008);
xor U14564 (N_14564,N_8425,N_10283);
nor U14565 (N_14565,N_9550,N_8300);
nor U14566 (N_14566,N_11400,N_8460);
nor U14567 (N_14567,N_6082,N_10265);
or U14568 (N_14568,N_9279,N_9516);
nor U14569 (N_14569,N_9923,N_8207);
nor U14570 (N_14570,N_11133,N_7358);
or U14571 (N_14571,N_10619,N_7190);
or U14572 (N_14572,N_7794,N_9646);
xnor U14573 (N_14573,N_11341,N_11857);
or U14574 (N_14574,N_6719,N_11306);
nor U14575 (N_14575,N_9850,N_10662);
nand U14576 (N_14576,N_10369,N_9963);
and U14577 (N_14577,N_9069,N_7425);
nor U14578 (N_14578,N_10786,N_10974);
nor U14579 (N_14579,N_9522,N_7235);
and U14580 (N_14580,N_10277,N_10122);
nand U14581 (N_14581,N_8366,N_7012);
and U14582 (N_14582,N_6599,N_6705);
nand U14583 (N_14583,N_11166,N_10079);
and U14584 (N_14584,N_10255,N_6454);
and U14585 (N_14585,N_9181,N_9164);
or U14586 (N_14586,N_7211,N_7999);
or U14587 (N_14587,N_6069,N_9592);
or U14588 (N_14588,N_9700,N_9196);
or U14589 (N_14589,N_10788,N_10323);
or U14590 (N_14590,N_9614,N_6882);
and U14591 (N_14591,N_8332,N_8483);
or U14592 (N_14592,N_7251,N_6668);
and U14593 (N_14593,N_6350,N_11631);
nor U14594 (N_14594,N_7077,N_11157);
and U14595 (N_14595,N_7458,N_7602);
or U14596 (N_14596,N_9747,N_6723);
or U14597 (N_14597,N_8492,N_8912);
xor U14598 (N_14598,N_10775,N_7924);
and U14599 (N_14599,N_9108,N_10068);
or U14600 (N_14600,N_11480,N_6814);
xor U14601 (N_14601,N_9995,N_9290);
or U14602 (N_14602,N_6308,N_10313);
nor U14603 (N_14603,N_7440,N_10647);
or U14604 (N_14604,N_11308,N_8352);
xor U14605 (N_14605,N_9458,N_8059);
nor U14606 (N_14606,N_7656,N_6952);
xnor U14607 (N_14607,N_8284,N_11261);
or U14608 (N_14608,N_11758,N_11834);
nor U14609 (N_14609,N_10755,N_7991);
or U14610 (N_14610,N_8921,N_6374);
or U14611 (N_14611,N_11993,N_11033);
nand U14612 (N_14612,N_11394,N_11580);
nand U14613 (N_14613,N_6794,N_6746);
nand U14614 (N_14614,N_7903,N_11818);
or U14615 (N_14615,N_7655,N_7402);
or U14616 (N_14616,N_9753,N_8426);
or U14617 (N_14617,N_11600,N_8654);
xor U14618 (N_14618,N_9025,N_7472);
nor U14619 (N_14619,N_7084,N_7299);
nor U14620 (N_14620,N_11550,N_11705);
or U14621 (N_14621,N_9339,N_9166);
or U14622 (N_14622,N_11925,N_7885);
or U14623 (N_14623,N_7810,N_10220);
xor U14624 (N_14624,N_8305,N_8976);
and U14625 (N_14625,N_11047,N_11132);
or U14626 (N_14626,N_10207,N_6681);
nor U14627 (N_14627,N_10132,N_11535);
nand U14628 (N_14628,N_6118,N_9672);
nor U14629 (N_14629,N_11473,N_8327);
and U14630 (N_14630,N_10025,N_8022);
or U14631 (N_14631,N_9771,N_10311);
and U14632 (N_14632,N_10397,N_8727);
nor U14633 (N_14633,N_7799,N_6836);
nand U14634 (N_14634,N_10683,N_11395);
nor U14635 (N_14635,N_11745,N_11688);
and U14636 (N_14636,N_9573,N_9353);
nor U14637 (N_14637,N_11876,N_10219);
nor U14638 (N_14638,N_10766,N_7104);
nor U14639 (N_14639,N_9882,N_7037);
and U14640 (N_14640,N_6445,N_10789);
and U14641 (N_14641,N_6367,N_6991);
nand U14642 (N_14642,N_10370,N_7983);
nor U14643 (N_14643,N_10129,N_6523);
xnor U14644 (N_14644,N_6855,N_8249);
nand U14645 (N_14645,N_10640,N_6130);
nand U14646 (N_14646,N_7940,N_8137);
and U14647 (N_14647,N_8966,N_10595);
xnor U14648 (N_14648,N_10694,N_9621);
and U14649 (N_14649,N_7283,N_6285);
xnor U14650 (N_14650,N_9649,N_8428);
xor U14651 (N_14651,N_9081,N_9848);
xor U14652 (N_14652,N_8072,N_10073);
xor U14653 (N_14653,N_9728,N_11873);
or U14654 (N_14654,N_8948,N_7255);
and U14655 (N_14655,N_7948,N_6099);
nor U14656 (N_14656,N_7462,N_9597);
nor U14657 (N_14657,N_9227,N_8640);
and U14658 (N_14658,N_10718,N_10155);
or U14659 (N_14659,N_8017,N_10092);
and U14660 (N_14660,N_9272,N_7552);
or U14661 (N_14661,N_8984,N_9063);
or U14662 (N_14662,N_7839,N_8451);
or U14663 (N_14663,N_11679,N_10098);
or U14664 (N_14664,N_6316,N_7534);
and U14665 (N_14665,N_8350,N_8760);
nand U14666 (N_14666,N_6269,N_9013);
and U14667 (N_14667,N_10156,N_6073);
nor U14668 (N_14668,N_6637,N_10884);
xor U14669 (N_14669,N_8224,N_8475);
nor U14670 (N_14670,N_7006,N_8788);
and U14671 (N_14671,N_7218,N_7137);
and U14672 (N_14672,N_8618,N_7747);
nand U14673 (N_14673,N_9921,N_10482);
or U14674 (N_14674,N_10965,N_7760);
and U14675 (N_14675,N_9334,N_8890);
or U14676 (N_14676,N_6254,N_7389);
or U14677 (N_14677,N_10652,N_8376);
or U14678 (N_14678,N_11052,N_8004);
or U14679 (N_14679,N_9357,N_8540);
and U14680 (N_14680,N_8044,N_8787);
nor U14681 (N_14681,N_8472,N_7902);
nand U14682 (N_14682,N_10047,N_8978);
and U14683 (N_14683,N_6158,N_8418);
and U14684 (N_14684,N_9559,N_6979);
and U14685 (N_14685,N_10065,N_10097);
xor U14686 (N_14686,N_11807,N_6042);
xor U14687 (N_14687,N_8667,N_8637);
and U14688 (N_14688,N_11833,N_9085);
and U14689 (N_14689,N_10878,N_8015);
xnor U14690 (N_14690,N_10935,N_7111);
or U14691 (N_14691,N_6524,N_8932);
nand U14692 (N_14692,N_7253,N_7912);
xor U14693 (N_14693,N_7174,N_8303);
nor U14694 (N_14694,N_11190,N_6593);
and U14695 (N_14695,N_7988,N_11491);
nor U14696 (N_14696,N_7931,N_11515);
xor U14697 (N_14697,N_7571,N_7823);
nand U14698 (N_14698,N_6075,N_9872);
nand U14699 (N_14699,N_6512,N_11836);
and U14700 (N_14700,N_8524,N_9149);
nand U14701 (N_14701,N_10322,N_6700);
xnor U14702 (N_14702,N_11263,N_8676);
xor U14703 (N_14703,N_10834,N_9035);
nand U14704 (N_14704,N_11093,N_8634);
nor U14705 (N_14705,N_7243,N_7797);
xor U14706 (N_14706,N_9794,N_9826);
or U14707 (N_14707,N_11070,N_10360);
nand U14708 (N_14708,N_8061,N_9692);
nand U14709 (N_14709,N_8164,N_11479);
nand U14710 (N_14710,N_7751,N_9297);
xnor U14711 (N_14711,N_7072,N_8834);
nor U14712 (N_14712,N_7350,N_6937);
nand U14713 (N_14713,N_9106,N_6310);
nand U14714 (N_14714,N_10565,N_8694);
nor U14715 (N_14715,N_9158,N_8496);
or U14716 (N_14716,N_10138,N_7814);
or U14717 (N_14717,N_8468,N_10495);
xnor U14718 (N_14718,N_9421,N_8987);
and U14719 (N_14719,N_8306,N_7834);
and U14720 (N_14720,N_7219,N_11095);
nand U14721 (N_14721,N_10780,N_10747);
and U14722 (N_14722,N_7566,N_11633);
nor U14723 (N_14723,N_10340,N_6610);
nand U14724 (N_14724,N_7863,N_6064);
nor U14725 (N_14725,N_6280,N_7943);
xnor U14726 (N_14726,N_6932,N_11673);
nand U14727 (N_14727,N_9571,N_11801);
nand U14728 (N_14728,N_9193,N_7573);
nor U14729 (N_14729,N_8585,N_11129);
xor U14730 (N_14730,N_11143,N_8811);
nor U14731 (N_14731,N_10616,N_10188);
nor U14732 (N_14732,N_11112,N_6608);
or U14733 (N_14733,N_11241,N_11312);
nor U14734 (N_14734,N_7427,N_7148);
nand U14735 (N_14735,N_11245,N_7787);
or U14736 (N_14736,N_9150,N_11626);
nor U14737 (N_14737,N_6718,N_10031);
or U14738 (N_14738,N_6586,N_11841);
and U14739 (N_14739,N_10457,N_10421);
and U14740 (N_14740,N_6196,N_6848);
nor U14741 (N_14741,N_7236,N_7518);
and U14742 (N_14742,N_6568,N_7296);
nor U14743 (N_14743,N_8342,N_9113);
or U14744 (N_14744,N_8259,N_7367);
nor U14745 (N_14745,N_6922,N_7116);
xnor U14746 (N_14746,N_6639,N_10405);
and U14747 (N_14747,N_11016,N_11390);
nor U14748 (N_14748,N_11270,N_8712);
and U14749 (N_14749,N_6507,N_7015);
and U14750 (N_14750,N_6683,N_6742);
nand U14751 (N_14751,N_8423,N_10902);
nand U14752 (N_14752,N_9537,N_8545);
nor U14753 (N_14753,N_11850,N_9089);
nor U14754 (N_14754,N_11822,N_6825);
or U14755 (N_14755,N_11054,N_9165);
nand U14756 (N_14756,N_9791,N_6071);
nor U14757 (N_14757,N_7735,N_9652);
xnor U14758 (N_14758,N_9820,N_10552);
or U14759 (N_14759,N_7635,N_8281);
xor U14760 (N_14760,N_9194,N_8517);
nor U14761 (N_14761,N_11030,N_11376);
or U14762 (N_14762,N_10203,N_9300);
xnor U14763 (N_14763,N_7163,N_6619);
xor U14764 (N_14764,N_7957,N_8689);
nor U14765 (N_14765,N_10907,N_7400);
nand U14766 (N_14766,N_8828,N_9466);
or U14767 (N_14767,N_7786,N_7698);
and U14768 (N_14768,N_11782,N_10712);
and U14769 (N_14769,N_7068,N_6884);
or U14770 (N_14770,N_11789,N_11606);
and U14771 (N_14771,N_8842,N_8444);
nand U14772 (N_14772,N_10839,N_10018);
nand U14773 (N_14773,N_8733,N_11806);
nor U14774 (N_14774,N_10665,N_9354);
nor U14775 (N_14775,N_11330,N_9464);
nand U14776 (N_14776,N_7613,N_7447);
xnor U14777 (N_14777,N_11598,N_8018);
nor U14778 (N_14778,N_8398,N_10465);
xor U14779 (N_14779,N_9183,N_10447);
xor U14780 (N_14780,N_8737,N_10684);
or U14781 (N_14781,N_9912,N_10888);
xor U14782 (N_14782,N_6175,N_8252);
nand U14783 (N_14783,N_7403,N_6800);
and U14784 (N_14784,N_11273,N_7765);
nor U14785 (N_14785,N_9998,N_9189);
nand U14786 (N_14786,N_9021,N_9801);
nand U14787 (N_14787,N_8195,N_8038);
nand U14788 (N_14788,N_9029,N_10572);
xor U14789 (N_14789,N_8632,N_7993);
nor U14790 (N_14790,N_10356,N_8141);
or U14791 (N_14791,N_7214,N_6015);
and U14792 (N_14792,N_8320,N_9479);
xor U14793 (N_14793,N_6085,N_9216);
xor U14794 (N_14794,N_11058,N_10288);
nor U14795 (N_14795,N_10720,N_8269);
and U14796 (N_14796,N_11408,N_8876);
nor U14797 (N_14797,N_7690,N_11647);
nor U14798 (N_14798,N_9008,N_11036);
and U14799 (N_14799,N_11618,N_8784);
xor U14800 (N_14800,N_9101,N_11504);
and U14801 (N_14801,N_8613,N_11372);
nand U14802 (N_14802,N_9434,N_8068);
nor U14803 (N_14803,N_10131,N_7672);
or U14804 (N_14804,N_10240,N_9174);
xor U14805 (N_14805,N_6859,N_11274);
and U14806 (N_14806,N_11418,N_9322);
nor U14807 (N_14807,N_9343,N_7248);
and U14808 (N_14808,N_11470,N_8457);
nor U14809 (N_14809,N_7639,N_7830);
xor U14810 (N_14810,N_9625,N_9388);
xnor U14811 (N_14811,N_8349,N_8085);
or U14812 (N_14812,N_10721,N_6982);
nor U14813 (N_14813,N_7580,N_9226);
and U14814 (N_14814,N_6878,N_8007);
or U14815 (N_14815,N_6459,N_9935);
nor U14816 (N_14816,N_11909,N_10135);
or U14817 (N_14817,N_10700,N_11082);
or U14818 (N_14818,N_11217,N_8505);
nor U14819 (N_14819,N_7921,N_9679);
and U14820 (N_14820,N_8365,N_8723);
nand U14821 (N_14821,N_9512,N_10762);
xnor U14822 (N_14822,N_6950,N_11374);
nor U14823 (N_14823,N_8478,N_11183);
nand U14824 (N_14824,N_7623,N_8539);
nand U14825 (N_14825,N_11639,N_7271);
and U14826 (N_14826,N_7191,N_9155);
nand U14827 (N_14827,N_8608,N_10914);
xnor U14828 (N_14828,N_8393,N_7213);
xor U14829 (N_14829,N_6314,N_7923);
or U14830 (N_14830,N_7558,N_10045);
and U14831 (N_14831,N_7741,N_8810);
nor U14832 (N_14832,N_10679,N_9561);
nand U14833 (N_14833,N_7356,N_8181);
nand U14834 (N_14834,N_8432,N_8997);
and U14835 (N_14835,N_8265,N_8805);
nor U14836 (N_14836,N_8914,N_11305);
nand U14837 (N_14837,N_10383,N_9982);
xnor U14838 (N_14838,N_9451,N_9784);
and U14839 (N_14839,N_7501,N_11123);
nand U14840 (N_14840,N_8543,N_10016);
or U14841 (N_14841,N_9762,N_6667);
nand U14842 (N_14842,N_10763,N_11276);
or U14843 (N_14843,N_8574,N_7728);
xnor U14844 (N_14844,N_8125,N_7262);
nand U14845 (N_14845,N_8652,N_10170);
xnor U14846 (N_14846,N_11226,N_7852);
nor U14847 (N_14847,N_10407,N_11698);
nand U14848 (N_14848,N_10361,N_11403);
nor U14849 (N_14849,N_11378,N_7119);
nor U14850 (N_14850,N_7339,N_10314);
nor U14851 (N_14851,N_10517,N_11997);
nand U14852 (N_14852,N_9582,N_6179);
xnor U14853 (N_14853,N_11055,N_9839);
or U14854 (N_14854,N_9028,N_6662);
xnor U14855 (N_14855,N_10948,N_10821);
xnor U14856 (N_14856,N_7035,N_6267);
nor U14857 (N_14857,N_11089,N_9071);
nor U14858 (N_14858,N_11923,N_7642);
nor U14859 (N_14859,N_11880,N_9064);
and U14860 (N_14860,N_7142,N_9298);
xnor U14861 (N_14861,N_8958,N_8527);
nor U14862 (N_14862,N_8319,N_6413);
nand U14863 (N_14863,N_6854,N_6252);
nor U14864 (N_14864,N_10512,N_8133);
or U14865 (N_14865,N_11988,N_6778);
and U14866 (N_14866,N_8915,N_8218);
or U14867 (N_14867,N_10624,N_8424);
nor U14868 (N_14868,N_9892,N_7811);
nand U14869 (N_14869,N_11960,N_6829);
nand U14870 (N_14870,N_10929,N_7216);
or U14871 (N_14871,N_10171,N_7156);
nor U14872 (N_14872,N_10833,N_7710);
or U14873 (N_14873,N_9994,N_7465);
nand U14874 (N_14874,N_10966,N_9946);
nor U14875 (N_14875,N_7662,N_8865);
nor U14876 (N_14876,N_7688,N_10388);
or U14877 (N_14877,N_8228,N_11657);
or U14878 (N_14878,N_7353,N_9897);
nor U14879 (N_14879,N_6238,N_6216);
nor U14880 (N_14880,N_9246,N_11370);
and U14881 (N_14881,N_6727,N_8037);
or U14882 (N_14882,N_11778,N_11087);
xnor U14883 (N_14883,N_10483,N_9012);
and U14884 (N_14884,N_6867,N_8276);
or U14885 (N_14885,N_6033,N_7105);
nand U14886 (N_14886,N_10927,N_8285);
or U14887 (N_14887,N_8573,N_9452);
nand U14888 (N_14888,N_9074,N_8189);
nor U14889 (N_14889,N_9969,N_7651);
nand U14890 (N_14890,N_7062,N_6694);
nor U14891 (N_14891,N_7510,N_10949);
nor U14892 (N_14892,N_8911,N_7395);
and U14893 (N_14893,N_6472,N_10108);
and U14894 (N_14894,N_11735,N_11819);
and U14895 (N_14895,N_11746,N_9913);
nor U14896 (N_14896,N_9970,N_9942);
and U14897 (N_14897,N_9110,N_9788);
and U14898 (N_14898,N_8462,N_8853);
and U14899 (N_14899,N_8905,N_6068);
nor U14900 (N_14900,N_11635,N_6635);
or U14901 (N_14901,N_8856,N_7753);
or U14902 (N_14902,N_6161,N_9523);
and U14903 (N_14903,N_10201,N_7980);
xor U14904 (N_14904,N_8677,N_9944);
nor U14905 (N_14905,N_8548,N_6062);
or U14906 (N_14906,N_8988,N_9020);
nor U14907 (N_14907,N_11803,N_10468);
and U14908 (N_14908,N_7461,N_10034);
nor U14909 (N_14909,N_11722,N_8454);
and U14910 (N_14910,N_9805,N_8612);
nand U14911 (N_14911,N_8666,N_7843);
nand U14912 (N_14912,N_9248,N_8337);
or U14913 (N_14913,N_6911,N_6747);
nor U14914 (N_14914,N_11456,N_10344);
nand U14915 (N_14915,N_10053,N_6750);
and U14916 (N_14916,N_9429,N_9005);
and U14917 (N_14917,N_7897,N_8767);
and U14918 (N_14918,N_9879,N_8882);
or U14919 (N_14919,N_9830,N_6327);
nor U14920 (N_14920,N_10770,N_10295);
nand U14921 (N_14921,N_11460,N_8506);
or U14922 (N_14922,N_10704,N_10614);
and U14923 (N_14923,N_7473,N_8730);
nor U14924 (N_14924,N_10214,N_10656);
or U14925 (N_14925,N_7971,N_7166);
nor U14926 (N_14926,N_8946,N_11740);
xor U14927 (N_14927,N_11573,N_7234);
nor U14928 (N_14928,N_8941,N_11875);
xor U14929 (N_14929,N_6857,N_7614);
or U14930 (N_14930,N_8369,N_7775);
or U14931 (N_14931,N_7298,N_6813);
nor U14932 (N_14932,N_6412,N_8032);
or U14933 (N_14933,N_8589,N_7221);
nand U14934 (N_14934,N_8096,N_10244);
and U14935 (N_14935,N_9179,N_8112);
or U14936 (N_14936,N_9217,N_9876);
or U14937 (N_14937,N_9188,N_11451);
or U14938 (N_14938,N_9361,N_7669);
nand U14939 (N_14939,N_6774,N_7990);
and U14940 (N_14940,N_10139,N_11099);
or U14941 (N_14941,N_6384,N_10408);
nor U14942 (N_14942,N_9239,N_8412);
nor U14943 (N_14943,N_9023,N_11022);
or U14944 (N_14944,N_11423,N_7290);
or U14945 (N_14945,N_8621,N_6219);
xor U14946 (N_14946,N_6039,N_7732);
xor U14947 (N_14947,N_11915,N_10711);
or U14948 (N_14948,N_11811,N_6724);
nor U14949 (N_14949,N_7588,N_6274);
nand U14950 (N_14950,N_9327,N_11167);
xor U14951 (N_14951,N_11324,N_8953);
xor U14952 (N_14952,N_6418,N_11503);
or U14953 (N_14953,N_8060,N_9669);
nor U14954 (N_14954,N_8770,N_6804);
xor U14955 (N_14955,N_9605,N_10411);
nand U14956 (N_14956,N_6261,N_11328);
and U14957 (N_14957,N_8501,N_8575);
nor U14958 (N_14958,N_11229,N_7738);
or U14959 (N_14959,N_10216,N_10930);
nor U14960 (N_14960,N_6944,N_6147);
nand U14961 (N_14961,N_9524,N_10235);
or U14962 (N_14962,N_8431,N_10807);
xnor U14963 (N_14963,N_7585,N_6014);
nor U14964 (N_14964,N_7210,N_8201);
and U14965 (N_14965,N_7399,N_9480);
and U14966 (N_14966,N_7112,N_9501);
or U14967 (N_14967,N_7469,N_8397);
nand U14968 (N_14968,N_10172,N_6215);
nor U14969 (N_14969,N_11065,N_10917);
nand U14970 (N_14970,N_9926,N_7648);
and U14971 (N_14971,N_9572,N_9477);
nor U14972 (N_14972,N_8333,N_7928);
xnor U14973 (N_14973,N_9238,N_6556);
nor U14974 (N_14974,N_6605,N_6543);
xnor U14975 (N_14975,N_8993,N_9566);
nand U14976 (N_14976,N_6478,N_6822);
xor U14977 (N_14977,N_6444,N_7724);
nand U14978 (N_14978,N_10868,N_9863);
or U14979 (N_14979,N_6388,N_9061);
nor U14980 (N_14980,N_6879,N_9589);
and U14981 (N_14981,N_7780,N_11406);
or U14982 (N_14982,N_10453,N_11405);
xnor U14983 (N_14983,N_8299,N_9168);
nand U14984 (N_14984,N_11018,N_11279);
nand U14985 (N_14985,N_11531,N_8740);
or U14986 (N_14986,N_10088,N_10500);
nor U14987 (N_14987,N_6924,N_11610);
xnor U14988 (N_14988,N_11985,N_11317);
xor U14989 (N_14989,N_10442,N_9888);
xnor U14990 (N_14990,N_6537,N_10580);
nor U14991 (N_14991,N_10223,N_6004);
nand U14992 (N_14992,N_8715,N_8186);
nand U14993 (N_14993,N_11974,N_8177);
and U14994 (N_14994,N_10695,N_9245);
nor U14995 (N_14995,N_11434,N_6546);
nand U14996 (N_14996,N_8508,N_11175);
and U14997 (N_14997,N_7475,N_6786);
nand U14998 (N_14998,N_10540,N_10690);
nor U14999 (N_14999,N_8741,N_7169);
nand U15000 (N_15000,N_11873,N_8761);
nor U15001 (N_15001,N_8600,N_7556);
nor U15002 (N_15002,N_6705,N_11332);
and U15003 (N_15003,N_6156,N_8048);
nand U15004 (N_15004,N_11244,N_10579);
nor U15005 (N_15005,N_9228,N_8169);
nand U15006 (N_15006,N_9120,N_9055);
nand U15007 (N_15007,N_11560,N_7888);
or U15008 (N_15008,N_11236,N_6566);
and U15009 (N_15009,N_10885,N_11044);
xor U15010 (N_15010,N_10738,N_10627);
xor U15011 (N_15011,N_9114,N_11573);
nand U15012 (N_15012,N_7129,N_9992);
xnor U15013 (N_15013,N_6962,N_8927);
or U15014 (N_15014,N_6457,N_10649);
nor U15015 (N_15015,N_6749,N_7419);
nand U15016 (N_15016,N_8632,N_7664);
nor U15017 (N_15017,N_9944,N_11412);
or U15018 (N_15018,N_9574,N_7266);
and U15019 (N_15019,N_10841,N_7704);
nor U15020 (N_15020,N_6956,N_11002);
nand U15021 (N_15021,N_7129,N_11260);
and U15022 (N_15022,N_6439,N_10748);
nand U15023 (N_15023,N_9527,N_9909);
or U15024 (N_15024,N_6977,N_6618);
xor U15025 (N_15025,N_6001,N_9515);
xnor U15026 (N_15026,N_11509,N_10925);
and U15027 (N_15027,N_8255,N_9366);
nor U15028 (N_15028,N_10427,N_10958);
or U15029 (N_15029,N_9363,N_10706);
nor U15030 (N_15030,N_11919,N_10090);
nor U15031 (N_15031,N_6421,N_10180);
and U15032 (N_15032,N_10094,N_7304);
nand U15033 (N_15033,N_11122,N_6405);
nand U15034 (N_15034,N_7905,N_8052);
nand U15035 (N_15035,N_9368,N_7011);
nor U15036 (N_15036,N_9495,N_11301);
or U15037 (N_15037,N_10621,N_9636);
and U15038 (N_15038,N_7736,N_9084);
xor U15039 (N_15039,N_10969,N_11522);
or U15040 (N_15040,N_7806,N_8072);
nand U15041 (N_15041,N_8977,N_8701);
xor U15042 (N_15042,N_8283,N_10466);
nand U15043 (N_15043,N_11059,N_9369);
nand U15044 (N_15044,N_11606,N_7165);
nor U15045 (N_15045,N_8553,N_10505);
nor U15046 (N_15046,N_10167,N_6861);
nand U15047 (N_15047,N_10584,N_9065);
and U15048 (N_15048,N_8498,N_6599);
nor U15049 (N_15049,N_7964,N_9760);
nor U15050 (N_15050,N_11839,N_6537);
nand U15051 (N_15051,N_7510,N_10104);
nor U15052 (N_15052,N_7304,N_7189);
nand U15053 (N_15053,N_9876,N_9485);
nor U15054 (N_15054,N_11915,N_7805);
and U15055 (N_15055,N_10933,N_9130);
xnor U15056 (N_15056,N_10733,N_10440);
and U15057 (N_15057,N_9958,N_11392);
and U15058 (N_15058,N_9758,N_7530);
nor U15059 (N_15059,N_7956,N_7416);
nor U15060 (N_15060,N_9774,N_6537);
and U15061 (N_15061,N_11727,N_6820);
or U15062 (N_15062,N_10592,N_11908);
nand U15063 (N_15063,N_6720,N_10550);
nand U15064 (N_15064,N_9234,N_7861);
nand U15065 (N_15065,N_7581,N_9582);
nor U15066 (N_15066,N_8598,N_7481);
and U15067 (N_15067,N_10287,N_8896);
xor U15068 (N_15068,N_11959,N_8310);
nand U15069 (N_15069,N_7586,N_6420);
and U15070 (N_15070,N_11076,N_6304);
nor U15071 (N_15071,N_9847,N_10898);
xnor U15072 (N_15072,N_10635,N_11688);
nand U15073 (N_15073,N_7073,N_7546);
xnor U15074 (N_15074,N_10318,N_9925);
and U15075 (N_15075,N_11612,N_9152);
xnor U15076 (N_15076,N_10472,N_8721);
nor U15077 (N_15077,N_7841,N_11424);
nor U15078 (N_15078,N_11212,N_11448);
or U15079 (N_15079,N_11315,N_7410);
or U15080 (N_15080,N_9939,N_8165);
and U15081 (N_15081,N_7368,N_10960);
or U15082 (N_15082,N_11979,N_9140);
nor U15083 (N_15083,N_6267,N_8859);
and U15084 (N_15084,N_10874,N_6649);
or U15085 (N_15085,N_8248,N_10339);
or U15086 (N_15086,N_11412,N_7816);
or U15087 (N_15087,N_8126,N_8202);
nand U15088 (N_15088,N_7680,N_10823);
nor U15089 (N_15089,N_11978,N_10522);
or U15090 (N_15090,N_9511,N_11621);
and U15091 (N_15091,N_7182,N_9502);
xor U15092 (N_15092,N_10792,N_7078);
xnor U15093 (N_15093,N_9253,N_6895);
and U15094 (N_15094,N_6940,N_9230);
xor U15095 (N_15095,N_7964,N_8042);
or U15096 (N_15096,N_11258,N_6982);
nor U15097 (N_15097,N_8100,N_10182);
nor U15098 (N_15098,N_10781,N_8719);
nand U15099 (N_15099,N_9145,N_10694);
xor U15100 (N_15100,N_9006,N_6951);
nor U15101 (N_15101,N_10213,N_8464);
xor U15102 (N_15102,N_8366,N_11159);
nand U15103 (N_15103,N_9172,N_8198);
nand U15104 (N_15104,N_7051,N_7439);
nand U15105 (N_15105,N_7483,N_8705);
nand U15106 (N_15106,N_6078,N_7350);
nor U15107 (N_15107,N_6033,N_7193);
nor U15108 (N_15108,N_6024,N_8498);
and U15109 (N_15109,N_8465,N_9840);
xnor U15110 (N_15110,N_6833,N_8152);
xor U15111 (N_15111,N_10134,N_9964);
xnor U15112 (N_15112,N_8669,N_11498);
nand U15113 (N_15113,N_7770,N_9238);
nor U15114 (N_15114,N_7632,N_10483);
or U15115 (N_15115,N_10192,N_8857);
or U15116 (N_15116,N_8101,N_11110);
xnor U15117 (N_15117,N_10358,N_11424);
and U15118 (N_15118,N_7638,N_7403);
or U15119 (N_15119,N_7131,N_11744);
nand U15120 (N_15120,N_9425,N_11899);
xor U15121 (N_15121,N_9016,N_6014);
nor U15122 (N_15122,N_8330,N_7624);
nand U15123 (N_15123,N_9780,N_9745);
nor U15124 (N_15124,N_8489,N_7525);
and U15125 (N_15125,N_10471,N_7491);
nand U15126 (N_15126,N_7622,N_8881);
and U15127 (N_15127,N_11723,N_10964);
nand U15128 (N_15128,N_6155,N_8107);
or U15129 (N_15129,N_7006,N_10425);
xor U15130 (N_15130,N_9727,N_6503);
nand U15131 (N_15131,N_7624,N_7801);
or U15132 (N_15132,N_7160,N_7171);
nor U15133 (N_15133,N_7519,N_11337);
and U15134 (N_15134,N_9260,N_8501);
and U15135 (N_15135,N_11355,N_7785);
nand U15136 (N_15136,N_9839,N_9228);
nor U15137 (N_15137,N_11348,N_10921);
nor U15138 (N_15138,N_8945,N_8185);
xor U15139 (N_15139,N_10337,N_7359);
nand U15140 (N_15140,N_10522,N_10554);
nor U15141 (N_15141,N_6700,N_8504);
or U15142 (N_15142,N_9004,N_11948);
nand U15143 (N_15143,N_6434,N_7412);
nor U15144 (N_15144,N_11804,N_9972);
nand U15145 (N_15145,N_7494,N_7866);
nor U15146 (N_15146,N_6648,N_6347);
xor U15147 (N_15147,N_7509,N_11781);
and U15148 (N_15148,N_6009,N_6476);
nand U15149 (N_15149,N_11623,N_6461);
nand U15150 (N_15150,N_8116,N_11027);
and U15151 (N_15151,N_8654,N_8229);
or U15152 (N_15152,N_10912,N_9670);
xor U15153 (N_15153,N_10917,N_7948);
nor U15154 (N_15154,N_7488,N_9057);
or U15155 (N_15155,N_8726,N_8379);
and U15156 (N_15156,N_10366,N_11288);
nor U15157 (N_15157,N_10612,N_6613);
nand U15158 (N_15158,N_7863,N_7816);
nand U15159 (N_15159,N_7447,N_8916);
or U15160 (N_15160,N_7218,N_9491);
or U15161 (N_15161,N_8181,N_9223);
nor U15162 (N_15162,N_7787,N_6264);
xor U15163 (N_15163,N_11785,N_9170);
or U15164 (N_15164,N_11571,N_10248);
and U15165 (N_15165,N_10549,N_10602);
nor U15166 (N_15166,N_11369,N_8269);
nor U15167 (N_15167,N_10623,N_10535);
or U15168 (N_15168,N_10086,N_7484);
and U15169 (N_15169,N_10195,N_6017);
and U15170 (N_15170,N_10308,N_6638);
nor U15171 (N_15171,N_8789,N_7689);
nand U15172 (N_15172,N_9701,N_9128);
xnor U15173 (N_15173,N_9318,N_11150);
nor U15174 (N_15174,N_6304,N_6190);
or U15175 (N_15175,N_8077,N_11768);
xnor U15176 (N_15176,N_10138,N_11875);
nor U15177 (N_15177,N_10675,N_10568);
nand U15178 (N_15178,N_7869,N_6060);
and U15179 (N_15179,N_8191,N_6425);
nand U15180 (N_15180,N_6796,N_9804);
nor U15181 (N_15181,N_10849,N_8016);
nand U15182 (N_15182,N_9291,N_6246);
or U15183 (N_15183,N_7221,N_11610);
and U15184 (N_15184,N_8262,N_6643);
nor U15185 (N_15185,N_8094,N_6358);
or U15186 (N_15186,N_11259,N_7619);
nand U15187 (N_15187,N_11340,N_9060);
and U15188 (N_15188,N_11375,N_9446);
and U15189 (N_15189,N_8233,N_6903);
xor U15190 (N_15190,N_9877,N_6830);
nand U15191 (N_15191,N_6175,N_11627);
or U15192 (N_15192,N_11812,N_9113);
xor U15193 (N_15193,N_7732,N_8975);
or U15194 (N_15194,N_10063,N_10457);
nor U15195 (N_15195,N_10978,N_6541);
nand U15196 (N_15196,N_6414,N_10872);
xnor U15197 (N_15197,N_10844,N_10975);
xnor U15198 (N_15198,N_10744,N_11041);
nand U15199 (N_15199,N_11021,N_6919);
nand U15200 (N_15200,N_7831,N_10773);
and U15201 (N_15201,N_6895,N_10784);
xor U15202 (N_15202,N_6421,N_8839);
or U15203 (N_15203,N_10233,N_10471);
nand U15204 (N_15204,N_10899,N_9857);
nand U15205 (N_15205,N_7954,N_9729);
nand U15206 (N_15206,N_9528,N_7068);
and U15207 (N_15207,N_8675,N_10421);
and U15208 (N_15208,N_6958,N_11971);
or U15209 (N_15209,N_7008,N_10850);
and U15210 (N_15210,N_10324,N_11900);
xnor U15211 (N_15211,N_6689,N_7403);
or U15212 (N_15212,N_10463,N_7971);
xnor U15213 (N_15213,N_8938,N_7784);
nand U15214 (N_15214,N_11590,N_6073);
nand U15215 (N_15215,N_7108,N_10452);
and U15216 (N_15216,N_9762,N_6140);
and U15217 (N_15217,N_10303,N_10443);
and U15218 (N_15218,N_11861,N_7684);
or U15219 (N_15219,N_11784,N_6345);
or U15220 (N_15220,N_6156,N_7051);
nand U15221 (N_15221,N_6658,N_9145);
nor U15222 (N_15222,N_7826,N_6598);
nor U15223 (N_15223,N_11615,N_7491);
nor U15224 (N_15224,N_11426,N_8393);
xor U15225 (N_15225,N_9233,N_9540);
nor U15226 (N_15226,N_10771,N_8473);
and U15227 (N_15227,N_7584,N_11793);
xor U15228 (N_15228,N_6370,N_8921);
nor U15229 (N_15229,N_8348,N_10399);
or U15230 (N_15230,N_8327,N_8718);
nor U15231 (N_15231,N_9243,N_7629);
xnor U15232 (N_15232,N_7528,N_8487);
and U15233 (N_15233,N_10415,N_10081);
xor U15234 (N_15234,N_6736,N_10251);
and U15235 (N_15235,N_6609,N_6475);
xnor U15236 (N_15236,N_8579,N_6264);
or U15237 (N_15237,N_8171,N_11241);
nor U15238 (N_15238,N_11116,N_11889);
nor U15239 (N_15239,N_9251,N_11212);
nor U15240 (N_15240,N_7673,N_10710);
nor U15241 (N_15241,N_8634,N_8182);
xnor U15242 (N_15242,N_7913,N_8900);
xor U15243 (N_15243,N_10282,N_9362);
and U15244 (N_15244,N_11059,N_10778);
nand U15245 (N_15245,N_6471,N_11434);
xor U15246 (N_15246,N_6028,N_7023);
nand U15247 (N_15247,N_7549,N_9632);
xnor U15248 (N_15248,N_11488,N_7939);
nand U15249 (N_15249,N_8404,N_7564);
and U15250 (N_15250,N_11801,N_7138);
and U15251 (N_15251,N_10573,N_9143);
nand U15252 (N_15252,N_11050,N_10250);
nand U15253 (N_15253,N_8797,N_8212);
nor U15254 (N_15254,N_7510,N_8466);
xnor U15255 (N_15255,N_7685,N_8138);
or U15256 (N_15256,N_8410,N_7092);
xor U15257 (N_15257,N_8286,N_7423);
nor U15258 (N_15258,N_9509,N_10305);
nand U15259 (N_15259,N_7775,N_11872);
or U15260 (N_15260,N_11223,N_7624);
or U15261 (N_15261,N_8622,N_6986);
and U15262 (N_15262,N_9044,N_9118);
nor U15263 (N_15263,N_6427,N_9312);
nor U15264 (N_15264,N_6480,N_9006);
and U15265 (N_15265,N_6616,N_6439);
and U15266 (N_15266,N_10065,N_7806);
and U15267 (N_15267,N_10524,N_11651);
xnor U15268 (N_15268,N_10517,N_9349);
xnor U15269 (N_15269,N_9054,N_7227);
xnor U15270 (N_15270,N_7701,N_9363);
nor U15271 (N_15271,N_6720,N_9581);
or U15272 (N_15272,N_8494,N_8997);
or U15273 (N_15273,N_11781,N_9332);
xor U15274 (N_15274,N_7119,N_10797);
and U15275 (N_15275,N_10553,N_6712);
or U15276 (N_15276,N_11254,N_11185);
nand U15277 (N_15277,N_10241,N_9053);
and U15278 (N_15278,N_9965,N_9790);
nand U15279 (N_15279,N_8886,N_8655);
nor U15280 (N_15280,N_9779,N_9342);
nor U15281 (N_15281,N_10927,N_8664);
or U15282 (N_15282,N_8119,N_9724);
and U15283 (N_15283,N_7406,N_8100);
nand U15284 (N_15284,N_6183,N_9543);
nand U15285 (N_15285,N_9041,N_9837);
or U15286 (N_15286,N_7290,N_8050);
and U15287 (N_15287,N_10029,N_11598);
nor U15288 (N_15288,N_7379,N_8085);
or U15289 (N_15289,N_11077,N_6028);
and U15290 (N_15290,N_6231,N_9758);
nor U15291 (N_15291,N_9577,N_6112);
nor U15292 (N_15292,N_7776,N_6885);
nor U15293 (N_15293,N_9993,N_10258);
and U15294 (N_15294,N_6965,N_9881);
nand U15295 (N_15295,N_6141,N_11734);
xnor U15296 (N_15296,N_7181,N_8007);
or U15297 (N_15297,N_10568,N_9044);
nand U15298 (N_15298,N_10277,N_9977);
xnor U15299 (N_15299,N_11944,N_8792);
nor U15300 (N_15300,N_6866,N_11904);
nor U15301 (N_15301,N_9477,N_9585);
xnor U15302 (N_15302,N_10598,N_10849);
nor U15303 (N_15303,N_10339,N_10299);
or U15304 (N_15304,N_11824,N_6642);
xor U15305 (N_15305,N_9349,N_8829);
nand U15306 (N_15306,N_10587,N_10865);
nor U15307 (N_15307,N_9117,N_11340);
and U15308 (N_15308,N_10777,N_10676);
or U15309 (N_15309,N_8890,N_7003);
xnor U15310 (N_15310,N_6273,N_10994);
xnor U15311 (N_15311,N_10767,N_7053);
or U15312 (N_15312,N_6777,N_10111);
xnor U15313 (N_15313,N_10219,N_7746);
nand U15314 (N_15314,N_10274,N_8098);
xnor U15315 (N_15315,N_10208,N_11782);
or U15316 (N_15316,N_7717,N_7167);
and U15317 (N_15317,N_7935,N_6574);
or U15318 (N_15318,N_11847,N_11285);
xnor U15319 (N_15319,N_11214,N_11141);
or U15320 (N_15320,N_11246,N_8943);
or U15321 (N_15321,N_10834,N_8009);
xnor U15322 (N_15322,N_7977,N_11060);
and U15323 (N_15323,N_9985,N_6381);
xnor U15324 (N_15324,N_9169,N_7577);
nand U15325 (N_15325,N_11360,N_11189);
xnor U15326 (N_15326,N_8925,N_11856);
xnor U15327 (N_15327,N_8078,N_10347);
xnor U15328 (N_15328,N_10722,N_7991);
or U15329 (N_15329,N_7347,N_11783);
nand U15330 (N_15330,N_9896,N_11554);
nor U15331 (N_15331,N_10603,N_8886);
and U15332 (N_15332,N_10384,N_8645);
or U15333 (N_15333,N_8801,N_6650);
and U15334 (N_15334,N_8359,N_11293);
nand U15335 (N_15335,N_9950,N_11310);
or U15336 (N_15336,N_6169,N_6072);
nand U15337 (N_15337,N_11389,N_11446);
nand U15338 (N_15338,N_10995,N_9299);
or U15339 (N_15339,N_8624,N_11167);
or U15340 (N_15340,N_7628,N_8746);
or U15341 (N_15341,N_6873,N_10311);
and U15342 (N_15342,N_8878,N_7749);
or U15343 (N_15343,N_6786,N_7304);
xnor U15344 (N_15344,N_10394,N_7829);
or U15345 (N_15345,N_8219,N_10636);
and U15346 (N_15346,N_7645,N_6726);
xnor U15347 (N_15347,N_7121,N_9494);
nor U15348 (N_15348,N_11961,N_6659);
xnor U15349 (N_15349,N_9711,N_10778);
nand U15350 (N_15350,N_8961,N_7502);
or U15351 (N_15351,N_9905,N_7816);
nor U15352 (N_15352,N_6103,N_7308);
nand U15353 (N_15353,N_8238,N_7359);
and U15354 (N_15354,N_9926,N_10737);
and U15355 (N_15355,N_6969,N_11133);
xor U15356 (N_15356,N_10241,N_7470);
and U15357 (N_15357,N_11080,N_8064);
nor U15358 (N_15358,N_6795,N_8767);
or U15359 (N_15359,N_6992,N_7642);
or U15360 (N_15360,N_9378,N_7655);
or U15361 (N_15361,N_6187,N_11783);
or U15362 (N_15362,N_6143,N_11957);
or U15363 (N_15363,N_9647,N_9561);
or U15364 (N_15364,N_9328,N_9225);
or U15365 (N_15365,N_10212,N_9555);
nor U15366 (N_15366,N_6099,N_8814);
or U15367 (N_15367,N_7034,N_7301);
or U15368 (N_15368,N_7704,N_9881);
xor U15369 (N_15369,N_6200,N_10468);
nor U15370 (N_15370,N_8564,N_9309);
nand U15371 (N_15371,N_10473,N_11932);
nand U15372 (N_15372,N_11507,N_7384);
nor U15373 (N_15373,N_6433,N_10894);
xor U15374 (N_15374,N_10410,N_6473);
nor U15375 (N_15375,N_10381,N_11818);
nor U15376 (N_15376,N_10939,N_7809);
nand U15377 (N_15377,N_6512,N_6372);
or U15378 (N_15378,N_11600,N_11179);
xnor U15379 (N_15379,N_7609,N_7316);
and U15380 (N_15380,N_6802,N_7955);
and U15381 (N_15381,N_11210,N_7351);
and U15382 (N_15382,N_11627,N_6945);
or U15383 (N_15383,N_6913,N_8379);
or U15384 (N_15384,N_6155,N_10858);
nand U15385 (N_15385,N_6272,N_6978);
xor U15386 (N_15386,N_7125,N_11337);
nor U15387 (N_15387,N_10665,N_7887);
or U15388 (N_15388,N_10597,N_7692);
or U15389 (N_15389,N_11955,N_7137);
or U15390 (N_15390,N_9606,N_10108);
and U15391 (N_15391,N_11593,N_6566);
and U15392 (N_15392,N_11095,N_11550);
xor U15393 (N_15393,N_11597,N_7769);
xor U15394 (N_15394,N_11136,N_9517);
nand U15395 (N_15395,N_8280,N_9791);
nand U15396 (N_15396,N_9849,N_8653);
nand U15397 (N_15397,N_11424,N_7634);
nor U15398 (N_15398,N_10796,N_8909);
nor U15399 (N_15399,N_6639,N_8056);
xor U15400 (N_15400,N_10820,N_10133);
or U15401 (N_15401,N_6646,N_8356);
and U15402 (N_15402,N_6845,N_6626);
nor U15403 (N_15403,N_8251,N_6508);
or U15404 (N_15404,N_6945,N_6465);
nor U15405 (N_15405,N_6057,N_6398);
or U15406 (N_15406,N_9161,N_9468);
nand U15407 (N_15407,N_10634,N_11171);
and U15408 (N_15408,N_8255,N_9567);
or U15409 (N_15409,N_6866,N_9012);
xor U15410 (N_15410,N_8702,N_11225);
nand U15411 (N_15411,N_6399,N_8291);
xnor U15412 (N_15412,N_7767,N_9720);
and U15413 (N_15413,N_9093,N_6489);
nor U15414 (N_15414,N_10190,N_11849);
and U15415 (N_15415,N_9726,N_9989);
xnor U15416 (N_15416,N_10509,N_10655);
nand U15417 (N_15417,N_8589,N_11791);
xor U15418 (N_15418,N_8501,N_9843);
and U15419 (N_15419,N_7435,N_10979);
nor U15420 (N_15420,N_10662,N_11863);
and U15421 (N_15421,N_10398,N_7545);
or U15422 (N_15422,N_9201,N_8623);
or U15423 (N_15423,N_8428,N_8001);
xnor U15424 (N_15424,N_8266,N_8753);
or U15425 (N_15425,N_8388,N_9968);
or U15426 (N_15426,N_7644,N_10933);
or U15427 (N_15427,N_9027,N_9084);
and U15428 (N_15428,N_7613,N_6983);
nor U15429 (N_15429,N_11256,N_9529);
and U15430 (N_15430,N_11806,N_9230);
or U15431 (N_15431,N_6146,N_6848);
or U15432 (N_15432,N_10528,N_9030);
nand U15433 (N_15433,N_9873,N_10297);
and U15434 (N_15434,N_8022,N_11928);
nor U15435 (N_15435,N_10616,N_9555);
or U15436 (N_15436,N_11860,N_10670);
xnor U15437 (N_15437,N_7433,N_10416);
and U15438 (N_15438,N_7573,N_11597);
nand U15439 (N_15439,N_6433,N_11761);
and U15440 (N_15440,N_6139,N_6082);
nor U15441 (N_15441,N_8040,N_6654);
xor U15442 (N_15442,N_8933,N_9910);
xnor U15443 (N_15443,N_7161,N_7113);
and U15444 (N_15444,N_8177,N_11999);
nor U15445 (N_15445,N_7036,N_10620);
nor U15446 (N_15446,N_8921,N_11410);
and U15447 (N_15447,N_7952,N_9318);
and U15448 (N_15448,N_8378,N_6263);
nand U15449 (N_15449,N_7793,N_7015);
or U15450 (N_15450,N_9883,N_10307);
nand U15451 (N_15451,N_6089,N_11718);
nand U15452 (N_15452,N_10508,N_7521);
or U15453 (N_15453,N_11833,N_8962);
xor U15454 (N_15454,N_6154,N_11963);
and U15455 (N_15455,N_8725,N_7401);
nand U15456 (N_15456,N_9676,N_10568);
or U15457 (N_15457,N_11858,N_9360);
and U15458 (N_15458,N_10250,N_10304);
xnor U15459 (N_15459,N_7237,N_10270);
or U15460 (N_15460,N_9701,N_6320);
xnor U15461 (N_15461,N_9263,N_6402);
or U15462 (N_15462,N_11247,N_11245);
nand U15463 (N_15463,N_9811,N_9974);
xor U15464 (N_15464,N_10814,N_8666);
and U15465 (N_15465,N_11000,N_9287);
and U15466 (N_15466,N_9187,N_9895);
nand U15467 (N_15467,N_6988,N_8074);
nor U15468 (N_15468,N_7329,N_6272);
nand U15469 (N_15469,N_8605,N_8122);
and U15470 (N_15470,N_11652,N_6454);
xor U15471 (N_15471,N_6730,N_10797);
xor U15472 (N_15472,N_7502,N_6510);
xnor U15473 (N_15473,N_9976,N_7951);
nand U15474 (N_15474,N_11364,N_8067);
nand U15475 (N_15475,N_11169,N_9540);
and U15476 (N_15476,N_7200,N_11020);
xor U15477 (N_15477,N_11956,N_6097);
nand U15478 (N_15478,N_8615,N_7754);
nand U15479 (N_15479,N_10511,N_9498);
nor U15480 (N_15480,N_7023,N_8475);
xnor U15481 (N_15481,N_7836,N_10912);
nand U15482 (N_15482,N_11316,N_9564);
or U15483 (N_15483,N_11241,N_11663);
nand U15484 (N_15484,N_8229,N_6153);
nor U15485 (N_15485,N_8873,N_7684);
xnor U15486 (N_15486,N_11011,N_10777);
or U15487 (N_15487,N_11108,N_8418);
nand U15488 (N_15488,N_7487,N_8858);
nor U15489 (N_15489,N_8325,N_10920);
nor U15490 (N_15490,N_6203,N_7772);
xnor U15491 (N_15491,N_11470,N_10245);
or U15492 (N_15492,N_9225,N_8420);
nand U15493 (N_15493,N_6415,N_9346);
xnor U15494 (N_15494,N_10707,N_10294);
or U15495 (N_15495,N_7069,N_10655);
and U15496 (N_15496,N_11205,N_9563);
or U15497 (N_15497,N_6329,N_10569);
or U15498 (N_15498,N_6089,N_9539);
or U15499 (N_15499,N_9449,N_11470);
nor U15500 (N_15500,N_8741,N_8195);
or U15501 (N_15501,N_8560,N_9202);
or U15502 (N_15502,N_7413,N_6003);
or U15503 (N_15503,N_7044,N_10349);
or U15504 (N_15504,N_7432,N_8997);
and U15505 (N_15505,N_9356,N_8320);
or U15506 (N_15506,N_9561,N_9628);
and U15507 (N_15507,N_11901,N_8485);
and U15508 (N_15508,N_9828,N_9444);
xnor U15509 (N_15509,N_10571,N_6673);
and U15510 (N_15510,N_7883,N_10625);
nor U15511 (N_15511,N_8971,N_11784);
or U15512 (N_15512,N_10905,N_6147);
or U15513 (N_15513,N_8167,N_10523);
nor U15514 (N_15514,N_8719,N_6738);
xor U15515 (N_15515,N_9799,N_8633);
xnor U15516 (N_15516,N_8324,N_9415);
nand U15517 (N_15517,N_11784,N_8862);
and U15518 (N_15518,N_6826,N_8169);
xor U15519 (N_15519,N_10726,N_8865);
nand U15520 (N_15520,N_6201,N_11225);
xor U15521 (N_15521,N_9613,N_10395);
or U15522 (N_15522,N_10209,N_7962);
nor U15523 (N_15523,N_6485,N_11908);
or U15524 (N_15524,N_10340,N_8413);
or U15525 (N_15525,N_9099,N_11088);
and U15526 (N_15526,N_10100,N_7775);
xnor U15527 (N_15527,N_6093,N_8263);
or U15528 (N_15528,N_11979,N_8573);
and U15529 (N_15529,N_8503,N_10050);
nor U15530 (N_15530,N_8853,N_10947);
xnor U15531 (N_15531,N_6482,N_6820);
xor U15532 (N_15532,N_6932,N_11744);
nor U15533 (N_15533,N_7611,N_7220);
and U15534 (N_15534,N_9724,N_9815);
or U15535 (N_15535,N_8908,N_10279);
xor U15536 (N_15536,N_6848,N_9916);
xnor U15537 (N_15537,N_6796,N_7847);
nand U15538 (N_15538,N_8841,N_9054);
or U15539 (N_15539,N_9565,N_7149);
and U15540 (N_15540,N_10735,N_8688);
nor U15541 (N_15541,N_9176,N_10109);
and U15542 (N_15542,N_11470,N_8772);
xor U15543 (N_15543,N_10267,N_9721);
or U15544 (N_15544,N_8619,N_10677);
xor U15545 (N_15545,N_7088,N_9337);
nand U15546 (N_15546,N_7731,N_7600);
or U15547 (N_15547,N_7759,N_8556);
nand U15548 (N_15548,N_8093,N_6071);
and U15549 (N_15549,N_10540,N_11088);
nand U15550 (N_15550,N_11578,N_6947);
nand U15551 (N_15551,N_7054,N_7015);
nand U15552 (N_15552,N_6616,N_10951);
nand U15553 (N_15553,N_8461,N_7377);
nand U15554 (N_15554,N_11543,N_10039);
nand U15555 (N_15555,N_9790,N_6612);
or U15556 (N_15556,N_11889,N_6616);
nor U15557 (N_15557,N_7588,N_9276);
nor U15558 (N_15558,N_8819,N_10358);
nand U15559 (N_15559,N_10650,N_9158);
or U15560 (N_15560,N_11791,N_7456);
xor U15561 (N_15561,N_9015,N_11420);
nor U15562 (N_15562,N_11566,N_9562);
and U15563 (N_15563,N_9768,N_6404);
nand U15564 (N_15564,N_10156,N_10898);
or U15565 (N_15565,N_8592,N_9045);
and U15566 (N_15566,N_8422,N_9834);
xor U15567 (N_15567,N_6196,N_10025);
or U15568 (N_15568,N_6486,N_10767);
xor U15569 (N_15569,N_7010,N_11824);
and U15570 (N_15570,N_7687,N_11766);
or U15571 (N_15571,N_6856,N_8780);
nor U15572 (N_15572,N_10204,N_11659);
or U15573 (N_15573,N_10615,N_11245);
xor U15574 (N_15574,N_6394,N_10303);
xnor U15575 (N_15575,N_9079,N_7297);
nand U15576 (N_15576,N_11851,N_11057);
nand U15577 (N_15577,N_7310,N_10010);
and U15578 (N_15578,N_8730,N_11983);
nor U15579 (N_15579,N_7125,N_7141);
and U15580 (N_15580,N_8836,N_6451);
nand U15581 (N_15581,N_6381,N_9244);
nand U15582 (N_15582,N_10396,N_7569);
nor U15583 (N_15583,N_6789,N_11510);
nor U15584 (N_15584,N_7111,N_7927);
or U15585 (N_15585,N_11133,N_7215);
nor U15586 (N_15586,N_10184,N_7099);
and U15587 (N_15587,N_8938,N_7755);
and U15588 (N_15588,N_7748,N_10962);
xor U15589 (N_15589,N_9708,N_10021);
nand U15590 (N_15590,N_9012,N_10077);
nand U15591 (N_15591,N_9757,N_8157);
and U15592 (N_15592,N_8932,N_6334);
xor U15593 (N_15593,N_11357,N_9543);
or U15594 (N_15594,N_6338,N_9672);
and U15595 (N_15595,N_11474,N_6406);
and U15596 (N_15596,N_10142,N_6828);
or U15597 (N_15597,N_11499,N_8975);
or U15598 (N_15598,N_6376,N_9964);
or U15599 (N_15599,N_9999,N_10467);
and U15600 (N_15600,N_8867,N_6058);
nor U15601 (N_15601,N_11110,N_9114);
and U15602 (N_15602,N_9589,N_9216);
or U15603 (N_15603,N_9109,N_10919);
nand U15604 (N_15604,N_9952,N_6070);
nand U15605 (N_15605,N_8500,N_6749);
xor U15606 (N_15606,N_11393,N_7108);
and U15607 (N_15607,N_8414,N_6211);
nand U15608 (N_15608,N_8575,N_9545);
or U15609 (N_15609,N_9079,N_8657);
nor U15610 (N_15610,N_8911,N_10205);
xnor U15611 (N_15611,N_11536,N_10461);
xor U15612 (N_15612,N_10084,N_10999);
xor U15613 (N_15613,N_11404,N_11337);
xnor U15614 (N_15614,N_9796,N_10106);
or U15615 (N_15615,N_11187,N_9130);
nor U15616 (N_15616,N_11335,N_11355);
nand U15617 (N_15617,N_9671,N_11952);
nor U15618 (N_15618,N_7189,N_8560);
xnor U15619 (N_15619,N_6211,N_11293);
nor U15620 (N_15620,N_8521,N_6454);
or U15621 (N_15621,N_10243,N_11206);
and U15622 (N_15622,N_9722,N_7349);
and U15623 (N_15623,N_8751,N_7685);
and U15624 (N_15624,N_9638,N_10931);
xnor U15625 (N_15625,N_7508,N_6125);
and U15626 (N_15626,N_7981,N_9314);
nand U15627 (N_15627,N_9519,N_8589);
xor U15628 (N_15628,N_10766,N_9633);
nand U15629 (N_15629,N_8389,N_8873);
nor U15630 (N_15630,N_11978,N_8438);
xnor U15631 (N_15631,N_11617,N_11701);
and U15632 (N_15632,N_7177,N_11523);
nor U15633 (N_15633,N_11856,N_11403);
and U15634 (N_15634,N_6120,N_8356);
and U15635 (N_15635,N_8617,N_8930);
nor U15636 (N_15636,N_9851,N_11710);
or U15637 (N_15637,N_11129,N_11136);
xor U15638 (N_15638,N_9590,N_7707);
xnor U15639 (N_15639,N_6892,N_11286);
xor U15640 (N_15640,N_9963,N_6830);
or U15641 (N_15641,N_6815,N_7791);
nand U15642 (N_15642,N_6237,N_8065);
and U15643 (N_15643,N_7722,N_11973);
nand U15644 (N_15644,N_8774,N_6024);
or U15645 (N_15645,N_8655,N_9328);
or U15646 (N_15646,N_7765,N_11285);
nand U15647 (N_15647,N_6111,N_11703);
or U15648 (N_15648,N_6317,N_10220);
nor U15649 (N_15649,N_10860,N_10002);
xor U15650 (N_15650,N_11828,N_10297);
nor U15651 (N_15651,N_6773,N_9108);
and U15652 (N_15652,N_6465,N_6677);
nand U15653 (N_15653,N_9485,N_6675);
xor U15654 (N_15654,N_6314,N_11422);
and U15655 (N_15655,N_10628,N_7347);
nand U15656 (N_15656,N_9350,N_9860);
xor U15657 (N_15657,N_9796,N_10587);
and U15658 (N_15658,N_6418,N_7447);
or U15659 (N_15659,N_10239,N_6342);
nor U15660 (N_15660,N_10670,N_9026);
nand U15661 (N_15661,N_9657,N_6319);
xnor U15662 (N_15662,N_6214,N_6853);
nand U15663 (N_15663,N_10487,N_10817);
nor U15664 (N_15664,N_11393,N_11874);
and U15665 (N_15665,N_11078,N_7176);
or U15666 (N_15666,N_11081,N_11228);
and U15667 (N_15667,N_9925,N_7413);
or U15668 (N_15668,N_10005,N_11494);
xnor U15669 (N_15669,N_8441,N_8385);
nor U15670 (N_15670,N_7662,N_11331);
nand U15671 (N_15671,N_10299,N_6011);
nor U15672 (N_15672,N_10958,N_8315);
xor U15673 (N_15673,N_8848,N_10290);
and U15674 (N_15674,N_11197,N_7337);
nor U15675 (N_15675,N_9693,N_10693);
nor U15676 (N_15676,N_10360,N_11941);
and U15677 (N_15677,N_10882,N_9525);
and U15678 (N_15678,N_10984,N_9602);
xnor U15679 (N_15679,N_6268,N_8467);
xnor U15680 (N_15680,N_11649,N_11329);
or U15681 (N_15681,N_6222,N_8789);
nand U15682 (N_15682,N_6836,N_11165);
or U15683 (N_15683,N_8292,N_9191);
and U15684 (N_15684,N_7903,N_9477);
xnor U15685 (N_15685,N_7726,N_10132);
nand U15686 (N_15686,N_9172,N_11272);
or U15687 (N_15687,N_7280,N_10940);
nand U15688 (N_15688,N_10223,N_6207);
or U15689 (N_15689,N_7403,N_8757);
nor U15690 (N_15690,N_9221,N_8752);
nor U15691 (N_15691,N_9491,N_8603);
and U15692 (N_15692,N_9427,N_9359);
nand U15693 (N_15693,N_10195,N_8947);
xor U15694 (N_15694,N_8666,N_6732);
xor U15695 (N_15695,N_9257,N_11394);
nor U15696 (N_15696,N_6471,N_9349);
nor U15697 (N_15697,N_9053,N_11852);
and U15698 (N_15698,N_9521,N_9258);
and U15699 (N_15699,N_6688,N_6493);
or U15700 (N_15700,N_11113,N_7796);
and U15701 (N_15701,N_7995,N_9362);
and U15702 (N_15702,N_7134,N_11581);
nand U15703 (N_15703,N_9152,N_9542);
or U15704 (N_15704,N_9881,N_6262);
nand U15705 (N_15705,N_6429,N_11469);
nand U15706 (N_15706,N_8089,N_7966);
and U15707 (N_15707,N_9991,N_6711);
nand U15708 (N_15708,N_10766,N_10920);
nor U15709 (N_15709,N_9485,N_8710);
nand U15710 (N_15710,N_6641,N_9980);
nor U15711 (N_15711,N_8352,N_6338);
xnor U15712 (N_15712,N_11526,N_8476);
and U15713 (N_15713,N_9406,N_11136);
nand U15714 (N_15714,N_6733,N_10033);
or U15715 (N_15715,N_7989,N_8117);
nand U15716 (N_15716,N_10167,N_6399);
xor U15717 (N_15717,N_8403,N_7412);
nand U15718 (N_15718,N_9088,N_9063);
and U15719 (N_15719,N_8864,N_7443);
xor U15720 (N_15720,N_7726,N_8479);
or U15721 (N_15721,N_9686,N_10713);
xnor U15722 (N_15722,N_9218,N_7847);
and U15723 (N_15723,N_10595,N_11341);
and U15724 (N_15724,N_11920,N_8013);
or U15725 (N_15725,N_8075,N_9315);
nor U15726 (N_15726,N_9412,N_6238);
nand U15727 (N_15727,N_8507,N_10525);
nand U15728 (N_15728,N_9108,N_6709);
or U15729 (N_15729,N_7994,N_6682);
xor U15730 (N_15730,N_10881,N_7815);
xnor U15731 (N_15731,N_8822,N_9890);
or U15732 (N_15732,N_7191,N_6091);
xnor U15733 (N_15733,N_9181,N_6939);
and U15734 (N_15734,N_9122,N_6547);
nor U15735 (N_15735,N_8971,N_8501);
and U15736 (N_15736,N_9683,N_11869);
nor U15737 (N_15737,N_6302,N_11699);
nor U15738 (N_15738,N_11220,N_9328);
and U15739 (N_15739,N_8087,N_10564);
nor U15740 (N_15740,N_11117,N_11368);
and U15741 (N_15741,N_11556,N_9991);
xor U15742 (N_15742,N_11075,N_11942);
xnor U15743 (N_15743,N_8721,N_9926);
or U15744 (N_15744,N_8393,N_6404);
and U15745 (N_15745,N_8398,N_11446);
xnor U15746 (N_15746,N_11105,N_8560);
nor U15747 (N_15747,N_11492,N_9148);
or U15748 (N_15748,N_11890,N_10044);
nor U15749 (N_15749,N_6988,N_10422);
xor U15750 (N_15750,N_9183,N_8057);
xnor U15751 (N_15751,N_6238,N_8225);
nand U15752 (N_15752,N_10207,N_8948);
xor U15753 (N_15753,N_10396,N_6316);
or U15754 (N_15754,N_6691,N_11709);
or U15755 (N_15755,N_6898,N_11266);
or U15756 (N_15756,N_11310,N_8305);
or U15757 (N_15757,N_8579,N_10421);
nor U15758 (N_15758,N_10291,N_6347);
and U15759 (N_15759,N_10477,N_10677);
nand U15760 (N_15760,N_8326,N_7120);
and U15761 (N_15761,N_8253,N_9918);
and U15762 (N_15762,N_9818,N_7670);
nor U15763 (N_15763,N_9050,N_9738);
and U15764 (N_15764,N_9666,N_9147);
xor U15765 (N_15765,N_10202,N_9296);
or U15766 (N_15766,N_6274,N_11896);
or U15767 (N_15767,N_6794,N_11375);
nor U15768 (N_15768,N_6417,N_10466);
or U15769 (N_15769,N_7117,N_6474);
or U15770 (N_15770,N_8167,N_10863);
nor U15771 (N_15771,N_11117,N_10194);
nor U15772 (N_15772,N_10327,N_6450);
and U15773 (N_15773,N_11390,N_8445);
or U15774 (N_15774,N_11032,N_7006);
xor U15775 (N_15775,N_10597,N_9098);
and U15776 (N_15776,N_7930,N_6000);
xor U15777 (N_15777,N_6346,N_11099);
xor U15778 (N_15778,N_7029,N_6359);
or U15779 (N_15779,N_6491,N_9543);
or U15780 (N_15780,N_8589,N_10163);
and U15781 (N_15781,N_11070,N_8036);
and U15782 (N_15782,N_10584,N_9202);
and U15783 (N_15783,N_6548,N_7331);
xnor U15784 (N_15784,N_11756,N_7134);
or U15785 (N_15785,N_9700,N_7563);
xnor U15786 (N_15786,N_9136,N_8721);
xor U15787 (N_15787,N_8020,N_7410);
xor U15788 (N_15788,N_9320,N_7359);
nor U15789 (N_15789,N_10404,N_6350);
and U15790 (N_15790,N_6840,N_9975);
xnor U15791 (N_15791,N_7569,N_6712);
and U15792 (N_15792,N_7226,N_8312);
xnor U15793 (N_15793,N_8000,N_9527);
nor U15794 (N_15794,N_8505,N_8284);
or U15795 (N_15795,N_7831,N_6150);
and U15796 (N_15796,N_11151,N_10725);
nor U15797 (N_15797,N_11060,N_9105);
or U15798 (N_15798,N_6543,N_9530);
xnor U15799 (N_15799,N_11748,N_7628);
nand U15800 (N_15800,N_11780,N_9887);
or U15801 (N_15801,N_10090,N_6752);
xnor U15802 (N_15802,N_8222,N_11060);
or U15803 (N_15803,N_6355,N_10536);
nand U15804 (N_15804,N_9730,N_6212);
xnor U15805 (N_15805,N_8499,N_9744);
and U15806 (N_15806,N_11930,N_7797);
nand U15807 (N_15807,N_10469,N_9324);
or U15808 (N_15808,N_7738,N_7049);
xor U15809 (N_15809,N_11879,N_7886);
xor U15810 (N_15810,N_9163,N_8582);
xor U15811 (N_15811,N_9133,N_10495);
and U15812 (N_15812,N_10994,N_7398);
or U15813 (N_15813,N_11542,N_9808);
or U15814 (N_15814,N_10979,N_6896);
nand U15815 (N_15815,N_8610,N_11903);
nor U15816 (N_15816,N_9287,N_8007);
nand U15817 (N_15817,N_6851,N_6066);
nor U15818 (N_15818,N_7000,N_10791);
or U15819 (N_15819,N_8370,N_10606);
and U15820 (N_15820,N_10878,N_7727);
and U15821 (N_15821,N_6265,N_11243);
nor U15822 (N_15822,N_9082,N_8164);
nand U15823 (N_15823,N_6232,N_7547);
nand U15824 (N_15824,N_7145,N_10396);
and U15825 (N_15825,N_9953,N_10616);
nand U15826 (N_15826,N_6720,N_6431);
xnor U15827 (N_15827,N_6524,N_11569);
xor U15828 (N_15828,N_7649,N_11428);
xnor U15829 (N_15829,N_9107,N_7373);
nor U15830 (N_15830,N_6082,N_7404);
xnor U15831 (N_15831,N_8724,N_11527);
nor U15832 (N_15832,N_11834,N_6345);
or U15833 (N_15833,N_8242,N_9737);
nand U15834 (N_15834,N_7785,N_9625);
nand U15835 (N_15835,N_10790,N_8505);
and U15836 (N_15836,N_7456,N_11129);
and U15837 (N_15837,N_7104,N_10924);
and U15838 (N_15838,N_9171,N_8153);
or U15839 (N_15839,N_7691,N_9478);
and U15840 (N_15840,N_9865,N_6775);
xnor U15841 (N_15841,N_6654,N_7433);
or U15842 (N_15842,N_8006,N_11630);
or U15843 (N_15843,N_10695,N_6609);
and U15844 (N_15844,N_11661,N_6965);
xnor U15845 (N_15845,N_9909,N_6064);
nand U15846 (N_15846,N_11026,N_11070);
nor U15847 (N_15847,N_7737,N_9564);
or U15848 (N_15848,N_6537,N_8976);
and U15849 (N_15849,N_8397,N_8783);
nand U15850 (N_15850,N_6105,N_6447);
nand U15851 (N_15851,N_9311,N_8612);
or U15852 (N_15852,N_11397,N_10592);
or U15853 (N_15853,N_10708,N_7197);
and U15854 (N_15854,N_7562,N_7374);
and U15855 (N_15855,N_8897,N_7293);
xnor U15856 (N_15856,N_10873,N_6262);
and U15857 (N_15857,N_7213,N_11343);
nand U15858 (N_15858,N_7879,N_10224);
and U15859 (N_15859,N_7550,N_6900);
xor U15860 (N_15860,N_9087,N_9038);
or U15861 (N_15861,N_7495,N_9930);
or U15862 (N_15862,N_7968,N_7313);
or U15863 (N_15863,N_8421,N_9775);
and U15864 (N_15864,N_7649,N_11274);
or U15865 (N_15865,N_8833,N_11569);
nor U15866 (N_15866,N_7440,N_7306);
xnor U15867 (N_15867,N_8340,N_9283);
nor U15868 (N_15868,N_10873,N_8892);
or U15869 (N_15869,N_8108,N_8041);
xnor U15870 (N_15870,N_11318,N_10720);
nor U15871 (N_15871,N_6149,N_6375);
or U15872 (N_15872,N_9565,N_10212);
or U15873 (N_15873,N_11544,N_6540);
or U15874 (N_15874,N_8469,N_8311);
or U15875 (N_15875,N_10212,N_11180);
and U15876 (N_15876,N_9271,N_8378);
and U15877 (N_15877,N_9707,N_9233);
nor U15878 (N_15878,N_7678,N_7110);
nor U15879 (N_15879,N_11013,N_9094);
or U15880 (N_15880,N_10576,N_8845);
nor U15881 (N_15881,N_9853,N_9546);
and U15882 (N_15882,N_7435,N_9657);
nand U15883 (N_15883,N_10455,N_11401);
nand U15884 (N_15884,N_10740,N_6672);
or U15885 (N_15885,N_10906,N_10834);
or U15886 (N_15886,N_7650,N_7783);
and U15887 (N_15887,N_6471,N_11631);
and U15888 (N_15888,N_9670,N_11622);
xnor U15889 (N_15889,N_11105,N_6173);
nor U15890 (N_15890,N_7636,N_11751);
nand U15891 (N_15891,N_8982,N_6532);
or U15892 (N_15892,N_8858,N_6907);
nor U15893 (N_15893,N_10822,N_9084);
nand U15894 (N_15894,N_7001,N_11641);
nand U15895 (N_15895,N_11214,N_6608);
or U15896 (N_15896,N_9523,N_11167);
xnor U15897 (N_15897,N_11166,N_7757);
nor U15898 (N_15898,N_9872,N_6357);
and U15899 (N_15899,N_6302,N_6316);
nand U15900 (N_15900,N_8811,N_9258);
or U15901 (N_15901,N_9347,N_10166);
and U15902 (N_15902,N_7149,N_10553);
or U15903 (N_15903,N_8451,N_7694);
nor U15904 (N_15904,N_8702,N_7123);
or U15905 (N_15905,N_11258,N_11598);
and U15906 (N_15906,N_7833,N_10068);
nand U15907 (N_15907,N_11056,N_6521);
and U15908 (N_15908,N_6740,N_11432);
nor U15909 (N_15909,N_10753,N_7749);
xor U15910 (N_15910,N_11244,N_9537);
nand U15911 (N_15911,N_10359,N_8241);
or U15912 (N_15912,N_11427,N_11138);
nor U15913 (N_15913,N_9543,N_10632);
nand U15914 (N_15914,N_7418,N_9751);
nand U15915 (N_15915,N_6037,N_7014);
or U15916 (N_15916,N_11432,N_9761);
or U15917 (N_15917,N_6806,N_9132);
nor U15918 (N_15918,N_11783,N_6734);
or U15919 (N_15919,N_9106,N_9027);
nand U15920 (N_15920,N_11791,N_6265);
and U15921 (N_15921,N_8667,N_9165);
and U15922 (N_15922,N_8509,N_8224);
xnor U15923 (N_15923,N_11646,N_7287);
xor U15924 (N_15924,N_8867,N_6519);
and U15925 (N_15925,N_11433,N_8445);
and U15926 (N_15926,N_11335,N_11855);
nor U15927 (N_15927,N_10329,N_7314);
nor U15928 (N_15928,N_6684,N_6662);
and U15929 (N_15929,N_8439,N_7008);
nor U15930 (N_15930,N_6165,N_11407);
xnor U15931 (N_15931,N_8286,N_7497);
nor U15932 (N_15932,N_9309,N_8692);
nand U15933 (N_15933,N_7155,N_11966);
nor U15934 (N_15934,N_11994,N_11933);
xnor U15935 (N_15935,N_11585,N_6481);
nand U15936 (N_15936,N_11951,N_11977);
nor U15937 (N_15937,N_11146,N_9143);
nand U15938 (N_15938,N_9570,N_7692);
and U15939 (N_15939,N_8649,N_9612);
and U15940 (N_15940,N_6155,N_8739);
and U15941 (N_15941,N_7612,N_11706);
nor U15942 (N_15942,N_10670,N_8042);
nor U15943 (N_15943,N_9721,N_10604);
xnor U15944 (N_15944,N_9778,N_9870);
nor U15945 (N_15945,N_10258,N_8433);
or U15946 (N_15946,N_6802,N_10839);
nand U15947 (N_15947,N_10034,N_11518);
or U15948 (N_15948,N_6635,N_9724);
nand U15949 (N_15949,N_7357,N_7729);
nand U15950 (N_15950,N_10853,N_8872);
nor U15951 (N_15951,N_7609,N_11788);
nand U15952 (N_15952,N_8372,N_6189);
and U15953 (N_15953,N_11943,N_10414);
nand U15954 (N_15954,N_6220,N_6469);
or U15955 (N_15955,N_6643,N_8887);
and U15956 (N_15956,N_11927,N_9493);
nor U15957 (N_15957,N_7327,N_7000);
nand U15958 (N_15958,N_10491,N_6077);
and U15959 (N_15959,N_6948,N_6084);
nand U15960 (N_15960,N_11003,N_6973);
nor U15961 (N_15961,N_7883,N_10276);
nand U15962 (N_15962,N_8676,N_8839);
xnor U15963 (N_15963,N_8435,N_11844);
xnor U15964 (N_15964,N_7439,N_11856);
nand U15965 (N_15965,N_9378,N_7149);
nand U15966 (N_15966,N_9856,N_8951);
and U15967 (N_15967,N_9333,N_10085);
xnor U15968 (N_15968,N_7304,N_7370);
nor U15969 (N_15969,N_11931,N_7502);
nand U15970 (N_15970,N_11003,N_9229);
and U15971 (N_15971,N_11465,N_6028);
or U15972 (N_15972,N_11186,N_9835);
nand U15973 (N_15973,N_8352,N_11413);
nand U15974 (N_15974,N_9707,N_11082);
nor U15975 (N_15975,N_9520,N_9542);
nand U15976 (N_15976,N_7455,N_7490);
xor U15977 (N_15977,N_6359,N_10635);
nand U15978 (N_15978,N_8200,N_9765);
xnor U15979 (N_15979,N_11942,N_10044);
and U15980 (N_15980,N_11400,N_6427);
and U15981 (N_15981,N_7879,N_9400);
nor U15982 (N_15982,N_9265,N_8700);
and U15983 (N_15983,N_6622,N_7041);
nand U15984 (N_15984,N_7158,N_6719);
or U15985 (N_15985,N_7578,N_9793);
or U15986 (N_15986,N_7904,N_11111);
xnor U15987 (N_15987,N_9979,N_9482);
xor U15988 (N_15988,N_6044,N_7691);
nand U15989 (N_15989,N_6902,N_8297);
xor U15990 (N_15990,N_11186,N_8997);
and U15991 (N_15991,N_9589,N_7669);
nand U15992 (N_15992,N_6410,N_11060);
or U15993 (N_15993,N_9610,N_7280);
or U15994 (N_15994,N_10060,N_7337);
nand U15995 (N_15995,N_6260,N_7421);
and U15996 (N_15996,N_8750,N_7086);
and U15997 (N_15997,N_9076,N_11709);
nand U15998 (N_15998,N_10987,N_10381);
nor U15999 (N_15999,N_9427,N_9680);
and U16000 (N_16000,N_8775,N_10527);
xnor U16001 (N_16001,N_6270,N_11580);
xor U16002 (N_16002,N_11813,N_9620);
xor U16003 (N_16003,N_6155,N_6781);
or U16004 (N_16004,N_11826,N_11383);
nor U16005 (N_16005,N_11320,N_10569);
nor U16006 (N_16006,N_11691,N_11365);
nand U16007 (N_16007,N_11797,N_6794);
or U16008 (N_16008,N_10678,N_6601);
xor U16009 (N_16009,N_9755,N_9959);
xnor U16010 (N_16010,N_11978,N_8099);
nand U16011 (N_16011,N_6902,N_6901);
or U16012 (N_16012,N_9283,N_8673);
nand U16013 (N_16013,N_10673,N_10771);
or U16014 (N_16014,N_8388,N_8609);
and U16015 (N_16015,N_7771,N_11732);
or U16016 (N_16016,N_6615,N_8588);
and U16017 (N_16017,N_11207,N_9802);
xnor U16018 (N_16018,N_9590,N_9195);
nor U16019 (N_16019,N_9401,N_8864);
nor U16020 (N_16020,N_10633,N_6822);
nand U16021 (N_16021,N_11662,N_7529);
xnor U16022 (N_16022,N_7621,N_11389);
nand U16023 (N_16023,N_9380,N_8557);
nand U16024 (N_16024,N_7559,N_9891);
or U16025 (N_16025,N_8431,N_6712);
nor U16026 (N_16026,N_8845,N_7886);
nor U16027 (N_16027,N_8855,N_7039);
and U16028 (N_16028,N_8023,N_11929);
or U16029 (N_16029,N_11937,N_8071);
xnor U16030 (N_16030,N_9821,N_9276);
nand U16031 (N_16031,N_11351,N_8736);
nand U16032 (N_16032,N_8419,N_7566);
nor U16033 (N_16033,N_9669,N_11859);
and U16034 (N_16034,N_7617,N_9263);
nand U16035 (N_16035,N_9379,N_9621);
and U16036 (N_16036,N_11116,N_11805);
nor U16037 (N_16037,N_8530,N_11793);
nand U16038 (N_16038,N_6662,N_8516);
xor U16039 (N_16039,N_7136,N_10355);
nor U16040 (N_16040,N_7098,N_9794);
nand U16041 (N_16041,N_11078,N_7192);
nand U16042 (N_16042,N_8650,N_10186);
and U16043 (N_16043,N_7181,N_10219);
nand U16044 (N_16044,N_8622,N_9009);
nor U16045 (N_16045,N_11409,N_11530);
nand U16046 (N_16046,N_10799,N_11473);
or U16047 (N_16047,N_10657,N_11884);
or U16048 (N_16048,N_7228,N_11802);
nand U16049 (N_16049,N_10927,N_8778);
and U16050 (N_16050,N_10075,N_7928);
xor U16051 (N_16051,N_11825,N_7899);
nand U16052 (N_16052,N_8602,N_6366);
nand U16053 (N_16053,N_7003,N_10594);
nor U16054 (N_16054,N_10739,N_7421);
and U16055 (N_16055,N_6262,N_6869);
xnor U16056 (N_16056,N_11551,N_8326);
xnor U16057 (N_16057,N_7094,N_8195);
xnor U16058 (N_16058,N_8978,N_9083);
and U16059 (N_16059,N_10004,N_11600);
nor U16060 (N_16060,N_7810,N_10161);
nor U16061 (N_16061,N_11179,N_6945);
or U16062 (N_16062,N_11107,N_6152);
xnor U16063 (N_16063,N_8213,N_8812);
and U16064 (N_16064,N_6873,N_7393);
xor U16065 (N_16065,N_10894,N_10586);
nand U16066 (N_16066,N_7477,N_7944);
or U16067 (N_16067,N_8375,N_6593);
and U16068 (N_16068,N_11115,N_8145);
nand U16069 (N_16069,N_7055,N_11285);
nand U16070 (N_16070,N_7651,N_11214);
or U16071 (N_16071,N_7330,N_7056);
nor U16072 (N_16072,N_7581,N_7886);
nand U16073 (N_16073,N_9942,N_6100);
nor U16074 (N_16074,N_8133,N_10779);
or U16075 (N_16075,N_7523,N_11894);
nand U16076 (N_16076,N_11540,N_8953);
nand U16077 (N_16077,N_10744,N_10537);
xnor U16078 (N_16078,N_8064,N_7028);
or U16079 (N_16079,N_10072,N_7190);
xor U16080 (N_16080,N_6383,N_7308);
or U16081 (N_16081,N_8134,N_6707);
and U16082 (N_16082,N_7091,N_8503);
xor U16083 (N_16083,N_7957,N_6041);
or U16084 (N_16084,N_10766,N_7847);
and U16085 (N_16085,N_10876,N_10944);
nand U16086 (N_16086,N_11630,N_10146);
and U16087 (N_16087,N_9051,N_10955);
nor U16088 (N_16088,N_11631,N_11392);
nand U16089 (N_16089,N_11100,N_8500);
xor U16090 (N_16090,N_6425,N_7356);
nand U16091 (N_16091,N_7602,N_11063);
nand U16092 (N_16092,N_9241,N_10875);
and U16093 (N_16093,N_8866,N_7169);
and U16094 (N_16094,N_8356,N_10008);
nand U16095 (N_16095,N_6935,N_9128);
or U16096 (N_16096,N_7561,N_7573);
nand U16097 (N_16097,N_7172,N_7910);
nor U16098 (N_16098,N_8257,N_6441);
and U16099 (N_16099,N_6626,N_9330);
xor U16100 (N_16100,N_9261,N_10594);
xnor U16101 (N_16101,N_8050,N_6188);
nand U16102 (N_16102,N_8579,N_7336);
and U16103 (N_16103,N_7675,N_7274);
and U16104 (N_16104,N_7760,N_9678);
xor U16105 (N_16105,N_8520,N_9477);
and U16106 (N_16106,N_9943,N_6730);
xnor U16107 (N_16107,N_6715,N_6538);
nand U16108 (N_16108,N_8173,N_10879);
or U16109 (N_16109,N_7415,N_9521);
and U16110 (N_16110,N_8601,N_9764);
nor U16111 (N_16111,N_8107,N_8901);
xnor U16112 (N_16112,N_6893,N_7331);
xor U16113 (N_16113,N_7370,N_7025);
or U16114 (N_16114,N_8808,N_6081);
or U16115 (N_16115,N_7650,N_6354);
or U16116 (N_16116,N_7051,N_6691);
nor U16117 (N_16117,N_10095,N_8395);
nand U16118 (N_16118,N_9042,N_10900);
or U16119 (N_16119,N_10383,N_10870);
nand U16120 (N_16120,N_7777,N_8591);
xnor U16121 (N_16121,N_8329,N_6886);
nand U16122 (N_16122,N_11054,N_8236);
or U16123 (N_16123,N_7896,N_10310);
nor U16124 (N_16124,N_8601,N_10073);
nand U16125 (N_16125,N_7987,N_10664);
or U16126 (N_16126,N_9731,N_11700);
and U16127 (N_16127,N_6896,N_10252);
nand U16128 (N_16128,N_8422,N_7224);
and U16129 (N_16129,N_7967,N_11719);
or U16130 (N_16130,N_8366,N_11824);
xor U16131 (N_16131,N_9939,N_9814);
and U16132 (N_16132,N_7939,N_6171);
and U16133 (N_16133,N_7633,N_7288);
nand U16134 (N_16134,N_10826,N_8795);
or U16135 (N_16135,N_11481,N_7876);
nand U16136 (N_16136,N_7240,N_10358);
or U16137 (N_16137,N_8844,N_8377);
and U16138 (N_16138,N_9695,N_8988);
nand U16139 (N_16139,N_7554,N_10373);
xor U16140 (N_16140,N_10665,N_10560);
nand U16141 (N_16141,N_10087,N_11036);
nand U16142 (N_16142,N_6532,N_10119);
nand U16143 (N_16143,N_10828,N_9163);
and U16144 (N_16144,N_9585,N_10383);
and U16145 (N_16145,N_6845,N_11202);
nand U16146 (N_16146,N_6882,N_10302);
or U16147 (N_16147,N_11809,N_8265);
and U16148 (N_16148,N_11416,N_8712);
and U16149 (N_16149,N_6815,N_11990);
xnor U16150 (N_16150,N_11617,N_11006);
xnor U16151 (N_16151,N_6130,N_6729);
nor U16152 (N_16152,N_11744,N_8042);
nor U16153 (N_16153,N_11616,N_11513);
nor U16154 (N_16154,N_6422,N_7928);
and U16155 (N_16155,N_8834,N_6760);
or U16156 (N_16156,N_11614,N_9958);
nor U16157 (N_16157,N_8778,N_6272);
nor U16158 (N_16158,N_6433,N_11827);
and U16159 (N_16159,N_11736,N_11333);
nor U16160 (N_16160,N_9728,N_10148);
nor U16161 (N_16161,N_8897,N_8909);
and U16162 (N_16162,N_11771,N_8594);
or U16163 (N_16163,N_6584,N_7053);
and U16164 (N_16164,N_7016,N_11779);
nand U16165 (N_16165,N_8749,N_10823);
and U16166 (N_16166,N_9133,N_9776);
nor U16167 (N_16167,N_8066,N_9263);
nor U16168 (N_16168,N_10766,N_9419);
or U16169 (N_16169,N_9674,N_7132);
xnor U16170 (N_16170,N_10396,N_7373);
or U16171 (N_16171,N_10460,N_10196);
xnor U16172 (N_16172,N_6744,N_6621);
xnor U16173 (N_16173,N_6052,N_6696);
or U16174 (N_16174,N_9369,N_10905);
or U16175 (N_16175,N_7937,N_8964);
xor U16176 (N_16176,N_9242,N_8263);
xnor U16177 (N_16177,N_9514,N_9606);
or U16178 (N_16178,N_7444,N_10988);
and U16179 (N_16179,N_8754,N_8514);
nor U16180 (N_16180,N_7262,N_7501);
xor U16181 (N_16181,N_6627,N_11737);
or U16182 (N_16182,N_9390,N_10787);
xor U16183 (N_16183,N_6010,N_8412);
nor U16184 (N_16184,N_11876,N_9928);
nand U16185 (N_16185,N_6918,N_8369);
xor U16186 (N_16186,N_10713,N_9310);
nand U16187 (N_16187,N_7998,N_11287);
and U16188 (N_16188,N_11377,N_9976);
xor U16189 (N_16189,N_9924,N_7016);
or U16190 (N_16190,N_9137,N_9543);
and U16191 (N_16191,N_8054,N_6545);
or U16192 (N_16192,N_9097,N_8863);
nand U16193 (N_16193,N_6243,N_10312);
and U16194 (N_16194,N_6380,N_11414);
and U16195 (N_16195,N_10558,N_9472);
or U16196 (N_16196,N_8376,N_10631);
or U16197 (N_16197,N_8684,N_9326);
or U16198 (N_16198,N_7605,N_8106);
and U16199 (N_16199,N_7179,N_6818);
or U16200 (N_16200,N_8514,N_8246);
and U16201 (N_16201,N_6531,N_8812);
or U16202 (N_16202,N_8992,N_10697);
or U16203 (N_16203,N_11218,N_10839);
or U16204 (N_16204,N_7605,N_11838);
xor U16205 (N_16205,N_10133,N_8693);
nor U16206 (N_16206,N_11265,N_7658);
nand U16207 (N_16207,N_11856,N_6524);
xor U16208 (N_16208,N_11898,N_9081);
nand U16209 (N_16209,N_6685,N_10335);
and U16210 (N_16210,N_9995,N_11849);
nor U16211 (N_16211,N_8184,N_7881);
and U16212 (N_16212,N_9874,N_11976);
nand U16213 (N_16213,N_8294,N_10435);
nand U16214 (N_16214,N_10067,N_7680);
nand U16215 (N_16215,N_7437,N_11921);
nand U16216 (N_16216,N_7354,N_10512);
or U16217 (N_16217,N_6312,N_11853);
xor U16218 (N_16218,N_8014,N_11558);
nand U16219 (N_16219,N_6273,N_11145);
and U16220 (N_16220,N_10909,N_11241);
nand U16221 (N_16221,N_8799,N_6210);
or U16222 (N_16222,N_11566,N_11351);
nand U16223 (N_16223,N_6943,N_10528);
nand U16224 (N_16224,N_9879,N_8076);
or U16225 (N_16225,N_9775,N_11341);
nand U16226 (N_16226,N_8922,N_8003);
nor U16227 (N_16227,N_7744,N_9901);
and U16228 (N_16228,N_8201,N_6264);
or U16229 (N_16229,N_9661,N_6415);
and U16230 (N_16230,N_7616,N_6721);
or U16231 (N_16231,N_6273,N_11094);
nand U16232 (N_16232,N_6526,N_10900);
and U16233 (N_16233,N_11564,N_7569);
or U16234 (N_16234,N_8093,N_9361);
or U16235 (N_16235,N_7389,N_10313);
or U16236 (N_16236,N_9721,N_11265);
nor U16237 (N_16237,N_11823,N_7985);
nor U16238 (N_16238,N_7729,N_7952);
and U16239 (N_16239,N_6952,N_10801);
and U16240 (N_16240,N_6659,N_11765);
xor U16241 (N_16241,N_11655,N_7080);
and U16242 (N_16242,N_7317,N_8344);
nand U16243 (N_16243,N_11233,N_9988);
and U16244 (N_16244,N_9022,N_11831);
or U16245 (N_16245,N_9887,N_11638);
nand U16246 (N_16246,N_8382,N_8249);
and U16247 (N_16247,N_11388,N_9782);
nor U16248 (N_16248,N_11432,N_10809);
and U16249 (N_16249,N_11809,N_10472);
and U16250 (N_16250,N_8117,N_8400);
and U16251 (N_16251,N_6365,N_7278);
nor U16252 (N_16252,N_8112,N_6565);
xor U16253 (N_16253,N_8240,N_8520);
nand U16254 (N_16254,N_9834,N_6998);
nand U16255 (N_16255,N_8216,N_10507);
xnor U16256 (N_16256,N_6737,N_6582);
and U16257 (N_16257,N_6326,N_8837);
xor U16258 (N_16258,N_11742,N_8191);
nand U16259 (N_16259,N_7385,N_9142);
nand U16260 (N_16260,N_6045,N_8865);
and U16261 (N_16261,N_11724,N_11831);
xnor U16262 (N_16262,N_9467,N_9991);
and U16263 (N_16263,N_11036,N_9124);
or U16264 (N_16264,N_10103,N_11133);
or U16265 (N_16265,N_8807,N_6553);
xnor U16266 (N_16266,N_8194,N_8376);
and U16267 (N_16267,N_10827,N_6586);
nand U16268 (N_16268,N_7162,N_8538);
nand U16269 (N_16269,N_10022,N_9820);
nor U16270 (N_16270,N_7793,N_10501);
and U16271 (N_16271,N_9162,N_9720);
nand U16272 (N_16272,N_8099,N_7345);
nand U16273 (N_16273,N_8871,N_6246);
nor U16274 (N_16274,N_6412,N_7974);
or U16275 (N_16275,N_6083,N_9043);
nand U16276 (N_16276,N_10912,N_8077);
nand U16277 (N_16277,N_9462,N_9913);
xnor U16278 (N_16278,N_6396,N_9540);
or U16279 (N_16279,N_8822,N_7922);
xnor U16280 (N_16280,N_6433,N_9801);
and U16281 (N_16281,N_7578,N_6096);
or U16282 (N_16282,N_11187,N_7873);
nor U16283 (N_16283,N_9383,N_8336);
nor U16284 (N_16284,N_9778,N_11686);
xnor U16285 (N_16285,N_7201,N_11002);
and U16286 (N_16286,N_10633,N_7151);
xor U16287 (N_16287,N_8401,N_11089);
nand U16288 (N_16288,N_11047,N_9026);
and U16289 (N_16289,N_6757,N_6423);
nand U16290 (N_16290,N_10059,N_6301);
xor U16291 (N_16291,N_7747,N_7516);
and U16292 (N_16292,N_6958,N_10419);
xnor U16293 (N_16293,N_9746,N_8149);
and U16294 (N_16294,N_11758,N_11946);
xor U16295 (N_16295,N_11851,N_7296);
nor U16296 (N_16296,N_8984,N_9025);
and U16297 (N_16297,N_6263,N_6444);
xnor U16298 (N_16298,N_10359,N_8534);
or U16299 (N_16299,N_6084,N_9898);
nand U16300 (N_16300,N_7838,N_6835);
xor U16301 (N_16301,N_8497,N_8122);
xnor U16302 (N_16302,N_7486,N_8961);
or U16303 (N_16303,N_6793,N_10173);
or U16304 (N_16304,N_8831,N_7837);
and U16305 (N_16305,N_7122,N_6524);
nand U16306 (N_16306,N_10050,N_8161);
and U16307 (N_16307,N_9240,N_8112);
xnor U16308 (N_16308,N_10354,N_10585);
nor U16309 (N_16309,N_10826,N_8769);
and U16310 (N_16310,N_9121,N_9029);
or U16311 (N_16311,N_8314,N_9591);
or U16312 (N_16312,N_9386,N_9431);
nand U16313 (N_16313,N_11030,N_8491);
and U16314 (N_16314,N_11431,N_10924);
xnor U16315 (N_16315,N_10559,N_6254);
nor U16316 (N_16316,N_6237,N_9206);
xnor U16317 (N_16317,N_9979,N_10471);
nor U16318 (N_16318,N_9848,N_6578);
nand U16319 (N_16319,N_8790,N_6346);
or U16320 (N_16320,N_11689,N_6658);
or U16321 (N_16321,N_8169,N_11984);
nand U16322 (N_16322,N_7382,N_11428);
and U16323 (N_16323,N_10779,N_11911);
nor U16324 (N_16324,N_11875,N_6722);
xor U16325 (N_16325,N_9116,N_11494);
or U16326 (N_16326,N_9180,N_6986);
nand U16327 (N_16327,N_6607,N_8452);
or U16328 (N_16328,N_7998,N_7555);
or U16329 (N_16329,N_7678,N_10863);
nor U16330 (N_16330,N_9535,N_8426);
and U16331 (N_16331,N_7201,N_8690);
xor U16332 (N_16332,N_11467,N_10051);
xnor U16333 (N_16333,N_11506,N_11847);
or U16334 (N_16334,N_11646,N_6665);
nand U16335 (N_16335,N_6427,N_7170);
nand U16336 (N_16336,N_6292,N_11270);
nor U16337 (N_16337,N_9049,N_9034);
xnor U16338 (N_16338,N_9886,N_8650);
nor U16339 (N_16339,N_9105,N_6643);
and U16340 (N_16340,N_8863,N_10772);
nand U16341 (N_16341,N_7540,N_9612);
xnor U16342 (N_16342,N_10100,N_9004);
or U16343 (N_16343,N_6940,N_8349);
nand U16344 (N_16344,N_9661,N_7845);
and U16345 (N_16345,N_11494,N_10316);
nand U16346 (N_16346,N_6555,N_7354);
nor U16347 (N_16347,N_10125,N_6477);
and U16348 (N_16348,N_8498,N_8593);
and U16349 (N_16349,N_9108,N_7609);
nor U16350 (N_16350,N_11277,N_8272);
or U16351 (N_16351,N_7326,N_7196);
nand U16352 (N_16352,N_9165,N_9559);
and U16353 (N_16353,N_6031,N_7393);
nor U16354 (N_16354,N_9031,N_9001);
xnor U16355 (N_16355,N_11405,N_8257);
xnor U16356 (N_16356,N_11325,N_10955);
xnor U16357 (N_16357,N_10312,N_6919);
nor U16358 (N_16358,N_9625,N_6825);
nor U16359 (N_16359,N_6009,N_8859);
or U16360 (N_16360,N_8973,N_9432);
or U16361 (N_16361,N_8692,N_6474);
nor U16362 (N_16362,N_8884,N_10523);
xor U16363 (N_16363,N_10598,N_7258);
nor U16364 (N_16364,N_9242,N_10001);
nand U16365 (N_16365,N_7425,N_10588);
xor U16366 (N_16366,N_6265,N_11767);
or U16367 (N_16367,N_9129,N_8373);
and U16368 (N_16368,N_8914,N_8008);
or U16369 (N_16369,N_8957,N_10365);
nor U16370 (N_16370,N_7602,N_9727);
nand U16371 (N_16371,N_11362,N_6238);
nor U16372 (N_16372,N_10367,N_7978);
nor U16373 (N_16373,N_10683,N_7040);
xnor U16374 (N_16374,N_11818,N_8873);
nor U16375 (N_16375,N_11646,N_11391);
or U16376 (N_16376,N_8659,N_7203);
and U16377 (N_16377,N_10353,N_9452);
xnor U16378 (N_16378,N_8938,N_6050);
xor U16379 (N_16379,N_11770,N_9600);
xnor U16380 (N_16380,N_9249,N_8852);
xnor U16381 (N_16381,N_7569,N_6926);
xor U16382 (N_16382,N_6722,N_6916);
nand U16383 (N_16383,N_10383,N_6833);
and U16384 (N_16384,N_11615,N_7451);
or U16385 (N_16385,N_8070,N_6135);
xnor U16386 (N_16386,N_8060,N_10774);
nor U16387 (N_16387,N_7504,N_11058);
and U16388 (N_16388,N_6223,N_8557);
or U16389 (N_16389,N_7343,N_11559);
and U16390 (N_16390,N_7727,N_10392);
nand U16391 (N_16391,N_7722,N_11312);
and U16392 (N_16392,N_7345,N_8487);
xor U16393 (N_16393,N_11219,N_7071);
or U16394 (N_16394,N_9682,N_10486);
xnor U16395 (N_16395,N_10108,N_9240);
or U16396 (N_16396,N_9851,N_11383);
nor U16397 (N_16397,N_11439,N_8825);
nor U16398 (N_16398,N_6379,N_6043);
nor U16399 (N_16399,N_6599,N_7825);
nand U16400 (N_16400,N_11915,N_11121);
nor U16401 (N_16401,N_7769,N_7772);
or U16402 (N_16402,N_7242,N_9302);
and U16403 (N_16403,N_8436,N_7229);
or U16404 (N_16404,N_7028,N_10574);
and U16405 (N_16405,N_6664,N_9758);
or U16406 (N_16406,N_11362,N_7236);
xnor U16407 (N_16407,N_7352,N_7042);
and U16408 (N_16408,N_11919,N_8684);
xnor U16409 (N_16409,N_7621,N_8288);
xnor U16410 (N_16410,N_7684,N_11264);
xnor U16411 (N_16411,N_11455,N_6553);
or U16412 (N_16412,N_10798,N_7065);
xor U16413 (N_16413,N_7629,N_9458);
or U16414 (N_16414,N_9087,N_9329);
and U16415 (N_16415,N_11046,N_6271);
or U16416 (N_16416,N_11010,N_10007);
xnor U16417 (N_16417,N_7454,N_11563);
or U16418 (N_16418,N_9488,N_8505);
and U16419 (N_16419,N_6301,N_8393);
nor U16420 (N_16420,N_10567,N_11991);
and U16421 (N_16421,N_6501,N_11653);
or U16422 (N_16422,N_8227,N_9817);
and U16423 (N_16423,N_7505,N_7089);
or U16424 (N_16424,N_9221,N_9013);
or U16425 (N_16425,N_6146,N_9221);
xor U16426 (N_16426,N_8028,N_10236);
xor U16427 (N_16427,N_11877,N_8149);
nor U16428 (N_16428,N_8765,N_8085);
or U16429 (N_16429,N_6478,N_7437);
or U16430 (N_16430,N_8490,N_6927);
nand U16431 (N_16431,N_10136,N_11760);
nand U16432 (N_16432,N_10647,N_7457);
xnor U16433 (N_16433,N_7910,N_7083);
or U16434 (N_16434,N_11302,N_6038);
nand U16435 (N_16435,N_11827,N_11583);
and U16436 (N_16436,N_6117,N_11936);
xnor U16437 (N_16437,N_6648,N_10219);
and U16438 (N_16438,N_10719,N_10050);
nor U16439 (N_16439,N_10972,N_10231);
nand U16440 (N_16440,N_9868,N_8296);
nand U16441 (N_16441,N_6894,N_8620);
xnor U16442 (N_16442,N_11038,N_9221);
nor U16443 (N_16443,N_8120,N_6022);
nand U16444 (N_16444,N_9026,N_11597);
nor U16445 (N_16445,N_9937,N_11758);
or U16446 (N_16446,N_11605,N_7400);
nor U16447 (N_16447,N_7714,N_10322);
and U16448 (N_16448,N_8748,N_9652);
or U16449 (N_16449,N_10903,N_7519);
xor U16450 (N_16450,N_8499,N_9086);
xor U16451 (N_16451,N_9301,N_8286);
nand U16452 (N_16452,N_8336,N_10143);
nand U16453 (N_16453,N_8855,N_6355);
or U16454 (N_16454,N_11675,N_10540);
or U16455 (N_16455,N_9950,N_7243);
nor U16456 (N_16456,N_10274,N_6632);
nor U16457 (N_16457,N_6979,N_9055);
and U16458 (N_16458,N_11373,N_11153);
or U16459 (N_16459,N_10151,N_10143);
nand U16460 (N_16460,N_6791,N_8210);
or U16461 (N_16461,N_6140,N_7633);
nand U16462 (N_16462,N_8837,N_10565);
xnor U16463 (N_16463,N_8067,N_6336);
xnor U16464 (N_16464,N_8083,N_10151);
nand U16465 (N_16465,N_10053,N_9937);
nand U16466 (N_16466,N_6135,N_8893);
and U16467 (N_16467,N_9101,N_6286);
nor U16468 (N_16468,N_6498,N_10755);
or U16469 (N_16469,N_10997,N_6523);
xor U16470 (N_16470,N_7094,N_9315);
nor U16471 (N_16471,N_9759,N_6180);
xnor U16472 (N_16472,N_8111,N_7886);
or U16473 (N_16473,N_7563,N_11391);
nand U16474 (N_16474,N_9986,N_8934);
or U16475 (N_16475,N_9393,N_9745);
and U16476 (N_16476,N_10786,N_9213);
and U16477 (N_16477,N_8392,N_11346);
and U16478 (N_16478,N_9933,N_8601);
or U16479 (N_16479,N_11054,N_10272);
or U16480 (N_16480,N_10064,N_7041);
xnor U16481 (N_16481,N_7924,N_9625);
xor U16482 (N_16482,N_7277,N_10680);
xnor U16483 (N_16483,N_9455,N_8372);
and U16484 (N_16484,N_10344,N_9050);
nand U16485 (N_16485,N_8615,N_10612);
xor U16486 (N_16486,N_9315,N_8438);
xor U16487 (N_16487,N_7707,N_11064);
nand U16488 (N_16488,N_9110,N_9853);
nor U16489 (N_16489,N_11329,N_10371);
xor U16490 (N_16490,N_9933,N_11722);
nor U16491 (N_16491,N_6971,N_8474);
nor U16492 (N_16492,N_6339,N_10211);
nor U16493 (N_16493,N_7025,N_9214);
and U16494 (N_16494,N_8666,N_8476);
and U16495 (N_16495,N_10991,N_7180);
nand U16496 (N_16496,N_11046,N_9365);
and U16497 (N_16497,N_8685,N_7981);
nand U16498 (N_16498,N_11942,N_11452);
xor U16499 (N_16499,N_10886,N_8811);
and U16500 (N_16500,N_9465,N_10005);
and U16501 (N_16501,N_10745,N_7599);
nor U16502 (N_16502,N_10092,N_8220);
and U16503 (N_16503,N_9771,N_10233);
or U16504 (N_16504,N_9789,N_8205);
nor U16505 (N_16505,N_7002,N_7994);
nand U16506 (N_16506,N_6537,N_6014);
xnor U16507 (N_16507,N_11408,N_11935);
nor U16508 (N_16508,N_6733,N_8612);
and U16509 (N_16509,N_10158,N_7090);
and U16510 (N_16510,N_7207,N_9436);
or U16511 (N_16511,N_9129,N_6081);
nor U16512 (N_16512,N_7982,N_11690);
nor U16513 (N_16513,N_9271,N_8285);
or U16514 (N_16514,N_6424,N_7826);
xor U16515 (N_16515,N_7090,N_9773);
or U16516 (N_16516,N_10473,N_8393);
or U16517 (N_16517,N_6477,N_9527);
nand U16518 (N_16518,N_6563,N_11479);
or U16519 (N_16519,N_10490,N_9329);
nor U16520 (N_16520,N_9117,N_10135);
nor U16521 (N_16521,N_6146,N_10456);
nor U16522 (N_16522,N_10841,N_11900);
and U16523 (N_16523,N_11196,N_7940);
nor U16524 (N_16524,N_6489,N_9385);
and U16525 (N_16525,N_8784,N_8458);
nand U16526 (N_16526,N_11655,N_9426);
and U16527 (N_16527,N_11883,N_9531);
or U16528 (N_16528,N_8893,N_9034);
nor U16529 (N_16529,N_7285,N_8027);
xor U16530 (N_16530,N_7885,N_6712);
xor U16531 (N_16531,N_6453,N_10661);
nor U16532 (N_16532,N_11671,N_9892);
or U16533 (N_16533,N_8041,N_6685);
nor U16534 (N_16534,N_8344,N_6580);
nand U16535 (N_16535,N_7265,N_8397);
and U16536 (N_16536,N_8280,N_10751);
or U16537 (N_16537,N_8839,N_8811);
or U16538 (N_16538,N_6426,N_11264);
nand U16539 (N_16539,N_9502,N_7469);
nor U16540 (N_16540,N_8929,N_7902);
and U16541 (N_16541,N_9117,N_7524);
xnor U16542 (N_16542,N_6525,N_8609);
xor U16543 (N_16543,N_8170,N_6675);
or U16544 (N_16544,N_9603,N_11062);
xor U16545 (N_16545,N_8330,N_10521);
xnor U16546 (N_16546,N_10566,N_11167);
or U16547 (N_16547,N_9755,N_10296);
xnor U16548 (N_16548,N_8335,N_9969);
xnor U16549 (N_16549,N_8477,N_11411);
xor U16550 (N_16550,N_11110,N_9986);
or U16551 (N_16551,N_11565,N_8890);
xnor U16552 (N_16552,N_8204,N_9683);
or U16553 (N_16553,N_6104,N_9959);
and U16554 (N_16554,N_11548,N_8396);
or U16555 (N_16555,N_7556,N_11883);
nor U16556 (N_16556,N_10624,N_6194);
nor U16557 (N_16557,N_10295,N_6028);
nor U16558 (N_16558,N_10646,N_11361);
and U16559 (N_16559,N_11085,N_10928);
nand U16560 (N_16560,N_6523,N_11849);
nor U16561 (N_16561,N_11766,N_7661);
xor U16562 (N_16562,N_7772,N_6240);
and U16563 (N_16563,N_10245,N_10645);
nor U16564 (N_16564,N_9294,N_8882);
xor U16565 (N_16565,N_7131,N_9609);
nand U16566 (N_16566,N_8305,N_8640);
nor U16567 (N_16567,N_9578,N_7256);
or U16568 (N_16568,N_6258,N_11003);
nand U16569 (N_16569,N_8674,N_7167);
nand U16570 (N_16570,N_11503,N_7809);
or U16571 (N_16571,N_8206,N_10921);
nor U16572 (N_16572,N_10570,N_11050);
or U16573 (N_16573,N_8438,N_6782);
and U16574 (N_16574,N_11154,N_10335);
nor U16575 (N_16575,N_9958,N_6786);
and U16576 (N_16576,N_6833,N_11413);
nor U16577 (N_16577,N_10748,N_10712);
nand U16578 (N_16578,N_11692,N_7053);
xor U16579 (N_16579,N_7063,N_11930);
nand U16580 (N_16580,N_10055,N_6939);
and U16581 (N_16581,N_9108,N_8740);
and U16582 (N_16582,N_11854,N_9624);
or U16583 (N_16583,N_7232,N_9469);
nand U16584 (N_16584,N_9890,N_9432);
nand U16585 (N_16585,N_8253,N_11073);
nand U16586 (N_16586,N_11156,N_6763);
and U16587 (N_16587,N_11838,N_8711);
or U16588 (N_16588,N_8565,N_7326);
and U16589 (N_16589,N_8504,N_8931);
nor U16590 (N_16590,N_9977,N_8075);
nor U16591 (N_16591,N_10124,N_11953);
or U16592 (N_16592,N_11259,N_10615);
xnor U16593 (N_16593,N_7417,N_11337);
nor U16594 (N_16594,N_11251,N_11956);
nor U16595 (N_16595,N_10412,N_9739);
nor U16596 (N_16596,N_6017,N_9376);
and U16597 (N_16597,N_11006,N_6344);
or U16598 (N_16598,N_11029,N_8605);
and U16599 (N_16599,N_7945,N_9359);
nor U16600 (N_16600,N_8458,N_7650);
xor U16601 (N_16601,N_10329,N_8591);
or U16602 (N_16602,N_8291,N_11312);
xor U16603 (N_16603,N_10110,N_9105);
nand U16604 (N_16604,N_8136,N_8745);
xor U16605 (N_16605,N_10598,N_7230);
and U16606 (N_16606,N_6527,N_6794);
nor U16607 (N_16607,N_6797,N_11281);
nand U16608 (N_16608,N_10852,N_9801);
nand U16609 (N_16609,N_7224,N_10235);
and U16610 (N_16610,N_11247,N_9565);
or U16611 (N_16611,N_10997,N_10483);
nand U16612 (N_16612,N_8688,N_9658);
xnor U16613 (N_16613,N_10094,N_10472);
nor U16614 (N_16614,N_11359,N_6968);
or U16615 (N_16615,N_9850,N_11381);
nand U16616 (N_16616,N_6174,N_8499);
and U16617 (N_16617,N_11680,N_7959);
or U16618 (N_16618,N_11560,N_7328);
or U16619 (N_16619,N_11895,N_9172);
and U16620 (N_16620,N_11941,N_8267);
xor U16621 (N_16621,N_10224,N_9069);
nand U16622 (N_16622,N_10750,N_9506);
nand U16623 (N_16623,N_11331,N_10268);
and U16624 (N_16624,N_11089,N_7469);
and U16625 (N_16625,N_9654,N_10059);
and U16626 (N_16626,N_10124,N_6378);
or U16627 (N_16627,N_7258,N_8245);
nor U16628 (N_16628,N_11600,N_8492);
nor U16629 (N_16629,N_11018,N_8369);
nand U16630 (N_16630,N_8009,N_9145);
or U16631 (N_16631,N_6192,N_10080);
or U16632 (N_16632,N_9409,N_11864);
xor U16633 (N_16633,N_6809,N_6892);
nand U16634 (N_16634,N_6674,N_10740);
nor U16635 (N_16635,N_7109,N_8394);
nor U16636 (N_16636,N_7298,N_7355);
nor U16637 (N_16637,N_8215,N_11046);
or U16638 (N_16638,N_9863,N_8384);
or U16639 (N_16639,N_8518,N_9957);
and U16640 (N_16640,N_11894,N_11095);
and U16641 (N_16641,N_8076,N_10824);
nand U16642 (N_16642,N_6510,N_7498);
nor U16643 (N_16643,N_7171,N_11216);
nor U16644 (N_16644,N_10148,N_8382);
and U16645 (N_16645,N_11755,N_11399);
or U16646 (N_16646,N_9854,N_7997);
and U16647 (N_16647,N_11276,N_6259);
or U16648 (N_16648,N_8031,N_6683);
nand U16649 (N_16649,N_7745,N_10842);
or U16650 (N_16650,N_6747,N_10188);
xnor U16651 (N_16651,N_11148,N_9806);
and U16652 (N_16652,N_6382,N_7764);
or U16653 (N_16653,N_7124,N_7708);
xor U16654 (N_16654,N_6446,N_7427);
xor U16655 (N_16655,N_9508,N_7980);
nor U16656 (N_16656,N_8723,N_9580);
nand U16657 (N_16657,N_8794,N_9919);
and U16658 (N_16658,N_11483,N_9512);
xor U16659 (N_16659,N_10698,N_8532);
nand U16660 (N_16660,N_11334,N_6381);
xor U16661 (N_16661,N_7699,N_9430);
xnor U16662 (N_16662,N_7087,N_9970);
xnor U16663 (N_16663,N_10001,N_6196);
xor U16664 (N_16664,N_11934,N_10163);
and U16665 (N_16665,N_11215,N_9328);
nand U16666 (N_16666,N_9305,N_9545);
and U16667 (N_16667,N_9220,N_8656);
or U16668 (N_16668,N_10059,N_7262);
nor U16669 (N_16669,N_9546,N_10427);
or U16670 (N_16670,N_10160,N_11893);
and U16671 (N_16671,N_8826,N_7935);
or U16672 (N_16672,N_10160,N_9893);
nand U16673 (N_16673,N_7100,N_8165);
and U16674 (N_16674,N_11090,N_8922);
nand U16675 (N_16675,N_6720,N_7767);
or U16676 (N_16676,N_7818,N_11709);
and U16677 (N_16677,N_9863,N_11711);
nand U16678 (N_16678,N_8685,N_11937);
and U16679 (N_16679,N_9858,N_7359);
nand U16680 (N_16680,N_10908,N_6268);
or U16681 (N_16681,N_11868,N_9862);
nand U16682 (N_16682,N_7482,N_11862);
nor U16683 (N_16683,N_9933,N_9163);
and U16684 (N_16684,N_7163,N_7825);
and U16685 (N_16685,N_7276,N_7855);
nand U16686 (N_16686,N_10577,N_6004);
xor U16687 (N_16687,N_8150,N_7439);
nand U16688 (N_16688,N_7799,N_6192);
nor U16689 (N_16689,N_10685,N_8479);
or U16690 (N_16690,N_8765,N_7869);
and U16691 (N_16691,N_6177,N_10707);
or U16692 (N_16692,N_9881,N_6511);
nor U16693 (N_16693,N_9379,N_8532);
nor U16694 (N_16694,N_9157,N_9678);
nor U16695 (N_16695,N_10903,N_11315);
nand U16696 (N_16696,N_9695,N_10888);
xor U16697 (N_16697,N_8825,N_8217);
or U16698 (N_16698,N_8325,N_8937);
nor U16699 (N_16699,N_9658,N_9373);
or U16700 (N_16700,N_11191,N_7755);
and U16701 (N_16701,N_11227,N_9960);
or U16702 (N_16702,N_7997,N_11273);
and U16703 (N_16703,N_11112,N_7866);
or U16704 (N_16704,N_8883,N_9716);
nor U16705 (N_16705,N_8414,N_10350);
xnor U16706 (N_16706,N_10938,N_7432);
nand U16707 (N_16707,N_10802,N_8541);
nand U16708 (N_16708,N_8861,N_9136);
nand U16709 (N_16709,N_9126,N_6551);
nand U16710 (N_16710,N_6098,N_8471);
and U16711 (N_16711,N_8244,N_8849);
nor U16712 (N_16712,N_7212,N_8466);
and U16713 (N_16713,N_8981,N_8406);
and U16714 (N_16714,N_10924,N_7684);
xor U16715 (N_16715,N_10888,N_11467);
nor U16716 (N_16716,N_8000,N_9314);
xnor U16717 (N_16717,N_6764,N_8727);
or U16718 (N_16718,N_6563,N_10462);
and U16719 (N_16719,N_8324,N_6594);
and U16720 (N_16720,N_8122,N_8024);
nand U16721 (N_16721,N_10493,N_10079);
or U16722 (N_16722,N_10242,N_7074);
nand U16723 (N_16723,N_10076,N_9148);
nor U16724 (N_16724,N_10025,N_10888);
xnor U16725 (N_16725,N_8818,N_9019);
xnor U16726 (N_16726,N_11708,N_11927);
nand U16727 (N_16727,N_8609,N_8135);
nor U16728 (N_16728,N_8119,N_8700);
nand U16729 (N_16729,N_7803,N_6167);
xnor U16730 (N_16730,N_7009,N_9723);
nor U16731 (N_16731,N_11872,N_11814);
xor U16732 (N_16732,N_8368,N_11805);
nor U16733 (N_16733,N_7989,N_10259);
nor U16734 (N_16734,N_10993,N_7063);
xor U16735 (N_16735,N_7775,N_8763);
and U16736 (N_16736,N_6755,N_6151);
nand U16737 (N_16737,N_7785,N_7067);
nor U16738 (N_16738,N_11973,N_6994);
nand U16739 (N_16739,N_6210,N_7616);
nand U16740 (N_16740,N_11780,N_10216);
or U16741 (N_16741,N_10768,N_8992);
xnor U16742 (N_16742,N_6244,N_11164);
nor U16743 (N_16743,N_6115,N_7452);
xnor U16744 (N_16744,N_6579,N_6114);
and U16745 (N_16745,N_9906,N_11503);
xnor U16746 (N_16746,N_10240,N_6509);
and U16747 (N_16747,N_11158,N_11650);
nand U16748 (N_16748,N_8840,N_11402);
nand U16749 (N_16749,N_10688,N_6484);
and U16750 (N_16750,N_8900,N_11033);
nor U16751 (N_16751,N_7901,N_7274);
nand U16752 (N_16752,N_11639,N_9316);
xor U16753 (N_16753,N_7672,N_6121);
or U16754 (N_16754,N_11630,N_7646);
nor U16755 (N_16755,N_6446,N_8138);
nand U16756 (N_16756,N_11441,N_7865);
nor U16757 (N_16757,N_6211,N_10259);
nand U16758 (N_16758,N_8886,N_7588);
nor U16759 (N_16759,N_6724,N_6614);
xnor U16760 (N_16760,N_7474,N_8256);
nor U16761 (N_16761,N_6545,N_11122);
nand U16762 (N_16762,N_7942,N_10092);
nor U16763 (N_16763,N_6945,N_6135);
nand U16764 (N_16764,N_7332,N_7115);
nand U16765 (N_16765,N_6740,N_7206);
or U16766 (N_16766,N_7453,N_10050);
xnor U16767 (N_16767,N_10370,N_8870);
and U16768 (N_16768,N_11168,N_10562);
and U16769 (N_16769,N_8609,N_10113);
nand U16770 (N_16770,N_8058,N_6980);
xor U16771 (N_16771,N_9626,N_6293);
or U16772 (N_16772,N_6899,N_10346);
nand U16773 (N_16773,N_11799,N_8595);
nor U16774 (N_16774,N_8223,N_6013);
nand U16775 (N_16775,N_9394,N_7912);
nor U16776 (N_16776,N_9312,N_10513);
nor U16777 (N_16777,N_6103,N_10346);
or U16778 (N_16778,N_9668,N_9677);
xor U16779 (N_16779,N_10852,N_9163);
and U16780 (N_16780,N_8421,N_8207);
nor U16781 (N_16781,N_10953,N_7394);
xnor U16782 (N_16782,N_9508,N_11869);
or U16783 (N_16783,N_9647,N_6041);
nor U16784 (N_16784,N_8138,N_9333);
or U16785 (N_16785,N_10908,N_7485);
nor U16786 (N_16786,N_11724,N_10196);
nor U16787 (N_16787,N_11024,N_11037);
nand U16788 (N_16788,N_7694,N_7830);
xor U16789 (N_16789,N_10859,N_8700);
nor U16790 (N_16790,N_10016,N_8880);
nor U16791 (N_16791,N_7733,N_10582);
nor U16792 (N_16792,N_9258,N_9654);
and U16793 (N_16793,N_6362,N_9090);
xnor U16794 (N_16794,N_11087,N_7293);
nor U16795 (N_16795,N_10242,N_7868);
xnor U16796 (N_16796,N_10445,N_8064);
nor U16797 (N_16797,N_8534,N_11766);
xor U16798 (N_16798,N_11513,N_8854);
and U16799 (N_16799,N_9619,N_10326);
xor U16800 (N_16800,N_8241,N_9467);
nor U16801 (N_16801,N_10254,N_11925);
nand U16802 (N_16802,N_10787,N_10474);
and U16803 (N_16803,N_11775,N_8537);
xnor U16804 (N_16804,N_7879,N_8510);
nor U16805 (N_16805,N_9103,N_6931);
xor U16806 (N_16806,N_7856,N_11616);
and U16807 (N_16807,N_10626,N_11285);
or U16808 (N_16808,N_11657,N_8190);
nor U16809 (N_16809,N_6634,N_10023);
nor U16810 (N_16810,N_11317,N_11981);
xnor U16811 (N_16811,N_7627,N_11069);
nand U16812 (N_16812,N_11956,N_6906);
nor U16813 (N_16813,N_10412,N_9366);
nor U16814 (N_16814,N_9490,N_6941);
xor U16815 (N_16815,N_9476,N_10112);
nand U16816 (N_16816,N_9095,N_6905);
and U16817 (N_16817,N_6027,N_10787);
xor U16818 (N_16818,N_8553,N_10805);
xnor U16819 (N_16819,N_6045,N_9252);
nand U16820 (N_16820,N_6480,N_7730);
nand U16821 (N_16821,N_6451,N_11555);
and U16822 (N_16822,N_7920,N_11645);
and U16823 (N_16823,N_7890,N_11138);
or U16824 (N_16824,N_9399,N_10480);
or U16825 (N_16825,N_7205,N_9736);
xor U16826 (N_16826,N_10170,N_9180);
nor U16827 (N_16827,N_10502,N_7685);
nand U16828 (N_16828,N_11353,N_8537);
xnor U16829 (N_16829,N_10167,N_6015);
nand U16830 (N_16830,N_8528,N_9365);
and U16831 (N_16831,N_7331,N_11839);
nor U16832 (N_16832,N_6608,N_7426);
or U16833 (N_16833,N_10183,N_8845);
xnor U16834 (N_16834,N_10389,N_9704);
nor U16835 (N_16835,N_8998,N_7708);
nor U16836 (N_16836,N_11376,N_10647);
xor U16837 (N_16837,N_6014,N_7328);
and U16838 (N_16838,N_7312,N_6135);
and U16839 (N_16839,N_8050,N_7070);
xnor U16840 (N_16840,N_11293,N_11066);
xnor U16841 (N_16841,N_11618,N_6905);
nor U16842 (N_16842,N_7657,N_10470);
or U16843 (N_16843,N_9794,N_9057);
and U16844 (N_16844,N_8738,N_11751);
nand U16845 (N_16845,N_8696,N_10416);
nand U16846 (N_16846,N_7433,N_9531);
nor U16847 (N_16847,N_10703,N_6033);
nor U16848 (N_16848,N_10854,N_9328);
and U16849 (N_16849,N_9843,N_11619);
xnor U16850 (N_16850,N_10812,N_9127);
or U16851 (N_16851,N_9960,N_7984);
xnor U16852 (N_16852,N_6232,N_9164);
nand U16853 (N_16853,N_7558,N_8804);
nand U16854 (N_16854,N_10412,N_11701);
xnor U16855 (N_16855,N_10717,N_11204);
and U16856 (N_16856,N_9100,N_8862);
nand U16857 (N_16857,N_9611,N_9953);
or U16858 (N_16858,N_7509,N_10384);
and U16859 (N_16859,N_8207,N_9988);
or U16860 (N_16860,N_10440,N_7761);
nand U16861 (N_16861,N_10457,N_7565);
and U16862 (N_16862,N_9273,N_8879);
nor U16863 (N_16863,N_10006,N_9054);
or U16864 (N_16864,N_6773,N_6632);
or U16865 (N_16865,N_8436,N_7331);
or U16866 (N_16866,N_11448,N_11421);
or U16867 (N_16867,N_11391,N_11685);
nor U16868 (N_16868,N_8966,N_7383);
nand U16869 (N_16869,N_8184,N_8443);
and U16870 (N_16870,N_8322,N_6615);
or U16871 (N_16871,N_8369,N_8168);
nand U16872 (N_16872,N_7331,N_11651);
and U16873 (N_16873,N_6835,N_8898);
or U16874 (N_16874,N_10919,N_7105);
nor U16875 (N_16875,N_7474,N_7200);
nor U16876 (N_16876,N_8997,N_11543);
nor U16877 (N_16877,N_10485,N_10091);
nor U16878 (N_16878,N_10491,N_11870);
xor U16879 (N_16879,N_7373,N_11041);
nor U16880 (N_16880,N_8523,N_9639);
nor U16881 (N_16881,N_11849,N_7160);
and U16882 (N_16882,N_8574,N_9378);
xnor U16883 (N_16883,N_10738,N_11041);
xor U16884 (N_16884,N_11664,N_9506);
or U16885 (N_16885,N_7032,N_8488);
nor U16886 (N_16886,N_7149,N_11094);
nor U16887 (N_16887,N_8127,N_11561);
nor U16888 (N_16888,N_8417,N_9612);
nor U16889 (N_16889,N_10406,N_6122);
nor U16890 (N_16890,N_8504,N_11546);
nand U16891 (N_16891,N_6038,N_11846);
or U16892 (N_16892,N_7390,N_8808);
xnor U16893 (N_16893,N_8415,N_8670);
and U16894 (N_16894,N_11865,N_10219);
or U16895 (N_16895,N_9051,N_7612);
or U16896 (N_16896,N_7790,N_7135);
or U16897 (N_16897,N_9873,N_7030);
and U16898 (N_16898,N_7723,N_9742);
nand U16899 (N_16899,N_10074,N_10627);
xor U16900 (N_16900,N_6323,N_6712);
nand U16901 (N_16901,N_9780,N_7610);
or U16902 (N_16902,N_8007,N_7267);
nand U16903 (N_16903,N_10748,N_7770);
and U16904 (N_16904,N_8641,N_9973);
and U16905 (N_16905,N_8644,N_9315);
nand U16906 (N_16906,N_11155,N_7465);
or U16907 (N_16907,N_9287,N_7258);
and U16908 (N_16908,N_11764,N_9681);
xnor U16909 (N_16909,N_8021,N_8200);
xnor U16910 (N_16910,N_8443,N_11080);
and U16911 (N_16911,N_9711,N_11239);
nand U16912 (N_16912,N_10212,N_9304);
nor U16913 (N_16913,N_7923,N_11949);
nor U16914 (N_16914,N_9211,N_6958);
and U16915 (N_16915,N_6330,N_11472);
nor U16916 (N_16916,N_6818,N_6549);
nor U16917 (N_16917,N_7077,N_6853);
nor U16918 (N_16918,N_6660,N_8744);
xor U16919 (N_16919,N_10687,N_6696);
nor U16920 (N_16920,N_9016,N_7047);
or U16921 (N_16921,N_9666,N_8087);
nor U16922 (N_16922,N_9143,N_6502);
and U16923 (N_16923,N_6015,N_6104);
nor U16924 (N_16924,N_10978,N_6606);
and U16925 (N_16925,N_7195,N_10134);
nand U16926 (N_16926,N_7492,N_11778);
xor U16927 (N_16927,N_9416,N_8895);
nand U16928 (N_16928,N_6924,N_11947);
nand U16929 (N_16929,N_7585,N_6136);
or U16930 (N_16930,N_7471,N_10024);
xor U16931 (N_16931,N_11515,N_10657);
or U16932 (N_16932,N_11268,N_10131);
or U16933 (N_16933,N_9907,N_10542);
or U16934 (N_16934,N_6475,N_11431);
xor U16935 (N_16935,N_8943,N_11209);
xor U16936 (N_16936,N_10200,N_11896);
nor U16937 (N_16937,N_11143,N_11738);
or U16938 (N_16938,N_8709,N_8873);
xnor U16939 (N_16939,N_11822,N_7267);
xor U16940 (N_16940,N_11358,N_9120);
xor U16941 (N_16941,N_9568,N_9390);
or U16942 (N_16942,N_9547,N_10525);
or U16943 (N_16943,N_11599,N_10055);
nor U16944 (N_16944,N_11345,N_9234);
nor U16945 (N_16945,N_9708,N_11946);
or U16946 (N_16946,N_7848,N_8596);
nand U16947 (N_16947,N_6542,N_8769);
nand U16948 (N_16948,N_8180,N_10546);
or U16949 (N_16949,N_11575,N_10095);
and U16950 (N_16950,N_6985,N_8476);
nand U16951 (N_16951,N_11172,N_10868);
nand U16952 (N_16952,N_7493,N_9364);
and U16953 (N_16953,N_9663,N_6418);
or U16954 (N_16954,N_8823,N_7906);
xnor U16955 (N_16955,N_10873,N_10931);
xor U16956 (N_16956,N_6098,N_10858);
nand U16957 (N_16957,N_9830,N_7509);
or U16958 (N_16958,N_6091,N_6172);
nor U16959 (N_16959,N_8364,N_10480);
and U16960 (N_16960,N_7639,N_6850);
xnor U16961 (N_16961,N_6736,N_6161);
nand U16962 (N_16962,N_7512,N_11062);
nor U16963 (N_16963,N_11769,N_8205);
and U16964 (N_16964,N_6867,N_8171);
xnor U16965 (N_16965,N_8001,N_7020);
nor U16966 (N_16966,N_7267,N_7206);
and U16967 (N_16967,N_11760,N_10140);
and U16968 (N_16968,N_8739,N_6998);
and U16969 (N_16969,N_6333,N_11068);
or U16970 (N_16970,N_11703,N_8327);
or U16971 (N_16971,N_9491,N_7994);
or U16972 (N_16972,N_10707,N_6541);
xnor U16973 (N_16973,N_11030,N_11988);
or U16974 (N_16974,N_8007,N_6811);
nand U16975 (N_16975,N_10955,N_10429);
or U16976 (N_16976,N_6706,N_10933);
nand U16977 (N_16977,N_6538,N_9477);
or U16978 (N_16978,N_6989,N_8570);
nor U16979 (N_16979,N_10335,N_9278);
or U16980 (N_16980,N_7454,N_10620);
or U16981 (N_16981,N_6833,N_11133);
and U16982 (N_16982,N_11486,N_11038);
nor U16983 (N_16983,N_8831,N_8435);
and U16984 (N_16984,N_8131,N_11004);
xnor U16985 (N_16985,N_11369,N_9982);
nor U16986 (N_16986,N_8203,N_10659);
and U16987 (N_16987,N_11404,N_8341);
and U16988 (N_16988,N_9777,N_7233);
xor U16989 (N_16989,N_9272,N_10230);
nand U16990 (N_16990,N_8503,N_11947);
nand U16991 (N_16991,N_10960,N_8985);
nand U16992 (N_16992,N_6419,N_10302);
nand U16993 (N_16993,N_8483,N_6330);
xnor U16994 (N_16994,N_11976,N_8713);
xnor U16995 (N_16995,N_6129,N_7522);
and U16996 (N_16996,N_6362,N_7118);
or U16997 (N_16997,N_7794,N_9068);
and U16998 (N_16998,N_8481,N_11817);
or U16999 (N_16999,N_10292,N_11464);
nor U17000 (N_17000,N_10662,N_10757);
nor U17001 (N_17001,N_6582,N_7595);
and U17002 (N_17002,N_7849,N_9866);
or U17003 (N_17003,N_6020,N_7186);
xor U17004 (N_17004,N_6149,N_10746);
xnor U17005 (N_17005,N_6843,N_6384);
xor U17006 (N_17006,N_8287,N_6362);
or U17007 (N_17007,N_9158,N_7229);
and U17008 (N_17008,N_7736,N_7041);
xor U17009 (N_17009,N_9443,N_6257);
nand U17010 (N_17010,N_8679,N_8801);
and U17011 (N_17011,N_11678,N_11558);
xnor U17012 (N_17012,N_11613,N_8185);
or U17013 (N_17013,N_6685,N_6214);
nor U17014 (N_17014,N_7340,N_8872);
or U17015 (N_17015,N_8909,N_7508);
and U17016 (N_17016,N_6220,N_7019);
nor U17017 (N_17017,N_7966,N_9940);
nor U17018 (N_17018,N_8591,N_7026);
xnor U17019 (N_17019,N_11046,N_6104);
or U17020 (N_17020,N_8630,N_9612);
or U17021 (N_17021,N_8884,N_7005);
nand U17022 (N_17022,N_6875,N_11737);
nor U17023 (N_17023,N_11086,N_9847);
nand U17024 (N_17024,N_11073,N_8980);
xnor U17025 (N_17025,N_8243,N_7646);
and U17026 (N_17026,N_10943,N_7994);
nand U17027 (N_17027,N_8842,N_8269);
or U17028 (N_17028,N_10441,N_9193);
nand U17029 (N_17029,N_11961,N_10713);
xor U17030 (N_17030,N_8755,N_8747);
xnor U17031 (N_17031,N_10603,N_10687);
nor U17032 (N_17032,N_11608,N_8943);
xnor U17033 (N_17033,N_7289,N_6213);
xnor U17034 (N_17034,N_8925,N_7020);
nand U17035 (N_17035,N_10957,N_7799);
nor U17036 (N_17036,N_8721,N_10349);
and U17037 (N_17037,N_8465,N_8558);
xor U17038 (N_17038,N_11648,N_9928);
nand U17039 (N_17039,N_7385,N_8714);
xor U17040 (N_17040,N_10808,N_7928);
and U17041 (N_17041,N_8186,N_9579);
or U17042 (N_17042,N_8057,N_7064);
nor U17043 (N_17043,N_8687,N_6007);
xor U17044 (N_17044,N_8895,N_8266);
xor U17045 (N_17045,N_11465,N_7609);
xnor U17046 (N_17046,N_7971,N_7076);
and U17047 (N_17047,N_7616,N_9937);
nand U17048 (N_17048,N_9458,N_8655);
nand U17049 (N_17049,N_8740,N_6102);
nor U17050 (N_17050,N_9079,N_9855);
nor U17051 (N_17051,N_10525,N_6888);
nor U17052 (N_17052,N_7477,N_6415);
xor U17053 (N_17053,N_10260,N_8713);
or U17054 (N_17054,N_8412,N_6299);
nand U17055 (N_17055,N_7642,N_9218);
xnor U17056 (N_17056,N_9040,N_8580);
and U17057 (N_17057,N_9457,N_7252);
nor U17058 (N_17058,N_10482,N_6632);
nor U17059 (N_17059,N_10979,N_9075);
nand U17060 (N_17060,N_9301,N_8736);
or U17061 (N_17061,N_9179,N_6896);
nand U17062 (N_17062,N_9535,N_10184);
or U17063 (N_17063,N_7030,N_8592);
or U17064 (N_17064,N_6293,N_8675);
and U17065 (N_17065,N_11134,N_7598);
nand U17066 (N_17066,N_7110,N_7247);
xor U17067 (N_17067,N_10761,N_9089);
xnor U17068 (N_17068,N_8416,N_8346);
or U17069 (N_17069,N_7726,N_11039);
nor U17070 (N_17070,N_11636,N_6230);
or U17071 (N_17071,N_11213,N_6902);
nor U17072 (N_17072,N_6178,N_6453);
and U17073 (N_17073,N_10176,N_10267);
nor U17074 (N_17074,N_10439,N_7746);
nand U17075 (N_17075,N_6264,N_6035);
nand U17076 (N_17076,N_10782,N_8636);
nor U17077 (N_17077,N_8939,N_7513);
or U17078 (N_17078,N_10514,N_11008);
or U17079 (N_17079,N_10638,N_10944);
or U17080 (N_17080,N_7156,N_10273);
and U17081 (N_17081,N_7905,N_7499);
or U17082 (N_17082,N_7123,N_7899);
or U17083 (N_17083,N_6299,N_6820);
nor U17084 (N_17084,N_8676,N_11530);
and U17085 (N_17085,N_6378,N_9390);
xnor U17086 (N_17086,N_11383,N_8214);
nand U17087 (N_17087,N_8599,N_9855);
or U17088 (N_17088,N_7104,N_10571);
nand U17089 (N_17089,N_7489,N_9506);
xor U17090 (N_17090,N_7206,N_6820);
and U17091 (N_17091,N_10703,N_8534);
and U17092 (N_17092,N_8469,N_8634);
nand U17093 (N_17093,N_6399,N_7426);
nor U17094 (N_17094,N_10876,N_11730);
nor U17095 (N_17095,N_9075,N_7286);
or U17096 (N_17096,N_8258,N_7404);
or U17097 (N_17097,N_6895,N_8994);
xor U17098 (N_17098,N_10879,N_6017);
xnor U17099 (N_17099,N_9308,N_8848);
nor U17100 (N_17100,N_7943,N_10133);
xnor U17101 (N_17101,N_6866,N_6760);
or U17102 (N_17102,N_8535,N_6170);
or U17103 (N_17103,N_7756,N_7636);
or U17104 (N_17104,N_6382,N_7006);
and U17105 (N_17105,N_8868,N_10334);
and U17106 (N_17106,N_11598,N_10488);
or U17107 (N_17107,N_9534,N_9252);
nor U17108 (N_17108,N_6768,N_9723);
or U17109 (N_17109,N_10844,N_10950);
and U17110 (N_17110,N_10781,N_11402);
nor U17111 (N_17111,N_9674,N_8939);
and U17112 (N_17112,N_7907,N_9692);
or U17113 (N_17113,N_6286,N_11656);
nand U17114 (N_17114,N_8155,N_6022);
and U17115 (N_17115,N_6393,N_9113);
nand U17116 (N_17116,N_7682,N_6674);
nor U17117 (N_17117,N_8109,N_6506);
nand U17118 (N_17118,N_6097,N_11171);
xor U17119 (N_17119,N_11886,N_11149);
and U17120 (N_17120,N_9117,N_11490);
nand U17121 (N_17121,N_9076,N_7879);
or U17122 (N_17122,N_6703,N_6605);
nor U17123 (N_17123,N_6684,N_7202);
nor U17124 (N_17124,N_6325,N_6826);
nor U17125 (N_17125,N_10202,N_9278);
nor U17126 (N_17126,N_11339,N_11253);
nor U17127 (N_17127,N_10550,N_10001);
nand U17128 (N_17128,N_9492,N_10866);
nor U17129 (N_17129,N_9919,N_8987);
and U17130 (N_17130,N_11868,N_10943);
xor U17131 (N_17131,N_8762,N_10721);
xnor U17132 (N_17132,N_9907,N_11066);
xnor U17133 (N_17133,N_11923,N_11752);
and U17134 (N_17134,N_6408,N_6501);
nand U17135 (N_17135,N_6864,N_6811);
nor U17136 (N_17136,N_7360,N_9815);
nand U17137 (N_17137,N_8348,N_8942);
nor U17138 (N_17138,N_10096,N_11522);
xor U17139 (N_17139,N_6595,N_8258);
xnor U17140 (N_17140,N_6762,N_6882);
and U17141 (N_17141,N_9937,N_7538);
and U17142 (N_17142,N_11029,N_6114);
or U17143 (N_17143,N_9695,N_9040);
nand U17144 (N_17144,N_7393,N_11334);
nor U17145 (N_17145,N_7847,N_9823);
and U17146 (N_17146,N_7925,N_11016);
xnor U17147 (N_17147,N_8274,N_7064);
and U17148 (N_17148,N_9627,N_8600);
nand U17149 (N_17149,N_6298,N_7122);
nand U17150 (N_17150,N_11907,N_10907);
or U17151 (N_17151,N_10373,N_7309);
xor U17152 (N_17152,N_10474,N_10828);
nand U17153 (N_17153,N_7996,N_9949);
nor U17154 (N_17154,N_6153,N_8639);
xnor U17155 (N_17155,N_6673,N_11799);
or U17156 (N_17156,N_8760,N_7462);
or U17157 (N_17157,N_8656,N_11459);
or U17158 (N_17158,N_11440,N_8004);
nor U17159 (N_17159,N_8279,N_10699);
nor U17160 (N_17160,N_7948,N_6469);
and U17161 (N_17161,N_6051,N_10168);
nor U17162 (N_17162,N_8248,N_9818);
or U17163 (N_17163,N_11008,N_11601);
nor U17164 (N_17164,N_10930,N_8674);
xor U17165 (N_17165,N_9095,N_11179);
or U17166 (N_17166,N_11713,N_10496);
nand U17167 (N_17167,N_6499,N_9834);
nand U17168 (N_17168,N_9862,N_6724);
nand U17169 (N_17169,N_9815,N_9258);
nand U17170 (N_17170,N_6146,N_7588);
and U17171 (N_17171,N_11124,N_10097);
and U17172 (N_17172,N_9401,N_11362);
and U17173 (N_17173,N_8945,N_7927);
or U17174 (N_17174,N_9648,N_11866);
nand U17175 (N_17175,N_10289,N_6716);
or U17176 (N_17176,N_6443,N_8683);
nand U17177 (N_17177,N_9222,N_9675);
nor U17178 (N_17178,N_10941,N_6896);
and U17179 (N_17179,N_10479,N_6248);
nand U17180 (N_17180,N_6210,N_8063);
and U17181 (N_17181,N_6041,N_6152);
or U17182 (N_17182,N_7484,N_8507);
nor U17183 (N_17183,N_6233,N_9679);
or U17184 (N_17184,N_8659,N_10185);
xor U17185 (N_17185,N_6420,N_11506);
nand U17186 (N_17186,N_7658,N_10001);
nor U17187 (N_17187,N_9079,N_7411);
nor U17188 (N_17188,N_9152,N_11623);
nor U17189 (N_17189,N_6742,N_6482);
and U17190 (N_17190,N_7622,N_10529);
nor U17191 (N_17191,N_7743,N_7861);
xor U17192 (N_17192,N_8889,N_7359);
and U17193 (N_17193,N_10838,N_9284);
nand U17194 (N_17194,N_6616,N_6243);
xnor U17195 (N_17195,N_8144,N_7178);
and U17196 (N_17196,N_6481,N_7496);
xor U17197 (N_17197,N_11617,N_6585);
and U17198 (N_17198,N_11728,N_7359);
nor U17199 (N_17199,N_11587,N_10975);
nor U17200 (N_17200,N_11797,N_9803);
nand U17201 (N_17201,N_11840,N_6782);
nand U17202 (N_17202,N_6191,N_8575);
nand U17203 (N_17203,N_8111,N_10112);
and U17204 (N_17204,N_6431,N_8462);
nor U17205 (N_17205,N_10160,N_6708);
nand U17206 (N_17206,N_8575,N_11216);
or U17207 (N_17207,N_7964,N_8212);
nor U17208 (N_17208,N_6089,N_11955);
nand U17209 (N_17209,N_10165,N_10912);
or U17210 (N_17210,N_11462,N_11702);
nor U17211 (N_17211,N_6069,N_6616);
nand U17212 (N_17212,N_10660,N_7425);
nor U17213 (N_17213,N_10045,N_11134);
nand U17214 (N_17214,N_7077,N_6187);
xnor U17215 (N_17215,N_8880,N_10340);
xnor U17216 (N_17216,N_11975,N_6316);
nor U17217 (N_17217,N_9178,N_8776);
and U17218 (N_17218,N_10927,N_10095);
nor U17219 (N_17219,N_10659,N_10474);
nor U17220 (N_17220,N_9638,N_9827);
or U17221 (N_17221,N_8727,N_6685);
nand U17222 (N_17222,N_11944,N_11795);
xor U17223 (N_17223,N_7666,N_9983);
xnor U17224 (N_17224,N_10936,N_10956);
nor U17225 (N_17225,N_9101,N_11681);
or U17226 (N_17226,N_7676,N_11285);
or U17227 (N_17227,N_11238,N_7424);
and U17228 (N_17228,N_8761,N_9520);
nand U17229 (N_17229,N_8067,N_11150);
nand U17230 (N_17230,N_6027,N_11100);
nor U17231 (N_17231,N_7250,N_9050);
nand U17232 (N_17232,N_7644,N_10400);
and U17233 (N_17233,N_11250,N_9623);
or U17234 (N_17234,N_8766,N_11728);
and U17235 (N_17235,N_9403,N_11017);
nor U17236 (N_17236,N_10577,N_10060);
xnor U17237 (N_17237,N_11848,N_10112);
nand U17238 (N_17238,N_9219,N_10312);
nor U17239 (N_17239,N_9615,N_10369);
nand U17240 (N_17240,N_6229,N_11588);
nand U17241 (N_17241,N_8376,N_8201);
xnor U17242 (N_17242,N_6161,N_7085);
xor U17243 (N_17243,N_11683,N_8060);
xor U17244 (N_17244,N_11921,N_11725);
or U17245 (N_17245,N_7954,N_11150);
nor U17246 (N_17246,N_6431,N_9495);
xor U17247 (N_17247,N_6752,N_8660);
xor U17248 (N_17248,N_11066,N_10696);
nand U17249 (N_17249,N_11790,N_9469);
and U17250 (N_17250,N_6813,N_7050);
nor U17251 (N_17251,N_6684,N_9097);
and U17252 (N_17252,N_7908,N_7197);
nor U17253 (N_17253,N_10480,N_6533);
nand U17254 (N_17254,N_10315,N_11824);
nand U17255 (N_17255,N_6978,N_9024);
and U17256 (N_17256,N_7778,N_11724);
and U17257 (N_17257,N_6719,N_11649);
nor U17258 (N_17258,N_7759,N_7448);
or U17259 (N_17259,N_8329,N_8279);
nor U17260 (N_17260,N_6351,N_10105);
or U17261 (N_17261,N_8763,N_9989);
nor U17262 (N_17262,N_6028,N_11356);
xor U17263 (N_17263,N_9488,N_9256);
and U17264 (N_17264,N_11224,N_7532);
nor U17265 (N_17265,N_10994,N_7361);
or U17266 (N_17266,N_11188,N_7118);
nor U17267 (N_17267,N_10814,N_7498);
xnor U17268 (N_17268,N_11285,N_9851);
and U17269 (N_17269,N_9837,N_11594);
and U17270 (N_17270,N_7688,N_6966);
and U17271 (N_17271,N_6603,N_8331);
or U17272 (N_17272,N_6022,N_7085);
nor U17273 (N_17273,N_6997,N_10758);
nor U17274 (N_17274,N_11730,N_9591);
xnor U17275 (N_17275,N_6651,N_7079);
nand U17276 (N_17276,N_9232,N_8916);
nand U17277 (N_17277,N_8376,N_10530);
and U17278 (N_17278,N_10498,N_10154);
or U17279 (N_17279,N_6679,N_11836);
xor U17280 (N_17280,N_7842,N_9932);
nor U17281 (N_17281,N_6429,N_10985);
nor U17282 (N_17282,N_6912,N_7239);
nand U17283 (N_17283,N_10064,N_10262);
xnor U17284 (N_17284,N_9244,N_10832);
and U17285 (N_17285,N_10311,N_10085);
nand U17286 (N_17286,N_9157,N_11627);
or U17287 (N_17287,N_6701,N_9949);
nor U17288 (N_17288,N_8789,N_7126);
nor U17289 (N_17289,N_9908,N_8110);
nand U17290 (N_17290,N_9557,N_6505);
nand U17291 (N_17291,N_10328,N_9445);
or U17292 (N_17292,N_7114,N_6087);
or U17293 (N_17293,N_10609,N_8668);
xor U17294 (N_17294,N_6959,N_7700);
xor U17295 (N_17295,N_11994,N_6117);
xnor U17296 (N_17296,N_11193,N_9255);
nor U17297 (N_17297,N_8218,N_11601);
and U17298 (N_17298,N_7096,N_7060);
nand U17299 (N_17299,N_7985,N_7546);
xor U17300 (N_17300,N_6674,N_7346);
nor U17301 (N_17301,N_10955,N_6219);
and U17302 (N_17302,N_7936,N_6009);
and U17303 (N_17303,N_11631,N_6178);
and U17304 (N_17304,N_8845,N_10878);
xnor U17305 (N_17305,N_7652,N_7914);
and U17306 (N_17306,N_7047,N_11390);
xnor U17307 (N_17307,N_8237,N_7176);
and U17308 (N_17308,N_10189,N_7334);
xnor U17309 (N_17309,N_9679,N_9032);
or U17310 (N_17310,N_8703,N_9926);
or U17311 (N_17311,N_9485,N_10295);
or U17312 (N_17312,N_8634,N_8049);
and U17313 (N_17313,N_8376,N_10642);
or U17314 (N_17314,N_9712,N_11100);
xor U17315 (N_17315,N_10133,N_6163);
xor U17316 (N_17316,N_10979,N_6329);
xor U17317 (N_17317,N_11204,N_8599);
xor U17318 (N_17318,N_7913,N_9451);
nor U17319 (N_17319,N_9128,N_11218);
and U17320 (N_17320,N_6246,N_8914);
nand U17321 (N_17321,N_8484,N_11621);
or U17322 (N_17322,N_9607,N_8259);
or U17323 (N_17323,N_10003,N_9362);
or U17324 (N_17324,N_11477,N_8218);
or U17325 (N_17325,N_8002,N_8972);
xor U17326 (N_17326,N_9642,N_7754);
nor U17327 (N_17327,N_8677,N_8079);
xor U17328 (N_17328,N_8527,N_10105);
nand U17329 (N_17329,N_11269,N_6268);
xnor U17330 (N_17330,N_10352,N_7322);
nor U17331 (N_17331,N_10906,N_11004);
and U17332 (N_17332,N_9261,N_7614);
nand U17333 (N_17333,N_11193,N_7562);
nand U17334 (N_17334,N_7605,N_9619);
nor U17335 (N_17335,N_7998,N_10805);
nand U17336 (N_17336,N_11122,N_8496);
xor U17337 (N_17337,N_9736,N_6334);
xnor U17338 (N_17338,N_7324,N_10034);
nor U17339 (N_17339,N_8874,N_10026);
nand U17340 (N_17340,N_8267,N_11962);
nor U17341 (N_17341,N_11785,N_10977);
or U17342 (N_17342,N_10352,N_11613);
and U17343 (N_17343,N_8734,N_11216);
and U17344 (N_17344,N_6421,N_9838);
xnor U17345 (N_17345,N_8629,N_11607);
nor U17346 (N_17346,N_10839,N_8687);
or U17347 (N_17347,N_7670,N_11840);
nor U17348 (N_17348,N_8424,N_11937);
or U17349 (N_17349,N_7357,N_7067);
nand U17350 (N_17350,N_6883,N_6044);
and U17351 (N_17351,N_10322,N_6489);
nand U17352 (N_17352,N_6160,N_8480);
nor U17353 (N_17353,N_11300,N_10450);
nor U17354 (N_17354,N_6266,N_10843);
xor U17355 (N_17355,N_10442,N_10448);
and U17356 (N_17356,N_6013,N_8092);
xnor U17357 (N_17357,N_6992,N_6886);
and U17358 (N_17358,N_8006,N_10676);
nor U17359 (N_17359,N_6687,N_10946);
xor U17360 (N_17360,N_11359,N_11286);
and U17361 (N_17361,N_7663,N_8324);
xor U17362 (N_17362,N_9717,N_8635);
or U17363 (N_17363,N_11732,N_10865);
nor U17364 (N_17364,N_8081,N_10968);
and U17365 (N_17365,N_10212,N_7714);
nor U17366 (N_17366,N_6697,N_7135);
and U17367 (N_17367,N_7092,N_10189);
and U17368 (N_17368,N_7891,N_8229);
or U17369 (N_17369,N_7261,N_9147);
or U17370 (N_17370,N_11021,N_7384);
nand U17371 (N_17371,N_9362,N_9780);
or U17372 (N_17372,N_8204,N_7259);
or U17373 (N_17373,N_11859,N_11652);
xnor U17374 (N_17374,N_11048,N_11186);
and U17375 (N_17375,N_6904,N_9933);
nand U17376 (N_17376,N_9872,N_8261);
nor U17377 (N_17377,N_10326,N_6732);
or U17378 (N_17378,N_11431,N_10933);
nor U17379 (N_17379,N_11332,N_11279);
or U17380 (N_17380,N_11218,N_6634);
nand U17381 (N_17381,N_7034,N_10723);
nor U17382 (N_17382,N_11939,N_7453);
nand U17383 (N_17383,N_6369,N_10965);
xnor U17384 (N_17384,N_7939,N_10992);
and U17385 (N_17385,N_10931,N_6929);
nor U17386 (N_17386,N_9140,N_8503);
and U17387 (N_17387,N_8436,N_8527);
or U17388 (N_17388,N_8692,N_8680);
xnor U17389 (N_17389,N_9060,N_11619);
and U17390 (N_17390,N_10175,N_11661);
nand U17391 (N_17391,N_7717,N_10400);
and U17392 (N_17392,N_7654,N_8119);
nand U17393 (N_17393,N_9737,N_8210);
or U17394 (N_17394,N_9867,N_8467);
xor U17395 (N_17395,N_11054,N_8857);
nor U17396 (N_17396,N_7735,N_8496);
or U17397 (N_17397,N_10236,N_11058);
nor U17398 (N_17398,N_9553,N_6268);
nand U17399 (N_17399,N_9238,N_9951);
nand U17400 (N_17400,N_9865,N_10986);
or U17401 (N_17401,N_7900,N_10960);
xor U17402 (N_17402,N_10259,N_7140);
or U17403 (N_17403,N_6387,N_9319);
xnor U17404 (N_17404,N_10727,N_6637);
and U17405 (N_17405,N_9177,N_9514);
nand U17406 (N_17406,N_8494,N_7343);
and U17407 (N_17407,N_10181,N_9856);
nor U17408 (N_17408,N_11554,N_10481);
and U17409 (N_17409,N_10056,N_6027);
xnor U17410 (N_17410,N_7262,N_6049);
and U17411 (N_17411,N_8817,N_9993);
or U17412 (N_17412,N_10568,N_10722);
xor U17413 (N_17413,N_7109,N_10911);
nor U17414 (N_17414,N_11507,N_10687);
and U17415 (N_17415,N_7262,N_11711);
nor U17416 (N_17416,N_11960,N_10465);
nor U17417 (N_17417,N_11905,N_7310);
and U17418 (N_17418,N_10948,N_11280);
or U17419 (N_17419,N_9811,N_11363);
nand U17420 (N_17420,N_7415,N_7972);
nand U17421 (N_17421,N_11313,N_10166);
nand U17422 (N_17422,N_9349,N_9481);
or U17423 (N_17423,N_6603,N_11401);
xnor U17424 (N_17424,N_7272,N_7858);
nor U17425 (N_17425,N_7462,N_11049);
or U17426 (N_17426,N_11133,N_6035);
xor U17427 (N_17427,N_11130,N_10315);
and U17428 (N_17428,N_7627,N_10076);
nor U17429 (N_17429,N_6639,N_10531);
xor U17430 (N_17430,N_10828,N_11706);
nor U17431 (N_17431,N_11405,N_11249);
or U17432 (N_17432,N_8502,N_9379);
xor U17433 (N_17433,N_7889,N_7368);
or U17434 (N_17434,N_9088,N_7537);
xnor U17435 (N_17435,N_8616,N_11348);
and U17436 (N_17436,N_9160,N_8333);
or U17437 (N_17437,N_7927,N_9278);
xnor U17438 (N_17438,N_11300,N_7773);
nand U17439 (N_17439,N_10093,N_6401);
nor U17440 (N_17440,N_10329,N_7997);
and U17441 (N_17441,N_9140,N_11393);
xor U17442 (N_17442,N_6148,N_9536);
nor U17443 (N_17443,N_10281,N_6583);
xor U17444 (N_17444,N_7748,N_8478);
nand U17445 (N_17445,N_8733,N_10529);
or U17446 (N_17446,N_7210,N_11635);
or U17447 (N_17447,N_6403,N_8777);
or U17448 (N_17448,N_7310,N_10610);
and U17449 (N_17449,N_6067,N_10237);
nand U17450 (N_17450,N_9783,N_8445);
nor U17451 (N_17451,N_9530,N_7505);
or U17452 (N_17452,N_9306,N_10071);
nor U17453 (N_17453,N_6187,N_7913);
xor U17454 (N_17454,N_6937,N_10932);
xor U17455 (N_17455,N_6298,N_10424);
and U17456 (N_17456,N_10076,N_9614);
xnor U17457 (N_17457,N_6216,N_7400);
nand U17458 (N_17458,N_7437,N_6154);
or U17459 (N_17459,N_8591,N_6582);
or U17460 (N_17460,N_9901,N_10239);
or U17461 (N_17461,N_8547,N_7544);
and U17462 (N_17462,N_7006,N_8614);
and U17463 (N_17463,N_11692,N_11502);
xor U17464 (N_17464,N_11717,N_8696);
nor U17465 (N_17465,N_10537,N_9715);
nor U17466 (N_17466,N_11776,N_7936);
and U17467 (N_17467,N_11843,N_9935);
nor U17468 (N_17468,N_7927,N_7990);
and U17469 (N_17469,N_9868,N_7112);
and U17470 (N_17470,N_11242,N_9631);
nor U17471 (N_17471,N_11688,N_11670);
xor U17472 (N_17472,N_8477,N_8210);
xor U17473 (N_17473,N_8936,N_7919);
and U17474 (N_17474,N_11526,N_11759);
and U17475 (N_17475,N_7440,N_8164);
or U17476 (N_17476,N_10075,N_6895);
or U17477 (N_17477,N_6381,N_9980);
nor U17478 (N_17478,N_11618,N_10557);
and U17479 (N_17479,N_10481,N_9719);
or U17480 (N_17480,N_10022,N_9988);
or U17481 (N_17481,N_8631,N_8697);
or U17482 (N_17482,N_6828,N_6380);
and U17483 (N_17483,N_11207,N_9269);
and U17484 (N_17484,N_6943,N_9089);
or U17485 (N_17485,N_7039,N_8593);
xnor U17486 (N_17486,N_6951,N_8362);
nor U17487 (N_17487,N_8562,N_9239);
xor U17488 (N_17488,N_10490,N_7973);
nor U17489 (N_17489,N_9865,N_11907);
and U17490 (N_17490,N_6248,N_8877);
nand U17491 (N_17491,N_10422,N_10262);
nor U17492 (N_17492,N_9184,N_9328);
and U17493 (N_17493,N_8088,N_10589);
and U17494 (N_17494,N_8911,N_8874);
nor U17495 (N_17495,N_11729,N_7106);
nor U17496 (N_17496,N_6442,N_11740);
nand U17497 (N_17497,N_9144,N_9050);
or U17498 (N_17498,N_8188,N_10859);
nor U17499 (N_17499,N_11578,N_10644);
xnor U17500 (N_17500,N_8870,N_6709);
and U17501 (N_17501,N_7125,N_7899);
or U17502 (N_17502,N_10916,N_9093);
and U17503 (N_17503,N_8711,N_11845);
or U17504 (N_17504,N_11261,N_8022);
nor U17505 (N_17505,N_7838,N_11428);
or U17506 (N_17506,N_10703,N_7745);
nand U17507 (N_17507,N_9485,N_7865);
or U17508 (N_17508,N_8914,N_11245);
and U17509 (N_17509,N_9032,N_6824);
nand U17510 (N_17510,N_8486,N_9402);
nand U17511 (N_17511,N_10749,N_7104);
nor U17512 (N_17512,N_7761,N_8973);
nor U17513 (N_17513,N_9042,N_6874);
nand U17514 (N_17514,N_9101,N_9358);
nor U17515 (N_17515,N_6078,N_9799);
or U17516 (N_17516,N_10020,N_8112);
xnor U17517 (N_17517,N_10147,N_8477);
xnor U17518 (N_17518,N_11905,N_8121);
or U17519 (N_17519,N_7595,N_8840);
or U17520 (N_17520,N_11319,N_10072);
and U17521 (N_17521,N_6111,N_11543);
xor U17522 (N_17522,N_8331,N_6346);
and U17523 (N_17523,N_10815,N_10093);
nand U17524 (N_17524,N_11906,N_9901);
and U17525 (N_17525,N_9748,N_10828);
nand U17526 (N_17526,N_9759,N_6249);
or U17527 (N_17527,N_8095,N_9143);
and U17528 (N_17528,N_9589,N_7294);
xnor U17529 (N_17529,N_10083,N_6907);
or U17530 (N_17530,N_10478,N_6079);
nand U17531 (N_17531,N_7308,N_6881);
nor U17532 (N_17532,N_10889,N_7034);
xor U17533 (N_17533,N_6761,N_6901);
nor U17534 (N_17534,N_10793,N_8627);
and U17535 (N_17535,N_9524,N_7613);
xor U17536 (N_17536,N_9330,N_7653);
nand U17537 (N_17537,N_6593,N_9710);
nor U17538 (N_17538,N_8984,N_7864);
xor U17539 (N_17539,N_9119,N_7198);
and U17540 (N_17540,N_11642,N_8894);
xor U17541 (N_17541,N_11828,N_7493);
nor U17542 (N_17542,N_6352,N_8196);
nor U17543 (N_17543,N_10229,N_6267);
nor U17544 (N_17544,N_10818,N_7140);
nand U17545 (N_17545,N_6184,N_8306);
and U17546 (N_17546,N_11943,N_8668);
xnor U17547 (N_17547,N_10898,N_7004);
nor U17548 (N_17548,N_10397,N_10725);
and U17549 (N_17549,N_8158,N_8470);
and U17550 (N_17550,N_11689,N_6638);
and U17551 (N_17551,N_9437,N_6036);
or U17552 (N_17552,N_10180,N_9676);
nand U17553 (N_17553,N_7462,N_6879);
or U17554 (N_17554,N_7970,N_10812);
nor U17555 (N_17555,N_9215,N_8452);
or U17556 (N_17556,N_8986,N_7844);
and U17557 (N_17557,N_9278,N_6732);
nor U17558 (N_17558,N_6950,N_7331);
nor U17559 (N_17559,N_10753,N_11486);
nand U17560 (N_17560,N_6485,N_8725);
nor U17561 (N_17561,N_10777,N_10805);
nor U17562 (N_17562,N_9626,N_8572);
nand U17563 (N_17563,N_7835,N_11253);
xor U17564 (N_17564,N_10622,N_7870);
xnor U17565 (N_17565,N_9915,N_7197);
nand U17566 (N_17566,N_11452,N_6834);
xor U17567 (N_17567,N_11923,N_11305);
nand U17568 (N_17568,N_11588,N_9667);
nand U17569 (N_17569,N_11613,N_7321);
xnor U17570 (N_17570,N_6040,N_7929);
and U17571 (N_17571,N_8108,N_9126);
or U17572 (N_17572,N_6437,N_8095);
and U17573 (N_17573,N_7639,N_11724);
xor U17574 (N_17574,N_8378,N_10643);
nor U17575 (N_17575,N_6475,N_11113);
nand U17576 (N_17576,N_11136,N_11158);
and U17577 (N_17577,N_8274,N_7372);
and U17578 (N_17578,N_6182,N_6886);
or U17579 (N_17579,N_11535,N_11303);
and U17580 (N_17580,N_9688,N_6394);
nor U17581 (N_17581,N_10250,N_8719);
nand U17582 (N_17582,N_6093,N_8109);
nand U17583 (N_17583,N_10032,N_9671);
or U17584 (N_17584,N_10033,N_11489);
or U17585 (N_17585,N_7294,N_11056);
xnor U17586 (N_17586,N_11692,N_11390);
xnor U17587 (N_17587,N_7630,N_11410);
xor U17588 (N_17588,N_7698,N_9036);
and U17589 (N_17589,N_7845,N_8937);
nand U17590 (N_17590,N_10547,N_6359);
or U17591 (N_17591,N_6305,N_8725);
nand U17592 (N_17592,N_10757,N_6426);
nand U17593 (N_17593,N_6332,N_6067);
or U17594 (N_17594,N_10842,N_11706);
and U17595 (N_17595,N_11911,N_11813);
and U17596 (N_17596,N_10791,N_8928);
nand U17597 (N_17597,N_8632,N_8166);
and U17598 (N_17598,N_7134,N_6407);
xnor U17599 (N_17599,N_8474,N_9836);
or U17600 (N_17600,N_11296,N_6255);
and U17601 (N_17601,N_6579,N_10952);
and U17602 (N_17602,N_8749,N_8707);
xnor U17603 (N_17603,N_8424,N_8561);
and U17604 (N_17604,N_7537,N_6905);
nor U17605 (N_17605,N_7661,N_11651);
or U17606 (N_17606,N_11048,N_11461);
and U17607 (N_17607,N_7649,N_6386);
nand U17608 (N_17608,N_11052,N_10308);
or U17609 (N_17609,N_6122,N_9619);
nand U17610 (N_17610,N_7981,N_11229);
nand U17611 (N_17611,N_11519,N_7302);
nand U17612 (N_17612,N_9801,N_10318);
nand U17613 (N_17613,N_6818,N_6591);
or U17614 (N_17614,N_7697,N_8209);
and U17615 (N_17615,N_10532,N_11791);
or U17616 (N_17616,N_8694,N_8561);
nand U17617 (N_17617,N_9654,N_7201);
and U17618 (N_17618,N_11075,N_9465);
nor U17619 (N_17619,N_10748,N_9545);
nand U17620 (N_17620,N_7133,N_10612);
nand U17621 (N_17621,N_7178,N_11779);
or U17622 (N_17622,N_7949,N_6500);
nand U17623 (N_17623,N_8211,N_8980);
or U17624 (N_17624,N_8271,N_7149);
and U17625 (N_17625,N_8152,N_11317);
nor U17626 (N_17626,N_10806,N_6858);
xor U17627 (N_17627,N_8081,N_11425);
nand U17628 (N_17628,N_9630,N_9790);
and U17629 (N_17629,N_11686,N_11189);
nor U17630 (N_17630,N_9760,N_10287);
xor U17631 (N_17631,N_8929,N_10062);
xor U17632 (N_17632,N_6951,N_11498);
xor U17633 (N_17633,N_11575,N_11976);
or U17634 (N_17634,N_8270,N_10070);
and U17635 (N_17635,N_11791,N_8545);
nand U17636 (N_17636,N_7019,N_9443);
nand U17637 (N_17637,N_6099,N_9513);
nand U17638 (N_17638,N_11825,N_6800);
or U17639 (N_17639,N_11380,N_10026);
and U17640 (N_17640,N_10146,N_11184);
nand U17641 (N_17641,N_11210,N_8065);
or U17642 (N_17642,N_6460,N_11249);
and U17643 (N_17643,N_7932,N_11001);
nor U17644 (N_17644,N_7987,N_10049);
and U17645 (N_17645,N_8139,N_7617);
xor U17646 (N_17646,N_6208,N_11932);
nor U17647 (N_17647,N_10686,N_11547);
nor U17648 (N_17648,N_11570,N_10167);
xor U17649 (N_17649,N_8611,N_6709);
nand U17650 (N_17650,N_9397,N_6819);
nor U17651 (N_17651,N_11670,N_7577);
or U17652 (N_17652,N_7205,N_11152);
nor U17653 (N_17653,N_9170,N_6712);
and U17654 (N_17654,N_10743,N_10448);
or U17655 (N_17655,N_6519,N_9959);
xor U17656 (N_17656,N_6715,N_10332);
and U17657 (N_17657,N_9247,N_6375);
xor U17658 (N_17658,N_10398,N_6670);
nor U17659 (N_17659,N_11608,N_6332);
xor U17660 (N_17660,N_7698,N_7198);
nand U17661 (N_17661,N_8857,N_7945);
nand U17662 (N_17662,N_7709,N_6423);
or U17663 (N_17663,N_8697,N_11884);
xor U17664 (N_17664,N_6093,N_8430);
xor U17665 (N_17665,N_10769,N_9823);
nor U17666 (N_17666,N_8746,N_6306);
nor U17667 (N_17667,N_8770,N_11862);
nand U17668 (N_17668,N_9196,N_9548);
nor U17669 (N_17669,N_10031,N_8683);
nor U17670 (N_17670,N_7828,N_7173);
nor U17671 (N_17671,N_10736,N_10900);
nand U17672 (N_17672,N_10014,N_6399);
and U17673 (N_17673,N_10849,N_9952);
and U17674 (N_17674,N_11334,N_8619);
nor U17675 (N_17675,N_8662,N_7074);
or U17676 (N_17676,N_9032,N_8785);
or U17677 (N_17677,N_7623,N_9380);
xnor U17678 (N_17678,N_6010,N_7953);
or U17679 (N_17679,N_10904,N_8113);
nand U17680 (N_17680,N_6021,N_7034);
and U17681 (N_17681,N_10315,N_10865);
nand U17682 (N_17682,N_8339,N_10460);
and U17683 (N_17683,N_7167,N_6016);
nand U17684 (N_17684,N_10003,N_8535);
or U17685 (N_17685,N_7885,N_6750);
nand U17686 (N_17686,N_10338,N_9963);
nor U17687 (N_17687,N_7039,N_6877);
nor U17688 (N_17688,N_7339,N_8074);
or U17689 (N_17689,N_6184,N_11070);
or U17690 (N_17690,N_6818,N_8904);
xor U17691 (N_17691,N_10255,N_6552);
and U17692 (N_17692,N_10345,N_6733);
xnor U17693 (N_17693,N_9981,N_10381);
and U17694 (N_17694,N_6007,N_7712);
nor U17695 (N_17695,N_10022,N_7072);
nand U17696 (N_17696,N_7675,N_11611);
nand U17697 (N_17697,N_7542,N_9392);
or U17698 (N_17698,N_6232,N_7411);
nand U17699 (N_17699,N_11405,N_7885);
nor U17700 (N_17700,N_9974,N_8047);
xor U17701 (N_17701,N_8643,N_9668);
nor U17702 (N_17702,N_6216,N_7000);
xnor U17703 (N_17703,N_6386,N_6227);
xor U17704 (N_17704,N_7928,N_11499);
nand U17705 (N_17705,N_7263,N_11005);
and U17706 (N_17706,N_10421,N_9726);
or U17707 (N_17707,N_9010,N_8057);
xor U17708 (N_17708,N_10730,N_9322);
xnor U17709 (N_17709,N_9329,N_11629);
or U17710 (N_17710,N_9097,N_8309);
and U17711 (N_17711,N_6948,N_11221);
and U17712 (N_17712,N_7027,N_11640);
xnor U17713 (N_17713,N_11662,N_10228);
or U17714 (N_17714,N_7057,N_6395);
nor U17715 (N_17715,N_11618,N_11590);
or U17716 (N_17716,N_6023,N_9633);
and U17717 (N_17717,N_7288,N_10676);
nand U17718 (N_17718,N_7459,N_6575);
nor U17719 (N_17719,N_11765,N_8035);
or U17720 (N_17720,N_6153,N_6423);
xor U17721 (N_17721,N_11141,N_6972);
xor U17722 (N_17722,N_9949,N_10470);
and U17723 (N_17723,N_6887,N_6000);
xor U17724 (N_17724,N_10411,N_7421);
nand U17725 (N_17725,N_6869,N_9923);
nor U17726 (N_17726,N_8136,N_11959);
or U17727 (N_17727,N_8950,N_10184);
xor U17728 (N_17728,N_9466,N_8840);
xnor U17729 (N_17729,N_6622,N_9988);
xnor U17730 (N_17730,N_6141,N_9851);
nand U17731 (N_17731,N_7328,N_11281);
nand U17732 (N_17732,N_9561,N_11179);
or U17733 (N_17733,N_10199,N_11427);
or U17734 (N_17734,N_6744,N_9992);
nor U17735 (N_17735,N_8187,N_9051);
or U17736 (N_17736,N_11699,N_6303);
or U17737 (N_17737,N_9988,N_9354);
or U17738 (N_17738,N_11347,N_9477);
nand U17739 (N_17739,N_6506,N_7845);
xnor U17740 (N_17740,N_6506,N_10516);
nor U17741 (N_17741,N_8331,N_10023);
xnor U17742 (N_17742,N_7146,N_6991);
nor U17743 (N_17743,N_8220,N_8789);
nand U17744 (N_17744,N_10445,N_10151);
or U17745 (N_17745,N_8947,N_8465);
nand U17746 (N_17746,N_8093,N_6803);
xnor U17747 (N_17747,N_8934,N_9384);
and U17748 (N_17748,N_10739,N_7746);
nor U17749 (N_17749,N_6622,N_6510);
xor U17750 (N_17750,N_7160,N_10621);
and U17751 (N_17751,N_9339,N_7121);
nor U17752 (N_17752,N_6048,N_6263);
nand U17753 (N_17753,N_9035,N_6216);
and U17754 (N_17754,N_8338,N_7140);
xor U17755 (N_17755,N_6422,N_11248);
nand U17756 (N_17756,N_9450,N_8501);
and U17757 (N_17757,N_6690,N_11204);
nand U17758 (N_17758,N_10083,N_10017);
nor U17759 (N_17759,N_8289,N_6670);
nand U17760 (N_17760,N_8732,N_9508);
xnor U17761 (N_17761,N_6375,N_6967);
or U17762 (N_17762,N_10364,N_11386);
nor U17763 (N_17763,N_9385,N_10319);
and U17764 (N_17764,N_11292,N_10162);
nor U17765 (N_17765,N_8660,N_6008);
or U17766 (N_17766,N_10176,N_7451);
xor U17767 (N_17767,N_11518,N_6792);
nand U17768 (N_17768,N_6638,N_11471);
nor U17769 (N_17769,N_7945,N_8565);
nor U17770 (N_17770,N_7957,N_9886);
xor U17771 (N_17771,N_9410,N_10420);
nor U17772 (N_17772,N_11833,N_6291);
nor U17773 (N_17773,N_7634,N_6854);
and U17774 (N_17774,N_6866,N_7228);
or U17775 (N_17775,N_10881,N_9621);
xnor U17776 (N_17776,N_9469,N_6663);
or U17777 (N_17777,N_11781,N_8321);
or U17778 (N_17778,N_10778,N_9174);
or U17779 (N_17779,N_8735,N_10231);
nand U17780 (N_17780,N_10455,N_10676);
nand U17781 (N_17781,N_8449,N_7222);
or U17782 (N_17782,N_11864,N_11390);
xor U17783 (N_17783,N_6233,N_10040);
xor U17784 (N_17784,N_9016,N_6861);
or U17785 (N_17785,N_7906,N_11306);
nand U17786 (N_17786,N_11578,N_11306);
and U17787 (N_17787,N_9956,N_11524);
nor U17788 (N_17788,N_11229,N_8132);
xor U17789 (N_17789,N_10049,N_6083);
nand U17790 (N_17790,N_7882,N_11479);
nand U17791 (N_17791,N_7680,N_10584);
nor U17792 (N_17792,N_6981,N_6357);
xor U17793 (N_17793,N_8774,N_10255);
nor U17794 (N_17794,N_8808,N_7017);
or U17795 (N_17795,N_6065,N_7798);
nand U17796 (N_17796,N_7324,N_10808);
nor U17797 (N_17797,N_6873,N_11770);
or U17798 (N_17798,N_9387,N_8660);
nand U17799 (N_17799,N_7740,N_11271);
nand U17800 (N_17800,N_7689,N_11718);
or U17801 (N_17801,N_9831,N_10354);
nand U17802 (N_17802,N_9750,N_10392);
nand U17803 (N_17803,N_7583,N_7098);
and U17804 (N_17804,N_11386,N_6571);
xor U17805 (N_17805,N_9968,N_8804);
nand U17806 (N_17806,N_9097,N_8809);
or U17807 (N_17807,N_8296,N_10251);
xor U17808 (N_17808,N_6846,N_7830);
nor U17809 (N_17809,N_6206,N_11271);
nand U17810 (N_17810,N_7029,N_8172);
or U17811 (N_17811,N_8152,N_10673);
nor U17812 (N_17812,N_6330,N_10223);
nand U17813 (N_17813,N_10959,N_7042);
or U17814 (N_17814,N_9776,N_10061);
or U17815 (N_17815,N_8004,N_8611);
xor U17816 (N_17816,N_9074,N_11404);
xnor U17817 (N_17817,N_9895,N_7689);
nor U17818 (N_17818,N_10017,N_10923);
nor U17819 (N_17819,N_6814,N_11850);
nor U17820 (N_17820,N_8911,N_10170);
and U17821 (N_17821,N_8558,N_6284);
and U17822 (N_17822,N_7686,N_8998);
nand U17823 (N_17823,N_9957,N_11257);
nand U17824 (N_17824,N_11942,N_11082);
nor U17825 (N_17825,N_10457,N_11943);
and U17826 (N_17826,N_7850,N_8339);
and U17827 (N_17827,N_9851,N_8452);
nand U17828 (N_17828,N_6818,N_9110);
nand U17829 (N_17829,N_7310,N_6400);
and U17830 (N_17830,N_11654,N_6267);
or U17831 (N_17831,N_7793,N_11190);
and U17832 (N_17832,N_6719,N_6881);
nor U17833 (N_17833,N_7307,N_9752);
nor U17834 (N_17834,N_8107,N_7887);
nand U17835 (N_17835,N_10159,N_8684);
and U17836 (N_17836,N_7004,N_6977);
nand U17837 (N_17837,N_9717,N_11526);
and U17838 (N_17838,N_9465,N_7787);
or U17839 (N_17839,N_10957,N_7625);
or U17840 (N_17840,N_11143,N_10882);
nor U17841 (N_17841,N_9613,N_11778);
nand U17842 (N_17842,N_9636,N_8304);
or U17843 (N_17843,N_10215,N_7113);
or U17844 (N_17844,N_6243,N_8919);
xor U17845 (N_17845,N_7715,N_11812);
or U17846 (N_17846,N_6055,N_7189);
nand U17847 (N_17847,N_7505,N_11995);
or U17848 (N_17848,N_9236,N_11837);
and U17849 (N_17849,N_9160,N_9880);
xor U17850 (N_17850,N_8763,N_8909);
or U17851 (N_17851,N_7287,N_10119);
xnor U17852 (N_17852,N_10474,N_11092);
or U17853 (N_17853,N_7985,N_9502);
nor U17854 (N_17854,N_11799,N_9914);
nand U17855 (N_17855,N_10386,N_7391);
nand U17856 (N_17856,N_8440,N_10049);
and U17857 (N_17857,N_9583,N_8031);
or U17858 (N_17858,N_11933,N_8157);
nand U17859 (N_17859,N_7805,N_8982);
and U17860 (N_17860,N_8364,N_9536);
nor U17861 (N_17861,N_10741,N_10075);
or U17862 (N_17862,N_8765,N_6224);
xnor U17863 (N_17863,N_10865,N_11387);
and U17864 (N_17864,N_7410,N_7090);
nand U17865 (N_17865,N_9562,N_8277);
nand U17866 (N_17866,N_6668,N_6664);
and U17867 (N_17867,N_7658,N_6884);
and U17868 (N_17868,N_6431,N_8623);
nand U17869 (N_17869,N_11288,N_11297);
nor U17870 (N_17870,N_10660,N_8987);
xnor U17871 (N_17871,N_6312,N_9806);
nand U17872 (N_17872,N_7966,N_8889);
or U17873 (N_17873,N_10295,N_9802);
xor U17874 (N_17874,N_7257,N_8996);
and U17875 (N_17875,N_8129,N_7570);
xnor U17876 (N_17876,N_11052,N_6798);
nand U17877 (N_17877,N_6676,N_9915);
nor U17878 (N_17878,N_7603,N_10856);
xor U17879 (N_17879,N_7205,N_7855);
or U17880 (N_17880,N_11722,N_9517);
or U17881 (N_17881,N_9605,N_9593);
nand U17882 (N_17882,N_8248,N_7925);
nand U17883 (N_17883,N_10948,N_9647);
xor U17884 (N_17884,N_6364,N_7760);
xor U17885 (N_17885,N_8189,N_7190);
and U17886 (N_17886,N_11675,N_11790);
nand U17887 (N_17887,N_10126,N_11197);
xnor U17888 (N_17888,N_7851,N_6020);
or U17889 (N_17889,N_9926,N_9814);
or U17890 (N_17890,N_10128,N_8520);
xnor U17891 (N_17891,N_6157,N_6290);
or U17892 (N_17892,N_8049,N_7059);
xnor U17893 (N_17893,N_9379,N_11353);
and U17894 (N_17894,N_11199,N_8705);
and U17895 (N_17895,N_7650,N_7504);
or U17896 (N_17896,N_9317,N_8532);
xnor U17897 (N_17897,N_9016,N_10706);
xnor U17898 (N_17898,N_6495,N_7099);
nand U17899 (N_17899,N_9517,N_9913);
and U17900 (N_17900,N_6102,N_9468);
and U17901 (N_17901,N_10616,N_9150);
nand U17902 (N_17902,N_10380,N_8295);
nand U17903 (N_17903,N_10405,N_10711);
nor U17904 (N_17904,N_7197,N_8730);
nand U17905 (N_17905,N_7322,N_8908);
nand U17906 (N_17906,N_7847,N_9683);
xor U17907 (N_17907,N_8774,N_10946);
or U17908 (N_17908,N_11155,N_9592);
nand U17909 (N_17909,N_10931,N_7192);
nand U17910 (N_17910,N_9302,N_10729);
and U17911 (N_17911,N_9164,N_9136);
or U17912 (N_17912,N_7094,N_11521);
and U17913 (N_17913,N_7260,N_7852);
nor U17914 (N_17914,N_11429,N_7026);
or U17915 (N_17915,N_6867,N_6687);
xnor U17916 (N_17916,N_7747,N_10345);
nor U17917 (N_17917,N_7130,N_10303);
nor U17918 (N_17918,N_7920,N_9705);
or U17919 (N_17919,N_6582,N_7021);
or U17920 (N_17920,N_9661,N_7256);
nor U17921 (N_17921,N_7059,N_9010);
and U17922 (N_17922,N_8827,N_8768);
xnor U17923 (N_17923,N_7337,N_7341);
nand U17924 (N_17924,N_9266,N_6438);
xor U17925 (N_17925,N_10745,N_9847);
nand U17926 (N_17926,N_7740,N_9532);
nor U17927 (N_17927,N_7011,N_9806);
nor U17928 (N_17928,N_8397,N_10399);
and U17929 (N_17929,N_11724,N_8931);
nand U17930 (N_17930,N_7990,N_6776);
nor U17931 (N_17931,N_10526,N_7517);
and U17932 (N_17932,N_10733,N_6554);
nor U17933 (N_17933,N_9227,N_7594);
and U17934 (N_17934,N_8204,N_8856);
xnor U17935 (N_17935,N_6945,N_9788);
and U17936 (N_17936,N_11753,N_6041);
xnor U17937 (N_17937,N_7299,N_11351);
and U17938 (N_17938,N_8912,N_10998);
xor U17939 (N_17939,N_7825,N_9646);
or U17940 (N_17940,N_6129,N_7347);
nand U17941 (N_17941,N_7004,N_9497);
or U17942 (N_17942,N_6182,N_8278);
or U17943 (N_17943,N_6292,N_6977);
nor U17944 (N_17944,N_10548,N_6253);
nor U17945 (N_17945,N_7769,N_8160);
and U17946 (N_17946,N_6950,N_6514);
nor U17947 (N_17947,N_11102,N_8787);
and U17948 (N_17948,N_10484,N_6465);
and U17949 (N_17949,N_9827,N_8006);
nand U17950 (N_17950,N_10872,N_7672);
or U17951 (N_17951,N_8149,N_10362);
or U17952 (N_17952,N_7572,N_6874);
nand U17953 (N_17953,N_9816,N_8343);
xnor U17954 (N_17954,N_9804,N_9258);
nand U17955 (N_17955,N_10268,N_7299);
xnor U17956 (N_17956,N_10977,N_8743);
or U17957 (N_17957,N_7347,N_7915);
nand U17958 (N_17958,N_8476,N_10963);
xnor U17959 (N_17959,N_9434,N_9337);
nand U17960 (N_17960,N_11339,N_6900);
nor U17961 (N_17961,N_11215,N_10664);
xor U17962 (N_17962,N_9550,N_11439);
or U17963 (N_17963,N_10741,N_11847);
nand U17964 (N_17964,N_7666,N_9833);
xnor U17965 (N_17965,N_11749,N_10501);
xor U17966 (N_17966,N_8076,N_9653);
or U17967 (N_17967,N_9803,N_6409);
and U17968 (N_17968,N_8281,N_11072);
or U17969 (N_17969,N_6629,N_10814);
nand U17970 (N_17970,N_6555,N_9351);
and U17971 (N_17971,N_6605,N_8994);
or U17972 (N_17972,N_10264,N_11875);
or U17973 (N_17973,N_7377,N_6486);
xor U17974 (N_17974,N_7629,N_6033);
nand U17975 (N_17975,N_7233,N_6802);
xor U17976 (N_17976,N_11765,N_11712);
nor U17977 (N_17977,N_10905,N_11057);
nand U17978 (N_17978,N_11425,N_6612);
nor U17979 (N_17979,N_9432,N_9645);
nor U17980 (N_17980,N_6242,N_9554);
and U17981 (N_17981,N_9402,N_6764);
and U17982 (N_17982,N_11805,N_8600);
nor U17983 (N_17983,N_10757,N_10340);
or U17984 (N_17984,N_8055,N_6058);
or U17985 (N_17985,N_6517,N_7732);
nor U17986 (N_17986,N_10283,N_11443);
and U17987 (N_17987,N_11388,N_9219);
and U17988 (N_17988,N_7232,N_6890);
nand U17989 (N_17989,N_8448,N_7052);
nand U17990 (N_17990,N_10841,N_11164);
nor U17991 (N_17991,N_6529,N_6743);
xor U17992 (N_17992,N_10744,N_9820);
xnor U17993 (N_17993,N_6544,N_8260);
xor U17994 (N_17994,N_10623,N_10601);
and U17995 (N_17995,N_6477,N_7767);
nor U17996 (N_17996,N_9860,N_11798);
xnor U17997 (N_17997,N_7990,N_7021);
nand U17998 (N_17998,N_11035,N_11134);
nand U17999 (N_17999,N_9899,N_10788);
nand U18000 (N_18000,N_16515,N_14874);
or U18001 (N_18001,N_13929,N_13877);
or U18002 (N_18002,N_16207,N_12848);
and U18003 (N_18003,N_16892,N_17938);
or U18004 (N_18004,N_13563,N_15695);
and U18005 (N_18005,N_15023,N_12839);
or U18006 (N_18006,N_14349,N_12739);
and U18007 (N_18007,N_13984,N_13123);
xor U18008 (N_18008,N_16930,N_17612);
and U18009 (N_18009,N_15222,N_14353);
or U18010 (N_18010,N_15152,N_15322);
nor U18011 (N_18011,N_12225,N_14794);
nor U18012 (N_18012,N_17196,N_14455);
nand U18013 (N_18013,N_14020,N_13257);
nor U18014 (N_18014,N_15821,N_16422);
nor U18015 (N_18015,N_14148,N_17897);
and U18016 (N_18016,N_14476,N_13934);
or U18017 (N_18017,N_12632,N_17604);
and U18018 (N_18018,N_14611,N_15318);
nand U18019 (N_18019,N_12933,N_13760);
and U18020 (N_18020,N_15382,N_14069);
or U18021 (N_18021,N_15301,N_12069);
and U18022 (N_18022,N_15334,N_13048);
and U18023 (N_18023,N_15542,N_13698);
nor U18024 (N_18024,N_17499,N_12418);
nor U18025 (N_18025,N_14593,N_14764);
xnor U18026 (N_18026,N_13358,N_15656);
nor U18027 (N_18027,N_16474,N_14809);
or U18028 (N_18028,N_14831,N_14294);
xnor U18029 (N_18029,N_17219,N_14852);
or U18030 (N_18030,N_13221,N_17703);
and U18031 (N_18031,N_15872,N_13819);
nor U18032 (N_18032,N_14670,N_15108);
xnor U18033 (N_18033,N_16224,N_14286);
xnor U18034 (N_18034,N_16925,N_16926);
or U18035 (N_18035,N_12108,N_16723);
or U18036 (N_18036,N_16480,N_16022);
xnor U18037 (N_18037,N_14782,N_16917);
and U18038 (N_18038,N_14696,N_16722);
xnor U18039 (N_18039,N_17632,N_13711);
and U18040 (N_18040,N_14521,N_15845);
nor U18041 (N_18041,N_14109,N_13979);
or U18042 (N_18042,N_14959,N_12858);
nor U18043 (N_18043,N_16913,N_16962);
and U18044 (N_18044,N_15983,N_17177);
or U18045 (N_18045,N_13655,N_14759);
nand U18046 (N_18046,N_15809,N_17186);
xor U18047 (N_18047,N_13443,N_17116);
or U18048 (N_18048,N_13441,N_12039);
xnor U18049 (N_18049,N_14549,N_17029);
nor U18050 (N_18050,N_17560,N_17583);
nor U18051 (N_18051,N_13611,N_16904);
nor U18052 (N_18052,N_14305,N_12977);
nand U18053 (N_18053,N_17137,N_14538);
nand U18054 (N_18054,N_17071,N_12321);
and U18055 (N_18055,N_15097,N_16237);
nand U18056 (N_18056,N_16487,N_14369);
nor U18057 (N_18057,N_17793,N_13779);
and U18058 (N_18058,N_14957,N_17153);
and U18059 (N_18059,N_12426,N_17496);
nor U18060 (N_18060,N_17718,N_17566);
and U18061 (N_18061,N_15618,N_15008);
xor U18062 (N_18062,N_17441,N_14882);
or U18063 (N_18063,N_14456,N_14773);
or U18064 (N_18064,N_13890,N_17143);
or U18065 (N_18065,N_14102,N_16510);
nor U18066 (N_18066,N_17643,N_13697);
nand U18067 (N_18067,N_16358,N_15242);
nor U18068 (N_18068,N_16730,N_16159);
and U18069 (N_18069,N_17966,N_12946);
and U18070 (N_18070,N_12608,N_16486);
or U18071 (N_18071,N_13116,N_12573);
nand U18072 (N_18072,N_16441,N_15364);
and U18073 (N_18073,N_17320,N_14560);
and U18074 (N_18074,N_12432,N_16184);
xnor U18075 (N_18075,N_17843,N_13456);
xnor U18076 (N_18076,N_16535,N_14311);
and U18077 (N_18077,N_15011,N_16217);
or U18078 (N_18078,N_15748,N_15466);
xor U18079 (N_18079,N_14139,N_16720);
nand U18080 (N_18080,N_16269,N_17809);
nand U18081 (N_18081,N_12835,N_13097);
nand U18082 (N_18082,N_14693,N_15243);
xnor U18083 (N_18083,N_13861,N_15250);
nor U18084 (N_18084,N_15615,N_13936);
nand U18085 (N_18085,N_14106,N_16130);
or U18086 (N_18086,N_13685,N_17651);
nor U18087 (N_18087,N_13504,N_17538);
nor U18088 (N_18088,N_16307,N_14453);
or U18089 (N_18089,N_15248,N_16910);
and U18090 (N_18090,N_13293,N_14376);
nand U18091 (N_18091,N_15525,N_16178);
nand U18092 (N_18092,N_13163,N_13206);
xor U18093 (N_18093,N_17865,N_13536);
and U18094 (N_18094,N_14184,N_15978);
xnor U18095 (N_18095,N_14884,N_13383);
nor U18096 (N_18096,N_13876,N_16861);
xor U18097 (N_18097,N_13962,N_16411);
xnor U18098 (N_18098,N_13332,N_16793);
or U18099 (N_18099,N_17311,N_15671);
nor U18100 (N_18100,N_15950,N_12097);
xnor U18101 (N_18101,N_12892,N_15811);
xor U18102 (N_18102,N_16079,N_14529);
nor U18103 (N_18103,N_14230,N_16779);
xor U18104 (N_18104,N_12054,N_14808);
nand U18105 (N_18105,N_12450,N_13408);
and U18106 (N_18106,N_12723,N_12491);
and U18107 (N_18107,N_16574,N_14027);
nor U18108 (N_18108,N_13609,N_17762);
nand U18109 (N_18109,N_16630,N_17147);
or U18110 (N_18110,N_15579,N_12184);
nand U18111 (N_18111,N_14394,N_17819);
or U18112 (N_18112,N_14598,N_17208);
nor U18113 (N_18113,N_13889,N_14997);
and U18114 (N_18114,N_14487,N_15981);
and U18115 (N_18115,N_16485,N_12076);
and U18116 (N_18116,N_12382,N_14200);
nor U18117 (N_18117,N_14144,N_17452);
nand U18118 (N_18118,N_17551,N_15054);
or U18119 (N_18119,N_15532,N_13136);
and U18120 (N_18120,N_15543,N_14741);
xnor U18121 (N_18121,N_17194,N_14480);
xnor U18122 (N_18122,N_12489,N_16238);
and U18123 (N_18123,N_15282,N_13532);
and U18124 (N_18124,N_14432,N_13676);
or U18125 (N_18125,N_12199,N_17711);
nor U18126 (N_18126,N_16335,N_14923);
nand U18127 (N_18127,N_15549,N_14012);
or U18128 (N_18128,N_14336,N_15733);
or U18129 (N_18129,N_12303,N_14071);
nor U18130 (N_18130,N_15649,N_12730);
nand U18131 (N_18131,N_12238,N_17038);
xor U18132 (N_18132,N_15269,N_12912);
nand U18133 (N_18133,N_15917,N_12697);
and U18134 (N_18134,N_16068,N_12319);
xnor U18135 (N_18135,N_17485,N_12618);
nand U18136 (N_18136,N_13510,N_13120);
and U18137 (N_18137,N_15782,N_16668);
or U18138 (N_18138,N_15094,N_12548);
nor U18139 (N_18139,N_16696,N_12127);
xnor U18140 (N_18140,N_17408,N_16653);
xor U18141 (N_18141,N_17122,N_17110);
or U18142 (N_18142,N_15799,N_14906);
and U18143 (N_18143,N_17430,N_16451);
nor U18144 (N_18144,N_17829,N_14338);
and U18145 (N_18145,N_16989,N_16518);
and U18146 (N_18146,N_17435,N_17201);
nor U18147 (N_18147,N_17719,N_16833);
nor U18148 (N_18148,N_13561,N_15345);
and U18149 (N_18149,N_13491,N_13498);
nor U18150 (N_18150,N_16349,N_12352);
or U18151 (N_18151,N_14779,N_15203);
nand U18152 (N_18152,N_13932,N_12711);
nor U18153 (N_18153,N_14373,N_16891);
and U18154 (N_18154,N_15701,N_16726);
and U18155 (N_18155,N_15149,N_16765);
or U18156 (N_18156,N_14424,N_17446);
and U18157 (N_18157,N_16885,N_15158);
nand U18158 (N_18158,N_16433,N_15425);
nand U18159 (N_18159,N_15463,N_15672);
nor U18160 (N_18160,N_12470,N_13952);
xnor U18161 (N_18161,N_15652,N_14155);
nand U18162 (N_18162,N_13864,N_14348);
nand U18163 (N_18163,N_15522,N_15472);
nand U18164 (N_18164,N_14697,N_14490);
xnor U18165 (N_18165,N_13964,N_17111);
nor U18166 (N_18166,N_14851,N_13066);
nand U18167 (N_18167,N_16658,N_17536);
nor U18168 (N_18168,N_17875,N_16967);
nand U18169 (N_18169,N_16368,N_16080);
nor U18170 (N_18170,N_13565,N_14592);
or U18171 (N_18171,N_17804,N_15766);
or U18172 (N_18172,N_16343,N_16923);
xor U18173 (N_18173,N_15370,N_17032);
xnor U18174 (N_18174,N_13114,N_14822);
nor U18175 (N_18175,N_12318,N_13201);
or U18176 (N_18176,N_16539,N_15412);
nand U18177 (N_18177,N_16119,N_15794);
or U18178 (N_18178,N_15187,N_15841);
nor U18179 (N_18179,N_14519,N_17306);
or U18180 (N_18180,N_12775,N_17624);
or U18181 (N_18181,N_16160,N_14534);
or U18182 (N_18182,N_13562,N_17973);
or U18183 (N_18183,N_16636,N_16203);
nand U18184 (N_18184,N_17146,N_14775);
or U18185 (N_18185,N_15637,N_14400);
nor U18186 (N_18186,N_12446,N_13807);
or U18187 (N_18187,N_17084,N_17205);
nand U18188 (N_18188,N_17689,N_12027);
or U18189 (N_18189,N_12278,N_15808);
xor U18190 (N_18190,N_13770,N_12003);
xnor U18191 (N_18191,N_15535,N_14352);
nand U18192 (N_18192,N_17813,N_14819);
nand U18193 (N_18193,N_17617,N_17217);
or U18194 (N_18194,N_17872,N_16573);
nor U18195 (N_18195,N_13720,N_14239);
nor U18196 (N_18196,N_15778,N_14335);
nor U18197 (N_18197,N_13037,N_16398);
nand U18198 (N_18198,N_17622,N_15868);
or U18199 (N_18199,N_13544,N_12999);
xnor U18200 (N_18200,N_16251,N_15600);
xor U18201 (N_18201,N_14416,N_12257);
and U18202 (N_18202,N_14772,N_16642);
nor U18203 (N_18203,N_13102,N_17357);
or U18204 (N_18204,N_15559,N_17789);
and U18205 (N_18205,N_17393,N_12226);
and U18206 (N_18206,N_14749,N_16645);
or U18207 (N_18207,N_12258,N_12824);
and U18208 (N_18208,N_17611,N_13212);
and U18209 (N_18209,N_17226,N_12733);
nor U18210 (N_18210,N_15531,N_17405);
xnor U18211 (N_18211,N_12164,N_17484);
xor U18212 (N_18212,N_13288,N_13714);
nand U18213 (N_18213,N_13618,N_16788);
xnor U18214 (N_18214,N_15586,N_16086);
nand U18215 (N_18215,N_13789,N_12411);
nor U18216 (N_18216,N_14440,N_17934);
xor U18217 (N_18217,N_14913,N_12520);
nand U18218 (N_18218,N_13260,N_12584);
nand U18219 (N_18219,N_12392,N_16694);
nand U18220 (N_18220,N_16135,N_13309);
or U18221 (N_18221,N_14327,N_13831);
nand U18222 (N_18222,N_13778,N_12659);
xnor U18223 (N_18223,N_14409,N_17045);
and U18224 (N_18224,N_15979,N_12563);
or U18225 (N_18225,N_15853,N_12991);
and U18226 (N_18226,N_12742,N_15046);
nand U18227 (N_18227,N_17886,N_15589);
and U18228 (N_18228,N_16186,N_12868);
xnor U18229 (N_18229,N_17746,N_12964);
nand U18230 (N_18230,N_17119,N_17106);
nor U18231 (N_18231,N_13080,N_13278);
nand U18232 (N_18232,N_12037,N_12098);
nand U18233 (N_18233,N_13673,N_17050);
and U18234 (N_18234,N_15914,N_13477);
xnor U18235 (N_18235,N_12201,N_14123);
and U18236 (N_18236,N_17817,N_15371);
nor U18237 (N_18237,N_12468,N_14131);
nor U18238 (N_18238,N_12102,N_17476);
nor U18239 (N_18239,N_16133,N_17531);
and U18240 (N_18240,N_14797,N_14663);
xnor U18241 (N_18241,N_17876,N_13166);
xnor U18242 (N_18242,N_14920,N_13208);
and U18243 (N_18243,N_14988,N_12908);
xnor U18244 (N_18244,N_16148,N_14499);
xor U18245 (N_18245,N_17782,N_13188);
or U18246 (N_18246,N_12431,N_12113);
xor U18247 (N_18247,N_14820,N_12645);
and U18248 (N_18248,N_14963,N_17572);
nand U18249 (N_18249,N_16226,N_13447);
xnor U18250 (N_18250,N_16836,N_13009);
xor U18251 (N_18251,N_13893,N_15066);
nand U18252 (N_18252,N_15747,N_14350);
and U18253 (N_18253,N_15373,N_13499);
nand U18254 (N_18254,N_12575,N_14934);
xnor U18255 (N_18255,N_15636,N_13853);
and U18256 (N_18256,N_14938,N_17915);
nand U18257 (N_18257,N_13574,N_15795);
xnor U18258 (N_18258,N_14583,N_14625);
xor U18259 (N_18259,N_14933,N_13560);
nor U18260 (N_18260,N_12528,N_16818);
and U18261 (N_18261,N_12081,N_14654);
xnor U18262 (N_18262,N_17928,N_16968);
nor U18263 (N_18263,N_14279,N_17607);
or U18264 (N_18264,N_15078,N_16084);
xnor U18265 (N_18265,N_13053,N_16428);
nor U18266 (N_18266,N_16562,N_13509);
nor U18267 (N_18267,N_14964,N_17343);
and U18268 (N_18268,N_16431,N_17362);
nand U18269 (N_18269,N_12911,N_14359);
nor U18270 (N_18270,N_13684,N_12245);
nand U18271 (N_18271,N_17418,N_13195);
xnor U18272 (N_18272,N_16718,N_14177);
xnor U18273 (N_18273,N_16240,N_12684);
nand U18274 (N_18274,N_16509,N_13549);
nand U18275 (N_18275,N_16382,N_15504);
xor U18276 (N_18276,N_13101,N_16544);
and U18277 (N_18277,N_17220,N_14763);
or U18278 (N_18278,N_15486,N_12228);
xnor U18279 (N_18279,N_13731,N_14580);
or U18280 (N_18280,N_13251,N_17675);
xor U18281 (N_18281,N_15278,N_17044);
nor U18282 (N_18282,N_15607,N_13223);
and U18283 (N_18283,N_16639,N_12409);
and U18284 (N_18284,N_12710,N_17302);
or U18285 (N_18285,N_17489,N_17274);
or U18286 (N_18286,N_12345,N_16969);
nand U18287 (N_18287,N_12276,N_16471);
xor U18288 (N_18288,N_13529,N_16258);
xnor U18289 (N_18289,N_13474,N_13911);
nor U18290 (N_18290,N_14040,N_14798);
and U18291 (N_18291,N_14126,N_15133);
xnor U18292 (N_18292,N_17682,N_12531);
nor U18293 (N_18293,N_13656,N_15698);
nand U18294 (N_18294,N_16511,N_15457);
xor U18295 (N_18295,N_15160,N_16704);
and U18296 (N_18296,N_16252,N_12793);
and U18297 (N_18297,N_12007,N_16513);
nand U18298 (N_18298,N_16475,N_14568);
or U18299 (N_18299,N_14304,N_16883);
nand U18300 (N_18300,N_14332,N_15319);
and U18301 (N_18301,N_17750,N_14950);
nor U18302 (N_18302,N_17558,N_12429);
and U18303 (N_18303,N_16834,N_15915);
and U18304 (N_18304,N_17814,N_13313);
xor U18305 (N_18305,N_14402,N_16193);
and U18306 (N_18306,N_17133,N_12815);
or U18307 (N_18307,N_12253,N_13977);
xnor U18308 (N_18308,N_14187,N_13143);
xor U18309 (N_18309,N_16927,N_13044);
and U18310 (N_18310,N_15424,N_16565);
and U18311 (N_18311,N_16303,N_16900);
and U18312 (N_18312,N_16586,N_13699);
nor U18313 (N_18313,N_15849,N_17664);
or U18314 (N_18314,N_13301,N_17327);
nor U18315 (N_18315,N_16152,N_15315);
or U18316 (N_18316,N_13997,N_15332);
xor U18317 (N_18317,N_15923,N_14823);
nor U18318 (N_18318,N_12328,N_17573);
and U18319 (N_18319,N_16609,N_14297);
or U18320 (N_18320,N_13868,N_15286);
nor U18321 (N_18321,N_13448,N_16255);
nand U18322 (N_18322,N_15602,N_12836);
xor U18323 (N_18323,N_15070,N_12100);
nand U18324 (N_18324,N_15837,N_13289);
nor U18325 (N_18325,N_17224,N_12072);
and U18326 (N_18326,N_14932,N_13949);
and U18327 (N_18327,N_12547,N_15302);
xnor U18328 (N_18328,N_17103,N_15040);
xor U18329 (N_18329,N_12546,N_16072);
nor U18330 (N_18330,N_16032,N_17591);
xnor U18331 (N_18331,N_17462,N_15650);
xnor U18332 (N_18332,N_16669,N_12699);
nand U18333 (N_18333,N_16634,N_12962);
or U18334 (N_18334,N_17169,N_17458);
and U18335 (N_18335,N_13969,N_15038);
nand U18336 (N_18336,N_12065,N_12654);
nor U18337 (N_18337,N_15729,N_17259);
and U18338 (N_18338,N_17975,N_15470);
nor U18339 (N_18339,N_15707,N_13394);
nand U18340 (N_18340,N_13083,N_12504);
or U18341 (N_18341,N_13087,N_13282);
or U18342 (N_18342,N_13700,N_14889);
xor U18343 (N_18343,N_15882,N_16447);
and U18344 (N_18344,N_12159,N_13571);
nand U18345 (N_18345,N_16626,N_15830);
or U18346 (N_18346,N_13464,N_16205);
nand U18347 (N_18347,N_17150,N_16289);
nand U18348 (N_18348,N_17370,N_12907);
nor U18349 (N_18349,N_14151,N_16014);
nor U18350 (N_18350,N_12634,N_16396);
nand U18351 (N_18351,N_16430,N_14385);
xnor U18352 (N_18352,N_15073,N_16602);
xor U18353 (N_18353,N_17922,N_12141);
nor U18354 (N_18354,N_15271,N_12362);
nor U18355 (N_18355,N_12840,N_13380);
or U18356 (N_18356,N_12168,N_17281);
and U18357 (N_18357,N_17982,N_14036);
or U18358 (N_18358,N_17200,N_15743);
or U18359 (N_18359,N_17830,N_13927);
and U18360 (N_18360,N_13060,N_15478);
nor U18361 (N_18361,N_17355,N_12623);
nor U18362 (N_18362,N_15590,N_15972);
xnor U18363 (N_18363,N_17542,N_12640);
nand U18364 (N_18364,N_15309,N_17473);
nor U18365 (N_18365,N_17047,N_17139);
xor U18366 (N_18366,N_14276,N_13356);
xnor U18367 (N_18367,N_17267,N_15376);
xnor U18368 (N_18368,N_16040,N_14472);
and U18369 (N_18369,N_12973,N_12348);
nand U18370 (N_18370,N_17248,N_12366);
nand U18371 (N_18371,N_13587,N_13903);
nor U18372 (N_18372,N_17545,N_15410);
or U18373 (N_18373,N_15014,N_15375);
xnor U18374 (N_18374,N_16204,N_17630);
xnor U18375 (N_18375,N_15280,N_17270);
or U18376 (N_18376,N_15349,N_14203);
xnor U18377 (N_18377,N_17881,N_17338);
xor U18378 (N_18378,N_12681,N_12811);
and U18379 (N_18379,N_17631,N_12901);
nor U18380 (N_18380,N_17190,N_13968);
nor U18381 (N_18381,N_14542,N_12187);
and U18382 (N_18382,N_15045,N_15694);
nor U18383 (N_18383,N_14209,N_14720);
xor U18384 (N_18384,N_17698,N_15047);
xor U18385 (N_18385,N_15735,N_13193);
nor U18386 (N_18386,N_13974,N_13526);
and U18387 (N_18387,N_17397,N_16651);
and U18388 (N_18388,N_17249,N_17176);
xnor U18389 (N_18389,N_13540,N_15886);
nand U18390 (N_18390,N_17697,N_13283);
or U18391 (N_18391,N_15227,N_14045);
or U18392 (N_18392,N_12286,N_12680);
xor U18393 (N_18393,N_13816,N_16675);
or U18394 (N_18394,N_16684,N_16286);
nor U18395 (N_18395,N_14674,N_12541);
nor U18396 (N_18396,N_16659,N_16473);
or U18397 (N_18397,N_14169,N_16108);
nor U18398 (N_18398,N_17135,N_13916);
xnor U18399 (N_18399,N_12261,N_16918);
xor U18400 (N_18400,N_15616,N_13866);
or U18401 (N_18401,N_12627,N_13459);
nor U18402 (N_18402,N_15666,N_16397);
xor U18403 (N_18403,N_13177,N_12262);
nand U18404 (N_18404,N_17810,N_16021);
nor U18405 (N_18405,N_13594,N_15580);
or U18406 (N_18406,N_15901,N_13125);
and U18407 (N_18407,N_16299,N_16019);
xnor U18408 (N_18408,N_15386,N_17594);
xor U18409 (N_18409,N_15477,N_13924);
and U18410 (N_18410,N_15894,N_14357);
and U18411 (N_18411,N_12604,N_17828);
xor U18412 (N_18412,N_13920,N_13096);
nor U18413 (N_18413,N_15138,N_17811);
xor U18414 (N_18414,N_14420,N_14632);
nand U18415 (N_18415,N_16886,N_16646);
and U18416 (N_18416,N_14965,N_16444);
and U18417 (N_18417,N_17507,N_14048);
xor U18418 (N_18418,N_13342,N_16106);
or U18419 (N_18419,N_16972,N_15814);
nand U18420 (N_18420,N_17969,N_13211);
nand U18421 (N_18421,N_13832,N_12974);
or U18422 (N_18422,N_17354,N_12255);
xor U18423 (N_18423,N_13295,N_13800);
or U18424 (N_18424,N_16373,N_12764);
nor U18425 (N_18425,N_13458,N_15564);
nor U18426 (N_18426,N_13763,N_16092);
nand U18427 (N_18427,N_15050,N_12967);
or U18428 (N_18428,N_13578,N_17204);
nor U18429 (N_18429,N_16782,N_14903);
nand U18430 (N_18430,N_12804,N_12306);
nand U18431 (N_18431,N_14367,N_17036);
nor U18432 (N_18432,N_17543,N_17300);
nand U18433 (N_18433,N_16667,N_14500);
nor U18434 (N_18434,N_16406,N_16421);
and U18435 (N_18435,N_14801,N_13390);
nand U18436 (N_18436,N_15180,N_14210);
xnor U18437 (N_18437,N_15102,N_15711);
and U18438 (N_18438,N_14642,N_15554);
nand U18439 (N_18439,N_14725,N_16994);
xnor U18440 (N_18440,N_13330,N_16557);
and U18441 (N_18441,N_14634,N_13658);
xor U18442 (N_18442,N_12246,N_12870);
and U18443 (N_18443,N_12736,N_17420);
or U18444 (N_18444,N_17506,N_16652);
nor U18445 (N_18445,N_12248,N_13186);
nor U18446 (N_18446,N_17957,N_16273);
xnor U18447 (N_18447,N_16144,N_12207);
xor U18448 (N_18448,N_17855,N_15132);
xnor U18449 (N_18449,N_13769,N_13967);
nand U18450 (N_18450,N_12929,N_13121);
xnor U18451 (N_18451,N_12674,N_14175);
and U18452 (N_18452,N_13735,N_14880);
nor U18453 (N_18453,N_14216,N_13200);
nand U18454 (N_18454,N_12828,N_17000);
nand U18455 (N_18455,N_13795,N_14661);
and U18456 (N_18456,N_16165,N_15864);
xnor U18457 (N_18457,N_16450,N_16915);
nor U18458 (N_18458,N_16619,N_13597);
xor U18459 (N_18459,N_14910,N_16052);
xnor U18460 (N_18460,N_16536,N_13228);
and U18461 (N_18461,N_16093,N_13384);
xor U18462 (N_18462,N_16976,N_16621);
or U18463 (N_18463,N_16414,N_15338);
and U18464 (N_18464,N_17563,N_12972);
nand U18465 (N_18465,N_14600,N_14980);
nor U18466 (N_18466,N_16437,N_12641);
or U18467 (N_18467,N_17223,N_13766);
xnor U18468 (N_18468,N_13294,N_14742);
xnor U18469 (N_18469,N_15274,N_13431);
and U18470 (N_18470,N_14493,N_12299);
or U18471 (N_18471,N_16033,N_13918);
nor U18472 (N_18472,N_12104,N_14262);
xnor U18473 (N_18473,N_12310,N_13183);
xor U18474 (N_18474,N_16666,N_14051);
nor U18475 (N_18475,N_14105,N_17619);
nand U18476 (N_18476,N_12337,N_12430);
xor U18477 (N_18477,N_17090,N_17062);
and U18478 (N_18478,N_14614,N_12358);
nand U18479 (N_18479,N_13272,N_16991);
nand U18480 (N_18480,N_17608,N_16256);
or U18481 (N_18481,N_13063,N_13256);
nor U18482 (N_18482,N_13848,N_14427);
nand U18483 (N_18483,N_12300,N_15523);
xor U18484 (N_18484,N_17539,N_15426);
nand U18485 (N_18485,N_15630,N_12052);
and U18486 (N_18486,N_17283,N_13803);
nor U18487 (N_18487,N_16048,N_14317);
nand U18488 (N_18488,N_15405,N_13273);
or U18489 (N_18489,N_12126,N_14288);
and U18490 (N_18490,N_14730,N_17599);
and U18491 (N_18491,N_12669,N_14842);
or U18492 (N_18492,N_15578,N_12878);
or U18493 (N_18493,N_13198,N_13151);
nor U18494 (N_18494,N_13019,N_15226);
nand U18495 (N_18495,N_17931,N_17896);
or U18496 (N_18496,N_12984,N_16377);
nand U18497 (N_18497,N_12668,N_13792);
and U18498 (N_18498,N_15755,N_15287);
xor U18499 (N_18499,N_14723,N_17237);
or U18500 (N_18500,N_13747,N_13745);
nand U18501 (N_18501,N_14452,N_16191);
nor U18502 (N_18502,N_13008,N_16379);
and U18503 (N_18503,N_14220,N_12580);
or U18504 (N_18504,N_13252,N_17760);
and U18505 (N_18505,N_13679,N_12073);
or U18506 (N_18506,N_16593,N_17402);
xor U18507 (N_18507,N_17268,N_15189);
nor U18508 (N_18508,N_16197,N_12646);
nor U18509 (N_18509,N_13031,N_15667);
xnor U18510 (N_18510,N_14438,N_14840);
xor U18511 (N_18511,N_14655,N_12445);
nand U18512 (N_18512,N_17033,N_13657);
or U18513 (N_18513,N_14095,N_17597);
nand U18514 (N_18514,N_16563,N_16825);
or U18515 (N_18515,N_16137,N_12761);
or U18516 (N_18516,N_16568,N_16483);
or U18517 (N_18517,N_17304,N_15880);
and U18518 (N_18518,N_16903,N_12189);
nand U18519 (N_18519,N_17880,N_13354);
or U18520 (N_18520,N_15496,N_14049);
xnor U18521 (N_18521,N_15548,N_13235);
nand U18522 (N_18522,N_14154,N_15705);
xor U18523 (N_18523,N_13403,N_12442);
xnor U18524 (N_18524,N_14011,N_14358);
xnor U18525 (N_18525,N_13497,N_16149);
and U18526 (N_18526,N_17126,N_17463);
nor U18527 (N_18527,N_13939,N_15460);
and U18528 (N_18528,N_12810,N_14866);
and U18529 (N_18529,N_15749,N_16678);
and U18530 (N_18530,N_13663,N_13219);
xnor U18531 (N_18531,N_16331,N_17455);
nand U18532 (N_18532,N_15774,N_13202);
or U18533 (N_18533,N_12791,N_17773);
nor U18534 (N_18534,N_14414,N_15439);
nand U18535 (N_18535,N_15856,N_15696);
nand U18536 (N_18536,N_12109,N_17693);
nand U18537 (N_18537,N_13122,N_14993);
nor U18538 (N_18538,N_16982,N_15604);
nand U18539 (N_18539,N_13218,N_15136);
or U18540 (N_18540,N_13247,N_14022);
and U18541 (N_18541,N_16374,N_15825);
xnor U18542 (N_18542,N_16440,N_16131);
or U18543 (N_18543,N_14992,N_13881);
and U18544 (N_18544,N_15290,N_17312);
and U18545 (N_18545,N_12402,N_17234);
or U18546 (N_18546,N_17278,N_17134);
xnor U18547 (N_18547,N_17015,N_14491);
and U18548 (N_18548,N_15943,N_12953);
nor U18549 (N_18549,N_14355,N_12373);
nand U18550 (N_18550,N_12656,N_12067);
nor U18551 (N_18551,N_14751,N_16713);
nand U18552 (N_18552,N_14242,N_15851);
or U18553 (N_18553,N_16039,N_17818);
xnor U18554 (N_18554,N_13018,N_17423);
nor U18555 (N_18555,N_17721,N_17785);
and U18556 (N_18556,N_12886,N_14059);
nor U18557 (N_18557,N_13215,N_14233);
or U18558 (N_18558,N_16742,N_16342);
nor U18559 (N_18559,N_17450,N_17740);
and U18560 (N_18560,N_15802,N_14213);
nand U18561 (N_18561,N_13035,N_17144);
or U18562 (N_18562,N_17264,N_15594);
nor U18563 (N_18563,N_14968,N_17694);
and U18564 (N_18564,N_14465,N_12148);
nor U18565 (N_18565,N_13243,N_17795);
nor U18566 (N_18566,N_13317,N_17580);
nand U18567 (N_18567,N_12036,N_16325);
and U18568 (N_18568,N_12401,N_15854);
or U18569 (N_18569,N_14029,N_16774);
nor U18570 (N_18570,N_14806,N_17731);
nor U18571 (N_18571,N_13472,N_15402);
nand U18572 (N_18572,N_15427,N_14621);
or U18573 (N_18573,N_17364,N_15498);
or U18574 (N_18574,N_13566,N_16244);
nand U18575 (N_18575,N_16791,N_16163);
and U18576 (N_18576,N_15858,N_16357);
or U18577 (N_18577,N_14743,N_15119);
or U18578 (N_18578,N_17082,N_13632);
and U18579 (N_18579,N_15305,N_15584);
nand U18580 (N_18580,N_16708,N_15713);
xor U18581 (N_18581,N_16959,N_16771);
nor U18582 (N_18582,N_14843,N_12157);
xor U18583 (N_18583,N_14316,N_13061);
nor U18584 (N_18584,N_17686,N_16465);
nor U18585 (N_18585,N_12727,N_17736);
xnor U18586 (N_18586,N_15758,N_17279);
nand U18587 (N_18587,N_16958,N_17188);
or U18588 (N_18588,N_17824,N_14941);
xor U18589 (N_18589,N_16839,N_17083);
and U18590 (N_18590,N_12722,N_17710);
and U18591 (N_18591,N_15710,N_17209);
nor U18592 (N_18592,N_17878,N_15777);
nor U18593 (N_18593,N_16749,N_12155);
and U18594 (N_18594,N_12591,N_15238);
nand U18595 (N_18595,N_17924,N_14306);
nand U18596 (N_18596,N_13450,N_17702);
nand U18597 (N_18597,N_17449,N_15860);
xnor U18598 (N_18598,N_16208,N_14667);
xnor U18599 (N_18599,N_16735,N_12251);
nor U18600 (N_18600,N_14167,N_16188);
or U18601 (N_18601,N_15398,N_13304);
nor U18602 (N_18602,N_13489,N_12260);
xnor U18603 (N_18603,N_12633,N_14867);
nand U18604 (N_18604,N_13805,N_16206);
nand U18605 (N_18605,N_13323,N_15002);
or U18606 (N_18606,N_16674,N_12706);
and U18607 (N_18607,N_17733,N_13538);
and U18608 (N_18608,N_16254,N_15257);
nor U18609 (N_18609,N_12380,N_12655);
and U18610 (N_18610,N_15022,N_12968);
nand U18611 (N_18611,N_14665,N_17687);
xnor U18612 (N_18612,N_13592,N_16724);
and U18613 (N_18613,N_12725,N_15714);
or U18614 (N_18614,N_16140,N_12182);
xor U18615 (N_18615,N_16580,N_12838);
xor U18616 (N_18616,N_14103,N_16446);
and U18617 (N_18617,N_15645,N_17744);
and U18618 (N_18618,N_14556,N_13802);
or U18619 (N_18619,N_12917,N_17947);
nand U18620 (N_18620,N_16202,N_14366);
xor U18621 (N_18621,N_15127,N_15381);
nor U18622 (N_18622,N_12652,N_14319);
nand U18623 (N_18623,N_13341,N_15988);
and U18624 (N_18624,N_14649,N_13569);
xnor U18625 (N_18625,N_12132,N_16425);
or U18626 (N_18626,N_13626,N_13882);
or U18627 (N_18627,N_17142,N_16321);
or U18628 (N_18628,N_15395,N_12265);
nand U18629 (N_18629,N_14044,N_14834);
or U18630 (N_18630,N_16493,N_16817);
nor U18631 (N_18631,N_17191,N_16291);
or U18632 (N_18632,N_16185,N_12585);
or U18633 (N_18633,N_15434,N_13664);
xnor U18634 (N_18634,N_17014,N_13869);
nor U18635 (N_18635,N_14532,N_15515);
or U18636 (N_18636,N_12956,N_14397);
and U18637 (N_18637,N_14285,N_15123);
nand U18638 (N_18638,N_12287,N_14464);
xnor U18639 (N_18639,N_17195,N_15184);
nand U18640 (N_18640,N_15260,N_15469);
nor U18641 (N_18641,N_12472,N_16504);
nor U18642 (N_18642,N_12570,N_15263);
xnor U18643 (N_18643,N_12313,N_12374);
or U18644 (N_18644,N_17492,N_17909);
nor U18645 (N_18645,N_17959,N_12790);
xnor U18646 (N_18646,N_17974,N_12927);
and U18647 (N_18647,N_17898,N_14739);
nor U18648 (N_18648,N_13501,N_13423);
xor U18649 (N_18649,N_14624,N_16823);
and U18650 (N_18650,N_13556,N_14517);
xnor U18651 (N_18651,N_14153,N_14684);
nor U18652 (N_18652,N_15331,N_17945);
or U18653 (N_18653,N_14707,N_12822);
nand U18654 (N_18654,N_12152,N_17004);
xnor U18655 (N_18655,N_13245,N_13788);
xnor U18656 (N_18656,N_17104,N_13988);
nand U18657 (N_18657,N_12378,N_17759);
nor U18658 (N_18658,N_14536,N_13065);
and U18659 (N_18659,N_12407,N_13303);
xnor U18660 (N_18660,N_14974,N_15644);
nor U18661 (N_18661,N_12215,N_16278);
xor U18662 (N_18662,N_14796,N_12297);
or U18663 (N_18663,N_13879,N_14246);
xnor U18664 (N_18664,N_13678,N_17447);
nand U18665 (N_18665,N_13173,N_12805);
nor U18666 (N_18666,N_14737,N_13214);
xnor U18667 (N_18667,N_12910,N_12149);
or U18668 (N_18668,N_16610,N_12008);
nor U18669 (N_18669,N_14236,N_14896);
nand U18670 (N_18670,N_14571,N_14486);
nor U18671 (N_18671,N_14443,N_13391);
nand U18672 (N_18672,N_17426,N_12320);
xor U18673 (N_18673,N_16043,N_16699);
and U18674 (N_18674,N_17299,N_12372);
or U18675 (N_18675,N_15763,N_13492);
nor U18676 (N_18676,N_16442,N_17403);
xor U18677 (N_18677,N_12863,N_16001);
nand U18678 (N_18678,N_17679,N_17858);
nand U18679 (N_18679,N_13170,N_17747);
nand U18680 (N_18680,N_15192,N_17232);
and U18681 (N_18681,N_13670,N_17568);
or U18682 (N_18682,N_17832,N_14792);
or U18683 (N_18683,N_15843,N_13479);
nor U18684 (N_18684,N_15569,N_15216);
or U18685 (N_18685,N_13998,N_14845);
or U18686 (N_18686,N_13012,N_17212);
xor U18687 (N_18687,N_14430,N_12213);
nor U18688 (N_18688,N_16089,N_16037);
nand U18689 (N_18689,N_14594,N_17018);
or U18690 (N_18690,N_15709,N_14735);
xor U18691 (N_18691,N_16220,N_13429);
xor U18692 (N_18692,N_17043,N_17319);
nor U18693 (N_18693,N_16897,N_12834);
xor U18694 (N_18694,N_16761,N_12740);
nor U18695 (N_18695,N_12556,N_16911);
nor U18696 (N_18696,N_13651,N_16596);
nor U18697 (N_18697,N_12347,N_16200);
and U18698 (N_18698,N_12125,N_15061);
xor U18699 (N_18699,N_17588,N_16871);
nor U18700 (N_18700,N_16378,N_13719);
nor U18701 (N_18701,N_14717,N_14116);
and U18702 (N_18702,N_12339,N_17633);
nand U18703 (N_18703,N_16992,N_14512);
nand U18704 (N_18704,N_17792,N_17498);
and U18705 (N_18705,N_16881,N_15333);
and U18706 (N_18706,N_14640,N_14237);
nand U18707 (N_18707,N_16796,N_14310);
nand U18708 (N_18708,N_12694,N_16169);
nor U18709 (N_18709,N_12648,N_16942);
nand U18710 (N_18710,N_15878,N_13387);
xnor U18711 (N_18711,N_13590,N_13671);
or U18712 (N_18712,N_15797,N_15327);
xor U18713 (N_18713,N_15682,N_16592);
nor U18714 (N_18714,N_13259,N_16218);
and U18715 (N_18715,N_12028,N_13768);
or U18716 (N_18716,N_16306,N_14447);
xor U18717 (N_18717,N_17554,N_13512);
nor U18718 (N_18718,N_17577,N_16427);
xor U18719 (N_18719,N_13548,N_14668);
or U18720 (N_18720,N_14434,N_13001);
nor U18721 (N_18721,N_17671,N_15582);
xnor U18722 (N_18722,N_12066,N_13942);
xor U18723 (N_18723,N_13261,N_17121);
xor U18724 (N_18724,N_17272,N_17753);
nor U18725 (N_18725,N_14870,N_17986);
or U18726 (N_18726,N_17108,N_15391);
nor U18727 (N_18727,N_12117,N_13424);
nand U18728 (N_18728,N_12642,N_16800);
or U18729 (N_18729,N_15818,N_12249);
or U18730 (N_18730,N_14482,N_15018);
and U18731 (N_18731,N_16481,N_17547);
nor U18732 (N_18732,N_15680,N_15473);
or U18733 (N_18733,N_14174,N_17788);
and U18734 (N_18734,N_16859,N_15081);
nor U18735 (N_18735,N_13191,N_16053);
xor U18736 (N_18736,N_13398,N_15400);
and U18737 (N_18737,N_14435,N_14835);
xnor U18738 (N_18738,N_15838,N_14198);
or U18739 (N_18739,N_16805,N_16582);
and U18740 (N_18740,N_12333,N_17087);
nand U18741 (N_18741,N_15279,N_16350);
and U18742 (N_18742,N_15708,N_14981);
nor U18743 (N_18743,N_12554,N_15389);
nor U18744 (N_18744,N_15629,N_17549);
nand U18745 (N_18745,N_12760,N_15429);
and U18746 (N_18746,N_12322,N_17522);
xor U18747 (N_18747,N_17109,N_17704);
nor U18748 (N_18748,N_13172,N_12507);
nand U18749 (N_18749,N_16405,N_17001);
and U18750 (N_18750,N_15497,N_15955);
xor U18751 (N_18751,N_15702,N_17921);
xnor U18752 (N_18752,N_17800,N_13158);
and U18753 (N_18753,N_16101,N_15730);
and U18754 (N_18754,N_14645,N_12511);
xnor U18755 (N_18755,N_12342,N_16112);
or U18756 (N_18756,N_16495,N_12211);
xor U18757 (N_18757,N_17318,N_14688);
or U18758 (N_18758,N_15320,N_14853);
nand U18759 (N_18759,N_15264,N_14342);
nor U18760 (N_18760,N_13002,N_13596);
nor U18761 (N_18761,N_14839,N_16051);
nand U18762 (N_18762,N_12140,N_12237);
nor U18763 (N_18763,N_12075,N_14628);
nor U18764 (N_18764,N_16187,N_17812);
and U18765 (N_18765,N_14972,N_15893);
nand U18766 (N_18766,N_12171,N_12252);
or U18767 (N_18767,N_15575,N_14518);
nand U18768 (N_18768,N_12644,N_16528);
or U18769 (N_18769,N_13591,N_16171);
and U18770 (N_18770,N_14562,N_14070);
and U18771 (N_18771,N_16531,N_13856);
and U18772 (N_18772,N_14879,N_15642);
or U18773 (N_18773,N_13781,N_15787);
or U18774 (N_18774,N_16514,N_16274);
nor U18775 (N_18775,N_12070,N_15019);
and U18776 (N_18776,N_15079,N_15458);
xor U18777 (N_18777,N_14633,N_15182);
nand U18778 (N_18778,N_16625,N_15910);
or U18779 (N_18779,N_17912,N_15655);
or U18780 (N_18780,N_15219,N_16896);
and U18781 (N_18781,N_17080,N_13014);
nand U18782 (N_18782,N_15664,N_14494);
or U18783 (N_18783,N_17317,N_15557);
and U18784 (N_18784,N_14838,N_17846);
xnor U18785 (N_18785,N_15217,N_15785);
xnor U18786 (N_18786,N_13858,N_16212);
nor U18787 (N_18787,N_17743,N_12068);
nor U18788 (N_18788,N_12079,N_15161);
xor U18789 (N_18789,N_12571,N_13445);
or U18790 (N_18790,N_14346,N_16837);
nor U18791 (N_18791,N_17433,N_16460);
and U18792 (N_18792,N_14145,N_12391);
nand U18793 (N_18793,N_17626,N_12731);
and U18794 (N_18794,N_14894,N_13922);
or U18795 (N_18795,N_15416,N_14620);
and U18796 (N_18796,N_14179,N_17401);
and U18797 (N_18797,N_16655,N_15686);
or U18798 (N_18798,N_17027,N_15233);
nor U18799 (N_18799,N_13649,N_14666);
xnor U18800 (N_18800,N_15143,N_13963);
nand U18801 (N_18801,N_12860,N_13055);
and U18802 (N_18802,N_15545,N_17303);
and U18803 (N_18803,N_14380,N_14446);
xnor U18804 (N_18804,N_13668,N_17030);
or U18805 (N_18805,N_17562,N_14470);
nand U18806 (N_18806,N_12460,N_14201);
nand U18807 (N_18807,N_12658,N_14282);
or U18808 (N_18808,N_16146,N_14951);
nand U18809 (N_18809,N_13614,N_17742);
nor U18810 (N_18810,N_15324,N_14927);
nand U18811 (N_18811,N_12561,N_16276);
or U18812 (N_18812,N_14229,N_12499);
or U18813 (N_18813,N_14524,N_16551);
and U18814 (N_18814,N_16380,N_14365);
nor U18815 (N_18815,N_13825,N_12406);
and U18816 (N_18816,N_13933,N_15307);
nand U18817 (N_18817,N_17953,N_15283);
xor U18818 (N_18818,N_13179,N_13425);
or U18819 (N_18819,N_16751,N_15683);
nand U18820 (N_18820,N_16272,N_12177);
xnor U18821 (N_18821,N_12587,N_14015);
xor U18822 (N_18822,N_15611,N_17064);
xnor U18823 (N_18823,N_12169,N_14565);
nor U18824 (N_18824,N_15240,N_14821);
or U18825 (N_18825,N_14716,N_17478);
nor U18826 (N_18826,N_13270,N_12368);
and U18827 (N_18827,N_12129,N_14962);
and U18828 (N_18828,N_14818,N_12357);
or U18829 (N_18829,N_14682,N_12166);
and U18830 (N_18830,N_17221,N_16277);
and U18831 (N_18831,N_12452,N_16745);
and U18832 (N_18832,N_12145,N_16963);
and U18833 (N_18833,N_13757,N_14596);
and U18834 (N_18834,N_12477,N_12759);
and U18835 (N_18835,N_12273,N_16640);
nand U18836 (N_18836,N_13606,N_17238);
or U18837 (N_18837,N_17275,N_16216);
and U18838 (N_18838,N_13551,N_17745);
or U18839 (N_18839,N_16710,N_16757);
nand U18840 (N_18840,N_17890,N_13264);
nor U18841 (N_18841,N_17431,N_16213);
nand U18842 (N_18842,N_14922,N_14979);
or U18843 (N_18843,N_12667,N_14727);
nor U18844 (N_18844,N_16558,N_14683);
and U18845 (N_18845,N_13249,N_15660);
nand U18846 (N_18846,N_15912,N_14644);
nor U18847 (N_18847,N_14858,N_16869);
xnor U18848 (N_18848,N_13442,N_14188);
nand U18849 (N_18849,N_15231,N_13812);
nand U18850 (N_18850,N_12370,N_16083);
and U18851 (N_18851,N_17888,N_14205);
and U18852 (N_18852,N_16066,N_12340);
xnor U18853 (N_18853,N_14007,N_13360);
xor U18854 (N_18854,N_14915,N_15124);
or U18855 (N_18855,N_12985,N_14766);
nand U18856 (N_18856,N_13025,N_16088);
xor U18857 (N_18857,N_16831,N_17326);
xnor U18858 (N_18858,N_17680,N_17331);
nand U18859 (N_18859,N_14115,N_15313);
and U18860 (N_18860,N_14729,N_15347);
xor U18861 (N_18861,N_14098,N_15210);
or U18862 (N_18862,N_13957,N_12926);
xor U18863 (N_18863,N_16756,N_15228);
or U18864 (N_18864,N_13137,N_16946);
xor U18865 (N_18865,N_13752,N_16546);
xor U18866 (N_18866,N_17101,N_17659);
nor U18867 (N_18867,N_12536,N_17749);
and U18868 (N_18868,N_12128,N_14032);
nor U18869 (N_18869,N_14289,N_14088);
or U18870 (N_18870,N_17381,N_14616);
nor U18871 (N_18871,N_15299,N_17206);
nand U18872 (N_18872,N_15157,N_16077);
and U18873 (N_18873,N_14646,N_13153);
or U18874 (N_18874,N_15346,N_13883);
nand U18875 (N_18875,N_17523,N_15967);
nor U18876 (N_18876,N_17672,N_16180);
and U18877 (N_18877,N_15064,N_14871);
xor U18878 (N_18878,N_12693,N_14047);
nand U18879 (N_18879,N_12614,N_15936);
xnor U18880 (N_18880,N_15392,N_13184);
xor U18881 (N_18881,N_13750,N_15421);
and U18882 (N_18882,N_12998,N_15632);
nand U18883 (N_18883,N_13003,N_12786);
nor U18884 (N_18884,N_17627,N_15715);
or U18885 (N_18885,N_17172,N_16182);
xnor U18886 (N_18886,N_13941,N_14631);
xnor U18887 (N_18887,N_13515,N_16890);
nand U18888 (N_18888,N_15903,N_17368);
and U18889 (N_18889,N_12712,N_15513);
or U18890 (N_18890,N_15296,N_12931);
xor U18891 (N_18891,N_16853,N_16100);
nor U18892 (N_18892,N_12721,N_15028);
and U18893 (N_18893,N_14572,N_15501);
or U18894 (N_18894,N_17942,N_14287);
xnor U18895 (N_18895,N_16769,N_16328);
nand U18896 (N_18896,N_17916,N_16633);
and U18897 (N_18897,N_12453,N_15016);
xor U18898 (N_18898,N_13178,N_16082);
and U18899 (N_18899,N_15842,N_12295);
or U18900 (N_18900,N_13537,N_12651);
nand U18901 (N_18901,N_14966,N_15517);
nor U18902 (N_18902,N_14573,N_16875);
nand U18903 (N_18903,N_15756,N_12662);
xor U18904 (N_18904,N_13762,N_12757);
xor U18905 (N_18905,N_14878,N_14900);
nor U18906 (N_18906,N_14168,N_16371);
xnor U18907 (N_18907,N_12930,N_13633);
nor U18908 (N_18908,N_13005,N_17028);
and U18909 (N_18909,N_12244,N_17464);
nor U18910 (N_18910,N_16585,N_13654);
nand U18911 (N_18911,N_14691,N_15027);
nor U18912 (N_18912,N_12376,N_12095);
or U18913 (N_18913,N_12481,N_14783);
nand U18914 (N_18914,N_17652,N_14445);
and U18915 (N_18915,N_15619,N_13845);
nand U18916 (N_18916,N_16005,N_12976);
xor U18917 (N_18917,N_12856,N_13854);
and U18918 (N_18918,N_14604,N_12613);
xnor U18919 (N_18919,N_13155,N_17256);
xnor U18920 (N_18920,N_14477,N_13016);
nor U18921 (N_18921,N_14158,N_15926);
and U18922 (N_18922,N_17124,N_15601);
nand U18923 (N_18923,N_15262,N_14211);
xnor U18924 (N_18924,N_14256,N_15946);
xnor U18925 (N_18925,N_12250,N_17948);
nand U18926 (N_18926,N_14599,N_13030);
or U18927 (N_18927,N_15166,N_12853);
nor U18928 (N_18928,N_17383,N_15071);
xor U18929 (N_18929,N_16403,N_17904);
nand U18930 (N_18930,N_15541,N_13134);
or U18931 (N_18931,N_16470,N_13267);
xnor U18932 (N_18932,N_15866,N_14263);
or U18933 (N_18933,N_15330,N_14629);
xor U18934 (N_18934,N_17836,N_17765);
nor U18935 (N_18935,N_17305,N_13335);
xor U18936 (N_18936,N_16211,N_15128);
xnor U18937 (N_18937,N_13475,N_15432);
nor U18938 (N_18938,N_15131,N_13508);
or U18939 (N_18939,N_15888,N_16170);
nand U18940 (N_18940,N_17067,N_13746);
xnor U18941 (N_18941,N_16351,N_16063);
nand U18942 (N_18942,N_15918,N_16570);
xor U18943 (N_18943,N_16550,N_17483);
xnor U18944 (N_18944,N_12796,N_15374);
and U18945 (N_18945,N_13995,N_12900);
and U18946 (N_18946,N_15049,N_16613);
and U18947 (N_18947,N_12459,N_12539);
or U18948 (N_18948,N_17055,N_13886);
and U18949 (N_18949,N_17990,N_16750);
nand U18950 (N_18950,N_13126,N_13986);
xor U18951 (N_18951,N_15775,N_13638);
nor U18952 (N_18952,N_17561,N_17665);
and U18953 (N_18953,N_13888,N_12405);
xor U18954 (N_18954,N_17037,N_15017);
or U18955 (N_18955,N_17166,N_14146);
and U18956 (N_18956,N_14046,N_12124);
nor U18957 (N_18957,N_16759,N_13434);
nand U18958 (N_18958,N_13471,N_15958);
xor U18959 (N_18959,N_14459,N_15881);
nor U18960 (N_18960,N_14270,N_14170);
xnor U18961 (N_18961,N_12090,N_15314);
xor U18962 (N_18962,N_14034,N_13994);
xnor U18963 (N_18963,N_17151,N_15104);
nor U18964 (N_18964,N_17722,N_13527);
xor U18965 (N_18965,N_13672,N_13534);
xor U18966 (N_18966,N_14615,N_13945);
or U18967 (N_18967,N_15436,N_16520);
xor U18968 (N_18968,N_16489,N_17363);
xnor U18969 (N_18969,N_16302,N_15328);
nor U18970 (N_18970,N_12394,N_14502);
nor U18971 (N_18971,N_15077,N_16768);
or U18972 (N_18972,N_12670,N_17376);
nand U18973 (N_18973,N_13739,N_16773);
nand U18974 (N_18974,N_13796,N_13705);
and U18975 (N_18975,N_16650,N_13318);
xnor U18976 (N_18976,N_16340,N_15390);
and U18977 (N_18977,N_14746,N_15962);
xor U18978 (N_18978,N_13473,N_16115);
nor U18979 (N_18979,N_12903,N_12865);
nand U18980 (N_18980,N_15030,N_14157);
or U18981 (N_18981,N_15606,N_13078);
nor U18982 (N_18982,N_16556,N_14419);
xor U18983 (N_18983,N_13131,N_14122);
xor U18984 (N_18984,N_15190,N_15092);
nor U18985 (N_18985,N_16503,N_13500);
or U18986 (N_18986,N_16257,N_14407);
and U18987 (N_18987,N_12565,N_16192);
or U18988 (N_18988,N_16363,N_13344);
nand U18989 (N_18989,N_17239,N_12924);
or U18990 (N_18990,N_15861,N_13849);
nor U18991 (N_18991,N_12151,N_17911);
xor U18992 (N_18992,N_14539,N_16827);
nor U18993 (N_18993,N_17096,N_13572);
or U18994 (N_18994,N_17998,N_15624);
nand U18995 (N_18995,N_13575,N_16271);
nor U18996 (N_18996,N_16741,N_14991);
nor U18997 (N_18997,N_16587,N_17603);
and U18998 (N_18998,N_13906,N_17870);
nand U18999 (N_18999,N_14613,N_13815);
nor U19000 (N_19000,N_12516,N_17469);
xnor U19001 (N_19001,N_15561,N_16056);
and U19002 (N_19002,N_14540,N_15508);
nand U19003 (N_19003,N_12420,N_14686);
nor U19004 (N_19004,N_12530,N_12700);
xor U19005 (N_19005,N_14982,N_15640);
xnor U19006 (N_19006,N_16183,N_15646);
or U19007 (N_19007,N_15206,N_14364);
nor U19008 (N_19008,N_14650,N_12144);
or U19009 (N_19009,N_13077,N_16198);
nand U19010 (N_19010,N_17026,N_13385);
nor U19011 (N_19011,N_12282,N_16223);
xnor U19012 (N_19012,N_17801,N_14384);
xnor U19013 (N_19013,N_17276,N_16177);
nor U19014 (N_19014,N_17734,N_12206);
and U19015 (N_19015,N_12043,N_12820);
and U19016 (N_19016,N_13983,N_17112);
xor U19017 (N_19017,N_14530,N_16458);
and U19018 (N_19018,N_17628,N_14120);
xnor U19019 (N_19019,N_13620,N_14561);
nor U19020 (N_19020,N_16851,N_16035);
and U19021 (N_19021,N_12535,N_16308);
nor U19022 (N_19022,N_17735,N_13742);
and U19023 (N_19023,N_17466,N_15112);
or U19024 (N_19024,N_14090,N_14485);
or U19025 (N_19025,N_12636,N_14769);
and U19026 (N_19026,N_17335,N_13042);
or U19027 (N_19027,N_16402,N_14501);
and U19028 (N_19028,N_15142,N_17849);
or U19029 (N_19029,N_15907,N_13161);
nor U19030 (N_19030,N_15595,N_16603);
nor U19031 (N_19031,N_15053,N_13150);
or U19032 (N_19032,N_12465,N_16054);
nor U19033 (N_19033,N_17107,N_12230);
nor U19034 (N_19034,N_17882,N_15172);
nor U19035 (N_19035,N_17225,N_12720);
nor U19036 (N_19036,N_14080,N_15176);
and U19037 (N_19037,N_13677,N_13598);
nor U19038 (N_19038,N_13427,N_16415);
or U19039 (N_19039,N_17460,N_15255);
xnor U19040 (N_19040,N_17352,N_17136);
or U19041 (N_19041,N_15221,N_15396);
or U19042 (N_19042,N_16388,N_13343);
or U19043 (N_19043,N_17535,N_14469);
or U19044 (N_19044,N_13791,N_14050);
or U19045 (N_19045,N_15183,N_16047);
or U19046 (N_19046,N_14503,N_14722);
nand U19047 (N_19047,N_15450,N_13368);
nand U19048 (N_19048,N_17163,N_15201);
nand U19049 (N_19049,N_14086,N_15712);
nor U19050 (N_19050,N_12485,N_17367);
xor U19051 (N_19051,N_13617,N_16590);
xnor U19052 (N_19052,N_17266,N_13899);
nand U19053 (N_19053,N_14186,N_15444);
and U19054 (N_19054,N_16496,N_15512);
or U19055 (N_19055,N_13359,N_12773);
and U19056 (N_19056,N_16599,N_14849);
and U19057 (N_19057,N_12523,N_16365);
or U19058 (N_19058,N_14601,N_15295);
nor U19059 (N_19059,N_14474,N_12061);
or U19060 (N_19060,N_12737,N_14360);
nand U19061 (N_19061,N_17779,N_16297);
xor U19062 (N_19062,N_17105,N_16194);
or U19063 (N_19063,N_15292,N_16283);
or U19064 (N_19064,N_15147,N_13959);
nand U19065 (N_19065,N_16932,N_14410);
nor U19066 (N_19066,N_15214,N_14676);
nand U19067 (N_19067,N_12506,N_15303);
and U19068 (N_19068,N_17419,N_16300);
and U19069 (N_19069,N_14273,N_12443);
nand U19070 (N_19070,N_14888,N_13068);
nor U19071 (N_19071,N_13020,N_17951);
nand U19072 (N_19072,N_15407,N_12508);
nand U19073 (N_19073,N_14704,N_16452);
nor U19074 (N_19074,N_14110,N_16392);
nand U19075 (N_19075,N_17884,N_14101);
nand U19076 (N_19076,N_17763,N_15352);
and U19077 (N_19077,N_13104,N_13240);
nand U19078 (N_19078,N_13411,N_13585);
and U19079 (N_19079,N_13377,N_13352);
or U19080 (N_19080,N_12387,N_13469);
xor U19081 (N_19081,N_12256,N_14940);
nand U19082 (N_19082,N_17802,N_16045);
nand U19083 (N_19083,N_15567,N_15750);
and U19084 (N_19084,N_13478,N_14507);
xor U19085 (N_19085,N_14030,N_16606);
or U19086 (N_19086,N_16057,N_14444);
or U19087 (N_19087,N_14128,N_14325);
and U19088 (N_19088,N_13246,N_16882);
xor U19089 (N_19089,N_15465,N_15990);
xor U19090 (N_19090,N_15798,N_15911);
xor U19091 (N_19091,N_16420,N_15126);
nor U19092 (N_19092,N_17211,N_12354);
or U19093 (N_19093,N_16329,N_13758);
and U19094 (N_19094,N_15697,N_13205);
and U19095 (N_19095,N_17786,N_15058);
and U19096 (N_19096,N_13971,N_16046);
and U19097 (N_19097,N_12234,N_13839);
or U19098 (N_19098,N_13297,N_14533);
and U19099 (N_19099,N_12346,N_14043);
nand U19100 (N_19100,N_16566,N_12861);
xor U19101 (N_19101,N_14113,N_13444);
xnor U19102 (N_19102,N_17339,N_14224);
xor U19103 (N_19103,N_14488,N_14162);
nand U19104 (N_19104,N_17941,N_12715);
and U19105 (N_19105,N_12107,N_12783);
nor U19106 (N_19106,N_14077,N_15443);
xnor U19107 (N_19107,N_14623,N_12696);
or U19108 (N_19108,N_12173,N_12809);
nand U19109 (N_19109,N_14166,N_15587);
nor U19110 (N_19110,N_13098,N_12649);
nor U19111 (N_19111,N_16790,N_15090);
nor U19112 (N_19112,N_17494,N_15527);
and U19113 (N_19113,N_17752,N_17493);
nor U19114 (N_19114,N_16820,N_17309);
and U19115 (N_19115,N_14314,N_17663);
nand U19116 (N_19116,N_16880,N_14226);
and U19117 (N_19117,N_16987,N_14546);
and U19118 (N_19118,N_13604,N_16236);
or U19119 (N_19119,N_12087,N_12880);
or U19120 (N_19120,N_15873,N_14509);
xor U19121 (N_19121,N_16426,N_16117);
or U19122 (N_19122,N_12454,N_17481);
and U19123 (N_19123,N_15834,N_13579);
xnor U19124 (N_19124,N_16941,N_13552);
or U19125 (N_19125,N_16929,N_12943);
or U19126 (N_19126,N_17860,N_16616);
nand U19127 (N_19127,N_13603,N_14828);
or U19128 (N_19128,N_12909,N_15409);
nand U19129 (N_19129,N_16243,N_17155);
and U19130 (N_19130,N_14899,N_12801);
nor U19131 (N_19131,N_12990,N_17548);
xnor U19132 (N_19132,N_12959,N_14347);
and U19133 (N_19133,N_13568,N_14075);
and U19134 (N_19134,N_15753,N_16588);
nor U19135 (N_19135,N_12198,N_15312);
nor U19136 (N_19136,N_14567,N_12396);
nand U19137 (N_19137,N_13253,N_15419);
nor U19138 (N_19138,N_16844,N_15122);
nor U19139 (N_19139,N_16799,N_15948);
nor U19140 (N_19140,N_16266,N_17766);
xor U19141 (N_19141,N_14904,N_13595);
nor U19142 (N_19142,N_13584,N_15399);
or U19143 (N_19143,N_16663,N_12270);
xnor U19144 (N_19144,N_12024,N_16372);
nor U19145 (N_19145,N_12588,N_16980);
and U19146 (N_19146,N_17060,N_14791);
nand U19147 (N_19147,N_14436,N_15850);
nand U19148 (N_19148,N_17646,N_12601);
nor U19149 (N_19149,N_12437,N_17621);
xor U19150 (N_19150,N_14089,N_15272);
and U19151 (N_19151,N_17516,N_13484);
nand U19152 (N_19152,N_17065,N_15765);
xor U19153 (N_19153,N_13627,N_17540);
nor U19154 (N_19154,N_13693,N_17235);
or U19155 (N_19155,N_13346,N_17427);
and U19156 (N_19156,N_12316,N_16219);
xor U19157 (N_19157,N_16716,N_12714);
or U19158 (N_19158,N_15961,N_12963);
nand U19159 (N_19159,N_17784,N_12769);
or U19160 (N_19160,N_12147,N_14140);
or U19161 (N_19161,N_13506,N_15767);
and U19162 (N_19162,N_14795,N_12116);
and U19163 (N_19163,N_17895,N_16912);
or U19164 (N_19164,N_15935,N_14147);
and U19165 (N_19165,N_12606,N_17831);
nand U19166 (N_19166,N_14208,N_14673);
nor U19167 (N_19167,N_13286,N_14698);
nand U19168 (N_19168,N_16157,N_15612);
nand U19169 (N_19169,N_16623,N_13794);
and U19170 (N_19170,N_13165,N_15989);
xor U19171 (N_19171,N_14543,N_12594);
nor U19172 (N_19172,N_16683,N_12572);
or U19173 (N_19173,N_17673,N_14214);
and U19174 (N_19174,N_12290,N_13040);
nor U19175 (N_19175,N_15736,N_17726);
nor U19176 (N_19176,N_13771,N_15963);
or U19177 (N_19177,N_12579,N_16067);
nor U19178 (N_19178,N_12557,N_12467);
nor U19179 (N_19179,N_16466,N_15001);
nand U19180 (N_19180,N_17685,N_16081);
xor U19181 (N_19181,N_15985,N_14868);
and U19182 (N_19182,N_17778,N_14526);
and U19183 (N_19183,N_16717,N_13734);
nor U19184 (N_19184,N_17524,N_13630);
xnor U19185 (N_19185,N_13152,N_13149);
xor U19186 (N_19186,N_13740,N_12495);
nand U19187 (N_19187,N_15052,N_14726);
or U19188 (N_19188,N_15091,N_17263);
xnor U19189 (N_19189,N_15906,N_15930);
or U19190 (N_19190,N_16118,N_13925);
and U19191 (N_19191,N_12231,N_17976);
or U19192 (N_19192,N_16449,N_12020);
xnor U19193 (N_19193,N_14280,N_16155);
xnor U19194 (N_19194,N_16581,N_15096);
and U19195 (N_19195,N_13109,N_17251);
nor U19196 (N_19196,N_15518,N_12476);
nor U19197 (N_19197,N_14732,N_15952);
and U19198 (N_19198,N_14066,N_13593);
nor U19199 (N_19199,N_15289,N_13234);
xnor U19200 (N_19200,N_12033,N_17906);
xor U19201 (N_19201,N_13488,N_17386);
and U19202 (N_19202,N_16895,N_15167);
or U19203 (N_19203,N_16097,N_12162);
nor U19204 (N_19204,N_17724,N_13366);
xor U19205 (N_19205,N_16416,N_15591);
nand U19206 (N_19206,N_13407,N_15746);
xnor U19207 (N_19207,N_17497,N_12509);
xnor U19208 (N_19208,N_12425,N_15093);
and U19209 (N_19209,N_17286,N_17454);
and U19210 (N_19210,N_13612,N_14245);
and U19211 (N_19211,N_13285,N_14947);
nor U19212 (N_19212,N_15852,N_16075);
nor U19213 (N_19213,N_16281,N_17442);
or U19214 (N_19214,N_15924,N_17322);
nand U19215 (N_19215,N_17764,N_17125);
nor U19216 (N_19216,N_13829,N_12898);
and U19217 (N_19217,N_13683,N_12462);
nor U19218 (N_19218,N_14037,N_12935);
nand U19219 (N_19219,N_12121,N_15411);
nor U19220 (N_19220,N_14510,N_12515);
or U19221 (N_19221,N_15169,N_17378);
xor U19222 (N_19222,N_12792,N_17094);
xor U19223 (N_19223,N_15562,N_15996);
and U19224 (N_19224,N_15365,N_15452);
xnor U19225 (N_19225,N_15488,N_17692);
or U19226 (N_19226,N_15482,N_15044);
xor U19227 (N_19227,N_17182,N_12381);
xor U19228 (N_19228,N_12114,N_15397);
and U19229 (N_19229,N_16931,N_12971);
and U19230 (N_19230,N_16709,N_13162);
nand U19231 (N_19231,N_12000,N_12208);
nand U19232 (N_19232,N_14221,N_17482);
and U19233 (N_19233,N_13738,N_17728);
xnor U19234 (N_19234,N_12752,N_16121);
and U19235 (N_19235,N_17013,N_15487);
nor U19236 (N_19236,N_15815,N_17255);
or U19237 (N_19237,N_14508,N_12315);
and U19238 (N_19238,N_14238,N_16725);
or U19239 (N_19239,N_14924,N_16492);
nand U19240 (N_19240,N_17606,N_15741);
nor U19241 (N_19241,N_15846,N_12800);
nand U19242 (N_19242,N_15111,N_12196);
and U19243 (N_19243,N_12922,N_13432);
nand U19244 (N_19244,N_16174,N_12267);
and U19245 (N_19245,N_16523,N_17372);
nor U19246 (N_19246,N_14659,N_14514);
or U19247 (N_19247,N_16816,N_16285);
xnor U19248 (N_19248,N_14608,N_17222);
and U19249 (N_19249,N_13281,N_17257);
and U19250 (N_19250,N_15806,N_13528);
and U19251 (N_19251,N_15140,N_17471);
or U19252 (N_19252,N_13522,N_15997);
or U19253 (N_19253,N_12896,N_12335);
and U19254 (N_19254,N_13690,N_13248);
nand U19255 (N_19255,N_15833,N_12032);
and U19256 (N_19256,N_15464,N_14907);
or U19257 (N_19257,N_12398,N_14939);
and U19258 (N_19258,N_15726,N_14602);
or U19259 (N_19259,N_12204,N_15035);
or U19260 (N_19260,N_12782,N_16614);
xor U19261 (N_19261,N_15012,N_13196);
xor U19262 (N_19262,N_14130,N_13582);
xor U19263 (N_19263,N_16006,N_16542);
xor U19264 (N_19264,N_13239,N_12209);
xor U19265 (N_19265,N_14413,N_16854);
nor U19266 (N_19266,N_15076,N_13072);
and U19267 (N_19267,N_12017,N_17165);
nor U19268 (N_19268,N_12361,N_16657);
nor U19269 (N_19269,N_13142,N_14361);
and U19270 (N_19270,N_16747,N_17950);
nand U19271 (N_19271,N_14429,N_17958);
nand U19272 (N_19272,N_15937,N_15139);
nand U19273 (N_19273,N_13577,N_17807);
nor U19274 (N_19274,N_13820,N_14958);
or U19275 (N_19275,N_17258,N_12025);
or U19276 (N_19276,N_15673,N_16235);
nand U19277 (N_19277,N_14936,N_13756);
xnor U19278 (N_19278,N_13857,N_14299);
and U19279 (N_19279,N_14844,N_17877);
nor U19280 (N_19280,N_15621,N_16961);
nor U19281 (N_19281,N_13646,N_16360);
nand U19282 (N_19282,N_13091,N_15121);
and U19283 (N_19283,N_15475,N_17021);
or U19284 (N_19284,N_17233,N_15087);
nor U19285 (N_19285,N_13570,N_16429);
or U19286 (N_19286,N_17207,N_15581);
nor U19287 (N_19287,N_17893,N_14378);
xor U19288 (N_19288,N_12471,N_17501);
and U19289 (N_19289,N_17244,N_17660);
or U19290 (N_19290,N_16315,N_12360);
xnor U19291 (N_19291,N_17871,N_14375);
nand U19292 (N_19292,N_15742,N_14117);
nand U19293 (N_19293,N_12867,N_14292);
or U19294 (N_19294,N_12513,N_14091);
nor U19295 (N_19295,N_15065,N_14234);
nor U19296 (N_19296,N_12219,N_17236);
xor U19297 (N_19297,N_17565,N_16122);
xor U19298 (N_19298,N_14570,N_16951);
and U19299 (N_19299,N_17358,N_14638);
and U19300 (N_19300,N_16059,N_16661);
nor U19301 (N_19301,N_17821,N_15484);
nor U19302 (N_19302,N_12083,N_17574);
nand U19303 (N_19303,N_14343,N_17504);
or U19304 (N_19304,N_16410,N_15209);
nor U19305 (N_19305,N_14761,N_15413);
xor U19306 (N_19306,N_12006,N_14829);
nor U19307 (N_19307,N_14949,N_14322);
or U19308 (N_19308,N_16162,N_13790);
nand U19309 (N_19309,N_12074,N_12160);
nor U19310 (N_19310,N_13111,N_13659);
nor U19311 (N_19311,N_13628,N_14555);
nor U19312 (N_19312,N_13209,N_17346);
or U19313 (N_19313,N_14622,N_15847);
or U19314 (N_19314,N_16622,N_16013);
and U19315 (N_19315,N_17161,N_14618);
xor U19316 (N_19316,N_14448,N_13872);
xnor U19317 (N_19317,N_16434,N_12705);
nor U19318 (N_19318,N_17154,N_15270);
or U19319 (N_19319,N_13324,N_13682);
xnor U19320 (N_19320,N_13287,N_13185);
nand U19321 (N_19321,N_12091,N_12367);
xor U19322 (N_19322,N_14987,N_16164);
xnor U19323 (N_19323,N_13130,N_15869);
nand U19324 (N_19324,N_12190,N_12010);
nand U19325 (N_19325,N_15377,N_15690);
nand U19326 (N_19326,N_17159,N_17991);
nand U19327 (N_19327,N_17944,N_15215);
nor U19328 (N_19328,N_15762,N_16353);
xnor U19329 (N_19329,N_15438,N_16943);
or U19330 (N_19330,N_14747,N_13824);
or U19331 (N_19331,N_12537,N_13325);
nand U19332 (N_19332,N_16841,N_15977);
nor U19333 (N_19333,N_13227,N_14859);
and U19334 (N_19334,N_12816,N_16988);
nand U19335 (N_19335,N_12524,N_16689);
and U19336 (N_19336,N_14038,N_15447);
xnor U19337 (N_19337,N_15141,N_16733);
nor U19338 (N_19338,N_13213,N_12592);
and U19339 (N_19339,N_12312,N_14557);
nor U19340 (N_19340,N_12913,N_15082);
xor U19341 (N_19341,N_14231,N_14405);
and U19342 (N_19342,N_16908,N_16819);
xnor U19343 (N_19343,N_16916,N_13931);
or U19344 (N_19344,N_16352,N_14333);
nand U19345 (N_19345,N_12650,N_12096);
nand U19346 (N_19346,N_15266,N_17852);
nand U19347 (N_19347,N_17864,N_15635);
and U19348 (N_19348,N_17550,N_15196);
nand U19349 (N_19349,N_14016,N_12795);
xnor U19350 (N_19350,N_17623,N_17157);
nor U19351 (N_19351,N_16516,N_13836);
and U19352 (N_19352,N_12188,N_15420);
nand U19353 (N_19353,N_13494,N_15737);
xnor U19354 (N_19354,N_13373,N_12647);
xnor U19355 (N_19355,N_12799,N_16974);
xnor U19356 (N_19356,N_16702,N_12543);
and U19357 (N_19357,N_13363,N_13232);
xnor U19358 (N_19358,N_15170,N_15191);
nor U19359 (N_19359,N_12205,N_17541);
and U19360 (N_19360,N_13299,N_16671);
xor U19361 (N_19361,N_16179,N_13776);
and U19362 (N_19362,N_12550,N_15676);
xnor U19363 (N_19363,N_14953,N_17723);
nand U19364 (N_19364,N_13006,N_12029);
nor U19365 (N_19365,N_16096,N_15446);
nand U19366 (N_19366,N_13463,N_12932);
xnor U19367 (N_19367,N_13306,N_14112);
and U19368 (N_19368,N_14467,N_16948);
nand U19369 (N_19369,N_14259,N_12156);
or U19370 (N_19370,N_16020,N_14374);
nand U19371 (N_19371,N_17853,N_12891);
or U19372 (N_19372,N_15883,N_14912);
nor U19373 (N_19373,N_15095,N_13843);
or U19374 (N_19374,N_13338,N_16628);
nand U19375 (N_19375,N_14994,N_15171);
nand U19376 (N_19376,N_16986,N_12015);
and U19377 (N_19377,N_13084,N_15941);
nand U19378 (N_19378,N_17717,N_14019);
or U19379 (N_19379,N_17977,N_16947);
nor U19380 (N_19380,N_12808,N_17350);
or U19381 (N_19381,N_12762,N_17553);
and U19382 (N_19382,N_16318,N_13581);
or U19383 (N_19383,N_13669,N_13644);
nand U19384 (N_19384,N_16953,N_12496);
xor U19385 (N_19385,N_13280,N_13483);
nand U19386 (N_19386,N_13513,N_14776);
nand U19387 (N_19387,N_15225,N_16849);
nand U19388 (N_19388,N_13576,N_16736);
nor U19389 (N_19389,N_16116,N_13466);
and U19390 (N_19390,N_17751,N_17187);
xor U19391 (N_19391,N_16359,N_12259);
xnor U19392 (N_19392,N_14767,N_15358);
xnor U19393 (N_19393,N_14160,N_12414);
xnor U19394 (N_19394,N_17641,N_15236);
and U19395 (N_19395,N_17413,N_12275);
and U19396 (N_19396,N_15435,N_13129);
or U19397 (N_19397,N_15974,N_17902);
xnor U19398 (N_19398,N_14687,N_13421);
xnor U19399 (N_19399,N_15417,N_14196);
nand U19400 (N_19400,N_15921,N_12936);
nor U19401 (N_19401,N_14114,N_15987);
xnor U19402 (N_19402,N_16810,N_16151);
nor U19403 (N_19403,N_13079,N_13749);
and U19404 (N_19404,N_14313,N_17253);
nor U19405 (N_19405,N_13007,N_13210);
or U19406 (N_19406,N_16323,N_14300);
or U19407 (N_19407,N_12326,N_17365);
nor U19408 (N_19408,N_14800,N_15716);
nor U19409 (N_19409,N_16413,N_17688);
nor U19410 (N_19410,N_16540,N_15234);
nor U19411 (N_19411,N_12041,N_13460);
or U19412 (N_19412,N_17647,N_15106);
or U19413 (N_19413,N_17310,N_15120);
or U19414 (N_19414,N_14498,N_15362);
or U19415 (N_19415,N_15144,N_16697);
nand U19416 (N_19416,N_16309,N_17620);
or U19417 (N_19417,N_12181,N_16843);
nor U19418 (N_19418,N_15288,N_13996);
and U19419 (N_19419,N_14021,N_12118);
or U19420 (N_19420,N_14141,N_14156);
or U19421 (N_19421,N_17532,N_16456);
and U19422 (N_19422,N_14195,N_13049);
xor U19423 (N_19423,N_14241,N_13830);
nor U19424 (N_19424,N_17412,N_16316);
xor U19425 (N_19425,N_17883,N_14108);
nand U19426 (N_19426,N_15253,N_15356);
nand U19427 (N_19427,N_12957,N_17669);
nor U19428 (N_19428,N_13786,N_14172);
or U19429 (N_19429,N_16239,N_16404);
nor U19430 (N_19430,N_13349,N_13583);
nand U19431 (N_19431,N_12307,N_12427);
and U19432 (N_19432,N_13242,N_12478);
xor U19433 (N_19433,N_16199,N_15193);
nor U19434 (N_19434,N_14522,N_12311);
or U19435 (N_19435,N_16828,N_15249);
and U19436 (N_19436,N_14886,N_13329);
xnor U19437 (N_19437,N_13036,N_15891);
and U19438 (N_19438,N_15445,N_14219);
and U19439 (N_19439,N_16387,N_13216);
nor U19440 (N_19440,N_15454,N_15453);
nand U19441 (N_19441,N_16439,N_14381);
and U19442 (N_19442,N_12223,N_14232);
and U19443 (N_19443,N_12612,N_17625);
nand U19444 (N_19444,N_12611,N_16949);
nand U19445 (N_19445,N_15528,N_13725);
nand U19446 (N_19446,N_16435,N_15029);
nor U19447 (N_19447,N_12277,N_12687);
or U19448 (N_19448,N_16038,N_15651);
or U19449 (N_19449,N_15675,N_15451);
xnor U19450 (N_19450,N_16094,N_14403);
and U19451 (N_19451,N_17653,N_12989);
xor U19452 (N_19452,N_15007,N_16401);
xor U19453 (N_19453,N_17039,N_12266);
and U19454 (N_19454,N_16785,N_17149);
xor U19455 (N_19455,N_15919,N_13897);
nand U19456 (N_19456,N_14826,N_16099);
or U19457 (N_19457,N_16250,N_15865);
and U19458 (N_19458,N_17277,N_13141);
xor U19459 (N_19459,N_14619,N_16098);
or U19460 (N_19460,N_13041,N_14999);
xor U19461 (N_19461,N_15471,N_17075);
or U19462 (N_19462,N_15783,N_13476);
or U19463 (N_19463,N_13862,N_13755);
xnor U19464 (N_19464,N_12167,N_13112);
or U19465 (N_19465,N_14679,N_12086);
or U19466 (N_19466,N_14321,N_12525);
xnor U19467 (N_19467,N_13650,N_16294);
nor U19468 (N_19468,N_13181,N_12919);
nor U19469 (N_19469,N_17589,N_14372);
or U19470 (N_19470,N_13082,N_12200);
nor U19471 (N_19471,N_17020,N_13027);
nor U19472 (N_19472,N_16488,N_15592);
xor U19473 (N_19473,N_17073,N_13784);
or U19474 (N_19474,N_12192,N_17716);
xor U19475 (N_19475,N_12434,N_13124);
nand U19476 (N_19476,N_14127,N_15807);
nand U19477 (N_19477,N_14511,N_15459);
xor U19478 (N_19478,N_17203,N_17336);
nor U19479 (N_19479,N_17715,N_12384);
nand U19480 (N_19480,N_15506,N_12600);
nor U19481 (N_19481,N_13308,N_14635);
nand U19482 (N_19482,N_17936,N_14475);
xnor U19483 (N_19483,N_14724,N_16049);
xor U19484 (N_19484,N_12503,N_13842);
nand U19485 (N_19485,N_15956,N_12864);
nor U19486 (N_19486,N_17041,N_14134);
and U19487 (N_19487,N_12671,N_14281);
nor U19488 (N_19488,N_16607,N_16766);
and U19489 (N_19489,N_14026,N_12802);
nor U19490 (N_19490,N_17410,N_16939);
xor U19491 (N_19491,N_15455,N_17696);
or U19492 (N_19492,N_15462,N_12847);
or U19493 (N_19493,N_12428,N_17648);
or U19494 (N_19494,N_12463,N_16436);
or U19495 (N_19495,N_15024,N_14793);
and U19496 (N_19496,N_12882,N_15335);
and U19497 (N_19497,N_17637,N_13026);
and U19498 (N_19498,N_12023,N_16850);
xnor U19499 (N_19499,N_17456,N_16336);
nor U19500 (N_19500,N_14185,N_16527);
xor U19501 (N_19501,N_15355,N_15776);
nor U19502 (N_19502,N_13182,N_14033);
and U19503 (N_19503,N_14132,N_16813);
and U19504 (N_19504,N_16505,N_12423);
nand U19505 (N_19505,N_15293,N_16499);
nand U19506 (N_19506,N_13884,N_16842);
or U19507 (N_19507,N_13319,N_13973);
xor U19508 (N_19508,N_13616,N_17923);
or U19509 (N_19509,N_16906,N_17042);
and U19510 (N_19510,N_13586,N_13231);
nand U19511 (N_19511,N_12728,N_16957);
nand U19512 (N_19512,N_15323,N_13396);
and U19513 (N_19513,N_14479,N_12574);
and U19514 (N_19514,N_16979,N_15826);
xor U19515 (N_19515,N_13333,N_13652);
nor U19516 (N_19516,N_13250,N_12436);
or U19517 (N_19517,N_17794,N_16649);
or U19518 (N_19518,N_16375,N_12009);
nor U19519 (N_19519,N_15115,N_17840);
nand U19520 (N_19520,N_12918,N_15075);
nor U19521 (N_19521,N_16301,N_15791);
nor U19522 (N_19522,N_15970,N_15285);
xnor U19523 (N_19523,N_16512,N_13692);
nor U19524 (N_19524,N_16209,N_16166);
or U19525 (N_19525,N_17230,N_15620);
xnor U19526 (N_19526,N_13328,N_17129);
nand U19527 (N_19527,N_14748,N_17670);
and U19528 (N_19528,N_13907,N_15403);
nor U19529 (N_19529,N_16002,N_13316);
xnor U19530 (N_19530,N_13470,N_16041);
or U19531 (N_19531,N_12987,N_15920);
xor U19532 (N_19532,N_14550,N_12560);
xor U19533 (N_19533,N_13645,N_15129);
xnor U19534 (N_19534,N_13361,N_15354);
nor U19535 (N_19535,N_17508,N_13691);
or U19536 (N_19536,N_13531,N_15784);
and U19537 (N_19537,N_12620,N_16921);
and U19538 (N_19538,N_12713,N_15530);
and U19539 (N_19539,N_16221,N_14218);
and U19540 (N_19540,N_14989,N_12222);
and U19541 (N_19541,N_17525,N_14003);
xnor U19542 (N_19542,N_13013,N_16559);
nor U19543 (N_19543,N_17380,N_15205);
xnor U19544 (N_19544,N_15839,N_17434);
and U19545 (N_19545,N_17175,N_12819);
nand U19546 (N_19546,N_14961,N_12603);
and U19547 (N_19547,N_15366,N_16677);
or U19548 (N_19548,N_16862,N_15235);
nand U19549 (N_19549,N_12797,N_17049);
or U19550 (N_19550,N_16025,N_13910);
nand U19551 (N_19551,N_16249,N_17377);
xor U19552 (N_19552,N_12897,N_17438);
and U19553 (N_19553,N_14265,N_12486);
nor U19554 (N_19554,N_16933,N_12329);
nor U19555 (N_19555,N_16110,N_17120);
and U19556 (N_19556,N_16526,N_14847);
and U19557 (N_19557,N_15015,N_14516);
nor U19558 (N_19558,N_14309,N_12031);
nand U19559 (N_19559,N_15728,N_12617);
nand U19560 (N_19560,N_17179,N_12894);
nor U19561 (N_19561,N_17382,N_17246);
nor U19562 (N_19562,N_17017,N_16830);
or U19563 (N_19563,N_14023,N_13514);
nor U19564 (N_19564,N_17964,N_12980);
nor U19565 (N_19565,N_13047,N_14389);
nor U19566 (N_19566,N_12638,N_12702);
and U19567 (N_19567,N_16381,N_14192);
or U19568 (N_19568,N_17899,N_14672);
or U19569 (N_19569,N_17349,N_12317);
nand U19570 (N_19570,N_14379,N_17040);
or U19571 (N_19571,N_16567,N_13621);
nor U19572 (N_19572,N_17231,N_14890);
nand U19573 (N_19573,N_17943,N_17127);
nor U19574 (N_19574,N_16287,N_16864);
nand U19575 (N_19575,N_15068,N_17240);
or U19576 (N_19576,N_12707,N_17555);
nand U19577 (N_19577,N_14354,N_17088);
or U19578 (N_19578,N_15552,N_13093);
nor U19579 (N_19579,N_12417,N_16914);
xor U19580 (N_19580,N_12279,N_15380);
and U19581 (N_19581,N_12105,N_16578);
xnor U19582 (N_19582,N_17424,N_15877);
nor U19583 (N_19583,N_15770,N_16484);
xor U19584 (N_19584,N_17850,N_12058);
or U19585 (N_19585,N_17873,N_16346);
or U19586 (N_19586,N_13439,N_15048);
and U19587 (N_19587,N_12676,N_12970);
xor U19588 (N_19588,N_13382,N_12293);
nor U19589 (N_19589,N_17213,N_15700);
nand U19590 (N_19590,N_16161,N_15819);
and U19591 (N_19591,N_17324,N_14093);
xnor U19592 (N_19592,N_14171,N_13292);
xnor U19593 (N_19593,N_16786,N_14329);
xnor U19594 (N_19594,N_16575,N_14193);
nor U19595 (N_19595,N_12842,N_15197);
nand U19596 (N_19596,N_16356,N_17521);
and U19597 (N_19597,N_14527,N_17509);
nor U19598 (N_19598,N_12493,N_16776);
or U19599 (N_19599,N_13461,N_16995);
or U19600 (N_19600,N_17012,N_15678);
and U19601 (N_19601,N_15114,N_12879);
and U19602 (N_19602,N_16924,N_13241);
nand U19603 (N_19603,N_16341,N_16789);
xor U19604 (N_19604,N_12843,N_16960);
and U19605 (N_19605,N_14892,N_12844);
xnor U19606 (N_19606,N_17406,N_12122);
nand U19607 (N_19607,N_14252,N_17429);
nor U19608 (N_19608,N_13347,N_16758);
nand U19609 (N_19609,N_17288,N_14576);
or U19610 (N_19610,N_16579,N_13355);
nor U19611 (N_19611,N_14462,N_13274);
nand U19612 (N_19612,N_13268,N_12683);
nand U19613 (N_19613,N_16832,N_17805);
and U19614 (N_19614,N_17437,N_15900);
xor U19615 (N_19615,N_15603,N_17913);
or U19616 (N_19616,N_12846,N_17293);
xnor U19617 (N_19617,N_16838,N_12751);
or U19618 (N_19618,N_12753,N_15277);
or U19619 (N_19619,N_16391,N_15490);
or U19620 (N_19620,N_12841,N_14612);
or U19621 (N_19621,N_14564,N_16901);
and U19622 (N_19622,N_12449,N_17054);
xor U19623 (N_19623,N_17210,N_12214);
nor U19624 (N_19624,N_16366,N_12247);
or U19625 (N_19625,N_17351,N_16966);
xor U19626 (N_19626,N_15663,N_13919);
nand U19627 (N_19627,N_13321,N_14119);
nand U19628 (N_19628,N_12235,N_15343);
xnor U19629 (N_19629,N_15423,N_17649);
or U19630 (N_19630,N_12893,N_16971);
nor U19631 (N_19631,N_12240,N_14952);
and U19632 (N_19632,N_13374,N_14547);
and U19633 (N_19633,N_15360,N_15113);
or U19634 (N_19634,N_14703,N_13828);
and U19635 (N_19635,N_15321,N_12763);
and U19636 (N_19636,N_15384,N_12390);
or U19637 (N_19637,N_13634,N_17009);
and U19638 (N_19638,N_17247,N_13961);
or U19639 (N_19639,N_12473,N_14948);
nor U19640 (N_19640,N_12743,N_13665);
nand U19641 (N_19641,N_13905,N_12881);
nand U19642 (N_19642,N_15574,N_17341);
or U19643 (N_19643,N_16326,N_17118);
nor U19644 (N_19644,N_17803,N_15933);
nand U19645 (N_19645,N_16824,N_12077);
or U19646 (N_19646,N_16364,N_17905);
nand U19647 (N_19647,N_13635,N_15538);
xnor U19648 (N_19648,N_16605,N_15722);
nor U19649 (N_19649,N_13573,N_13976);
and U19650 (N_19650,N_14864,N_12042);
or U19651 (N_19651,N_16259,N_12784);
nand U19652 (N_19652,N_12048,N_14553);
xnor U19653 (N_19653,N_13801,N_15751);
or U19654 (N_19654,N_13926,N_14052);
and U19655 (N_19655,N_13000,N_13351);
nor U19656 (N_19656,N_17148,N_12035);
or U19657 (N_19657,N_17480,N_12527);
nand U19658 (N_19658,N_13870,N_14425);
or U19659 (N_19659,N_16964,N_14100);
nor U19660 (N_19660,N_17706,N_14771);
and U19661 (N_19661,N_12758,N_13015);
xnor U19662 (N_19662,N_17683,N_14648);
xnor U19663 (N_19663,N_15544,N_13533);
xnor U19664 (N_19664,N_16549,N_16464);
xnor U19665 (N_19665,N_17360,N_14496);
xor U19666 (N_19666,N_15033,N_14700);
xor U19667 (N_19667,N_12050,N_15039);
or U19668 (N_19668,N_16507,N_12657);
xor U19669 (N_19669,N_17443,N_16981);
xnor U19670 (N_19670,N_14558,N_14944);
xnor U19671 (N_19671,N_17907,N_17031);
or U19672 (N_19672,N_16113,N_13639);
and U19673 (N_19673,N_14194,N_14308);
and U19674 (N_19674,N_16879,N_17214);
xor U19675 (N_19675,N_15241,N_12616);
and U19676 (N_19676,N_14001,N_12637);
nand U19677 (N_19677,N_12708,N_16423);
and U19678 (N_19678,N_17707,N_16246);
or U19679 (N_19679,N_12532,N_17421);
xor U19680 (N_19680,N_17737,N_17477);
and U19681 (N_19681,N_12291,N_12379);
and U19682 (N_19682,N_13326,N_16288);
xnor U19683 (N_19683,N_14861,N_12022);
nand U19684 (N_19684,N_14223,N_13467);
nand U19685 (N_19685,N_13999,N_14848);
or U19686 (N_19686,N_13667,N_13422);
nand U19687 (N_19687,N_13947,N_16345);
nand U19688 (N_19688,N_12660,N_12455);
nand U19689 (N_19689,N_17025,N_17407);
nor U19690 (N_19690,N_17316,N_12060);
nand U19691 (N_19691,N_12833,N_12517);
nand U19692 (N_19692,N_16270,N_12709);
xnor U19693 (N_19693,N_15185,N_14671);
nor U19694 (N_19694,N_16627,N_15654);
nor U19695 (N_19695,N_15693,N_12071);
and U19696 (N_19696,N_16457,N_14396);
and U19697 (N_19697,N_17167,N_17772);
nor U19698 (N_19698,N_15199,N_16432);
or U19699 (N_19699,N_16091,N_14862);
and U19700 (N_19700,N_13495,N_13718);
nor U19701 (N_19701,N_12103,N_14802);
and U19702 (N_19702,N_12873,N_14345);
xnor U19703 (N_19703,N_13440,N_15089);
or U19704 (N_19704,N_15085,N_14072);
and U19705 (N_19705,N_17366,N_14525);
xnor U19706 (N_19706,N_12457,N_12538);
nor U19707 (N_19707,N_15928,N_17051);
or U19708 (N_19708,N_15577,N_15608);
and U19709 (N_19709,N_13863,N_12635);
nand U19710 (N_19710,N_13117,N_14370);
or U19711 (N_19711,N_13978,N_17791);
nor U19712 (N_19712,N_16327,N_13144);
xor U19713 (N_19713,N_13045,N_15369);
xor U19714 (N_19714,N_14609,N_14421);
xor U19715 (N_19715,N_15134,N_16158);
or U19716 (N_19716,N_12887,N_15641);
xnor U19717 (N_19717,N_14307,N_14437);
xor U19718 (N_19718,N_16230,N_17593);
and U19719 (N_19719,N_12268,N_12883);
xor U19720 (N_19720,N_17436,N_14528);
xnor U19721 (N_19721,N_17399,N_17815);
nor U19722 (N_19722,N_12047,N_14257);
nand U19723 (N_19723,N_17243,N_12663);
xor U19724 (N_19724,N_17439,N_15353);
and U19725 (N_19725,N_17970,N_14911);
and U19726 (N_19726,N_12343,N_16783);
or U19727 (N_19727,N_15968,N_12923);
xor U19728 (N_19728,N_12518,N_16692);
and U19729 (N_19729,N_12400,N_12851);
nand U19730 (N_19730,N_17461,N_12233);
xnor U19731 (N_19731,N_12274,N_12175);
and U19732 (N_19732,N_16656,N_17841);
nand U19733 (N_19733,N_12937,N_15980);
or U19734 (N_19734,N_17984,N_16660);
or U19735 (N_19735,N_14789,N_15422);
or U19736 (N_19736,N_14149,N_15622);
nand U19737 (N_19737,N_15107,N_14489);
nand U19738 (N_19738,N_12399,N_13449);
xnor U19739 (N_19739,N_15489,N_13992);
nand U19740 (N_19740,N_12451,N_12220);
xor U19741 (N_19741,N_13372,N_13717);
or U19742 (N_19742,N_15430,N_15072);
nor U19743 (N_19743,N_16934,N_12363);
xnor U19744 (N_19744,N_16552,N_15164);
nand U19745 (N_19745,N_15687,N_17862);
nor U19746 (N_19746,N_16015,N_16632);
or U19747 (N_19747,N_15558,N_15298);
nor U19748 (N_19748,N_17488,N_14097);
or U19749 (N_19749,N_12665,N_16954);
and U19750 (N_19750,N_13694,N_17511);
nor U19751 (N_19751,N_17301,N_13039);
xor U19752 (N_19752,N_15524,N_17962);
nor U19753 (N_19753,N_14137,N_15218);
nand U19754 (N_19754,N_12193,N_15163);
and U19755 (N_19755,N_17375,N_16295);
nor U19756 (N_19756,N_12830,N_13176);
nand U19757 (N_19757,N_16109,N_14770);
xor U19758 (N_19758,N_12094,N_16031);
nand U19759 (N_19759,N_12735,N_13076);
nor U19760 (N_19760,N_12698,N_17586);
nor U19761 (N_19761,N_15275,N_17798);
nand U19762 (N_19762,N_13841,N_15689);
nand U19763 (N_19763,N_12057,N_17556);
nor U19764 (N_19764,N_15895,N_12837);
nor U19765 (N_19765,N_12947,N_17640);
nor U19766 (N_19766,N_17956,N_16695);
and U19767 (N_19767,N_15945,N_13365);
or U19768 (N_19768,N_17559,N_14805);
nand U19769 (N_19769,N_16314,N_12850);
and U19770 (N_19770,N_13090,N_16055);
or U19771 (N_19771,N_17374,N_12049);
nor U19772 (N_19772,N_14377,N_16624);
or U19773 (N_19773,N_13965,N_16577);
nand U19774 (N_19774,N_12772,N_13765);
xor U19775 (N_19775,N_16732,N_12174);
xnor U19776 (N_19776,N_16909,N_14125);
nand U19777 (N_19777,N_17323,N_15060);
and U19778 (N_19778,N_14014,N_17385);
nand U19779 (N_19779,N_13736,N_15526);
and U19780 (N_19780,N_13728,N_16754);
nor U19781 (N_19781,N_17874,N_13190);
nand U19782 (N_19782,N_12688,N_15929);
nor U19783 (N_19783,N_12788,N_17005);
xnor U19784 (N_19784,N_14428,N_16344);
xor U19785 (N_19785,N_15281,N_12551);
nand U19786 (N_19786,N_15173,N_17168);
nand U19787 (N_19787,N_13822,N_16234);
or U19788 (N_19788,N_15125,N_15316);
nor U19789 (N_19789,N_12578,N_14846);
and U19790 (N_19790,N_17972,N_12944);
nor U19791 (N_19791,N_13647,N_17512);
nor U19792 (N_19792,N_14505,N_14393);
nor U19793 (N_19793,N_17834,N_12336);
nor U19794 (N_19794,N_16608,N_17690);
nand U19795 (N_19795,N_15020,N_16322);
nor U19796 (N_19796,N_14606,N_15633);
and U19797 (N_19797,N_12664,N_15625);
and U19798 (N_19798,N_12419,N_15159);
and U19799 (N_19799,N_12895,N_14921);
nor U19800 (N_19800,N_17639,N_17002);
xnor U19801 (N_19801,N_13751,N_12803);
nand U19802 (N_19802,N_15151,N_17552);
nor U19803 (N_19803,N_13914,N_17359);
or U19804 (N_19804,N_12040,N_17010);
nor U19805 (N_19805,N_17919,N_12356);
nor U19806 (N_19806,N_12180,N_13823);
or U19807 (N_19807,N_13271,N_13951);
nand U19808 (N_19808,N_15805,N_13029);
nand U19809 (N_19809,N_16555,N_15100);
or U19810 (N_19810,N_12088,N_15634);
or U19811 (N_19811,N_15605,N_14630);
or U19812 (N_19812,N_13902,N_12589);
nor U19813 (N_19813,N_16638,N_14278);
nand U19814 (N_19814,N_15037,N_13687);
nand U19815 (N_19815,N_13230,N_17582);
and U19816 (N_19816,N_16524,N_13455);
and U19817 (N_19817,N_16715,N_17069);
nand U19818 (N_19818,N_14099,N_17914);
nor U19819 (N_19819,N_12653,N_16073);
xor U19820 (N_19820,N_16635,N_16139);
and U19821 (N_19821,N_17575,N_13511);
xnor U19822 (N_19822,N_15976,N_14607);
and U19823 (N_19823,N_16195,N_13081);
or U19824 (N_19824,N_16298,N_17298);
xor U19825 (N_19825,N_15884,N_15385);
nor U19826 (N_19826,N_13833,N_17289);
nor U19827 (N_19827,N_14254,N_15551);
or U19828 (N_19828,N_13712,N_14824);
nor U19829 (N_19829,N_13783,N_14368);
or U19830 (N_19830,N_17530,N_15674);
nand U19831 (N_19831,N_15229,N_12978);
nand U19832 (N_19832,N_14260,N_17885);
xnor U19833 (N_19833,N_12939,N_13225);
xor U19834 (N_19834,N_13913,N_16743);
xnor U19835 (N_19835,N_14872,N_16313);
or U19836 (N_19836,N_16026,N_12216);
xnor U19837 (N_19837,N_17394,N_12995);
and U19838 (N_19838,N_13937,N_15297);
nor U19839 (N_19839,N_14695,N_14323);
nand U19840 (N_19840,N_12823,N_15691);
nand U19841 (N_19841,N_13542,N_13199);
or U19842 (N_19842,N_15195,N_12982);
nand U19843 (N_19843,N_17334,N_15659);
xnor U19844 (N_19844,N_15239,N_12332);
xnor U19845 (N_19845,N_12941,N_13010);
or U19846 (N_19846,N_13192,N_13605);
nor U19847 (N_19847,N_13092,N_14909);
and U19848 (N_19848,N_17519,N_16894);
and U19849 (N_19849,N_16394,N_16647);
nor U19850 (N_19850,N_16348,N_13367);
or U19851 (N_19851,N_17448,N_16132);
nor U19852 (N_19852,N_13164,N_12288);
or U19853 (N_19853,N_12369,N_13613);
and U19854 (N_19854,N_13827,N_13412);
and U19855 (N_19855,N_15610,N_16320);
nor U19856 (N_19856,N_16985,N_12334);
nand U19857 (N_19857,N_13516,N_15156);
xor U19858 (N_19858,N_17768,N_16589);
xor U19859 (N_19859,N_15896,N_14298);
nor U19860 (N_19860,N_15609,N_17657);
and U19861 (N_19861,N_14545,N_12202);
nand U19862 (N_19862,N_14404,N_16455);
and U19863 (N_19863,N_17428,N_14295);
or U19864 (N_19864,N_12777,N_14222);
xor U19865 (N_19865,N_16018,N_14176);
xnor U19866 (N_19866,N_16835,N_16795);
nand U19867 (N_19867,N_15055,N_12940);
nor U19868 (N_19868,N_14689,N_17173);
or U19869 (N_19869,N_17459,N_14651);
nand U19870 (N_19870,N_15268,N_12872);
and U19871 (N_19871,N_12988,N_15898);
xor U19872 (N_19872,N_12217,N_16030);
or U19873 (N_19873,N_15960,N_15661);
xor U19874 (N_19874,N_13993,N_15306);
nand U19875 (N_19875,N_17598,N_12899);
and U19876 (N_19876,N_14495,N_12053);
nor U19877 (N_19877,N_17092,N_15560);
nand U19878 (N_19878,N_15879,N_15116);
xor U19879 (N_19879,N_14986,N_13386);
nor U19880 (N_19880,N_14678,N_12482);
nor U19881 (N_19881,N_12619,N_13375);
or U19882 (N_19882,N_12371,N_15146);
nor U19883 (N_19883,N_12408,N_17445);
xnor U19884 (N_19884,N_17838,N_16746);
xnor U19885 (N_19885,N_14092,N_13662);
xor U19886 (N_19886,N_13846,N_14973);
nor U19887 (N_19887,N_16691,N_13530);
nor U19888 (N_19888,N_13420,N_13437);
nor U19889 (N_19889,N_17425,N_13970);
and U19890 (N_19890,N_17837,N_16332);
or U19891 (N_19891,N_16873,N_12331);
and U19892 (N_19892,N_14977,N_13539);
nand U19893 (N_19893,N_14983,N_17102);
xor U19894 (N_19894,N_13865,N_12172);
nor U19895 (N_19895,N_15437,N_17918);
nor U19896 (N_19896,N_16898,N_16424);
xor U19897 (N_19897,N_12502,N_17908);
xor U19898 (N_19898,N_15021,N_16760);
nor U19899 (N_19899,N_12271,N_12704);
and U19900 (N_19900,N_14143,N_17892);
xor U19901 (N_19901,N_17954,N_14873);
nor U19902 (N_19902,N_17422,N_14212);
and U19903 (N_19903,N_14382,N_13944);
or U19904 (N_19904,N_15583,N_15638);
or U19905 (N_19905,N_12745,N_15208);
nor U19906 (N_19906,N_16714,N_12678);
or U19907 (N_19907,N_16545,N_14087);
nand U19908 (N_19908,N_14662,N_13774);
nand U19909 (N_19909,N_17569,N_17714);
xor U19910 (N_19910,N_13043,N_13194);
nor U19911 (N_19911,N_15628,N_13972);
xnor U19912 (N_19912,N_16637,N_13787);
and U19913 (N_19913,N_15177,N_16459);
or U19914 (N_19914,N_14758,N_12338);
nand U19915 (N_19915,N_12544,N_14856);
xor U19916 (N_19916,N_13233,N_15703);
or U19917 (N_19917,N_16482,N_16062);
xnor U19918 (N_19918,N_14094,N_12170);
and U19919 (N_19919,N_17537,N_14774);
and U19920 (N_19920,N_12082,N_16173);
nor U19921 (N_19921,N_17269,N_12916);
nor U19922 (N_19922,N_14031,N_17979);
or U19923 (N_19923,N_13222,N_15493);
nor U19924 (N_19924,N_16784,N_14249);
and U19925 (N_19925,N_17758,N_17823);
and U19926 (N_19926,N_16560,N_17337);
xor U19927 (N_19927,N_13350,N_12416);
nor U19928 (N_19928,N_15951,N_14713);
nand U19929 (N_19929,N_13452,N_17738);
and U19930 (N_19930,N_16215,N_13277);
xor U19931 (N_19931,N_15614,N_15051);
and U19932 (N_19932,N_15481,N_13255);
xor U19933 (N_19933,N_12631,N_12344);
nor U19934 (N_19934,N_13564,N_15662);
or U19935 (N_19935,N_15734,N_17342);
and U19936 (N_19936,N_12154,N_17502);
nand U19937 (N_19937,N_12925,N_13543);
nand U19938 (N_19938,N_12115,N_14591);
xnor U19939 (N_19939,N_14275,N_15934);
nand U19940 (N_19940,N_15118,N_12483);
nor U19941 (N_19941,N_13401,N_13878);
and U19942 (N_19942,N_16395,N_14261);
nand U19943 (N_19943,N_16983,N_14908);
or U19944 (N_19944,N_14152,N_14587);
nand U19945 (N_19945,N_16028,N_13764);
or U19946 (N_19946,N_14811,N_17727);
nand U19947 (N_19947,N_17250,N_13132);
xnor U19948 (N_19948,N_14142,N_13395);
xor U19949 (N_19949,N_14253,N_17371);
or U19950 (N_19950,N_17379,N_15491);
xnor U19951 (N_19951,N_16537,N_13311);
xnor U19952 (N_19952,N_16009,N_14978);
and U19953 (N_19953,N_16150,N_17297);
nand U19954 (N_19954,N_16594,N_17546);
nor U19955 (N_19955,N_15394,N_17457);
xnor U19956 (N_19956,N_13110,N_12533);
nand U19957 (N_19957,N_16803,N_15230);
nand U19958 (N_19958,N_17453,N_17614);
nor U19959 (N_19959,N_15086,N_15088);
nor U19960 (N_19960,N_12510,N_13946);
nand U19961 (N_19961,N_12415,N_14523);
nand U19962 (N_19962,N_15105,N_13057);
nand U19963 (N_19963,N_13785,N_12002);
and U19964 (N_19964,N_13520,N_16775);
or U19965 (N_19965,N_17520,N_15720);
nor U19966 (N_19966,N_13607,N_15006);
nand U19967 (N_19967,N_16975,N_16738);
nor U19968 (N_19968,N_17925,N_13320);
nor U19969 (N_19969,N_17866,N_12691);
or U19970 (N_19970,N_15110,N_14589);
nor U19971 (N_19971,N_12724,N_17797);
nand U19972 (N_19972,N_17292,N_16978);
nand U19973 (N_19973,N_17968,N_16061);
and U19974 (N_19974,N_16547,N_12403);
xnor U19975 (N_19975,N_13811,N_16253);
xnor U19976 (N_19976,N_13465,N_14386);
xnor U19977 (N_19977,N_15004,N_13602);
and U19978 (N_19978,N_14832,N_13737);
xnor U19979 (N_19979,N_12120,N_14919);
nor U19980 (N_19980,N_13716,N_13103);
nand U19981 (N_19981,N_12979,N_13954);
nor U19982 (N_19982,N_15657,N_16777);
or U19983 (N_19983,N_12490,N_17691);
xnor U19984 (N_19984,N_12441,N_15479);
xor U19985 (N_19985,N_13558,N_13237);
or U19986 (N_19986,N_14484,N_14339);
nor U19987 (N_19987,N_14401,N_12774);
nor U19988 (N_19988,N_13535,N_12602);
or U19989 (N_19989,N_17391,N_16553);
nor U19990 (N_19990,N_14076,N_16232);
xor U19991 (N_19991,N_16731,N_16463);
and U19992 (N_19992,N_17189,N_16384);
nand U19993 (N_19993,N_17528,N_15908);
nand U19994 (N_19994,N_13298,N_14740);
nor U19995 (N_19995,N_15503,N_13759);
nand U19996 (N_19996,N_14180,N_13557);
nor U19997 (N_19997,N_14255,N_12595);
nand U19998 (N_19998,N_17282,N_16330);
nor U19999 (N_19999,N_17940,N_14085);
xnor U20000 (N_20000,N_12194,N_15761);
and U20001 (N_20001,N_17720,N_13011);
and U20002 (N_20002,N_15940,N_16290);
nand U20003 (N_20003,N_15032,N_14133);
and U20004 (N_20004,N_17291,N_13559);
and U20005 (N_20005,N_13753,N_15223);
and U20006 (N_20006,N_15835,N_14028);
nand U20007 (N_20007,N_15494,N_14041);
nand U20008 (N_20008,N_13619,N_16687);
xor U20009 (N_20009,N_13935,N_15200);
nand U20010 (N_20010,N_13928,N_13900);
xor U20011 (N_20011,N_14513,N_17980);
nor U20012 (N_20012,N_15294,N_13220);
or U20013 (N_20013,N_13837,N_17725);
or U20014 (N_20014,N_12854,N_12243);
nor U20015 (N_20015,N_12150,N_17117);
xnor U20016 (N_20016,N_12365,N_14930);
nand U20017 (N_20017,N_14096,N_14164);
nor U20018 (N_20018,N_15174,N_13397);
xor U20019 (N_20019,N_17929,N_14320);
xnor U20020 (N_20020,N_12540,N_16154);
xor U20021 (N_20021,N_15725,N_13426);
nor U20022 (N_20022,N_15339,N_14857);
xor U20023 (N_20023,N_14575,N_17046);
nor U20024 (N_20024,N_17409,N_16706);
nor U20025 (N_20025,N_16263,N_17086);
nor U20026 (N_20026,N_16965,N_12133);
or U20027 (N_20027,N_17451,N_12951);
nor U20028 (N_20028,N_17011,N_14068);
or U20029 (N_20029,N_13302,N_17295);
xor U20030 (N_20030,N_14461,N_15537);
or U20031 (N_20031,N_16584,N_17254);
and U20032 (N_20032,N_16134,N_15668);
nand U20033 (N_20033,N_16770,N_13541);
nand U20034 (N_20034,N_14869,N_15836);
and U20035 (N_20035,N_14925,N_17662);
xor U20036 (N_20036,N_13487,N_16685);
nor U20037 (N_20037,N_17681,N_14217);
nand U20038 (N_20038,N_12330,N_13064);
and U20039 (N_20039,N_17833,N_12280);
and U20040 (N_20040,N_15109,N_17325);
and U20041 (N_20041,N_14637,N_13428);
nand U20042 (N_20042,N_17174,N_17063);
and U20043 (N_20043,N_14757,N_12610);
and U20044 (N_20044,N_15553,N_13547);
nor U20045 (N_20045,N_14392,N_16794);
nand U20046 (N_20046,N_14581,N_16337);
nor U20047 (N_20047,N_13519,N_12857);
nand U20048 (N_20048,N_12438,N_12005);
nor U20049 (N_20049,N_17868,N_14902);
and U20050 (N_20050,N_16846,N_13923);
and U20051 (N_20051,N_14905,N_12433);
or U20052 (N_20052,N_14004,N_14669);
or U20053 (N_20053,N_14617,N_16620);
nor U20054 (N_20054,N_15670,N_16847);
nor U20055 (N_20055,N_15817,N_15237);
xnor U20056 (N_20056,N_17835,N_14876);
or U20057 (N_20057,N_17806,N_14898);
or U20058 (N_20058,N_15653,N_17775);
nor U20059 (N_20059,N_13269,N_14551);
nand U20060 (N_20060,N_15565,N_15507);
nand U20061 (N_20061,N_16069,N_17414);
nand U20062 (N_20062,N_15957,N_14647);
or U20063 (N_20063,N_16127,N_17930);
xor U20064 (N_20064,N_17983,N_14627);
and U20065 (N_20065,N_12178,N_17822);
nand U20066 (N_20066,N_16945,N_12779);
nor U20067 (N_20067,N_16284,N_16125);
nand U20068 (N_20068,N_12719,N_17158);
or U20069 (N_20069,N_12609,N_13229);
nand U20070 (N_20070,N_13265,N_14442);
nand U20071 (N_20071,N_12553,N_16973);
and U20072 (N_20072,N_14340,N_13904);
nand U20073 (N_20073,N_17193,N_17910);
and U20074 (N_20074,N_17903,N_13312);
nand U20075 (N_20075,N_14548,N_13675);
nand U20076 (N_20076,N_14163,N_16902);
nand U20077 (N_20077,N_13726,N_12741);
nor U20078 (N_20078,N_12210,N_16468);
nor U20079 (N_20079,N_12599,N_13610);
xnor U20080 (N_20080,N_17059,N_17003);
and U20081 (N_20081,N_17677,N_17099);
and U20082 (N_20082,N_16654,N_14411);
nor U20083 (N_20083,N_13204,N_12229);
nor U20084 (N_20084,N_13189,N_15627);
and U20085 (N_20085,N_13262,N_13892);
or U20086 (N_20086,N_16662,N_16543);
nand U20087 (N_20087,N_12062,N_13767);
and U20088 (N_20088,N_14165,N_17638);
nor U20089 (N_20089,N_15804,N_13169);
and U20090 (N_20090,N_15224,N_13340);
xor U20091 (N_20091,N_15597,N_12787);
or U20092 (N_20092,N_13414,N_16445);
nor U20093 (N_20093,N_15406,N_12359);
xor U20094 (N_20094,N_14643,N_17307);
or U20095 (N_20095,N_15461,N_17491);
nand U20096 (N_20096,N_14269,N_12583);
nor U20097 (N_20097,N_17993,N_16105);
or U20098 (N_20098,N_13405,N_16175);
nand U20099 (N_20099,N_14129,N_15859);
and U20100 (N_20100,N_15372,N_16522);
xor U20101 (N_20101,N_16597,N_15790);
xor U20102 (N_20102,N_12488,N_13028);
nor U20103 (N_20103,N_14863,N_14161);
or U20104 (N_20104,N_13203,N_15658);
nand U20105 (N_20105,N_12388,N_15613);
nand U20106 (N_20106,N_15768,N_17658);
and U20107 (N_20107,N_12624,N_13038);
and U20108 (N_20108,N_17271,N_16008);
and U20109 (N_20109,N_13709,N_14657);
nor U20110 (N_20110,N_14264,N_17218);
or U20111 (N_20111,N_16705,N_14356);
or U20112 (N_20112,N_15599,N_16899);
or U20113 (N_20113,N_17770,N_15771);
and U20114 (N_20114,N_12011,N_14191);
xnor U20115 (N_20115,N_14318,N_14719);
and U20116 (N_20116,N_12013,N_17988);
nor U20117 (N_20117,N_17949,N_13024);
xnor U20118 (N_20118,N_14303,N_14481);
and U20119 (N_20119,N_13608,N_13503);
xor U20120 (N_20120,N_12375,N_12914);
xnor U20121 (N_20121,N_13835,N_13838);
xnor U20122 (N_20122,N_14733,N_14468);
xnor U20123 (N_20123,N_16922,N_15772);
xnor U20124 (N_20124,N_13388,N_16376);
xor U20125 (N_20125,N_14074,N_13254);
nand U20126 (N_20126,N_13748,N_14010);
nor U20127 (N_20127,N_13545,N_16727);
xor U20128 (N_20128,N_13930,N_13631);
and U20129 (N_20129,N_17078,N_12227);
xor U20130 (N_20130,N_12123,N_17035);
or U20131 (N_20131,N_17160,N_14945);
nand U20132 (N_20132,N_13336,N_16370);
nand U20133 (N_20133,N_12626,N_16201);
nand U20134 (N_20134,N_12666,N_16454);
or U20135 (N_20135,N_14854,N_12325);
and U20136 (N_20136,N_15953,N_15340);
nor U20137 (N_20137,N_16065,N_17654);
nor U20138 (N_20138,N_13860,N_16490);
or U20139 (N_20139,N_17308,N_12685);
nor U20140 (N_20140,N_12165,N_16029);
nand U20141 (N_20141,N_14118,N_13732);
xor U20142 (N_20142,N_12915,N_17052);
xor U20143 (N_20143,N_14681,N_13032);
or U20144 (N_20144,N_13099,N_16279);
nor U20145 (N_20145,N_15827,N_14653);
or U20146 (N_20146,N_16940,N_15414);
or U20147 (N_20147,N_12866,N_17595);
nor U20148 (N_20148,N_14754,N_16595);
or U20149 (N_20149,N_16242,N_15480);
or U20150 (N_20150,N_16517,N_14431);
or U20151 (N_20151,N_14433,N_12958);
nand U20152 (N_20152,N_16950,N_17384);
nand U20153 (N_20153,N_12439,N_14535);
nand U20154 (N_20154,N_15534,N_13168);
nand U20155 (N_20155,N_12301,N_14664);
xor U20156 (N_20156,N_16767,N_16190);
and U20157 (N_20157,N_17034,N_12263);
nand U20158 (N_20158,N_16729,N_12862);
nor U20159 (N_20159,N_12018,N_12993);
or U20160 (N_20160,N_13798,N_12292);
xor U20161 (N_20161,N_17995,N_15862);
and U20162 (N_20162,N_17100,N_12078);
and U20163 (N_20163,N_15492,N_13686);
nor U20164 (N_20164,N_12661,N_15732);
or U20165 (N_20165,N_16058,N_13873);
and U20166 (N_20166,N_13987,N_12826);
nor U20167 (N_20167,N_13840,N_16129);
and U20168 (N_20168,N_13174,N_14850);
xor U20169 (N_20169,N_16797,N_16538);
and U20170 (N_20170,N_13707,N_16920);
xnor U20171 (N_20171,N_15154,N_15803);
and U20172 (N_20172,N_13086,N_15995);
xor U20173 (N_20173,N_17348,N_16787);
or U20174 (N_20174,N_12890,N_13381);
nor U20175 (N_20175,N_17170,N_16938);
xor U20176 (N_20176,N_14266,N_17989);
xor U20177 (N_20177,N_14680,N_16044);
nor U20178 (N_20178,N_12106,N_12875);
xnor U20179 (N_20179,N_14457,N_17668);
nor U20180 (N_20180,N_12966,N_12484);
nor U20181 (N_20181,N_14967,N_17192);
or U20182 (N_20182,N_16347,N_16601);
xor U20183 (N_20183,N_15969,N_13955);
and U20184 (N_20184,N_17570,N_15254);
nand U20185 (N_20185,N_17089,N_15408);
xor U20186 (N_20186,N_15773,N_17503);
and U20187 (N_20187,N_13480,N_15148);
or U20188 (N_20188,N_14054,N_16479);
and U20189 (N_20189,N_15739,N_15456);
xnor U20190 (N_20190,N_13680,N_13724);
nor U20191 (N_20191,N_17215,N_15909);
and U20192 (N_20192,N_14351,N_17867);
and U20193 (N_20193,N_12143,N_17008);
nand U20194 (N_20194,N_17114,N_17140);
nor U20195 (N_20195,N_14463,N_12264);
nor U20196 (N_20196,N_16564,N_15026);
nand U20197 (N_20197,N_14541,N_12458);
xnor U20198 (N_20198,N_15796,N_15175);
nor U20199 (N_20199,N_16778,N_15786);
nand U20200 (N_20200,N_15573,N_15669);
xnor U20201 (N_20201,N_12689,N_16631);
xnor U20202 (N_20202,N_16629,N_14181);
and U20203 (N_20203,N_14712,N_12545);
nor U20204 (N_20204,N_13943,N_17981);
nor U20205 (N_20205,N_17757,N_12732);
nor U20206 (N_20206,N_14833,N_15626);
and U20207 (N_20207,N_16907,N_13982);
or U20208 (N_20208,N_16554,N_16740);
or U20209 (N_20209,N_13451,N_16138);
nor U20210 (N_20210,N_16070,N_16711);
xor U20211 (N_20211,N_12965,N_17389);
xor U20212 (N_20212,N_12158,N_13345);
and U20213 (N_20213,N_16707,N_15145);
xnor U20214 (N_20214,N_14277,N_17844);
xnor U20215 (N_20215,N_12101,N_17629);
nand U20216 (N_20216,N_16618,N_16867);
nand U20217 (N_20217,N_14750,N_17252);
or U20218 (N_20218,N_15155,N_14588);
nor U20219 (N_20219,N_14415,N_13648);
or U20220 (N_20220,N_17344,N_13446);
or U20221 (N_20221,N_13909,N_16798);
nand U20222 (N_20222,N_17856,N_15792);
or U20223 (N_20223,N_14390,N_17610);
xor U20224 (N_20224,N_16023,N_15361);
nor U20225 (N_20225,N_13486,N_12056);
xor U20226 (N_20226,N_15964,N_17500);
nand U20227 (N_20227,N_16107,N_16467);
nand U20228 (N_20228,N_16060,N_12395);
xnor U20229 (N_20229,N_16147,N_16693);
or U20230 (N_20230,N_15570,N_14636);
or U20231 (N_20231,N_16469,N_15533);
or U20232 (N_20232,N_15718,N_15207);
xnor U20233 (N_20233,N_14417,N_13023);
and U20234 (N_20234,N_14331,N_13075);
xnor U20235 (N_20235,N_14056,N_14752);
and U20236 (N_20236,N_12566,N_15010);
or U20237 (N_20237,N_13818,N_13417);
or U20238 (N_20238,N_15563,N_16399);
nor U20239 (N_20239,N_15198,N_14885);
and U20240 (N_20240,N_15857,N_12131);
or U20241 (N_20241,N_17946,N_15211);
and U20242 (N_20242,N_15300,N_17022);
and U20243 (N_20243,N_14138,N_15485);
nor U20244 (N_20244,N_14078,N_17613);
or U20245 (N_20245,N_14701,N_14928);
nor U20246 (N_20246,N_13793,N_14324);
xnor U20247 (N_20247,N_15848,N_14692);
and U20248 (N_20248,N_12456,N_12734);
nor U20249 (N_20249,N_17616,N_17557);
and U20250 (N_20250,N_16644,N_14002);
or U20251 (N_20251,N_12904,N_15367);
or U20252 (N_20252,N_17171,N_13279);
and U20253 (N_20253,N_15813,N_12749);
and U20254 (N_20254,N_16648,N_12855);
xnor U20255 (N_20255,N_16956,N_17113);
and U20256 (N_20256,N_14084,N_16541);
xor U20257 (N_20257,N_15137,N_12232);
xnor U20258 (N_20258,N_16111,N_15704);
and U20259 (N_20259,N_13106,N_13400);
nand U20260 (N_20260,N_12832,N_15348);
or U20261 (N_20261,N_14597,N_12176);
nor U20262 (N_20262,N_14887,N_15994);
and U20263 (N_20263,N_16214,N_14816);
nor U20264 (N_20264,N_16120,N_13418);
xnor U20265 (N_20265,N_14865,N_15350);
and U20266 (N_20266,N_12692,N_14362);
or U20267 (N_20267,N_15904,N_16521);
and U20268 (N_20268,N_13088,N_13761);
xnor U20269 (N_20269,N_12139,N_17474);
xor U20270 (N_20270,N_16017,N_17790);
nor U20271 (N_20271,N_16293,N_16095);
nand U20272 (N_20272,N_16003,N_17152);
or U20273 (N_20273,N_14005,N_17859);
and U20274 (N_20274,N_12950,N_13073);
or U20275 (N_20275,N_17756,N_15529);
nand U20276 (N_20276,N_14579,N_17847);
xor U20277 (N_20277,N_17048,N_17845);
or U20278 (N_20278,N_17518,N_17185);
or U20279 (N_20279,N_15179,N_13275);
nand U20280 (N_20280,N_13772,N_12254);
nand U20281 (N_20281,N_14931,N_15499);
and U20282 (N_20282,N_15467,N_16548);
and U20283 (N_20283,N_13912,N_17952);
or U20284 (N_20284,N_13171,N_12888);
nand U20285 (N_20285,N_16700,N_16780);
and U20286 (N_20286,N_12552,N_17296);
nor U20287 (N_20287,N_13490,N_16261);
nor U20288 (N_20288,N_17329,N_17294);
nand U20289 (N_20289,N_17245,N_17198);
or U20290 (N_20290,N_13453,N_16304);
and U20291 (N_20291,N_16104,N_12942);
xor U20292 (N_20292,N_12492,N_13898);
nand U20293 (N_20293,N_17644,N_14753);
nand U20294 (N_20294,N_17705,N_16984);
and U20295 (N_20295,N_15991,N_13688);
or U20296 (N_20296,N_13896,N_13744);
nor U20297 (N_20297,N_16888,N_17181);
and U20298 (N_20298,N_15310,N_16826);
and U20299 (N_20299,N_16282,N_14017);
or U20300 (N_20300,N_14765,N_13071);
nand U20301 (N_20301,N_14715,N_16324);
xnor U20302 (N_20302,N_12586,N_12341);
nand U20303 (N_20303,N_17678,N_14603);
nor U20304 (N_20304,N_14079,N_17996);
or U20305 (N_20305,N_13307,N_17085);
or U20306 (N_20306,N_13804,N_14699);
or U20307 (N_20307,N_13138,N_14399);
nand U20308 (N_20308,N_17963,N_16997);
and U20309 (N_20309,N_17415,N_16050);
or U20310 (N_20310,N_17581,N_15939);
xnor U20311 (N_20311,N_17058,N_15393);
nand U20312 (N_20312,N_17138,N_12386);
xor U20313 (N_20313,N_13291,N_14268);
and U20314 (N_20314,N_16569,N_16872);
nand U20315 (N_20315,N_13624,N_14985);
or U20316 (N_20316,N_16448,N_17332);
or U20317 (N_20317,N_13875,N_13507);
or U20318 (N_20318,N_16822,N_15252);
nor U20319 (N_20319,N_13135,N_17340);
nor U20320 (N_20320,N_15520,N_12884);
and U20321 (N_20321,N_15874,N_15999);
nand U20322 (N_20322,N_13553,N_15779);
or U20323 (N_20323,N_16275,N_17416);
nor U20324 (N_20324,N_12349,N_13851);
nand U20325 (N_20325,N_15308,N_15942);
nand U20326 (N_20326,N_12064,N_13482);
or U20327 (N_20327,N_15329,N_17072);
xor U20328 (N_20328,N_16811,N_12576);
and U20329 (N_20329,N_14586,N_14675);
or U20330 (N_20330,N_15831,N_13867);
xnor U20331 (N_20331,N_13305,N_17709);
nand U20332 (N_20332,N_17162,N_12643);
nand U20333 (N_20333,N_13689,N_14449);
nor U20334 (N_20334,N_17444,N_14258);
nor U20335 (N_20335,N_13871,N_14734);
nand U20336 (N_20336,N_12289,N_12994);
nand U20337 (N_20337,N_15351,N_17007);
or U20338 (N_20338,N_16856,N_16764);
nor U20339 (N_20339,N_16408,N_16612);
and U20340 (N_20340,N_14283,N_15514);
nand U20341 (N_20341,N_13917,N_12045);
nand U20342 (N_20342,N_16367,N_15631);
nor U20343 (N_20343,N_16698,N_16919);
nor U20344 (N_20344,N_12323,N_13826);
nand U20345 (N_20345,N_12738,N_15311);
nor U20346 (N_20346,N_15034,N_16393);
xor U20347 (N_20347,N_16296,N_13140);
or U20348 (N_20348,N_14660,N_16561);
nand U20349 (N_20349,N_12377,N_13364);
and U20350 (N_20350,N_12781,N_12996);
and U20351 (N_20351,N_15194,N_13119);
nor U20352 (N_20352,N_17961,N_14694);
or U20353 (N_20353,N_14121,N_13314);
xnor U20354 (N_20354,N_12298,N_13901);
nand U20355 (N_20355,N_12038,N_12353);
xnor U20356 (N_20356,N_14439,N_12019);
nand U20357 (N_20357,N_15441,N_16248);
and U20358 (N_20358,N_14159,N_16807);
or U20359 (N_20359,N_13133,N_15738);
nor U20360 (N_20360,N_15665,N_13674);
nand U20361 (N_20361,N_13402,N_15168);
nand U20362 (N_20362,N_12928,N_13052);
nand U20363 (N_20363,N_13160,N_14235);
nand U20364 (N_20364,N_17164,N_14901);
xor U20365 (N_20365,N_14935,N_13410);
nor U20366 (N_20366,N_15793,N_12615);
nand U20367 (N_20367,N_17527,N_14057);
and U20368 (N_20368,N_15973,N_12063);
nand U20369 (N_20369,N_14762,N_15648);
or U20370 (N_20370,N_12014,N_13601);
xnor U20371 (N_20371,N_16874,N_15643);
or U20372 (N_20372,N_15692,N_15975);
and U20373 (N_20373,N_15889,N_15284);
and U20374 (N_20374,N_12806,N_15378);
nor U20375 (N_20375,N_13810,N_17799);
or U20376 (N_20376,N_14566,N_15617);
xor U20377 (N_20377,N_17345,N_14929);
nor U20378 (N_20378,N_17290,N_16310);
nor U20379 (N_20379,N_13915,N_12448);
nor U20380 (N_20380,N_16168,N_13266);
nand U20381 (N_20381,N_13413,N_15723);
and U20382 (N_20382,N_16497,N_17787);
xnor U20383 (N_20383,N_17634,N_17517);
or U20384 (N_20384,N_16993,N_12153);
nor U20385 (N_20385,N_16845,N_12849);
nor U20386 (N_20386,N_13399,N_17130);
nor U20387 (N_20387,N_14207,N_14423);
xnor U20388 (N_20388,N_12505,N_13852);
nor U20389 (N_20389,N_16664,N_13885);
or U20390 (N_20390,N_13369,N_13550);
and U20391 (N_20391,N_14942,N_12955);
and U20392 (N_20392,N_13502,N_12997);
and U20393 (N_20393,N_13100,N_14471);
nand U20394 (N_20394,N_17879,N_14247);
xor U20395 (N_20395,N_15938,N_12986);
or U20396 (N_20396,N_14136,N_12981);
xor U20397 (N_20397,N_16319,N_15468);
and U20398 (N_20398,N_12718,N_12921);
nand U20399 (N_20399,N_14291,N_15744);
nor U20400 (N_20400,N_15916,N_15431);
nand U20401 (N_20401,N_12080,N_13046);
and U20402 (N_20402,N_14554,N_16478);
and U20403 (N_20403,N_16500,N_17261);
nor U20404 (N_20404,N_16389,N_13070);
nand U20405 (N_20405,N_14721,N_15769);
and U20406 (N_20406,N_14107,N_12542);
nand U20407 (N_20407,N_13721,N_15647);
nor U20408 (N_20408,N_17315,N_13339);
or U20409 (N_20409,N_17861,N_13085);
and U20410 (N_20410,N_15500,N_12519);
and U20411 (N_20411,N_13695,N_17997);
or U20412 (N_20412,N_14916,N_17479);
xor U20413 (N_20413,N_13989,N_14009);
nor U20414 (N_20414,N_17676,N_15387);
and U20415 (N_20415,N_15754,N_13154);
nand U20416 (N_20416,N_14228,N_16870);
or U20417 (N_20417,N_15925,N_15556);
and U20418 (N_20418,N_17825,N_17684);
and U20419 (N_20419,N_15550,N_13817);
and U20420 (N_20420,N_14605,N_14584);
nand U20421 (N_20421,N_14690,N_12562);
xnor U20422 (N_20422,N_17141,N_15025);
and U20423 (N_20423,N_17330,N_14458);
nand U20424 (N_20424,N_17369,N_14881);
nand U20425 (N_20425,N_14067,N_15781);
nand U20426 (N_20426,N_17280,N_15598);
nor U20427 (N_20427,N_15502,N_12628);
and U20428 (N_20428,N_14656,N_14124);
nor U20429 (N_20429,N_15546,N_17411);
and U20430 (N_20430,N_12568,N_16090);
or U20431 (N_20431,N_17926,N_17605);
and U20432 (N_20432,N_14937,N_14652);
and U20433 (N_20433,N_12327,N_14055);
nor U20434 (N_20434,N_16792,N_17068);
nand U20435 (N_20435,N_13108,N_17769);
nand U20436 (N_20436,N_16262,N_14267);
and U20437 (N_20437,N_17285,N_16877);
xnor U20438 (N_20438,N_15571,N_13636);
xor U20439 (N_20439,N_12920,N_14240);
xor U20440 (N_20440,N_12983,N_14875);
nand U20441 (N_20441,N_15511,N_15041);
nand U20442 (N_20442,N_17353,N_15685);
xor U20443 (N_20443,N_13908,N_14227);
and U20444 (N_20444,N_13599,N_12059);
nor U20445 (N_20445,N_16354,N_12389);
nand U20446 (N_20446,N_14760,N_14708);
nand U20447 (N_20447,N_16887,N_15576);
nand U20448 (N_20448,N_17091,N_16889);
nand U20449 (N_20449,N_15036,N_12089);
nand U20450 (N_20450,N_16000,N_13703);
and U20451 (N_20451,N_15905,N_12593);
and U20452 (N_20452,N_13034,N_14460);
or U20453 (N_20453,N_14183,N_16576);
nor U20454 (N_20454,N_15913,N_14202);
and U20455 (N_20455,N_17978,N_12283);
nand U20456 (N_20456,N_16734,N_13331);
nor U20457 (N_20457,N_15922,N_12703);
xnor U20458 (N_20458,N_15516,N_16145);
nand U20459 (N_20459,N_15304,N_12021);
or U20460 (N_20460,N_17887,N_14877);
nor U20461 (N_20461,N_13416,N_12827);
nor U20462 (N_20462,N_17123,N_17699);
and U20463 (N_20463,N_13555,N_13710);
xnor U20464 (N_20464,N_16571,N_13625);
and U20465 (N_20465,N_15337,N_14714);
xnor U20466 (N_20466,N_16519,N_12221);
or U20467 (N_20467,N_17816,N_14956);
xnor U20468 (N_20468,N_16231,N_12130);
and U20469 (N_20469,N_15359,N_14926);
nand U20470 (N_20470,N_12567,N_15982);
or U20471 (N_20471,N_14271,N_17321);
and U20472 (N_20472,N_14810,N_12085);
nand U20473 (N_20473,N_14777,N_12776);
nand U20474 (N_20474,N_14918,N_12768);
and U20475 (N_20475,N_13392,N_13834);
or U20476 (N_20476,N_12241,N_13637);
nand U20477 (N_20477,N_14827,N_13159);
or U20478 (N_20478,N_15752,N_17571);
nor U20479 (N_20479,N_12770,N_16311);
nor U20480 (N_20480,N_15181,N_14641);
nor U20481 (N_20481,N_16762,N_16763);
nand U20482 (N_20482,N_16944,N_17729);
and U20483 (N_20483,N_12785,N_13145);
nor U20484 (N_20484,N_16935,N_14595);
nor U20485 (N_20485,N_13921,N_13438);
or U20486 (N_20486,N_13643,N_14969);
or U20487 (N_20487,N_13435,N_16362);
xnor U20488 (N_20488,N_12577,N_15256);
nand U20489 (N_20489,N_14710,N_13207);
and U20490 (N_20490,N_12163,N_17732);
and U20491 (N_20491,N_14395,N_13217);
xnor U20492 (N_20492,N_14135,N_14422);
xnor U20493 (N_20493,N_13094,N_15336);
xnor U20494 (N_20494,N_16673,N_16228);
nor U20495 (N_20495,N_14976,N_12497);
and U20496 (N_20496,N_16878,N_15074);
xnor U20497 (N_20497,N_17475,N_14296);
or U20498 (N_20498,N_14860,N_12569);
or U20499 (N_20499,N_15043,N_16999);
xnor U20500 (N_20500,N_14341,N_14897);
or U20501 (N_20501,N_17701,N_16508);
xnor U20502 (N_20502,N_17183,N_13389);
nand U20503 (N_20503,N_16812,N_16443);
xor U20504 (N_20504,N_14790,N_12798);
or U20505 (N_20505,N_15428,N_15899);
and U20506 (N_20506,N_16604,N_16027);
or U20507 (N_20507,N_17767,N_14328);
xor U20508 (N_20508,N_15954,N_12494);
nand U20509 (N_20509,N_17754,N_17132);
nand U20510 (N_20510,N_13702,N_14454);
and U20511 (N_20511,N_14784,N_12767);
or U20512 (N_20512,N_12203,N_17016);
nor U20513 (N_20513,N_16412,N_13887);
nand U20514 (N_20514,N_16476,N_14042);
or U20515 (N_20515,N_13990,N_17515);
and U20516 (N_20516,N_14334,N_13244);
or U20517 (N_20517,N_13485,N_12564);
nand U20518 (N_20518,N_17667,N_12134);
nor U20519 (N_20519,N_16739,N_13462);
xnor U20520 (N_20520,N_16808,N_14371);
nand U20521 (N_20521,N_13322,N_13069);
xor U20522 (N_20522,N_13334,N_17006);
and U20523 (N_20523,N_16502,N_15810);
xor U20524 (N_20524,N_16868,N_14391);
and U20525 (N_20525,N_12807,N_16012);
xor U20526 (N_20526,N_17774,N_14473);
xor U20527 (N_20527,N_14225,N_16809);
nand U20528 (N_20528,N_14590,N_12825);
xor U20529 (N_20529,N_15947,N_14825);
xnor U20530 (N_20530,N_15971,N_13940);
xnor U20531 (N_20531,N_12948,N_16172);
nand U20532 (N_20532,N_12529,N_13580);
or U20533 (N_20533,N_14173,N_15679);
or U20534 (N_20534,N_14024,N_16680);
and U20535 (N_20535,N_13180,N_14061);
nand U20536 (N_20536,N_13404,N_12514);
or U20537 (N_20537,N_14582,N_16728);
nor U20538 (N_20538,N_16977,N_13187);
nor U20539 (N_20539,N_15555,N_13115);
and U20540 (N_20540,N_15800,N_13855);
nor U20541 (N_20541,N_17564,N_17356);
and U20542 (N_20542,N_17854,N_17645);
or U20543 (N_20543,N_12142,N_17851);
nand U20544 (N_20544,N_16317,N_16305);
nor U20545 (N_20545,N_15568,N_13821);
and U20546 (N_20546,N_12501,N_12487);
or U20547 (N_20547,N_17241,N_15731);
xnor U20548 (N_20548,N_14830,N_12239);
nor U20549 (N_20549,N_15062,N_14585);
and U20550 (N_20550,N_13310,N_12906);
nor U20551 (N_20551,N_14506,N_14073);
nor U20552 (N_20552,N_12480,N_12197);
xor U20553 (N_20553,N_12975,N_16501);
and U20554 (N_20554,N_12195,N_17585);
and U20555 (N_20555,N_17074,N_14841);
nand U20556 (N_20556,N_16438,N_15326);
and U20557 (N_20557,N_12945,N_15764);
xnor U20558 (N_20558,N_17863,N_14478);
xor U20559 (N_20559,N_14451,N_15273);
or U20560 (N_20560,N_16071,N_12639);
nand U20561 (N_20561,N_16525,N_17495);
and U20562 (N_20562,N_16866,N_14284);
nor U20563 (N_20563,N_17533,N_16181);
and U20564 (N_20564,N_13642,N_14466);
or U20565 (N_20565,N_17761,N_16905);
xnor U20566 (N_20566,N_16074,N_14197);
or U20567 (N_20567,N_13808,N_16222);
xor U20568 (N_20568,N_16533,N_12526);
nor U20569 (N_20569,N_13661,N_14914);
and U20570 (N_20570,N_15013,N_12992);
nand U20571 (N_20571,N_16407,N_14883);
nor U20572 (N_20572,N_16004,N_13723);
or U20573 (N_20573,N_15521,N_14035);
nor U20574 (N_20574,N_13729,N_17513);
nand U20575 (N_20575,N_14008,N_17960);
xor U20576 (N_20576,N_13554,N_12812);
nand U20577 (N_20577,N_16712,N_17796);
nand U20578 (N_20578,N_13113,N_13895);
and U20579 (N_20579,N_16355,N_13775);
nand U20580 (N_20580,N_12305,N_14781);
or U20581 (N_20581,N_14412,N_12771);
nor U20582 (N_20582,N_14104,N_15688);
and U20583 (N_20583,N_12512,N_12625);
or U20584 (N_20584,N_17490,N_15135);
xor U20585 (N_20585,N_15801,N_15449);
and U20586 (N_20586,N_14946,N_13782);
or U20587 (N_20587,N_14426,N_12596);
and U20588 (N_20588,N_15959,N_12350);
xor U20589 (N_20589,N_14786,N_15699);
xor U20590 (N_20590,N_17505,N_13468);
xnor U20591 (N_20591,N_17901,N_16690);
nand U20592 (N_20592,N_14408,N_17578);
and U20593 (N_20593,N_17287,N_15265);
nor U20594 (N_20594,N_14504,N_17650);
xnor U20595 (N_20595,N_16123,N_14817);
and U20596 (N_20596,N_16085,N_13353);
nor U20597 (N_20597,N_12949,N_17057);
nor U20598 (N_20598,N_17095,N_16681);
nand U20599 (N_20599,N_14190,N_17618);
xor U20600 (N_20600,N_12475,N_14315);
or U20601 (N_20601,N_17848,N_16128);
and U20602 (N_20602,N_13600,N_17999);
or U20603 (N_20603,N_15897,N_14744);
xor U20604 (N_20604,N_17216,N_14814);
xor U20605 (N_20605,N_16821,N_15325);
and U20606 (N_20606,N_16572,N_17842);
or U20607 (N_20607,N_15745,N_16753);
and U20608 (N_20608,N_17827,N_13118);
nand U20609 (N_20609,N_17070,N_12597);
nor U20610 (N_20610,N_12136,N_15966);
nand U20611 (N_20611,N_14984,N_17939);
and U20612 (N_20612,N_17145,N_15816);
and U20613 (N_20613,N_15213,N_16701);
or U20614 (N_20614,N_12479,N_13960);
or U20615 (N_20615,N_14891,N_15099);
or U20616 (N_20616,N_15993,N_16333);
xor U20617 (N_20617,N_15357,N_15840);
nor U20618 (N_20618,N_17713,N_17932);
nor U20619 (N_20619,N_15080,N_12393);
or U20620 (N_20620,N_13666,N_15870);
xor U20621 (N_20621,N_16167,N_14018);
nand U20622 (N_20622,N_14060,N_13147);
xnor U20623 (N_20623,N_15031,N_12954);
and U20624 (N_20624,N_15684,N_12859);
nor U20625 (N_20625,N_15220,N_17199);
nand U20626 (N_20626,N_12185,N_16241);
nand U20627 (N_20627,N_16860,N_17053);
or U20628 (N_20628,N_14768,N_14199);
and U20629 (N_20629,N_17400,N_13521);
and U20630 (N_20630,N_16400,N_13496);
xor U20631 (N_20631,N_17468,N_16016);
nor U20632 (N_20632,N_16076,N_15887);
xnor U20633 (N_20633,N_16928,N_17398);
and U20634 (N_20634,N_14738,N_13074);
xor U20635 (N_20635,N_13806,N_12435);
or U20636 (N_20636,N_12084,N_13615);
xnor U20637 (N_20637,N_14736,N_15788);
or U20638 (N_20638,N_15483,N_16386);
nand U20639 (N_20639,N_17937,N_14063);
nand U20640 (N_20640,N_14344,N_12871);
nand U20641 (N_20641,N_14062,N_17695);
nand U20642 (N_20642,N_17642,N_13981);
nand U20643 (N_20643,N_16643,N_15165);
or U20644 (N_20644,N_12522,N_14559);
and U20645 (N_20645,N_16686,N_15780);
xor U20646 (N_20646,N_13948,N_12682);
nand U20647 (N_20647,N_15998,N_13966);
xor U20648 (N_20648,N_17388,N_12701);
or U20649 (N_20649,N_14807,N_14971);
nor U20650 (N_20650,N_15593,N_12092);
nand U20651 (N_20651,N_13059,N_13799);
nor U20652 (N_20652,N_13641,N_13156);
nand U20653 (N_20653,N_17197,N_12111);
nand U20654 (N_20654,N_12630,N_16865);
nand U20655 (N_20655,N_12672,N_14745);
xnor U20656 (N_20656,N_17700,N_15379);
and U20657 (N_20657,N_13371,N_15267);
nor U20658 (N_20658,N_15448,N_17992);
nor U20659 (N_20659,N_15383,N_12869);
nor U20660 (N_20660,N_13226,N_17602);
and U20661 (N_20661,N_12555,N_15000);
or U20662 (N_20662,N_14025,N_13128);
and U20663 (N_20663,N_13730,N_16210);
or U20664 (N_20664,N_15363,N_13850);
nand U20665 (N_20665,N_12905,N_14406);
xnor U20666 (N_20666,N_16136,N_14398);
and U20667 (N_20667,N_17674,N_13567);
or U20668 (N_20668,N_17387,N_15871);
nor U20669 (N_20669,N_16814,N_12690);
xnor U20670 (N_20670,N_17079,N_16385);
xor U20671 (N_20671,N_17228,N_15547);
nand U20672 (N_20672,N_15418,N_17730);
nand U20673 (N_20673,N_15540,N_16721);
or U20674 (N_20674,N_16532,N_15536);
nand U20675 (N_20675,N_15539,N_12324);
xnor U20676 (N_20676,N_14387,N_14626);
xor U20677 (N_20677,N_16703,N_17601);
or U20678 (N_20678,N_13696,N_12952);
nor U20679 (N_20679,N_13589,N_16042);
and U20680 (N_20680,N_16970,N_17262);
or U20681 (N_20681,N_16679,N_12212);
and U20682 (N_20682,N_15681,N_14685);
and U20683 (N_20683,N_15677,N_17985);
xnor U20684 (N_20684,N_17894,N_13430);
nand U20685 (N_20685,N_14718,N_17056);
and U20686 (N_20686,N_17131,N_17260);
nor U20687 (N_20687,N_17656,N_17712);
nand U20688 (N_20688,N_17596,N_15415);
xor U20689 (N_20689,N_12351,N_16858);
nand U20690 (N_20690,N_16829,N_16126);
xnor U20691 (N_20691,N_13139,N_13157);
and U20692 (N_20692,N_16087,N_12474);
and U20693 (N_20693,N_12598,N_14705);
xor U20694 (N_20694,N_12677,N_14756);
or U20695 (N_20695,N_14520,N_14244);
or U20696 (N_20696,N_12304,N_13894);
xor U20697 (N_20697,N_12498,N_16893);
xnor U20698 (N_20698,N_17857,N_14388);
nor U20699 (N_20699,N_14450,N_17576);
and U20700 (N_20700,N_17635,N_14337);
and U20701 (N_20701,N_14799,N_15984);
xor U20702 (N_20702,N_13393,N_17741);
or U20703 (N_20703,N_16036,N_17178);
nand U20704 (N_20704,N_15056,N_14960);
or U20705 (N_20705,N_13021,N_15344);
or U20706 (N_20706,N_17965,N_15986);
or U20707 (N_20707,N_15098,N_14996);
nand U20708 (N_20708,N_15291,N_16247);
nand U20709 (N_20709,N_17927,N_15890);
nor U20710 (N_20710,N_17529,N_15117);
nor U20711 (N_20711,N_17242,N_17333);
or U20712 (N_20712,N_14383,N_14274);
or U20713 (N_20713,N_12410,N_12030);
xor U20714 (N_20714,N_13296,N_16840);
xnor U20715 (N_20715,N_13236,N_16124);
xor U20716 (N_20716,N_12889,N_15823);
nand U20717 (N_20717,N_12729,N_16227);
nor U20718 (N_20718,N_13708,N_13809);
nor U20719 (N_20719,N_12218,N_16755);
or U20720 (N_20720,N_13985,N_13224);
nand U20721 (N_20721,N_14658,N_14803);
nand U20722 (N_20722,N_12285,N_13436);
nand U20723 (N_20723,N_15246,N_16142);
xnor U20724 (N_20724,N_13148,N_12469);
nor U20725 (N_20725,N_17900,N_13370);
or U20726 (N_20726,N_15623,N_16955);
xor U20727 (N_20727,N_14000,N_12747);
nor U20728 (N_20728,N_15812,N_14064);
xnor U20729 (N_20729,N_16472,N_17780);
or U20730 (N_20730,N_13847,N_14639);
nand U20731 (N_20731,N_16280,N_15519);
nor U20732 (N_20732,N_17510,N_17600);
nand U20733 (N_20733,N_13493,N_16802);
nand U20734 (N_20734,N_12093,N_12179);
or U20735 (N_20735,N_13715,N_14998);
or U20736 (N_20736,N_16801,N_12558);
and U20737 (N_20737,N_14787,N_17392);
nand U20738 (N_20738,N_14248,N_16369);
or U20739 (N_20739,N_13950,N_15510);
or U20740 (N_20740,N_17023,N_17708);
xnor U20741 (N_20741,N_16312,N_12605);
or U20742 (N_20742,N_17347,N_12679);
or U20743 (N_20743,N_16670,N_16245);
nand U20744 (N_20744,N_16781,N_15992);
and U20745 (N_20745,N_12521,N_14178);
and U20746 (N_20746,N_14975,N_17592);
nor U20747 (N_20747,N_16530,N_17534);
xor U20748 (N_20748,N_14836,N_13067);
nand U20749 (N_20749,N_13033,N_15057);
nor U20750 (N_20750,N_12934,N_16176);
nand U20751 (N_20751,N_15101,N_12284);
xor U20752 (N_20752,N_12440,N_16665);
or U20753 (N_20753,N_16676,N_12814);
and U20754 (N_20754,N_16010,N_16996);
nand U20755 (N_20755,N_16855,N_14272);
and U20756 (N_20756,N_17748,N_16034);
xor U20757 (N_20757,N_16078,N_17066);
nand U20758 (N_20758,N_17655,N_17465);
nor U20759 (N_20759,N_13975,N_17781);
xor U20760 (N_20760,N_13958,N_15186);
xor U20761 (N_20761,N_13050,N_12191);
or U20762 (N_20762,N_13089,N_13415);
nor U20763 (N_20763,N_14990,N_15204);
or U20764 (N_20764,N_16141,N_17202);
nand U20765 (N_20765,N_15232,N_17098);
xnor U20766 (N_20766,N_14497,N_15067);
nor U20767 (N_20767,N_12422,N_16102);
or U20768 (N_20768,N_12756,N_13054);
nand U20769 (N_20769,N_15244,N_13741);
nor U20770 (N_20770,N_14302,N_12269);
or U20771 (N_20771,N_14577,N_12242);
nor U20772 (N_20772,N_16617,N_16852);
and U20773 (N_20773,N_12146,N_13197);
nor U20774 (N_20774,N_16848,N_13175);
nor U20775 (N_20775,N_16114,N_16143);
nand U20776 (N_20776,N_17115,N_15202);
nor U20777 (N_20777,N_14788,N_12272);
nand U20778 (N_20778,N_17373,N_12051);
nand U20779 (N_20779,N_14728,N_17777);
and U20780 (N_20780,N_12765,N_14206);
nand U20781 (N_20781,N_13681,N_12397);
nor U20782 (N_20782,N_14150,N_17024);
or U20783 (N_20783,N_17440,N_13524);
or U20784 (N_20784,N_14755,N_17487);
nor U20785 (N_20785,N_12099,N_15317);
xnor U20786 (N_20786,N_16806,N_16153);
and U20787 (N_20787,N_15931,N_15258);
nand U20788 (N_20788,N_13523,N_14363);
nand U20789 (N_20789,N_14780,N_15009);
and U20790 (N_20790,N_13127,N_13704);
and U20791 (N_20791,N_15059,N_14804);
nor U20792 (N_20792,N_12138,N_16672);
xnor U20793 (N_20793,N_15433,N_15721);
nand U20794 (N_20794,N_14531,N_15719);
xnor U20795 (N_20795,N_15585,N_16772);
and U20796 (N_20796,N_16267,N_12135);
nor U20797 (N_20797,N_16752,N_14215);
and U20798 (N_20798,N_15717,N_12877);
xor U20799 (N_20799,N_12581,N_16583);
nand U20800 (N_20800,N_13653,N_12876);
nand U20801 (N_20801,N_13623,N_16857);
or U20802 (N_20802,N_14569,N_12412);
or U20803 (N_20803,N_17987,N_12582);
nor U20804 (N_20804,N_17081,N_13062);
or U20805 (N_20805,N_16863,N_12821);
nor U20806 (N_20806,N_12186,N_16529);
or U20807 (N_20807,N_16268,N_13713);
xnor U20808 (N_20808,N_13891,N_17184);
and U20809 (N_20809,N_15892,N_12026);
nand U20810 (N_20810,N_13348,N_12817);
nor U20811 (N_20811,N_14081,N_14778);
and U20812 (N_20812,N_14013,N_14702);
and U20813 (N_20813,N_17666,N_13722);
nand U20814 (N_20814,N_17579,N_15476);
nor U20815 (N_20815,N_17955,N_15965);
or U20816 (N_20816,N_16719,N_14970);
nand U20817 (N_20817,N_12461,N_15440);
nand U20818 (N_20818,N_16419,N_14301);
and U20819 (N_20819,N_15083,N_13546);
nand U20820 (N_20820,N_13518,N_15588);
and U20821 (N_20821,N_15368,N_16534);
nand U20822 (N_20822,N_13276,N_12778);
or U20823 (N_20823,N_14250,N_16361);
nor U20824 (N_20824,N_14243,N_15188);
nand U20825 (N_20825,N_13640,N_14917);
or U20826 (N_20826,N_16233,N_14706);
xor U20827 (N_20827,N_17661,N_12413);
or U20828 (N_20828,N_13051,N_14552);
nor U20829 (N_20829,N_17891,N_17808);
xnor U20830 (N_20830,N_12766,N_17839);
nand U20831 (N_20831,N_16815,N_12789);
and U20832 (N_20832,N_12161,N_13588);
xnor U20833 (N_20833,N_12607,N_17404);
nand U20834 (N_20834,N_14053,N_15944);
or U20835 (N_20835,N_12726,N_17097);
or U20836 (N_20836,N_15832,N_17609);
nand U20837 (N_20837,N_17567,N_17771);
nor U20838 (N_20838,N_15932,N_17971);
or U20839 (N_20839,N_15342,N_15927);
nand U20840 (N_20840,N_12559,N_12885);
nand U20841 (N_20841,N_13263,N_12119);
xnor U20842 (N_20842,N_17826,N_15084);
and U20843 (N_20843,N_17128,N_17917);
xor U20844 (N_20844,N_12622,N_17284);
and U20845 (N_20845,N_17472,N_16952);
xnor U20846 (N_20846,N_13406,N_15727);
and U20847 (N_20847,N_17933,N_17776);
and U20848 (N_20848,N_15760,N_17180);
and U20849 (N_20849,N_13956,N_15949);
and U20850 (N_20850,N_17783,N_15902);
nor U20851 (N_20851,N_14711,N_12813);
and U20852 (N_20852,N_15003,N_16682);
nand U20853 (N_20853,N_12055,N_15824);
nand U20854 (N_20854,N_14039,N_13146);
and U20855 (N_20855,N_14813,N_12831);
and U20856 (N_20856,N_13880,N_17755);
nor U20857 (N_20857,N_16418,N_15509);
and U20858 (N_20858,N_12686,N_15724);
nor U20859 (N_20859,N_13813,N_17935);
and U20860 (N_20860,N_12309,N_16600);
xor U20861 (N_20861,N_12294,N_12717);
and U20862 (N_20862,N_12938,N_12852);
nand U20863 (N_20863,N_12780,N_15855);
xnor U20864 (N_20864,N_15566,N_15505);
xnor U20865 (N_20865,N_15572,N_13362);
and U20866 (N_20866,N_17227,N_16265);
and U20867 (N_20867,N_15757,N_16477);
nor U20868 (N_20868,N_16196,N_14578);
nand U20869 (N_20869,N_16744,N_14251);
nand U20870 (N_20870,N_17156,N_15401);
xnor U20871 (N_20871,N_13284,N_13056);
nor U20872 (N_20872,N_17526,N_12302);
nand U20873 (N_20873,N_12829,N_16936);
xor U20874 (N_20874,N_16884,N_15759);
xnor U20875 (N_20875,N_15844,N_17920);
or U20876 (N_20876,N_17361,N_17432);
xnor U20877 (N_20877,N_17467,N_17615);
and U20878 (N_20878,N_15596,N_16506);
xor U20879 (N_20879,N_16024,N_15341);
nand U20880 (N_20880,N_12746,N_16615);
and U20881 (N_20881,N_14855,N_16598);
or U20882 (N_20882,N_12110,N_14111);
and U20883 (N_20883,N_13814,N_17544);
xor U20884 (N_20884,N_15706,N_14515);
or U20885 (N_20885,N_13433,N_15251);
nand U20886 (N_20886,N_14483,N_16748);
and U20887 (N_20887,N_15876,N_13357);
xnor U20888 (N_20888,N_15875,N_15153);
and U20889 (N_20889,N_15178,N_15276);
or U20890 (N_20890,N_17019,N_16937);
xor U20891 (N_20891,N_16103,N_13300);
xnor U20892 (N_20892,N_13419,N_14189);
and U20893 (N_20893,N_12355,N_14330);
and U20894 (N_20894,N_13525,N_14895);
xor U20895 (N_20895,N_16417,N_17061);
or U20896 (N_20896,N_16339,N_16264);
xnor U20897 (N_20897,N_13517,N_13167);
nor U20898 (N_20898,N_12001,N_13376);
and U20899 (N_20899,N_14955,N_16804);
nor U20900 (N_20900,N_12383,N_12385);
and U20901 (N_20901,N_17076,N_15261);
or U20902 (N_20902,N_12549,N_12444);
nand U20903 (N_20903,N_15474,N_16409);
nand U20904 (N_20904,N_12424,N_16641);
xor U20905 (N_20905,N_14082,N_16461);
nor U20906 (N_20906,N_13454,N_13953);
nor U20907 (N_20907,N_12794,N_12046);
or U20908 (N_20908,N_16462,N_16292);
and U20909 (N_20909,N_12314,N_13327);
or U20910 (N_20910,N_12421,N_16494);
xnor U20911 (N_20911,N_15885,N_13379);
xor U20912 (N_20912,N_17820,N_17514);
nand U20913 (N_20913,N_12112,N_14812);
or U20914 (N_20914,N_12016,N_14544);
or U20915 (N_20915,N_16491,N_14731);
or U20916 (N_20916,N_13290,N_15042);
nor U20917 (N_20917,N_16156,N_12404);
or U20918 (N_20918,N_16338,N_14563);
and U20919 (N_20919,N_13315,N_16007);
nor U20920 (N_20920,N_13733,N_17889);
nor U20921 (N_20921,N_14204,N_17869);
nand U20922 (N_20922,N_17739,N_15404);
nand U20923 (N_20923,N_17273,N_14785);
nor U20924 (N_20924,N_12675,N_17314);
and U20925 (N_20925,N_13622,N_12308);
xnor U20926 (N_20926,N_12961,N_15829);
xnor U20927 (N_20927,N_14954,N_16453);
and U20928 (N_20928,N_17967,N_17390);
or U20929 (N_20929,N_13859,N_12754);
and U20930 (N_20930,N_15063,N_12534);
or U20931 (N_20931,N_14058,N_12236);
nand U20932 (N_20932,N_14893,N_17077);
nand U20933 (N_20933,N_13727,N_12281);
nor U20934 (N_20934,N_13095,N_12969);
and U20935 (N_20935,N_13058,N_12748);
or U20936 (N_20936,N_17328,N_13457);
nor U20937 (N_20937,N_17229,N_17994);
or U20938 (N_20938,N_15247,N_15863);
xor U20939 (N_20939,N_15069,N_12296);
nor U20940 (N_20940,N_13797,N_17486);
nor U20941 (N_20941,N_14574,N_14312);
or U20942 (N_20942,N_12183,N_13780);
nor U20943 (N_20943,N_17636,N_13754);
or U20944 (N_20944,N_12224,N_15442);
nand U20945 (N_20945,N_13004,N_16591);
nand U20946 (N_20946,N_13706,N_13378);
xnor U20947 (N_20947,N_16998,N_15130);
and U20948 (N_20948,N_14418,N_13409);
or U20949 (N_20949,N_15005,N_13105);
or U20950 (N_20950,N_15867,N_15245);
nor U20951 (N_20951,N_13337,N_15162);
or U20952 (N_20952,N_15789,N_15639);
nand U20953 (N_20953,N_17093,N_16011);
nand U20954 (N_20954,N_13743,N_17587);
and U20955 (N_20955,N_12845,N_16260);
or U20956 (N_20956,N_12364,N_17265);
xor U20957 (N_20957,N_17417,N_16611);
or U20958 (N_20958,N_12960,N_15259);
xor U20959 (N_20959,N_16064,N_16498);
and U20960 (N_20960,N_12137,N_15820);
nand U20961 (N_20961,N_17584,N_15740);
nand U20962 (N_20962,N_13980,N_12874);
xor U20963 (N_20963,N_16225,N_13629);
nand U20964 (N_20964,N_13777,N_12466);
nand U20965 (N_20965,N_14182,N_14065);
xor U20966 (N_20966,N_12012,N_14492);
or U20967 (N_20967,N_14083,N_13874);
or U20968 (N_20968,N_12818,N_13017);
nor U20969 (N_20969,N_12044,N_16876);
nand U20970 (N_20970,N_12464,N_12590);
nand U20971 (N_20971,N_13107,N_12621);
nor U20972 (N_20972,N_15212,N_14995);
or U20973 (N_20973,N_15388,N_17590);
and U20974 (N_20974,N_17470,N_14709);
nor U20975 (N_20975,N_16229,N_13481);
and U20976 (N_20976,N_12034,N_13660);
xor U20977 (N_20977,N_16390,N_12500);
or U20978 (N_20978,N_17395,N_12716);
and U20979 (N_20979,N_12902,N_15103);
nand U20980 (N_20980,N_13238,N_14943);
nand U20981 (N_20981,N_14610,N_14815);
nor U20982 (N_20982,N_13938,N_15150);
nor U20983 (N_20983,N_15822,N_16189);
or U20984 (N_20984,N_12673,N_14441);
and U20985 (N_20985,N_13844,N_14006);
xnor U20986 (N_20986,N_13022,N_13505);
xnor U20987 (N_20987,N_16688,N_12695);
nor U20988 (N_20988,N_15828,N_14326);
nor U20989 (N_20989,N_17396,N_12755);
nand U20990 (N_20990,N_13773,N_12004);
nor U20991 (N_20991,N_12750,N_14293);
xnor U20992 (N_20992,N_13991,N_14537);
and U20993 (N_20993,N_12629,N_14677);
and U20994 (N_20994,N_13701,N_16383);
or U20995 (N_20995,N_12744,N_12447);
nand U20996 (N_20996,N_16334,N_17313);
xor U20997 (N_20997,N_16990,N_16737);
xnor U20998 (N_20998,N_13258,N_14290);
xor U20999 (N_20999,N_15495,N_14837);
xnor U21000 (N_21000,N_14665,N_13978);
nand U21001 (N_21001,N_14030,N_12513);
and U21002 (N_21002,N_12163,N_13709);
or U21003 (N_21003,N_17841,N_13237);
xor U21004 (N_21004,N_17358,N_12446);
nor U21005 (N_21005,N_14260,N_15970);
or U21006 (N_21006,N_14515,N_12447);
nand U21007 (N_21007,N_14811,N_13438);
nand U21008 (N_21008,N_12072,N_12519);
or U21009 (N_21009,N_15410,N_17795);
xnor U21010 (N_21010,N_13256,N_12808);
and U21011 (N_21011,N_17175,N_17270);
nand U21012 (N_21012,N_12390,N_17698);
nor U21013 (N_21013,N_13343,N_15732);
nor U21014 (N_21014,N_17771,N_12218);
and U21015 (N_21015,N_15364,N_15633);
nand U21016 (N_21016,N_16579,N_14743);
and U21017 (N_21017,N_16985,N_13498);
and U21018 (N_21018,N_16355,N_14016);
xnor U21019 (N_21019,N_14132,N_16601);
nand U21020 (N_21020,N_14271,N_15139);
nor U21021 (N_21021,N_12297,N_13673);
nor U21022 (N_21022,N_13525,N_17922);
xnor U21023 (N_21023,N_16058,N_16910);
nand U21024 (N_21024,N_16577,N_15766);
xor U21025 (N_21025,N_14825,N_17287);
xnor U21026 (N_21026,N_17351,N_15586);
and U21027 (N_21027,N_15923,N_13393);
and U21028 (N_21028,N_17412,N_12290);
xnor U21029 (N_21029,N_15781,N_12034);
nand U21030 (N_21030,N_16644,N_13389);
nand U21031 (N_21031,N_12265,N_17319);
xnor U21032 (N_21032,N_13507,N_14250);
and U21033 (N_21033,N_16412,N_15586);
and U21034 (N_21034,N_15472,N_15099);
xor U21035 (N_21035,N_16575,N_12905);
or U21036 (N_21036,N_17405,N_15259);
xor U21037 (N_21037,N_14489,N_14437);
and U21038 (N_21038,N_14832,N_14359);
or U21039 (N_21039,N_14943,N_14208);
and U21040 (N_21040,N_15047,N_13034);
or U21041 (N_21041,N_13127,N_16745);
nor U21042 (N_21042,N_14798,N_15717);
and U21043 (N_21043,N_16052,N_14639);
xor U21044 (N_21044,N_14531,N_15467);
and U21045 (N_21045,N_17993,N_17316);
nand U21046 (N_21046,N_15343,N_12491);
and U21047 (N_21047,N_17416,N_14238);
nand U21048 (N_21048,N_17707,N_13952);
or U21049 (N_21049,N_13879,N_14832);
nand U21050 (N_21050,N_17869,N_14093);
and U21051 (N_21051,N_14794,N_13986);
and U21052 (N_21052,N_17934,N_17061);
nor U21053 (N_21053,N_15437,N_12205);
nand U21054 (N_21054,N_12406,N_14436);
and U21055 (N_21055,N_14509,N_16101);
nor U21056 (N_21056,N_13859,N_15920);
and U21057 (N_21057,N_12123,N_14832);
nor U21058 (N_21058,N_14629,N_13365);
nor U21059 (N_21059,N_13423,N_12563);
nor U21060 (N_21060,N_17927,N_17250);
or U21061 (N_21061,N_13735,N_15414);
or U21062 (N_21062,N_14337,N_13909);
or U21063 (N_21063,N_14379,N_12565);
nand U21064 (N_21064,N_17509,N_13272);
and U21065 (N_21065,N_16207,N_13962);
or U21066 (N_21066,N_15307,N_12540);
nor U21067 (N_21067,N_13054,N_15568);
nor U21068 (N_21068,N_15284,N_15202);
xor U21069 (N_21069,N_12477,N_14546);
xor U21070 (N_21070,N_13117,N_12382);
or U21071 (N_21071,N_15445,N_12032);
or U21072 (N_21072,N_17703,N_17038);
xnor U21073 (N_21073,N_13342,N_16745);
xor U21074 (N_21074,N_14971,N_13100);
xnor U21075 (N_21075,N_16466,N_17741);
nor U21076 (N_21076,N_14181,N_12517);
nand U21077 (N_21077,N_13651,N_16436);
or U21078 (N_21078,N_13365,N_14689);
nand U21079 (N_21079,N_15797,N_15545);
nand U21080 (N_21080,N_16847,N_17890);
nand U21081 (N_21081,N_14127,N_17126);
and U21082 (N_21082,N_17567,N_13913);
nand U21083 (N_21083,N_17887,N_14631);
nand U21084 (N_21084,N_14024,N_17172);
nor U21085 (N_21085,N_12150,N_13312);
or U21086 (N_21086,N_12810,N_13523);
and U21087 (N_21087,N_14593,N_14005);
nor U21088 (N_21088,N_17777,N_15580);
nor U21089 (N_21089,N_13268,N_13510);
and U21090 (N_21090,N_17012,N_17714);
xnor U21091 (N_21091,N_13166,N_17878);
nand U21092 (N_21092,N_13810,N_13726);
xnor U21093 (N_21093,N_17342,N_14369);
nand U21094 (N_21094,N_17799,N_17540);
nand U21095 (N_21095,N_14844,N_16441);
nand U21096 (N_21096,N_15334,N_13583);
nand U21097 (N_21097,N_13689,N_17732);
xnor U21098 (N_21098,N_16193,N_14374);
nor U21099 (N_21099,N_15062,N_14264);
nand U21100 (N_21100,N_12277,N_14698);
nor U21101 (N_21101,N_13454,N_13699);
and U21102 (N_21102,N_13087,N_17123);
nand U21103 (N_21103,N_15576,N_16214);
nor U21104 (N_21104,N_14875,N_14599);
nand U21105 (N_21105,N_16535,N_16219);
and U21106 (N_21106,N_16582,N_14366);
nor U21107 (N_21107,N_13409,N_13473);
nand U21108 (N_21108,N_17004,N_12231);
nand U21109 (N_21109,N_12024,N_17493);
xor U21110 (N_21110,N_12461,N_15066);
xor U21111 (N_21111,N_12841,N_17686);
xnor U21112 (N_21112,N_16008,N_13895);
nand U21113 (N_21113,N_12773,N_15066);
nor U21114 (N_21114,N_16884,N_15194);
and U21115 (N_21115,N_17799,N_14800);
nand U21116 (N_21116,N_15568,N_13313);
and U21117 (N_21117,N_17442,N_13715);
or U21118 (N_21118,N_14236,N_12200);
xnor U21119 (N_21119,N_13151,N_13948);
or U21120 (N_21120,N_13273,N_13833);
or U21121 (N_21121,N_12603,N_14195);
or U21122 (N_21122,N_12458,N_14798);
and U21123 (N_21123,N_15481,N_17532);
nand U21124 (N_21124,N_15133,N_15095);
nand U21125 (N_21125,N_13776,N_14220);
nand U21126 (N_21126,N_14603,N_16305);
nand U21127 (N_21127,N_14720,N_14221);
and U21128 (N_21128,N_13779,N_15291);
nor U21129 (N_21129,N_15635,N_16605);
or U21130 (N_21130,N_16258,N_16764);
or U21131 (N_21131,N_17703,N_15580);
nand U21132 (N_21132,N_14375,N_14873);
and U21133 (N_21133,N_15881,N_15385);
nand U21134 (N_21134,N_17596,N_14723);
or U21135 (N_21135,N_12786,N_17115);
nand U21136 (N_21136,N_16751,N_14071);
xnor U21137 (N_21137,N_12788,N_14994);
or U21138 (N_21138,N_17763,N_12476);
or U21139 (N_21139,N_14493,N_17728);
nor U21140 (N_21140,N_13351,N_14984);
or U21141 (N_21141,N_14579,N_12317);
and U21142 (N_21142,N_15396,N_16730);
xnor U21143 (N_21143,N_13910,N_14191);
or U21144 (N_21144,N_13293,N_17377);
and U21145 (N_21145,N_15777,N_16446);
nand U21146 (N_21146,N_15685,N_15219);
nor U21147 (N_21147,N_13823,N_16534);
nand U21148 (N_21148,N_13556,N_17044);
or U21149 (N_21149,N_15584,N_14192);
nand U21150 (N_21150,N_13520,N_17084);
or U21151 (N_21151,N_15290,N_16559);
or U21152 (N_21152,N_15453,N_14280);
xor U21153 (N_21153,N_14053,N_14327);
and U21154 (N_21154,N_17843,N_15839);
nor U21155 (N_21155,N_16706,N_12481);
and U21156 (N_21156,N_13324,N_14755);
nand U21157 (N_21157,N_16929,N_17674);
or U21158 (N_21158,N_13663,N_12162);
xor U21159 (N_21159,N_14206,N_16312);
and U21160 (N_21160,N_13366,N_14633);
xnor U21161 (N_21161,N_14424,N_15610);
or U21162 (N_21162,N_16095,N_14777);
or U21163 (N_21163,N_14695,N_16215);
and U21164 (N_21164,N_16953,N_15780);
and U21165 (N_21165,N_16201,N_16254);
or U21166 (N_21166,N_15693,N_14953);
xnor U21167 (N_21167,N_12220,N_12798);
and U21168 (N_21168,N_12947,N_17578);
or U21169 (N_21169,N_13522,N_15965);
or U21170 (N_21170,N_15024,N_15853);
xor U21171 (N_21171,N_12941,N_16630);
nor U21172 (N_21172,N_16890,N_15235);
or U21173 (N_21173,N_14383,N_15414);
or U21174 (N_21174,N_12689,N_13150);
and U21175 (N_21175,N_13454,N_16485);
and U21176 (N_21176,N_15147,N_14287);
nand U21177 (N_21177,N_13186,N_12066);
xor U21178 (N_21178,N_13145,N_14407);
and U21179 (N_21179,N_16619,N_14061);
xnor U21180 (N_21180,N_12916,N_12471);
nor U21181 (N_21181,N_12226,N_12467);
nor U21182 (N_21182,N_15526,N_12089);
nor U21183 (N_21183,N_14280,N_17307);
or U21184 (N_21184,N_16656,N_14349);
nand U21185 (N_21185,N_15702,N_14494);
nor U21186 (N_21186,N_17788,N_15559);
nor U21187 (N_21187,N_14911,N_16929);
xor U21188 (N_21188,N_13876,N_17453);
nor U21189 (N_21189,N_12071,N_15144);
nand U21190 (N_21190,N_13623,N_16622);
and U21191 (N_21191,N_13573,N_14849);
nor U21192 (N_21192,N_15617,N_16771);
nand U21193 (N_21193,N_15718,N_13445);
xnor U21194 (N_21194,N_15300,N_17708);
or U21195 (N_21195,N_14261,N_15070);
and U21196 (N_21196,N_12257,N_17300);
nor U21197 (N_21197,N_12165,N_14351);
and U21198 (N_21198,N_14461,N_17389);
xor U21199 (N_21199,N_15730,N_16622);
and U21200 (N_21200,N_12141,N_17709);
or U21201 (N_21201,N_16210,N_17024);
and U21202 (N_21202,N_16162,N_16786);
and U21203 (N_21203,N_16824,N_16153);
xnor U21204 (N_21204,N_13200,N_14623);
xnor U21205 (N_21205,N_15414,N_15686);
nor U21206 (N_21206,N_17575,N_12429);
xnor U21207 (N_21207,N_13406,N_16388);
and U21208 (N_21208,N_13128,N_17479);
nor U21209 (N_21209,N_14500,N_15267);
xnor U21210 (N_21210,N_12270,N_17112);
or U21211 (N_21211,N_15935,N_12954);
nor U21212 (N_21212,N_15677,N_16792);
and U21213 (N_21213,N_17602,N_14994);
and U21214 (N_21214,N_13330,N_13026);
xor U21215 (N_21215,N_16436,N_12985);
or U21216 (N_21216,N_16869,N_16089);
xor U21217 (N_21217,N_17313,N_17149);
xnor U21218 (N_21218,N_12393,N_15660);
nor U21219 (N_21219,N_15206,N_16005);
and U21220 (N_21220,N_12725,N_12896);
or U21221 (N_21221,N_15275,N_14393);
or U21222 (N_21222,N_12689,N_15306);
or U21223 (N_21223,N_16722,N_12083);
nand U21224 (N_21224,N_13182,N_12720);
nand U21225 (N_21225,N_14464,N_13918);
nand U21226 (N_21226,N_14971,N_14956);
nor U21227 (N_21227,N_13147,N_13879);
or U21228 (N_21228,N_15519,N_14636);
or U21229 (N_21229,N_16082,N_15801);
or U21230 (N_21230,N_17604,N_15294);
xor U21231 (N_21231,N_13769,N_13898);
nor U21232 (N_21232,N_13789,N_17783);
nor U21233 (N_21233,N_13664,N_17683);
nor U21234 (N_21234,N_13911,N_12386);
xor U21235 (N_21235,N_12545,N_14699);
nor U21236 (N_21236,N_13617,N_12018);
xor U21237 (N_21237,N_17816,N_14733);
and U21238 (N_21238,N_15560,N_17390);
xnor U21239 (N_21239,N_12053,N_16720);
and U21240 (N_21240,N_16377,N_12519);
and U21241 (N_21241,N_17032,N_17925);
xor U21242 (N_21242,N_16469,N_17222);
nor U21243 (N_21243,N_12649,N_12859);
and U21244 (N_21244,N_12836,N_16612);
nand U21245 (N_21245,N_15542,N_12131);
or U21246 (N_21246,N_12537,N_14518);
or U21247 (N_21247,N_16823,N_16585);
nor U21248 (N_21248,N_14701,N_14390);
and U21249 (N_21249,N_12969,N_17459);
nand U21250 (N_21250,N_15967,N_15857);
nor U21251 (N_21251,N_13675,N_13965);
and U21252 (N_21252,N_17060,N_17144);
or U21253 (N_21253,N_16364,N_12015);
nor U21254 (N_21254,N_13769,N_13501);
and U21255 (N_21255,N_14386,N_13273);
or U21256 (N_21256,N_16165,N_17681);
or U21257 (N_21257,N_14449,N_12875);
or U21258 (N_21258,N_16014,N_14254);
and U21259 (N_21259,N_15199,N_17122);
xnor U21260 (N_21260,N_12266,N_15226);
and U21261 (N_21261,N_17242,N_13299);
or U21262 (N_21262,N_17383,N_16016);
and U21263 (N_21263,N_16228,N_14201);
or U21264 (N_21264,N_17543,N_12788);
nor U21265 (N_21265,N_13333,N_16055);
xnor U21266 (N_21266,N_12295,N_15554);
xnor U21267 (N_21267,N_15341,N_14599);
nand U21268 (N_21268,N_17186,N_13597);
xor U21269 (N_21269,N_15437,N_13764);
xnor U21270 (N_21270,N_13390,N_17799);
xnor U21271 (N_21271,N_16331,N_14434);
nand U21272 (N_21272,N_15048,N_16889);
and U21273 (N_21273,N_17536,N_13914);
or U21274 (N_21274,N_12190,N_13673);
xnor U21275 (N_21275,N_13658,N_17330);
nand U21276 (N_21276,N_15260,N_16748);
and U21277 (N_21277,N_17571,N_17770);
nor U21278 (N_21278,N_12270,N_17474);
and U21279 (N_21279,N_12564,N_13131);
nand U21280 (N_21280,N_12296,N_12857);
nor U21281 (N_21281,N_15485,N_15162);
or U21282 (N_21282,N_12414,N_13637);
nor U21283 (N_21283,N_16269,N_12797);
and U21284 (N_21284,N_14219,N_16157);
and U21285 (N_21285,N_14442,N_13753);
xnor U21286 (N_21286,N_16538,N_17890);
nor U21287 (N_21287,N_12967,N_15078);
xnor U21288 (N_21288,N_14861,N_16722);
nor U21289 (N_21289,N_13244,N_12698);
xor U21290 (N_21290,N_16152,N_12660);
nor U21291 (N_21291,N_14944,N_14197);
xnor U21292 (N_21292,N_12861,N_14238);
nand U21293 (N_21293,N_15127,N_17463);
nor U21294 (N_21294,N_15216,N_16911);
or U21295 (N_21295,N_16228,N_12543);
nor U21296 (N_21296,N_15241,N_14723);
xor U21297 (N_21297,N_14829,N_14287);
xnor U21298 (N_21298,N_14496,N_12032);
nor U21299 (N_21299,N_15685,N_15345);
and U21300 (N_21300,N_16761,N_12474);
xor U21301 (N_21301,N_13366,N_15868);
xor U21302 (N_21302,N_16812,N_13826);
nor U21303 (N_21303,N_13317,N_13693);
or U21304 (N_21304,N_12388,N_15817);
nor U21305 (N_21305,N_15926,N_14111);
nor U21306 (N_21306,N_13884,N_14680);
and U21307 (N_21307,N_15129,N_13118);
xor U21308 (N_21308,N_12956,N_15807);
or U21309 (N_21309,N_17836,N_17699);
or U21310 (N_21310,N_17453,N_12481);
or U21311 (N_21311,N_14806,N_14420);
and U21312 (N_21312,N_16100,N_12180);
nor U21313 (N_21313,N_12455,N_13946);
nor U21314 (N_21314,N_15285,N_13218);
xnor U21315 (N_21315,N_14076,N_16775);
and U21316 (N_21316,N_17585,N_15311);
nand U21317 (N_21317,N_17978,N_12632);
nand U21318 (N_21318,N_15992,N_14454);
or U21319 (N_21319,N_16853,N_14221);
nand U21320 (N_21320,N_12122,N_17636);
or U21321 (N_21321,N_14747,N_13179);
nand U21322 (N_21322,N_16257,N_14141);
nor U21323 (N_21323,N_17628,N_15840);
and U21324 (N_21324,N_13144,N_16400);
and U21325 (N_21325,N_16009,N_12905);
nor U21326 (N_21326,N_17289,N_17348);
xnor U21327 (N_21327,N_15355,N_13569);
and U21328 (N_21328,N_14469,N_15232);
nor U21329 (N_21329,N_15224,N_14463);
xnor U21330 (N_21330,N_14200,N_17346);
nand U21331 (N_21331,N_17577,N_14933);
and U21332 (N_21332,N_16431,N_14876);
xor U21333 (N_21333,N_16303,N_12687);
nor U21334 (N_21334,N_13326,N_15290);
and U21335 (N_21335,N_16346,N_16197);
and U21336 (N_21336,N_15892,N_15061);
xnor U21337 (N_21337,N_12940,N_13703);
nand U21338 (N_21338,N_13018,N_13588);
and U21339 (N_21339,N_16800,N_15699);
and U21340 (N_21340,N_16536,N_13951);
or U21341 (N_21341,N_16810,N_12678);
nor U21342 (N_21342,N_16399,N_16042);
nand U21343 (N_21343,N_16398,N_13445);
nand U21344 (N_21344,N_17965,N_13546);
and U21345 (N_21345,N_16346,N_16568);
nor U21346 (N_21346,N_13676,N_13856);
nand U21347 (N_21347,N_16270,N_17957);
nor U21348 (N_21348,N_17682,N_17587);
and U21349 (N_21349,N_14238,N_17936);
and U21350 (N_21350,N_14741,N_14754);
nor U21351 (N_21351,N_13955,N_15697);
nand U21352 (N_21352,N_12975,N_17697);
and U21353 (N_21353,N_12517,N_13914);
nor U21354 (N_21354,N_14373,N_14743);
nor U21355 (N_21355,N_13762,N_16438);
and U21356 (N_21356,N_13791,N_14101);
or U21357 (N_21357,N_14241,N_16626);
or U21358 (N_21358,N_12356,N_16610);
and U21359 (N_21359,N_12028,N_16543);
and U21360 (N_21360,N_15599,N_17121);
nand U21361 (N_21361,N_15583,N_14563);
nand U21362 (N_21362,N_12557,N_17005);
and U21363 (N_21363,N_14022,N_17239);
nor U21364 (N_21364,N_13486,N_16270);
xnor U21365 (N_21365,N_12586,N_15876);
nand U21366 (N_21366,N_12217,N_12382);
nor U21367 (N_21367,N_14024,N_17411);
nand U21368 (N_21368,N_14582,N_15073);
nor U21369 (N_21369,N_12049,N_15062);
and U21370 (N_21370,N_13299,N_16724);
or U21371 (N_21371,N_16580,N_17550);
or U21372 (N_21372,N_12584,N_13809);
or U21373 (N_21373,N_13067,N_17217);
xor U21374 (N_21374,N_15904,N_12635);
xnor U21375 (N_21375,N_12591,N_13607);
nor U21376 (N_21376,N_15347,N_12151);
and U21377 (N_21377,N_12541,N_15979);
or U21378 (N_21378,N_12717,N_13086);
nor U21379 (N_21379,N_16732,N_17237);
and U21380 (N_21380,N_12920,N_13671);
xnor U21381 (N_21381,N_12801,N_12321);
or U21382 (N_21382,N_15681,N_15810);
nand U21383 (N_21383,N_13563,N_17404);
nor U21384 (N_21384,N_17230,N_15953);
nand U21385 (N_21385,N_15271,N_16959);
and U21386 (N_21386,N_13492,N_16903);
xor U21387 (N_21387,N_13908,N_15638);
nor U21388 (N_21388,N_15091,N_12227);
xnor U21389 (N_21389,N_14570,N_13084);
nand U21390 (N_21390,N_16203,N_14520);
and U21391 (N_21391,N_17901,N_13085);
and U21392 (N_21392,N_16194,N_13112);
and U21393 (N_21393,N_16996,N_12265);
and U21394 (N_21394,N_12642,N_12327);
nand U21395 (N_21395,N_17994,N_17949);
or U21396 (N_21396,N_17540,N_15897);
nor U21397 (N_21397,N_14148,N_14183);
nor U21398 (N_21398,N_14283,N_15042);
and U21399 (N_21399,N_17365,N_15101);
nor U21400 (N_21400,N_16623,N_15425);
nand U21401 (N_21401,N_12709,N_13952);
xnor U21402 (N_21402,N_12810,N_13455);
nor U21403 (N_21403,N_12423,N_15080);
xor U21404 (N_21404,N_13562,N_17088);
nand U21405 (N_21405,N_12691,N_16220);
nand U21406 (N_21406,N_17874,N_15192);
nand U21407 (N_21407,N_15121,N_13557);
or U21408 (N_21408,N_14737,N_13097);
xor U21409 (N_21409,N_17114,N_15743);
xnor U21410 (N_21410,N_17973,N_13089);
nor U21411 (N_21411,N_16667,N_12884);
nor U21412 (N_21412,N_14646,N_14772);
nand U21413 (N_21413,N_15909,N_16725);
nor U21414 (N_21414,N_14383,N_15358);
or U21415 (N_21415,N_15174,N_17200);
xnor U21416 (N_21416,N_13291,N_14594);
and U21417 (N_21417,N_12337,N_17619);
and U21418 (N_21418,N_16253,N_12694);
and U21419 (N_21419,N_15675,N_16019);
nand U21420 (N_21420,N_17444,N_17837);
nor U21421 (N_21421,N_13749,N_17189);
xor U21422 (N_21422,N_15146,N_16865);
nand U21423 (N_21423,N_14829,N_14226);
xor U21424 (N_21424,N_16027,N_15487);
nand U21425 (N_21425,N_12215,N_14116);
or U21426 (N_21426,N_14139,N_12684);
nand U21427 (N_21427,N_13017,N_12011);
nand U21428 (N_21428,N_17320,N_17724);
xor U21429 (N_21429,N_17028,N_14506);
nor U21430 (N_21430,N_15349,N_15933);
nor U21431 (N_21431,N_16753,N_17410);
and U21432 (N_21432,N_12655,N_12014);
xnor U21433 (N_21433,N_14554,N_17272);
and U21434 (N_21434,N_15614,N_17730);
xor U21435 (N_21435,N_16782,N_14719);
and U21436 (N_21436,N_16331,N_12410);
or U21437 (N_21437,N_13958,N_17190);
nor U21438 (N_21438,N_17276,N_14230);
or U21439 (N_21439,N_12761,N_17824);
xor U21440 (N_21440,N_12526,N_12294);
nand U21441 (N_21441,N_13761,N_16684);
nand U21442 (N_21442,N_16549,N_17924);
nor U21443 (N_21443,N_12190,N_15183);
nor U21444 (N_21444,N_17686,N_16846);
or U21445 (N_21445,N_15098,N_14913);
and U21446 (N_21446,N_17677,N_15389);
or U21447 (N_21447,N_17181,N_15327);
xor U21448 (N_21448,N_14970,N_14291);
nor U21449 (N_21449,N_15620,N_14451);
or U21450 (N_21450,N_16256,N_17279);
xnor U21451 (N_21451,N_13168,N_15308);
and U21452 (N_21452,N_12754,N_12473);
xnor U21453 (N_21453,N_15704,N_17866);
and U21454 (N_21454,N_16640,N_13261);
and U21455 (N_21455,N_13260,N_16917);
xnor U21456 (N_21456,N_13316,N_17393);
or U21457 (N_21457,N_17795,N_14275);
xnor U21458 (N_21458,N_12197,N_12767);
nand U21459 (N_21459,N_13126,N_17713);
nand U21460 (N_21460,N_13667,N_13686);
or U21461 (N_21461,N_17796,N_13612);
and U21462 (N_21462,N_12224,N_14436);
or U21463 (N_21463,N_14393,N_17827);
or U21464 (N_21464,N_17020,N_17792);
or U21465 (N_21465,N_15281,N_12360);
or U21466 (N_21466,N_13539,N_16189);
or U21467 (N_21467,N_15661,N_14430);
and U21468 (N_21468,N_16510,N_16350);
nand U21469 (N_21469,N_17690,N_17937);
nor U21470 (N_21470,N_12635,N_14613);
xnor U21471 (N_21471,N_12509,N_15848);
or U21472 (N_21472,N_12373,N_14420);
nand U21473 (N_21473,N_14440,N_16345);
or U21474 (N_21474,N_12347,N_15977);
nor U21475 (N_21475,N_17457,N_12525);
nand U21476 (N_21476,N_13759,N_16488);
and U21477 (N_21477,N_13450,N_17738);
nand U21478 (N_21478,N_15838,N_15805);
and U21479 (N_21479,N_14519,N_17730);
nand U21480 (N_21480,N_15885,N_12467);
or U21481 (N_21481,N_17235,N_12444);
or U21482 (N_21482,N_16884,N_13167);
or U21483 (N_21483,N_13611,N_17750);
nand U21484 (N_21484,N_15016,N_15306);
and U21485 (N_21485,N_12254,N_17777);
nand U21486 (N_21486,N_14328,N_17249);
nand U21487 (N_21487,N_17786,N_16767);
and U21488 (N_21488,N_15910,N_16102);
and U21489 (N_21489,N_14623,N_13450);
xor U21490 (N_21490,N_15408,N_14119);
xnor U21491 (N_21491,N_16864,N_13923);
xor U21492 (N_21492,N_16611,N_12369);
and U21493 (N_21493,N_12017,N_14327);
or U21494 (N_21494,N_13403,N_12373);
or U21495 (N_21495,N_12500,N_12675);
xor U21496 (N_21496,N_12480,N_13424);
and U21497 (N_21497,N_16463,N_13696);
xor U21498 (N_21498,N_17685,N_13735);
xnor U21499 (N_21499,N_13858,N_16191);
xnor U21500 (N_21500,N_13118,N_16324);
xnor U21501 (N_21501,N_12652,N_16083);
or U21502 (N_21502,N_13305,N_15323);
xnor U21503 (N_21503,N_13266,N_13751);
nor U21504 (N_21504,N_14252,N_16802);
or U21505 (N_21505,N_13278,N_14989);
nand U21506 (N_21506,N_15265,N_12011);
xnor U21507 (N_21507,N_12753,N_15046);
xnor U21508 (N_21508,N_12083,N_13256);
nor U21509 (N_21509,N_15684,N_15328);
or U21510 (N_21510,N_13356,N_15461);
or U21511 (N_21511,N_17866,N_17532);
or U21512 (N_21512,N_17306,N_15798);
and U21513 (N_21513,N_16276,N_15087);
nor U21514 (N_21514,N_14418,N_13761);
and U21515 (N_21515,N_15632,N_12120);
or U21516 (N_21516,N_15827,N_13418);
and U21517 (N_21517,N_17987,N_15819);
nor U21518 (N_21518,N_15900,N_15295);
or U21519 (N_21519,N_16096,N_13187);
nand U21520 (N_21520,N_12521,N_17176);
nor U21521 (N_21521,N_15173,N_17751);
xnor U21522 (N_21522,N_16437,N_16268);
nand U21523 (N_21523,N_14775,N_13518);
nand U21524 (N_21524,N_16286,N_16334);
and U21525 (N_21525,N_17085,N_17171);
nand U21526 (N_21526,N_15316,N_16132);
nand U21527 (N_21527,N_16750,N_14850);
and U21528 (N_21528,N_15357,N_14531);
or U21529 (N_21529,N_14455,N_12348);
xnor U21530 (N_21530,N_17577,N_14585);
nor U21531 (N_21531,N_14117,N_15784);
or U21532 (N_21532,N_14185,N_13732);
xnor U21533 (N_21533,N_16677,N_17476);
xor U21534 (N_21534,N_16795,N_13608);
xnor U21535 (N_21535,N_12823,N_12676);
xor U21536 (N_21536,N_17161,N_17381);
or U21537 (N_21537,N_14279,N_12125);
or U21538 (N_21538,N_17269,N_12166);
nand U21539 (N_21539,N_14092,N_13362);
and U21540 (N_21540,N_15043,N_17869);
and U21541 (N_21541,N_14783,N_17275);
nand U21542 (N_21542,N_13229,N_13384);
or U21543 (N_21543,N_16839,N_14436);
xnor U21544 (N_21544,N_13361,N_14601);
nor U21545 (N_21545,N_17589,N_14057);
xor U21546 (N_21546,N_17920,N_15259);
xor U21547 (N_21547,N_13854,N_13614);
and U21548 (N_21548,N_14868,N_15970);
and U21549 (N_21549,N_14138,N_17701);
or U21550 (N_21550,N_17791,N_12901);
and U21551 (N_21551,N_13644,N_13578);
nand U21552 (N_21552,N_14526,N_16143);
and U21553 (N_21553,N_17705,N_17303);
and U21554 (N_21554,N_16415,N_15976);
nor U21555 (N_21555,N_17648,N_12234);
nand U21556 (N_21556,N_12944,N_16432);
or U21557 (N_21557,N_12441,N_16626);
nand U21558 (N_21558,N_16512,N_16389);
nor U21559 (N_21559,N_17662,N_13524);
and U21560 (N_21560,N_17986,N_13031);
or U21561 (N_21561,N_16081,N_15171);
and U21562 (N_21562,N_12311,N_16196);
nand U21563 (N_21563,N_17181,N_13781);
and U21564 (N_21564,N_16228,N_15474);
nor U21565 (N_21565,N_16517,N_15477);
nor U21566 (N_21566,N_12060,N_12249);
nand U21567 (N_21567,N_16284,N_16793);
nor U21568 (N_21568,N_14051,N_17744);
xnor U21569 (N_21569,N_13771,N_12705);
or U21570 (N_21570,N_14974,N_12717);
nand U21571 (N_21571,N_17230,N_16720);
nor U21572 (N_21572,N_12280,N_15628);
nor U21573 (N_21573,N_17572,N_17427);
or U21574 (N_21574,N_13007,N_14525);
or U21575 (N_21575,N_13729,N_13512);
and U21576 (N_21576,N_14693,N_14472);
and U21577 (N_21577,N_12731,N_17797);
nor U21578 (N_21578,N_17070,N_16864);
nor U21579 (N_21579,N_15573,N_14144);
nor U21580 (N_21580,N_17819,N_13355);
and U21581 (N_21581,N_16164,N_17314);
xor U21582 (N_21582,N_16225,N_15840);
nor U21583 (N_21583,N_13593,N_13162);
nand U21584 (N_21584,N_15547,N_16309);
and U21585 (N_21585,N_13846,N_16977);
xor U21586 (N_21586,N_13124,N_16932);
nor U21587 (N_21587,N_17191,N_13391);
or U21588 (N_21588,N_14205,N_12732);
or U21589 (N_21589,N_13575,N_17810);
nand U21590 (N_21590,N_15587,N_12966);
and U21591 (N_21591,N_13344,N_17955);
nor U21592 (N_21592,N_15882,N_16516);
or U21593 (N_21593,N_12554,N_17746);
nand U21594 (N_21594,N_16413,N_13083);
or U21595 (N_21595,N_12998,N_13054);
or U21596 (N_21596,N_13166,N_14741);
nor U21597 (N_21597,N_12863,N_14878);
and U21598 (N_21598,N_17488,N_14677);
and U21599 (N_21599,N_16290,N_17623);
nand U21600 (N_21600,N_16170,N_16158);
or U21601 (N_21601,N_17251,N_12984);
xnor U21602 (N_21602,N_12688,N_15920);
and U21603 (N_21603,N_14286,N_16368);
nor U21604 (N_21604,N_14939,N_17667);
nand U21605 (N_21605,N_16571,N_14025);
nor U21606 (N_21606,N_14186,N_12398);
xnor U21607 (N_21607,N_13036,N_17357);
or U21608 (N_21608,N_12182,N_15966);
xnor U21609 (N_21609,N_13697,N_12135);
xor U21610 (N_21610,N_13586,N_15132);
nor U21611 (N_21611,N_14338,N_17572);
or U21612 (N_21612,N_15854,N_15557);
and U21613 (N_21613,N_13591,N_17426);
and U21614 (N_21614,N_14722,N_13107);
and U21615 (N_21615,N_13829,N_14420);
nor U21616 (N_21616,N_15009,N_16864);
or U21617 (N_21617,N_17983,N_12721);
and U21618 (N_21618,N_14187,N_16951);
and U21619 (N_21619,N_16960,N_17649);
or U21620 (N_21620,N_14961,N_13011);
xor U21621 (N_21621,N_16865,N_13815);
xnor U21622 (N_21622,N_15343,N_13937);
or U21623 (N_21623,N_15074,N_15079);
or U21624 (N_21624,N_15959,N_15212);
and U21625 (N_21625,N_15260,N_17667);
and U21626 (N_21626,N_15333,N_17365);
and U21627 (N_21627,N_15199,N_14204);
or U21628 (N_21628,N_13058,N_17432);
or U21629 (N_21629,N_17978,N_16086);
nand U21630 (N_21630,N_13125,N_14565);
and U21631 (N_21631,N_15606,N_13401);
nor U21632 (N_21632,N_14753,N_14265);
nor U21633 (N_21633,N_13209,N_13172);
or U21634 (N_21634,N_17606,N_13306);
xnor U21635 (N_21635,N_17507,N_16035);
nor U21636 (N_21636,N_15911,N_17899);
nand U21637 (N_21637,N_17069,N_12284);
or U21638 (N_21638,N_14713,N_15602);
nand U21639 (N_21639,N_14891,N_12155);
or U21640 (N_21640,N_14496,N_17157);
or U21641 (N_21641,N_17323,N_17394);
nand U21642 (N_21642,N_17003,N_15865);
or U21643 (N_21643,N_17225,N_17210);
or U21644 (N_21644,N_16000,N_12200);
nand U21645 (N_21645,N_12988,N_13668);
or U21646 (N_21646,N_13831,N_12245);
nor U21647 (N_21647,N_14073,N_14124);
or U21648 (N_21648,N_13666,N_14647);
xor U21649 (N_21649,N_17147,N_12336);
xnor U21650 (N_21650,N_16630,N_12141);
xor U21651 (N_21651,N_15102,N_13596);
and U21652 (N_21652,N_15432,N_14535);
or U21653 (N_21653,N_15128,N_17586);
nand U21654 (N_21654,N_14939,N_15414);
or U21655 (N_21655,N_14723,N_17321);
xnor U21656 (N_21656,N_12915,N_15151);
and U21657 (N_21657,N_14031,N_13992);
nand U21658 (N_21658,N_15126,N_14369);
xnor U21659 (N_21659,N_15057,N_14724);
nand U21660 (N_21660,N_17748,N_13287);
nor U21661 (N_21661,N_16897,N_16523);
or U21662 (N_21662,N_14834,N_13022);
or U21663 (N_21663,N_15327,N_15611);
or U21664 (N_21664,N_17073,N_16071);
xnor U21665 (N_21665,N_15597,N_13429);
nor U21666 (N_21666,N_14475,N_17112);
nor U21667 (N_21667,N_14927,N_14912);
nor U21668 (N_21668,N_12028,N_14679);
xnor U21669 (N_21669,N_16690,N_17144);
xnor U21670 (N_21670,N_12147,N_15190);
or U21671 (N_21671,N_13164,N_14935);
or U21672 (N_21672,N_14061,N_15391);
and U21673 (N_21673,N_17270,N_14404);
or U21674 (N_21674,N_16688,N_14340);
and U21675 (N_21675,N_12920,N_16638);
nor U21676 (N_21676,N_12988,N_13620);
nor U21677 (N_21677,N_14297,N_16771);
nand U21678 (N_21678,N_16367,N_16333);
nand U21679 (N_21679,N_14167,N_16359);
xor U21680 (N_21680,N_14242,N_13582);
xor U21681 (N_21681,N_15497,N_15078);
nor U21682 (N_21682,N_16528,N_12797);
nand U21683 (N_21683,N_17180,N_17026);
and U21684 (N_21684,N_15821,N_17600);
xor U21685 (N_21685,N_13637,N_15017);
nor U21686 (N_21686,N_15786,N_12174);
and U21687 (N_21687,N_12231,N_14016);
or U21688 (N_21688,N_14049,N_12824);
xor U21689 (N_21689,N_17983,N_14234);
or U21690 (N_21690,N_13093,N_17922);
and U21691 (N_21691,N_14871,N_16123);
xnor U21692 (N_21692,N_14145,N_13543);
and U21693 (N_21693,N_15139,N_14140);
nor U21694 (N_21694,N_16274,N_14238);
xor U21695 (N_21695,N_14600,N_16924);
or U21696 (N_21696,N_17958,N_14997);
and U21697 (N_21697,N_13351,N_17440);
xnor U21698 (N_21698,N_14423,N_15461);
nor U21699 (N_21699,N_13643,N_12175);
xnor U21700 (N_21700,N_12834,N_14494);
nand U21701 (N_21701,N_16726,N_13640);
nor U21702 (N_21702,N_16088,N_13934);
nor U21703 (N_21703,N_16796,N_13872);
xnor U21704 (N_21704,N_16358,N_17626);
nand U21705 (N_21705,N_12876,N_13629);
nor U21706 (N_21706,N_16168,N_14991);
nand U21707 (N_21707,N_16740,N_16766);
or U21708 (N_21708,N_13574,N_14434);
and U21709 (N_21709,N_17358,N_12175);
nand U21710 (N_21710,N_14868,N_12660);
and U21711 (N_21711,N_13285,N_15412);
or U21712 (N_21712,N_12223,N_15176);
nor U21713 (N_21713,N_13347,N_15821);
or U21714 (N_21714,N_16464,N_17630);
or U21715 (N_21715,N_14132,N_15031);
nor U21716 (N_21716,N_17070,N_15119);
and U21717 (N_21717,N_12886,N_13698);
nand U21718 (N_21718,N_15616,N_14361);
xnor U21719 (N_21719,N_14910,N_13835);
nand U21720 (N_21720,N_15504,N_17624);
or U21721 (N_21721,N_14488,N_16249);
or U21722 (N_21722,N_13767,N_15122);
xnor U21723 (N_21723,N_16854,N_13521);
xnor U21724 (N_21724,N_17241,N_17165);
nand U21725 (N_21725,N_17313,N_17263);
nand U21726 (N_21726,N_12818,N_16545);
or U21727 (N_21727,N_15527,N_15105);
nor U21728 (N_21728,N_13682,N_12903);
or U21729 (N_21729,N_17115,N_14116);
or U21730 (N_21730,N_17741,N_12569);
nand U21731 (N_21731,N_13071,N_16040);
nand U21732 (N_21732,N_14157,N_14958);
nor U21733 (N_21733,N_13080,N_13786);
xor U21734 (N_21734,N_16476,N_17257);
or U21735 (N_21735,N_12359,N_14253);
and U21736 (N_21736,N_12780,N_16075);
xor U21737 (N_21737,N_16332,N_15866);
xnor U21738 (N_21738,N_17668,N_14569);
nor U21739 (N_21739,N_15613,N_15075);
nor U21740 (N_21740,N_17592,N_17868);
xnor U21741 (N_21741,N_14589,N_16703);
nand U21742 (N_21742,N_12073,N_15830);
or U21743 (N_21743,N_16735,N_15796);
nand U21744 (N_21744,N_14742,N_16042);
xnor U21745 (N_21745,N_15747,N_12718);
and U21746 (N_21746,N_16782,N_12735);
xnor U21747 (N_21747,N_14848,N_15410);
xor U21748 (N_21748,N_16714,N_15098);
or U21749 (N_21749,N_12045,N_17892);
xnor U21750 (N_21750,N_15173,N_17036);
or U21751 (N_21751,N_12395,N_15138);
nand U21752 (N_21752,N_13166,N_13657);
or U21753 (N_21753,N_14885,N_14671);
or U21754 (N_21754,N_13387,N_15855);
nor U21755 (N_21755,N_16503,N_12885);
nand U21756 (N_21756,N_14220,N_13275);
nand U21757 (N_21757,N_14975,N_13549);
nor U21758 (N_21758,N_16177,N_12142);
xor U21759 (N_21759,N_15857,N_16850);
xor U21760 (N_21760,N_17670,N_17181);
nor U21761 (N_21761,N_12356,N_13893);
nand U21762 (N_21762,N_12917,N_13796);
nand U21763 (N_21763,N_16516,N_17542);
nand U21764 (N_21764,N_14603,N_16945);
and U21765 (N_21765,N_12039,N_13494);
xnor U21766 (N_21766,N_13561,N_17684);
nor U21767 (N_21767,N_13502,N_12169);
nor U21768 (N_21768,N_13205,N_17657);
xor U21769 (N_21769,N_17005,N_15312);
nand U21770 (N_21770,N_15995,N_14426);
nor U21771 (N_21771,N_17608,N_15011);
and U21772 (N_21772,N_14383,N_13685);
nor U21773 (N_21773,N_15055,N_13638);
nor U21774 (N_21774,N_12869,N_15983);
or U21775 (N_21775,N_12156,N_17102);
or U21776 (N_21776,N_15655,N_12977);
nand U21777 (N_21777,N_17248,N_15818);
nand U21778 (N_21778,N_17455,N_12639);
or U21779 (N_21779,N_17083,N_15862);
nand U21780 (N_21780,N_14376,N_17763);
and U21781 (N_21781,N_13545,N_16102);
nand U21782 (N_21782,N_16284,N_12956);
nor U21783 (N_21783,N_17734,N_17181);
xnor U21784 (N_21784,N_16990,N_15253);
and U21785 (N_21785,N_14364,N_16224);
xor U21786 (N_21786,N_15518,N_12762);
nand U21787 (N_21787,N_13590,N_12468);
or U21788 (N_21788,N_16205,N_14868);
nor U21789 (N_21789,N_14819,N_15777);
nand U21790 (N_21790,N_16728,N_14221);
xnor U21791 (N_21791,N_12447,N_15976);
xnor U21792 (N_21792,N_16694,N_12212);
nand U21793 (N_21793,N_13169,N_12505);
xnor U21794 (N_21794,N_13194,N_17715);
or U21795 (N_21795,N_14742,N_14558);
and U21796 (N_21796,N_16655,N_14953);
or U21797 (N_21797,N_17176,N_15121);
nand U21798 (N_21798,N_13608,N_16960);
nand U21799 (N_21799,N_17933,N_14038);
and U21800 (N_21800,N_16517,N_17211);
or U21801 (N_21801,N_12814,N_13552);
and U21802 (N_21802,N_13293,N_14384);
or U21803 (N_21803,N_16137,N_15665);
or U21804 (N_21804,N_17406,N_12293);
nand U21805 (N_21805,N_13187,N_12440);
nand U21806 (N_21806,N_12691,N_15896);
nand U21807 (N_21807,N_15263,N_15019);
or U21808 (N_21808,N_15319,N_14929);
and U21809 (N_21809,N_12647,N_13522);
and U21810 (N_21810,N_12919,N_16362);
nand U21811 (N_21811,N_14739,N_15860);
xnor U21812 (N_21812,N_15635,N_14979);
and U21813 (N_21813,N_13436,N_14248);
or U21814 (N_21814,N_12386,N_12684);
and U21815 (N_21815,N_14188,N_16211);
or U21816 (N_21816,N_17045,N_15864);
and U21817 (N_21817,N_14775,N_16874);
and U21818 (N_21818,N_16899,N_14183);
xnor U21819 (N_21819,N_14190,N_15814);
and U21820 (N_21820,N_17949,N_16119);
or U21821 (N_21821,N_14530,N_16833);
nand U21822 (N_21822,N_13839,N_15996);
and U21823 (N_21823,N_12312,N_16632);
or U21824 (N_21824,N_15669,N_13692);
or U21825 (N_21825,N_13795,N_13283);
xor U21826 (N_21826,N_15010,N_13115);
or U21827 (N_21827,N_17611,N_15149);
nand U21828 (N_21828,N_14676,N_15418);
and U21829 (N_21829,N_14294,N_13081);
or U21830 (N_21830,N_17531,N_13075);
xor U21831 (N_21831,N_13456,N_12058);
nand U21832 (N_21832,N_14072,N_14618);
nor U21833 (N_21833,N_14773,N_13709);
and U21834 (N_21834,N_12002,N_13833);
and U21835 (N_21835,N_14207,N_13368);
nand U21836 (N_21836,N_13999,N_15340);
or U21837 (N_21837,N_14220,N_13790);
nand U21838 (N_21838,N_12077,N_15978);
nand U21839 (N_21839,N_12540,N_13881);
and U21840 (N_21840,N_14360,N_15259);
and U21841 (N_21841,N_13226,N_17220);
and U21842 (N_21842,N_17223,N_14756);
or U21843 (N_21843,N_12593,N_14185);
or U21844 (N_21844,N_13288,N_17131);
xor U21845 (N_21845,N_12582,N_13198);
nor U21846 (N_21846,N_12725,N_13903);
nor U21847 (N_21847,N_14841,N_13639);
and U21848 (N_21848,N_14873,N_12654);
or U21849 (N_21849,N_14536,N_16630);
xor U21850 (N_21850,N_16237,N_12030);
nor U21851 (N_21851,N_14853,N_16820);
nor U21852 (N_21852,N_16778,N_15296);
nor U21853 (N_21853,N_14490,N_13808);
xor U21854 (N_21854,N_17362,N_15975);
xor U21855 (N_21855,N_17876,N_16812);
nand U21856 (N_21856,N_14543,N_14707);
xnor U21857 (N_21857,N_12210,N_13468);
nand U21858 (N_21858,N_17728,N_13277);
nor U21859 (N_21859,N_14872,N_17185);
xor U21860 (N_21860,N_14577,N_16451);
or U21861 (N_21861,N_16224,N_17105);
nor U21862 (N_21862,N_14613,N_12979);
nor U21863 (N_21863,N_17910,N_14008);
xnor U21864 (N_21864,N_16032,N_16253);
xnor U21865 (N_21865,N_14337,N_13592);
or U21866 (N_21866,N_14806,N_16002);
or U21867 (N_21867,N_14050,N_13675);
or U21868 (N_21868,N_14602,N_17893);
and U21869 (N_21869,N_15461,N_13171);
nor U21870 (N_21870,N_14697,N_12500);
nor U21871 (N_21871,N_17245,N_16476);
nand U21872 (N_21872,N_16844,N_13320);
xnor U21873 (N_21873,N_14335,N_12970);
and U21874 (N_21874,N_16863,N_12617);
xnor U21875 (N_21875,N_17228,N_17416);
xnor U21876 (N_21876,N_12446,N_14219);
or U21877 (N_21877,N_14262,N_12977);
xnor U21878 (N_21878,N_14548,N_13037);
or U21879 (N_21879,N_12391,N_14152);
nand U21880 (N_21880,N_13120,N_16484);
xor U21881 (N_21881,N_12083,N_14590);
xor U21882 (N_21882,N_17677,N_13168);
or U21883 (N_21883,N_15573,N_17870);
nand U21884 (N_21884,N_16407,N_14093);
and U21885 (N_21885,N_16953,N_14030);
xnor U21886 (N_21886,N_12364,N_15677);
xnor U21887 (N_21887,N_16800,N_14117);
and U21888 (N_21888,N_13293,N_16709);
and U21889 (N_21889,N_12866,N_17222);
or U21890 (N_21890,N_17846,N_12439);
and U21891 (N_21891,N_12055,N_15020);
or U21892 (N_21892,N_12196,N_17589);
nand U21893 (N_21893,N_14515,N_13683);
nand U21894 (N_21894,N_17561,N_14492);
or U21895 (N_21895,N_15283,N_12275);
or U21896 (N_21896,N_16477,N_14326);
and U21897 (N_21897,N_14952,N_13902);
nor U21898 (N_21898,N_15566,N_17440);
nand U21899 (N_21899,N_15144,N_12147);
xor U21900 (N_21900,N_17580,N_13504);
nor U21901 (N_21901,N_16861,N_14425);
and U21902 (N_21902,N_16712,N_17932);
nand U21903 (N_21903,N_13980,N_17197);
nor U21904 (N_21904,N_17313,N_17588);
or U21905 (N_21905,N_17585,N_12617);
or U21906 (N_21906,N_14581,N_17770);
nand U21907 (N_21907,N_15637,N_14102);
or U21908 (N_21908,N_17267,N_14063);
or U21909 (N_21909,N_16620,N_15909);
nor U21910 (N_21910,N_16759,N_13663);
or U21911 (N_21911,N_12750,N_17360);
and U21912 (N_21912,N_15706,N_13329);
or U21913 (N_21913,N_17693,N_14789);
nor U21914 (N_21914,N_13049,N_17387);
and U21915 (N_21915,N_15626,N_13541);
or U21916 (N_21916,N_14657,N_16591);
or U21917 (N_21917,N_16253,N_17967);
or U21918 (N_21918,N_14325,N_17779);
xor U21919 (N_21919,N_13281,N_12152);
and U21920 (N_21920,N_17280,N_12116);
nor U21921 (N_21921,N_16466,N_13827);
xnor U21922 (N_21922,N_13889,N_14331);
xor U21923 (N_21923,N_12815,N_12516);
nand U21924 (N_21924,N_15772,N_17679);
nand U21925 (N_21925,N_17902,N_14782);
or U21926 (N_21926,N_14898,N_16243);
nor U21927 (N_21927,N_13009,N_12394);
and U21928 (N_21928,N_14304,N_16860);
xnor U21929 (N_21929,N_12872,N_12129);
nor U21930 (N_21930,N_16768,N_17211);
nand U21931 (N_21931,N_15288,N_16002);
and U21932 (N_21932,N_14544,N_14900);
and U21933 (N_21933,N_17711,N_15957);
or U21934 (N_21934,N_17813,N_15381);
xor U21935 (N_21935,N_12126,N_16693);
or U21936 (N_21936,N_15270,N_13361);
and U21937 (N_21937,N_13569,N_12191);
xnor U21938 (N_21938,N_16229,N_14828);
and U21939 (N_21939,N_16765,N_13483);
nand U21940 (N_21940,N_12849,N_17717);
nand U21941 (N_21941,N_16298,N_14464);
or U21942 (N_21942,N_17640,N_12024);
and U21943 (N_21943,N_17937,N_14454);
nand U21944 (N_21944,N_14279,N_15399);
and U21945 (N_21945,N_13661,N_13342);
xor U21946 (N_21946,N_15916,N_16896);
nand U21947 (N_21947,N_17234,N_16472);
nor U21948 (N_21948,N_15633,N_15691);
or U21949 (N_21949,N_12068,N_12751);
or U21950 (N_21950,N_17113,N_12412);
nor U21951 (N_21951,N_15377,N_13858);
xor U21952 (N_21952,N_14278,N_15848);
nor U21953 (N_21953,N_13406,N_13107);
and U21954 (N_21954,N_15138,N_12724);
and U21955 (N_21955,N_15999,N_14501);
nor U21956 (N_21956,N_12577,N_13687);
and U21957 (N_21957,N_16395,N_14836);
nor U21958 (N_21958,N_13890,N_14731);
nand U21959 (N_21959,N_13926,N_16839);
nor U21960 (N_21960,N_13432,N_14751);
nor U21961 (N_21961,N_12972,N_12304);
nand U21962 (N_21962,N_13008,N_13428);
and U21963 (N_21963,N_16002,N_12078);
nand U21964 (N_21964,N_12267,N_17090);
and U21965 (N_21965,N_15379,N_17528);
nand U21966 (N_21966,N_12875,N_13198);
nand U21967 (N_21967,N_12336,N_12615);
xnor U21968 (N_21968,N_17713,N_17728);
and U21969 (N_21969,N_14106,N_12565);
nor U21970 (N_21970,N_15263,N_15434);
nand U21971 (N_21971,N_17987,N_17464);
and U21972 (N_21972,N_15850,N_17648);
and U21973 (N_21973,N_14087,N_12275);
xnor U21974 (N_21974,N_17728,N_13998);
or U21975 (N_21975,N_13246,N_17556);
and U21976 (N_21976,N_13225,N_12515);
nor U21977 (N_21977,N_12974,N_14091);
nand U21978 (N_21978,N_16165,N_17207);
nand U21979 (N_21979,N_17475,N_13647);
xnor U21980 (N_21980,N_15368,N_12465);
xor U21981 (N_21981,N_17561,N_12042);
or U21982 (N_21982,N_16210,N_13920);
xor U21983 (N_21983,N_17936,N_17032);
xnor U21984 (N_21984,N_16498,N_16995);
xor U21985 (N_21985,N_14963,N_17832);
nand U21986 (N_21986,N_17938,N_13977);
nor U21987 (N_21987,N_15563,N_12575);
or U21988 (N_21988,N_12153,N_15584);
nand U21989 (N_21989,N_17317,N_14469);
nand U21990 (N_21990,N_16045,N_12327);
and U21991 (N_21991,N_13619,N_13488);
or U21992 (N_21992,N_17499,N_16932);
xor U21993 (N_21993,N_13140,N_12358);
xnor U21994 (N_21994,N_14680,N_14572);
and U21995 (N_21995,N_13605,N_13594);
or U21996 (N_21996,N_15928,N_16012);
nor U21997 (N_21997,N_13943,N_15934);
nand U21998 (N_21998,N_14905,N_13761);
nor U21999 (N_21999,N_14318,N_12208);
and U22000 (N_22000,N_14645,N_14635);
xor U22001 (N_22001,N_16431,N_15694);
and U22002 (N_22002,N_14829,N_17312);
nand U22003 (N_22003,N_14738,N_17579);
and U22004 (N_22004,N_13880,N_14428);
nand U22005 (N_22005,N_13818,N_13628);
and U22006 (N_22006,N_12138,N_17614);
and U22007 (N_22007,N_13073,N_16139);
and U22008 (N_22008,N_15116,N_17421);
nor U22009 (N_22009,N_14724,N_15164);
and U22010 (N_22010,N_12427,N_14491);
or U22011 (N_22011,N_17147,N_16727);
nor U22012 (N_22012,N_12750,N_16768);
or U22013 (N_22013,N_15472,N_12066);
nand U22014 (N_22014,N_17997,N_14566);
nor U22015 (N_22015,N_12020,N_15234);
nor U22016 (N_22016,N_15160,N_16774);
nand U22017 (N_22017,N_16396,N_16919);
or U22018 (N_22018,N_14928,N_14444);
and U22019 (N_22019,N_12108,N_17121);
nor U22020 (N_22020,N_17246,N_15476);
and U22021 (N_22021,N_13635,N_16110);
and U22022 (N_22022,N_17918,N_15583);
and U22023 (N_22023,N_15807,N_12877);
or U22024 (N_22024,N_12590,N_12834);
nand U22025 (N_22025,N_16744,N_12829);
and U22026 (N_22026,N_17331,N_15693);
and U22027 (N_22027,N_17090,N_15302);
nand U22028 (N_22028,N_13757,N_16930);
xnor U22029 (N_22029,N_15228,N_17429);
and U22030 (N_22030,N_13831,N_15440);
nor U22031 (N_22031,N_12811,N_15060);
nor U22032 (N_22032,N_14273,N_15102);
nand U22033 (N_22033,N_12954,N_15627);
and U22034 (N_22034,N_13811,N_15538);
and U22035 (N_22035,N_13838,N_12521);
nand U22036 (N_22036,N_17475,N_17395);
xor U22037 (N_22037,N_14650,N_15850);
nor U22038 (N_22038,N_17712,N_15643);
nand U22039 (N_22039,N_16087,N_14680);
nand U22040 (N_22040,N_14690,N_12714);
and U22041 (N_22041,N_13840,N_14593);
or U22042 (N_22042,N_15201,N_17027);
nor U22043 (N_22043,N_16105,N_14024);
or U22044 (N_22044,N_14579,N_17013);
and U22045 (N_22045,N_12873,N_16808);
or U22046 (N_22046,N_16894,N_13150);
nand U22047 (N_22047,N_14352,N_16092);
nand U22048 (N_22048,N_13459,N_15301);
or U22049 (N_22049,N_15953,N_15241);
and U22050 (N_22050,N_16903,N_13360);
or U22051 (N_22051,N_15903,N_12250);
nor U22052 (N_22052,N_15315,N_15973);
nor U22053 (N_22053,N_13826,N_14198);
or U22054 (N_22054,N_12395,N_13140);
nor U22055 (N_22055,N_14632,N_14534);
nor U22056 (N_22056,N_13283,N_15300);
xnor U22057 (N_22057,N_13969,N_14929);
nand U22058 (N_22058,N_13245,N_13883);
or U22059 (N_22059,N_12958,N_15166);
nor U22060 (N_22060,N_13434,N_12062);
nand U22061 (N_22061,N_15514,N_16063);
nand U22062 (N_22062,N_17794,N_15519);
xnor U22063 (N_22063,N_13961,N_14810);
xor U22064 (N_22064,N_12689,N_16685);
and U22065 (N_22065,N_14604,N_12083);
nand U22066 (N_22066,N_13486,N_15075);
nor U22067 (N_22067,N_17795,N_12759);
nor U22068 (N_22068,N_15256,N_16734);
and U22069 (N_22069,N_13797,N_15117);
nand U22070 (N_22070,N_15011,N_12396);
or U22071 (N_22071,N_17963,N_15902);
xnor U22072 (N_22072,N_15179,N_15259);
nor U22073 (N_22073,N_13733,N_17688);
nor U22074 (N_22074,N_16817,N_14882);
and U22075 (N_22075,N_14939,N_16832);
xor U22076 (N_22076,N_17453,N_13661);
or U22077 (N_22077,N_16021,N_14458);
or U22078 (N_22078,N_16238,N_14166);
nand U22079 (N_22079,N_17168,N_17973);
nor U22080 (N_22080,N_15021,N_13833);
and U22081 (N_22081,N_17921,N_13926);
or U22082 (N_22082,N_15944,N_13577);
or U22083 (N_22083,N_15107,N_13638);
and U22084 (N_22084,N_13611,N_12018);
xnor U22085 (N_22085,N_13217,N_15855);
nand U22086 (N_22086,N_15392,N_16535);
xnor U22087 (N_22087,N_12089,N_17530);
nor U22088 (N_22088,N_14479,N_14798);
or U22089 (N_22089,N_17924,N_17653);
nand U22090 (N_22090,N_14811,N_15780);
nand U22091 (N_22091,N_17898,N_12514);
nand U22092 (N_22092,N_17759,N_16957);
xnor U22093 (N_22093,N_14596,N_15657);
or U22094 (N_22094,N_15909,N_16638);
nor U22095 (N_22095,N_12744,N_17897);
nor U22096 (N_22096,N_16735,N_13832);
and U22097 (N_22097,N_15431,N_13061);
nor U22098 (N_22098,N_14034,N_15633);
or U22099 (N_22099,N_15492,N_16106);
or U22100 (N_22100,N_15171,N_13094);
xnor U22101 (N_22101,N_16813,N_13051);
nand U22102 (N_22102,N_17089,N_13840);
nor U22103 (N_22103,N_14597,N_15177);
nor U22104 (N_22104,N_14751,N_14391);
or U22105 (N_22105,N_15502,N_13160);
nor U22106 (N_22106,N_15557,N_13253);
or U22107 (N_22107,N_17879,N_13486);
xor U22108 (N_22108,N_14313,N_14216);
nor U22109 (N_22109,N_12419,N_14423);
or U22110 (N_22110,N_14687,N_17189);
or U22111 (N_22111,N_13165,N_16898);
and U22112 (N_22112,N_14180,N_15730);
and U22113 (N_22113,N_14735,N_15881);
xor U22114 (N_22114,N_17760,N_15825);
nand U22115 (N_22115,N_14250,N_17860);
nand U22116 (N_22116,N_17330,N_14721);
xor U22117 (N_22117,N_13083,N_16324);
nor U22118 (N_22118,N_16558,N_14689);
nand U22119 (N_22119,N_13708,N_15319);
xor U22120 (N_22120,N_12780,N_14180);
and U22121 (N_22121,N_13475,N_15690);
nor U22122 (N_22122,N_15864,N_15729);
or U22123 (N_22123,N_13872,N_17518);
and U22124 (N_22124,N_15607,N_12301);
or U22125 (N_22125,N_16722,N_16405);
nor U22126 (N_22126,N_14294,N_14111);
nor U22127 (N_22127,N_17998,N_12572);
xor U22128 (N_22128,N_16693,N_14963);
and U22129 (N_22129,N_13690,N_16678);
or U22130 (N_22130,N_12499,N_17116);
nor U22131 (N_22131,N_15922,N_16486);
and U22132 (N_22132,N_15002,N_15202);
nand U22133 (N_22133,N_15200,N_13754);
or U22134 (N_22134,N_17123,N_14064);
nand U22135 (N_22135,N_12656,N_17197);
xor U22136 (N_22136,N_12550,N_17575);
nor U22137 (N_22137,N_13294,N_15500);
nor U22138 (N_22138,N_15989,N_12834);
and U22139 (N_22139,N_16181,N_15911);
xnor U22140 (N_22140,N_14876,N_17750);
or U22141 (N_22141,N_12670,N_13711);
nand U22142 (N_22142,N_15362,N_12389);
xnor U22143 (N_22143,N_12992,N_14100);
or U22144 (N_22144,N_14122,N_15758);
or U22145 (N_22145,N_14107,N_14105);
nor U22146 (N_22146,N_17475,N_12728);
and U22147 (N_22147,N_13304,N_14692);
nor U22148 (N_22148,N_14747,N_12442);
nand U22149 (N_22149,N_15177,N_17567);
nand U22150 (N_22150,N_16824,N_16357);
nor U22151 (N_22151,N_12629,N_15579);
nor U22152 (N_22152,N_15420,N_16359);
or U22153 (N_22153,N_17916,N_12725);
nand U22154 (N_22154,N_13038,N_16297);
or U22155 (N_22155,N_14998,N_12392);
and U22156 (N_22156,N_13205,N_13548);
or U22157 (N_22157,N_12014,N_15178);
nand U22158 (N_22158,N_12481,N_12286);
nand U22159 (N_22159,N_13584,N_13228);
xor U22160 (N_22160,N_15293,N_12847);
or U22161 (N_22161,N_17652,N_13582);
nor U22162 (N_22162,N_17430,N_12799);
or U22163 (N_22163,N_17774,N_15364);
nor U22164 (N_22164,N_16628,N_15981);
nor U22165 (N_22165,N_15120,N_16387);
or U22166 (N_22166,N_14373,N_14342);
nor U22167 (N_22167,N_16052,N_13319);
and U22168 (N_22168,N_12149,N_14928);
and U22169 (N_22169,N_17795,N_17981);
nor U22170 (N_22170,N_14392,N_13962);
or U22171 (N_22171,N_13372,N_16790);
and U22172 (N_22172,N_14586,N_16854);
and U22173 (N_22173,N_13365,N_15078);
xnor U22174 (N_22174,N_17280,N_12763);
or U22175 (N_22175,N_13714,N_13940);
xnor U22176 (N_22176,N_12350,N_16303);
nor U22177 (N_22177,N_12344,N_14358);
or U22178 (N_22178,N_14296,N_15480);
nor U22179 (N_22179,N_12250,N_14938);
nand U22180 (N_22180,N_16277,N_16346);
xnor U22181 (N_22181,N_16723,N_12799);
nor U22182 (N_22182,N_12347,N_17303);
nand U22183 (N_22183,N_17803,N_17691);
nor U22184 (N_22184,N_13052,N_12277);
and U22185 (N_22185,N_12929,N_15234);
or U22186 (N_22186,N_15305,N_15868);
nor U22187 (N_22187,N_13299,N_14129);
nor U22188 (N_22188,N_16457,N_14865);
nor U22189 (N_22189,N_12883,N_15581);
nor U22190 (N_22190,N_17675,N_13260);
nand U22191 (N_22191,N_12436,N_15008);
or U22192 (N_22192,N_16938,N_16495);
nor U22193 (N_22193,N_16669,N_14627);
nand U22194 (N_22194,N_14464,N_17112);
nor U22195 (N_22195,N_13600,N_13201);
xor U22196 (N_22196,N_15418,N_13938);
xor U22197 (N_22197,N_13027,N_17861);
nand U22198 (N_22198,N_16647,N_14481);
or U22199 (N_22199,N_12240,N_16360);
nor U22200 (N_22200,N_12734,N_12768);
and U22201 (N_22201,N_12049,N_12558);
nor U22202 (N_22202,N_13665,N_16215);
xnor U22203 (N_22203,N_14711,N_16705);
and U22204 (N_22204,N_17148,N_13269);
xor U22205 (N_22205,N_15803,N_17984);
xnor U22206 (N_22206,N_15715,N_17011);
or U22207 (N_22207,N_15524,N_13087);
or U22208 (N_22208,N_12709,N_12965);
nand U22209 (N_22209,N_12335,N_14865);
or U22210 (N_22210,N_13011,N_16681);
and U22211 (N_22211,N_14889,N_16768);
xnor U22212 (N_22212,N_17124,N_13443);
nor U22213 (N_22213,N_15831,N_12136);
or U22214 (N_22214,N_16849,N_12480);
and U22215 (N_22215,N_14894,N_17503);
nor U22216 (N_22216,N_12139,N_14030);
or U22217 (N_22217,N_17262,N_17446);
nand U22218 (N_22218,N_17191,N_17139);
and U22219 (N_22219,N_15693,N_12313);
or U22220 (N_22220,N_17444,N_13154);
and U22221 (N_22221,N_14205,N_12092);
xor U22222 (N_22222,N_16886,N_13726);
xnor U22223 (N_22223,N_14101,N_17539);
nand U22224 (N_22224,N_15631,N_17122);
and U22225 (N_22225,N_14392,N_13895);
nand U22226 (N_22226,N_12640,N_15556);
xnor U22227 (N_22227,N_16769,N_15223);
or U22228 (N_22228,N_14474,N_15011);
and U22229 (N_22229,N_12360,N_14500);
nor U22230 (N_22230,N_17080,N_16168);
xor U22231 (N_22231,N_16077,N_14161);
and U22232 (N_22232,N_13792,N_13202);
nand U22233 (N_22233,N_13193,N_12362);
xor U22234 (N_22234,N_14518,N_13462);
nand U22235 (N_22235,N_17713,N_16159);
xor U22236 (N_22236,N_16800,N_17710);
or U22237 (N_22237,N_15936,N_13414);
and U22238 (N_22238,N_17774,N_15010);
or U22239 (N_22239,N_17940,N_15831);
xnor U22240 (N_22240,N_13884,N_13926);
xor U22241 (N_22241,N_13120,N_17800);
xor U22242 (N_22242,N_16737,N_14767);
and U22243 (N_22243,N_15480,N_13654);
or U22244 (N_22244,N_15096,N_13317);
nor U22245 (N_22245,N_13455,N_14099);
nor U22246 (N_22246,N_14121,N_17058);
or U22247 (N_22247,N_15836,N_13437);
or U22248 (N_22248,N_17700,N_13941);
or U22249 (N_22249,N_16822,N_14217);
or U22250 (N_22250,N_16158,N_12028);
nor U22251 (N_22251,N_15463,N_12101);
or U22252 (N_22252,N_13065,N_17044);
xor U22253 (N_22253,N_14342,N_12864);
nor U22254 (N_22254,N_16049,N_12645);
or U22255 (N_22255,N_14323,N_13061);
or U22256 (N_22256,N_17685,N_14562);
and U22257 (N_22257,N_14878,N_13600);
xnor U22258 (N_22258,N_15101,N_17267);
or U22259 (N_22259,N_12878,N_14414);
and U22260 (N_22260,N_14056,N_14042);
and U22261 (N_22261,N_14518,N_12025);
or U22262 (N_22262,N_14507,N_14021);
nand U22263 (N_22263,N_12066,N_17520);
or U22264 (N_22264,N_14983,N_17505);
or U22265 (N_22265,N_12108,N_12495);
nor U22266 (N_22266,N_15646,N_17597);
and U22267 (N_22267,N_14447,N_14621);
nand U22268 (N_22268,N_13648,N_13230);
nand U22269 (N_22269,N_13379,N_17265);
nor U22270 (N_22270,N_13570,N_13601);
or U22271 (N_22271,N_12729,N_17112);
nor U22272 (N_22272,N_16640,N_14637);
xor U22273 (N_22273,N_13009,N_12487);
nand U22274 (N_22274,N_12142,N_14433);
and U22275 (N_22275,N_17070,N_16936);
xor U22276 (N_22276,N_16863,N_16888);
xnor U22277 (N_22277,N_17510,N_15144);
nor U22278 (N_22278,N_15133,N_16931);
and U22279 (N_22279,N_13259,N_12855);
nand U22280 (N_22280,N_16369,N_12969);
nand U22281 (N_22281,N_16617,N_15048);
and U22282 (N_22282,N_15768,N_14839);
or U22283 (N_22283,N_17499,N_14847);
and U22284 (N_22284,N_16038,N_16495);
or U22285 (N_22285,N_15610,N_14827);
nor U22286 (N_22286,N_12853,N_14609);
or U22287 (N_22287,N_16609,N_14122);
and U22288 (N_22288,N_15405,N_14620);
xor U22289 (N_22289,N_12124,N_14766);
or U22290 (N_22290,N_16974,N_12036);
nand U22291 (N_22291,N_14681,N_15999);
nand U22292 (N_22292,N_13109,N_14375);
nor U22293 (N_22293,N_17704,N_17720);
and U22294 (N_22294,N_14582,N_13228);
or U22295 (N_22295,N_16767,N_15300);
nor U22296 (N_22296,N_12675,N_14431);
nor U22297 (N_22297,N_16877,N_17391);
nand U22298 (N_22298,N_13234,N_17620);
or U22299 (N_22299,N_13039,N_14883);
or U22300 (N_22300,N_17701,N_17983);
nor U22301 (N_22301,N_14593,N_15003);
nand U22302 (N_22302,N_12344,N_15826);
and U22303 (N_22303,N_17361,N_12820);
nand U22304 (N_22304,N_13499,N_14597);
xor U22305 (N_22305,N_17268,N_13006);
or U22306 (N_22306,N_14964,N_16132);
or U22307 (N_22307,N_16563,N_16146);
xnor U22308 (N_22308,N_14025,N_13554);
or U22309 (N_22309,N_17080,N_16919);
nand U22310 (N_22310,N_17342,N_12208);
and U22311 (N_22311,N_13396,N_14431);
and U22312 (N_22312,N_16721,N_12510);
xnor U22313 (N_22313,N_13438,N_14930);
and U22314 (N_22314,N_12441,N_15101);
xnor U22315 (N_22315,N_13531,N_15407);
or U22316 (N_22316,N_17649,N_15328);
xnor U22317 (N_22317,N_15967,N_13040);
nand U22318 (N_22318,N_15057,N_15541);
or U22319 (N_22319,N_13008,N_15206);
or U22320 (N_22320,N_12803,N_17370);
nand U22321 (N_22321,N_13906,N_16785);
nor U22322 (N_22322,N_15477,N_15239);
nand U22323 (N_22323,N_17428,N_12035);
nand U22324 (N_22324,N_13231,N_12889);
or U22325 (N_22325,N_12131,N_12121);
xnor U22326 (N_22326,N_16084,N_16276);
nor U22327 (N_22327,N_17513,N_12157);
nand U22328 (N_22328,N_13973,N_14877);
nor U22329 (N_22329,N_17611,N_14872);
or U22330 (N_22330,N_12704,N_13409);
nand U22331 (N_22331,N_12220,N_17378);
and U22332 (N_22332,N_16182,N_13783);
or U22333 (N_22333,N_17161,N_14468);
and U22334 (N_22334,N_17160,N_17567);
or U22335 (N_22335,N_12759,N_13575);
nand U22336 (N_22336,N_15274,N_17892);
nor U22337 (N_22337,N_12139,N_16383);
and U22338 (N_22338,N_13384,N_17162);
nor U22339 (N_22339,N_14515,N_14406);
and U22340 (N_22340,N_16288,N_14395);
or U22341 (N_22341,N_14856,N_13331);
xor U22342 (N_22342,N_17233,N_14998);
nor U22343 (N_22343,N_14510,N_15396);
nor U22344 (N_22344,N_14488,N_12511);
xnor U22345 (N_22345,N_17059,N_14451);
or U22346 (N_22346,N_14809,N_13158);
or U22347 (N_22347,N_12239,N_14470);
nand U22348 (N_22348,N_17266,N_15811);
or U22349 (N_22349,N_12782,N_14366);
and U22350 (N_22350,N_13911,N_17306);
nor U22351 (N_22351,N_17506,N_16733);
xnor U22352 (N_22352,N_16663,N_13541);
xnor U22353 (N_22353,N_14336,N_14654);
or U22354 (N_22354,N_14764,N_15899);
nor U22355 (N_22355,N_16285,N_15298);
or U22356 (N_22356,N_16965,N_16927);
or U22357 (N_22357,N_16422,N_15503);
or U22358 (N_22358,N_15098,N_15335);
nand U22359 (N_22359,N_13084,N_14862);
nand U22360 (N_22360,N_14273,N_12034);
nor U22361 (N_22361,N_13304,N_14971);
and U22362 (N_22362,N_15262,N_15897);
nand U22363 (N_22363,N_17533,N_13483);
nor U22364 (N_22364,N_17631,N_12693);
xor U22365 (N_22365,N_12488,N_13343);
xor U22366 (N_22366,N_16419,N_13806);
xnor U22367 (N_22367,N_12729,N_12713);
and U22368 (N_22368,N_14547,N_16015);
and U22369 (N_22369,N_16913,N_15439);
nor U22370 (N_22370,N_16587,N_13288);
xnor U22371 (N_22371,N_17795,N_14465);
nor U22372 (N_22372,N_13014,N_16618);
nor U22373 (N_22373,N_15781,N_12246);
nor U22374 (N_22374,N_17542,N_14784);
or U22375 (N_22375,N_15000,N_16809);
nand U22376 (N_22376,N_15584,N_16934);
xor U22377 (N_22377,N_13060,N_15802);
nand U22378 (N_22378,N_12346,N_16544);
xor U22379 (N_22379,N_15781,N_14588);
nand U22380 (N_22380,N_14760,N_16809);
nand U22381 (N_22381,N_12011,N_15223);
or U22382 (N_22382,N_12176,N_14913);
and U22383 (N_22383,N_13769,N_17582);
nand U22384 (N_22384,N_13899,N_12767);
and U22385 (N_22385,N_16481,N_14027);
and U22386 (N_22386,N_12668,N_15947);
xnor U22387 (N_22387,N_15808,N_16919);
xnor U22388 (N_22388,N_13861,N_17665);
nand U22389 (N_22389,N_16411,N_14506);
nand U22390 (N_22390,N_16370,N_12543);
and U22391 (N_22391,N_13926,N_13224);
nor U22392 (N_22392,N_16500,N_12367);
xnor U22393 (N_22393,N_13675,N_14860);
nor U22394 (N_22394,N_15486,N_15425);
or U22395 (N_22395,N_16381,N_15117);
nand U22396 (N_22396,N_12476,N_16057);
nand U22397 (N_22397,N_17629,N_15111);
or U22398 (N_22398,N_15525,N_13805);
nand U22399 (N_22399,N_16269,N_12691);
or U22400 (N_22400,N_17478,N_13578);
nand U22401 (N_22401,N_13784,N_16898);
nor U22402 (N_22402,N_15429,N_17659);
or U22403 (N_22403,N_17661,N_16340);
nor U22404 (N_22404,N_15037,N_13480);
or U22405 (N_22405,N_16386,N_13483);
nor U22406 (N_22406,N_14074,N_14873);
xnor U22407 (N_22407,N_15141,N_17439);
xor U22408 (N_22408,N_12726,N_13120);
nor U22409 (N_22409,N_16879,N_15939);
xnor U22410 (N_22410,N_15102,N_15010);
xnor U22411 (N_22411,N_15683,N_12609);
or U22412 (N_22412,N_14854,N_17634);
or U22413 (N_22413,N_15540,N_15158);
nand U22414 (N_22414,N_17797,N_13033);
or U22415 (N_22415,N_14967,N_16348);
and U22416 (N_22416,N_17509,N_15235);
nor U22417 (N_22417,N_12750,N_16827);
xor U22418 (N_22418,N_15143,N_12446);
or U22419 (N_22419,N_17889,N_14997);
or U22420 (N_22420,N_14733,N_15541);
nand U22421 (N_22421,N_13049,N_17755);
xor U22422 (N_22422,N_14524,N_17955);
nand U22423 (N_22423,N_16251,N_15943);
or U22424 (N_22424,N_15689,N_13482);
and U22425 (N_22425,N_13978,N_12445);
nor U22426 (N_22426,N_15952,N_13469);
and U22427 (N_22427,N_13478,N_14234);
nand U22428 (N_22428,N_15576,N_13347);
and U22429 (N_22429,N_15421,N_17495);
and U22430 (N_22430,N_13641,N_15334);
and U22431 (N_22431,N_17310,N_16251);
xor U22432 (N_22432,N_17915,N_15362);
xnor U22433 (N_22433,N_15319,N_17281);
nand U22434 (N_22434,N_13841,N_17543);
nor U22435 (N_22435,N_13550,N_14254);
nor U22436 (N_22436,N_14542,N_14198);
xnor U22437 (N_22437,N_13243,N_16618);
nand U22438 (N_22438,N_17900,N_16153);
nor U22439 (N_22439,N_17876,N_13643);
nand U22440 (N_22440,N_17716,N_17707);
xnor U22441 (N_22441,N_16378,N_12881);
and U22442 (N_22442,N_16339,N_13081);
and U22443 (N_22443,N_14411,N_13250);
or U22444 (N_22444,N_16937,N_15072);
nor U22445 (N_22445,N_16347,N_13375);
and U22446 (N_22446,N_15844,N_12008);
nand U22447 (N_22447,N_16237,N_17640);
and U22448 (N_22448,N_16987,N_14773);
nor U22449 (N_22449,N_17354,N_13693);
or U22450 (N_22450,N_12925,N_14391);
or U22451 (N_22451,N_14987,N_14148);
nand U22452 (N_22452,N_15759,N_16390);
xnor U22453 (N_22453,N_12262,N_12040);
and U22454 (N_22454,N_13165,N_14555);
and U22455 (N_22455,N_13614,N_12609);
and U22456 (N_22456,N_15289,N_15904);
xnor U22457 (N_22457,N_14601,N_16120);
or U22458 (N_22458,N_14101,N_15776);
nor U22459 (N_22459,N_12719,N_13244);
or U22460 (N_22460,N_16821,N_12354);
or U22461 (N_22461,N_13413,N_14126);
xnor U22462 (N_22462,N_14680,N_12341);
nor U22463 (N_22463,N_16769,N_16868);
xnor U22464 (N_22464,N_16906,N_13158);
and U22465 (N_22465,N_17570,N_16888);
xor U22466 (N_22466,N_15040,N_12057);
xnor U22467 (N_22467,N_12103,N_15035);
nand U22468 (N_22468,N_16284,N_13675);
nand U22469 (N_22469,N_12416,N_15270);
and U22470 (N_22470,N_15349,N_12136);
or U22471 (N_22471,N_17669,N_16188);
or U22472 (N_22472,N_15241,N_16992);
nor U22473 (N_22473,N_15000,N_13975);
xor U22474 (N_22474,N_16278,N_15229);
xnor U22475 (N_22475,N_12659,N_13637);
or U22476 (N_22476,N_16203,N_15251);
xor U22477 (N_22477,N_15895,N_15206);
nand U22478 (N_22478,N_14159,N_16126);
or U22479 (N_22479,N_15400,N_12174);
nor U22480 (N_22480,N_17398,N_14482);
or U22481 (N_22481,N_13974,N_14946);
nand U22482 (N_22482,N_12891,N_15226);
and U22483 (N_22483,N_14787,N_12069);
and U22484 (N_22484,N_14450,N_15225);
nand U22485 (N_22485,N_12109,N_12195);
nor U22486 (N_22486,N_14013,N_12034);
nor U22487 (N_22487,N_16105,N_14704);
xnor U22488 (N_22488,N_14450,N_12791);
or U22489 (N_22489,N_16917,N_14476);
nand U22490 (N_22490,N_15525,N_12845);
nor U22491 (N_22491,N_12975,N_16668);
nor U22492 (N_22492,N_12907,N_15494);
nand U22493 (N_22493,N_17195,N_16783);
or U22494 (N_22494,N_13655,N_13923);
nor U22495 (N_22495,N_12009,N_12153);
xor U22496 (N_22496,N_15034,N_12643);
xor U22497 (N_22497,N_17804,N_13100);
nand U22498 (N_22498,N_14270,N_14608);
xnor U22499 (N_22499,N_12107,N_14799);
nor U22500 (N_22500,N_17395,N_15556);
xor U22501 (N_22501,N_13488,N_12242);
nand U22502 (N_22502,N_16576,N_12649);
and U22503 (N_22503,N_14564,N_12004);
and U22504 (N_22504,N_12761,N_15079);
or U22505 (N_22505,N_15954,N_13073);
xor U22506 (N_22506,N_12433,N_12883);
or U22507 (N_22507,N_15748,N_15497);
nand U22508 (N_22508,N_14949,N_16151);
nor U22509 (N_22509,N_16510,N_14049);
and U22510 (N_22510,N_13944,N_17924);
or U22511 (N_22511,N_14856,N_15283);
xnor U22512 (N_22512,N_15969,N_14468);
xnor U22513 (N_22513,N_17831,N_14299);
nor U22514 (N_22514,N_17728,N_12507);
nor U22515 (N_22515,N_17177,N_13636);
nand U22516 (N_22516,N_12548,N_16953);
nand U22517 (N_22517,N_14786,N_14718);
nor U22518 (N_22518,N_15247,N_14316);
and U22519 (N_22519,N_14789,N_15281);
nor U22520 (N_22520,N_15669,N_17528);
or U22521 (N_22521,N_15961,N_16522);
and U22522 (N_22522,N_13611,N_12436);
or U22523 (N_22523,N_15051,N_12091);
nand U22524 (N_22524,N_14281,N_12725);
or U22525 (N_22525,N_15207,N_13193);
nand U22526 (N_22526,N_13894,N_14398);
and U22527 (N_22527,N_13427,N_13823);
xor U22528 (N_22528,N_15446,N_16834);
and U22529 (N_22529,N_12182,N_13957);
nor U22530 (N_22530,N_12756,N_12542);
or U22531 (N_22531,N_14525,N_16487);
xnor U22532 (N_22532,N_14815,N_12801);
nand U22533 (N_22533,N_14587,N_12025);
nand U22534 (N_22534,N_12978,N_15451);
xnor U22535 (N_22535,N_17728,N_13358);
nand U22536 (N_22536,N_17303,N_13066);
nand U22537 (N_22537,N_16153,N_15764);
nor U22538 (N_22538,N_12685,N_16053);
nor U22539 (N_22539,N_14992,N_13773);
nor U22540 (N_22540,N_14138,N_16146);
nand U22541 (N_22541,N_17509,N_17766);
nor U22542 (N_22542,N_12572,N_12507);
nor U22543 (N_22543,N_13667,N_15594);
nor U22544 (N_22544,N_13876,N_16978);
or U22545 (N_22545,N_12753,N_14875);
and U22546 (N_22546,N_17604,N_15986);
nor U22547 (N_22547,N_13137,N_16788);
and U22548 (N_22548,N_13719,N_17738);
or U22549 (N_22549,N_13533,N_14287);
nand U22550 (N_22550,N_14348,N_15995);
nor U22551 (N_22551,N_16109,N_14245);
nor U22552 (N_22552,N_12712,N_15110);
xor U22553 (N_22553,N_17141,N_12710);
nand U22554 (N_22554,N_16102,N_15824);
and U22555 (N_22555,N_17491,N_12907);
nand U22556 (N_22556,N_16125,N_17365);
or U22557 (N_22557,N_12077,N_15918);
or U22558 (N_22558,N_12118,N_15324);
xor U22559 (N_22559,N_14448,N_15666);
and U22560 (N_22560,N_17428,N_15274);
xor U22561 (N_22561,N_14141,N_16309);
or U22562 (N_22562,N_17361,N_12397);
nand U22563 (N_22563,N_15866,N_12187);
nor U22564 (N_22564,N_16786,N_12070);
nand U22565 (N_22565,N_14967,N_17796);
nor U22566 (N_22566,N_13809,N_15798);
and U22567 (N_22567,N_13850,N_14471);
or U22568 (N_22568,N_13544,N_12658);
nor U22569 (N_22569,N_15639,N_13225);
or U22570 (N_22570,N_16990,N_16520);
xnor U22571 (N_22571,N_12401,N_15595);
and U22572 (N_22572,N_15366,N_14964);
and U22573 (N_22573,N_13717,N_14221);
or U22574 (N_22574,N_13109,N_17492);
or U22575 (N_22575,N_16991,N_14505);
or U22576 (N_22576,N_15002,N_16044);
xor U22577 (N_22577,N_16529,N_12569);
nor U22578 (N_22578,N_17369,N_13465);
nand U22579 (N_22579,N_13211,N_12011);
nand U22580 (N_22580,N_17294,N_14616);
or U22581 (N_22581,N_14355,N_12960);
or U22582 (N_22582,N_14330,N_15041);
or U22583 (N_22583,N_17604,N_16197);
nor U22584 (N_22584,N_16700,N_16513);
nor U22585 (N_22585,N_15978,N_12951);
and U22586 (N_22586,N_16456,N_14654);
and U22587 (N_22587,N_14126,N_17589);
nor U22588 (N_22588,N_17310,N_15646);
xnor U22589 (N_22589,N_13016,N_15906);
nand U22590 (N_22590,N_16248,N_13662);
nor U22591 (N_22591,N_14226,N_12367);
and U22592 (N_22592,N_15561,N_12049);
xor U22593 (N_22593,N_17497,N_16030);
or U22594 (N_22594,N_17861,N_15957);
nor U22595 (N_22595,N_14278,N_17948);
and U22596 (N_22596,N_17841,N_14498);
and U22597 (N_22597,N_17117,N_14231);
and U22598 (N_22598,N_12756,N_17268);
and U22599 (N_22599,N_17798,N_13621);
nand U22600 (N_22600,N_14556,N_16003);
or U22601 (N_22601,N_14398,N_17071);
xnor U22602 (N_22602,N_12867,N_16887);
xnor U22603 (N_22603,N_16815,N_15211);
and U22604 (N_22604,N_16562,N_15107);
xor U22605 (N_22605,N_17157,N_13850);
xor U22606 (N_22606,N_16503,N_16340);
or U22607 (N_22607,N_16027,N_14182);
nor U22608 (N_22608,N_14649,N_13981);
xor U22609 (N_22609,N_17257,N_14692);
nor U22610 (N_22610,N_16197,N_16451);
xnor U22611 (N_22611,N_16193,N_14328);
nand U22612 (N_22612,N_17754,N_12899);
and U22613 (N_22613,N_13379,N_12599);
or U22614 (N_22614,N_16355,N_15660);
nor U22615 (N_22615,N_14218,N_17459);
nand U22616 (N_22616,N_15522,N_17206);
xor U22617 (N_22617,N_13133,N_16187);
or U22618 (N_22618,N_17560,N_13063);
xnor U22619 (N_22619,N_15201,N_15401);
xnor U22620 (N_22620,N_16009,N_15952);
or U22621 (N_22621,N_15849,N_14485);
xnor U22622 (N_22622,N_15882,N_15935);
nor U22623 (N_22623,N_17486,N_13835);
xor U22624 (N_22624,N_15531,N_16685);
nand U22625 (N_22625,N_17087,N_16050);
xnor U22626 (N_22626,N_14007,N_14712);
xnor U22627 (N_22627,N_15604,N_17284);
and U22628 (N_22628,N_17624,N_15410);
nor U22629 (N_22629,N_17288,N_14018);
xnor U22630 (N_22630,N_13581,N_12822);
or U22631 (N_22631,N_16378,N_14562);
nand U22632 (N_22632,N_16048,N_15540);
and U22633 (N_22633,N_17691,N_14381);
or U22634 (N_22634,N_13411,N_17800);
nor U22635 (N_22635,N_15074,N_12231);
xor U22636 (N_22636,N_12329,N_17521);
nand U22637 (N_22637,N_12298,N_16993);
xor U22638 (N_22638,N_14811,N_15296);
nand U22639 (N_22639,N_14160,N_12368);
and U22640 (N_22640,N_13260,N_14838);
nand U22641 (N_22641,N_14478,N_15637);
or U22642 (N_22642,N_17713,N_12422);
nor U22643 (N_22643,N_15529,N_15793);
xor U22644 (N_22644,N_15266,N_13638);
xor U22645 (N_22645,N_17764,N_13635);
xnor U22646 (N_22646,N_17406,N_15696);
or U22647 (N_22647,N_16970,N_12901);
or U22648 (N_22648,N_17681,N_15265);
and U22649 (N_22649,N_13365,N_16828);
or U22650 (N_22650,N_17962,N_14844);
nor U22651 (N_22651,N_12149,N_17618);
nand U22652 (N_22652,N_17650,N_16112);
nor U22653 (N_22653,N_15577,N_16923);
nor U22654 (N_22654,N_14511,N_15398);
nor U22655 (N_22655,N_13077,N_16902);
or U22656 (N_22656,N_15361,N_13730);
xor U22657 (N_22657,N_16244,N_14522);
nor U22658 (N_22658,N_16383,N_12458);
xor U22659 (N_22659,N_16445,N_14309);
nand U22660 (N_22660,N_12916,N_12851);
nor U22661 (N_22661,N_15718,N_15972);
or U22662 (N_22662,N_17621,N_13113);
nand U22663 (N_22663,N_12057,N_16738);
nor U22664 (N_22664,N_14347,N_15680);
nor U22665 (N_22665,N_15218,N_14917);
nor U22666 (N_22666,N_12524,N_16037);
xor U22667 (N_22667,N_17632,N_12508);
xnor U22668 (N_22668,N_13075,N_12559);
and U22669 (N_22669,N_15070,N_16582);
nor U22670 (N_22670,N_14046,N_15567);
xnor U22671 (N_22671,N_12057,N_14719);
xnor U22672 (N_22672,N_14240,N_14287);
and U22673 (N_22673,N_15185,N_17527);
nor U22674 (N_22674,N_14252,N_17121);
nor U22675 (N_22675,N_16414,N_16146);
or U22676 (N_22676,N_15907,N_13436);
and U22677 (N_22677,N_17457,N_12267);
nor U22678 (N_22678,N_16785,N_13059);
and U22679 (N_22679,N_17587,N_15447);
and U22680 (N_22680,N_15030,N_14250);
or U22681 (N_22681,N_12761,N_13210);
nor U22682 (N_22682,N_14372,N_14397);
nand U22683 (N_22683,N_14106,N_12456);
or U22684 (N_22684,N_13697,N_16296);
nand U22685 (N_22685,N_15332,N_14352);
nand U22686 (N_22686,N_15959,N_17567);
and U22687 (N_22687,N_13439,N_15016);
or U22688 (N_22688,N_16673,N_15068);
and U22689 (N_22689,N_16151,N_17068);
nand U22690 (N_22690,N_15976,N_17295);
nand U22691 (N_22691,N_14064,N_12800);
and U22692 (N_22692,N_12979,N_12683);
xor U22693 (N_22693,N_16507,N_12204);
nand U22694 (N_22694,N_17804,N_13814);
and U22695 (N_22695,N_15657,N_12223);
nand U22696 (N_22696,N_17174,N_14489);
nor U22697 (N_22697,N_12373,N_12327);
or U22698 (N_22698,N_14197,N_14179);
nor U22699 (N_22699,N_12670,N_14551);
nand U22700 (N_22700,N_15276,N_16271);
and U22701 (N_22701,N_17782,N_17835);
and U22702 (N_22702,N_12746,N_17844);
and U22703 (N_22703,N_12300,N_12213);
nor U22704 (N_22704,N_14768,N_15608);
and U22705 (N_22705,N_17784,N_13610);
xor U22706 (N_22706,N_15517,N_12489);
or U22707 (N_22707,N_14001,N_17575);
nor U22708 (N_22708,N_12193,N_13966);
nor U22709 (N_22709,N_12937,N_17036);
and U22710 (N_22710,N_12593,N_17195);
or U22711 (N_22711,N_17087,N_14113);
nor U22712 (N_22712,N_15177,N_12015);
and U22713 (N_22713,N_14251,N_16160);
xor U22714 (N_22714,N_13035,N_16426);
or U22715 (N_22715,N_14131,N_13978);
xor U22716 (N_22716,N_14511,N_14479);
nor U22717 (N_22717,N_12664,N_12295);
or U22718 (N_22718,N_15379,N_12008);
and U22719 (N_22719,N_15543,N_15411);
xnor U22720 (N_22720,N_13275,N_14922);
xnor U22721 (N_22721,N_13387,N_13671);
and U22722 (N_22722,N_14763,N_13933);
nand U22723 (N_22723,N_14441,N_13094);
xor U22724 (N_22724,N_12634,N_14048);
nor U22725 (N_22725,N_14974,N_15482);
xor U22726 (N_22726,N_16767,N_12846);
nand U22727 (N_22727,N_12343,N_16764);
nor U22728 (N_22728,N_15538,N_13257);
or U22729 (N_22729,N_16967,N_12037);
xor U22730 (N_22730,N_17024,N_14497);
or U22731 (N_22731,N_13956,N_17944);
and U22732 (N_22732,N_14411,N_17434);
nand U22733 (N_22733,N_17313,N_16881);
or U22734 (N_22734,N_16747,N_13466);
xor U22735 (N_22735,N_16452,N_14309);
and U22736 (N_22736,N_17636,N_17391);
xnor U22737 (N_22737,N_15159,N_16110);
nand U22738 (N_22738,N_17605,N_12539);
and U22739 (N_22739,N_17202,N_14950);
or U22740 (N_22740,N_15300,N_13652);
and U22741 (N_22741,N_16452,N_16041);
or U22742 (N_22742,N_15646,N_17236);
nand U22743 (N_22743,N_13429,N_16373);
or U22744 (N_22744,N_15807,N_17938);
or U22745 (N_22745,N_16950,N_12221);
or U22746 (N_22746,N_15918,N_13755);
or U22747 (N_22747,N_12283,N_16696);
nand U22748 (N_22748,N_13606,N_15823);
and U22749 (N_22749,N_16056,N_17712);
and U22750 (N_22750,N_13226,N_15777);
nor U22751 (N_22751,N_17114,N_13498);
nor U22752 (N_22752,N_14170,N_15498);
nor U22753 (N_22753,N_12099,N_16970);
nor U22754 (N_22754,N_14197,N_17770);
xnor U22755 (N_22755,N_16135,N_17864);
xnor U22756 (N_22756,N_14204,N_16978);
nand U22757 (N_22757,N_12486,N_15524);
nand U22758 (N_22758,N_13957,N_13106);
and U22759 (N_22759,N_16436,N_17618);
nand U22760 (N_22760,N_13935,N_13086);
nand U22761 (N_22761,N_17931,N_14360);
or U22762 (N_22762,N_13004,N_16919);
nor U22763 (N_22763,N_17216,N_12138);
nor U22764 (N_22764,N_12199,N_17173);
nor U22765 (N_22765,N_16221,N_16136);
xor U22766 (N_22766,N_15607,N_12092);
nand U22767 (N_22767,N_13667,N_17824);
nor U22768 (N_22768,N_15831,N_14662);
xor U22769 (N_22769,N_14874,N_14462);
nand U22770 (N_22770,N_17935,N_13368);
and U22771 (N_22771,N_14451,N_16162);
xnor U22772 (N_22772,N_14923,N_14120);
xnor U22773 (N_22773,N_14949,N_13856);
xor U22774 (N_22774,N_14749,N_14540);
nor U22775 (N_22775,N_17565,N_17162);
nor U22776 (N_22776,N_14057,N_14548);
xnor U22777 (N_22777,N_15692,N_12640);
and U22778 (N_22778,N_16880,N_16306);
and U22779 (N_22779,N_16225,N_14455);
nor U22780 (N_22780,N_15896,N_14634);
and U22781 (N_22781,N_17979,N_15355);
nor U22782 (N_22782,N_17178,N_15047);
or U22783 (N_22783,N_12102,N_16014);
xnor U22784 (N_22784,N_15587,N_15561);
and U22785 (N_22785,N_13335,N_17854);
xor U22786 (N_22786,N_17779,N_13009);
or U22787 (N_22787,N_12679,N_13051);
and U22788 (N_22788,N_14569,N_16342);
nand U22789 (N_22789,N_12167,N_14132);
and U22790 (N_22790,N_13597,N_15504);
xnor U22791 (N_22791,N_15045,N_12914);
nand U22792 (N_22792,N_12877,N_15424);
and U22793 (N_22793,N_12227,N_13049);
xnor U22794 (N_22794,N_16848,N_12412);
nor U22795 (N_22795,N_13428,N_14509);
nand U22796 (N_22796,N_12230,N_14997);
nand U22797 (N_22797,N_15093,N_16297);
xor U22798 (N_22798,N_14198,N_13856);
xor U22799 (N_22799,N_14301,N_17028);
nor U22800 (N_22800,N_14583,N_12194);
and U22801 (N_22801,N_15293,N_17764);
nor U22802 (N_22802,N_16720,N_17694);
nand U22803 (N_22803,N_15054,N_12765);
nand U22804 (N_22804,N_17362,N_16407);
or U22805 (N_22805,N_16284,N_12401);
or U22806 (N_22806,N_14548,N_12562);
nand U22807 (N_22807,N_13640,N_13004);
or U22808 (N_22808,N_12108,N_17090);
nand U22809 (N_22809,N_16021,N_16649);
nor U22810 (N_22810,N_17532,N_15679);
nand U22811 (N_22811,N_17809,N_12502);
xor U22812 (N_22812,N_17323,N_13994);
or U22813 (N_22813,N_15505,N_15814);
or U22814 (N_22814,N_14883,N_13830);
nor U22815 (N_22815,N_14156,N_14334);
and U22816 (N_22816,N_12926,N_15452);
xor U22817 (N_22817,N_16663,N_16024);
nand U22818 (N_22818,N_13398,N_16296);
or U22819 (N_22819,N_17970,N_17001);
or U22820 (N_22820,N_15911,N_12719);
or U22821 (N_22821,N_15181,N_13108);
xnor U22822 (N_22822,N_16935,N_12387);
and U22823 (N_22823,N_16582,N_14002);
nand U22824 (N_22824,N_14326,N_15955);
and U22825 (N_22825,N_15564,N_13778);
nand U22826 (N_22826,N_15274,N_17039);
nand U22827 (N_22827,N_17612,N_13410);
and U22828 (N_22828,N_14249,N_17773);
and U22829 (N_22829,N_13262,N_16646);
or U22830 (N_22830,N_16865,N_17352);
nand U22831 (N_22831,N_17947,N_13812);
or U22832 (N_22832,N_13497,N_14722);
nor U22833 (N_22833,N_14040,N_17648);
and U22834 (N_22834,N_14610,N_16927);
or U22835 (N_22835,N_13981,N_15308);
xor U22836 (N_22836,N_12210,N_12129);
and U22837 (N_22837,N_13240,N_14789);
and U22838 (N_22838,N_16568,N_14465);
xnor U22839 (N_22839,N_15250,N_12624);
xor U22840 (N_22840,N_16933,N_14916);
or U22841 (N_22841,N_13113,N_16420);
and U22842 (N_22842,N_14728,N_12474);
nor U22843 (N_22843,N_13887,N_12585);
nor U22844 (N_22844,N_17543,N_16429);
nor U22845 (N_22845,N_15866,N_13901);
and U22846 (N_22846,N_12420,N_17131);
and U22847 (N_22847,N_15867,N_14453);
nand U22848 (N_22848,N_12148,N_12769);
xnor U22849 (N_22849,N_14721,N_16116);
xor U22850 (N_22850,N_15505,N_17131);
nand U22851 (N_22851,N_14056,N_13296);
or U22852 (N_22852,N_14354,N_17597);
and U22853 (N_22853,N_12446,N_12675);
nand U22854 (N_22854,N_13921,N_12510);
xnor U22855 (N_22855,N_15688,N_15344);
nor U22856 (N_22856,N_15555,N_16225);
nand U22857 (N_22857,N_17387,N_16074);
or U22858 (N_22858,N_13716,N_12328);
and U22859 (N_22859,N_12501,N_16345);
or U22860 (N_22860,N_16155,N_14591);
nand U22861 (N_22861,N_12555,N_14422);
nand U22862 (N_22862,N_17487,N_12907);
nor U22863 (N_22863,N_12724,N_12063);
nand U22864 (N_22864,N_14997,N_14672);
and U22865 (N_22865,N_17231,N_17616);
nand U22866 (N_22866,N_12723,N_15795);
xor U22867 (N_22867,N_17454,N_13518);
nor U22868 (N_22868,N_16349,N_13277);
or U22869 (N_22869,N_12730,N_14332);
nor U22870 (N_22870,N_16027,N_14786);
or U22871 (N_22871,N_13595,N_14194);
or U22872 (N_22872,N_12117,N_13353);
nor U22873 (N_22873,N_15724,N_17826);
and U22874 (N_22874,N_16751,N_17695);
or U22875 (N_22875,N_17557,N_17191);
and U22876 (N_22876,N_12062,N_14983);
nand U22877 (N_22877,N_14372,N_14080);
or U22878 (N_22878,N_17375,N_14016);
or U22879 (N_22879,N_16138,N_17275);
nor U22880 (N_22880,N_16897,N_12850);
nor U22881 (N_22881,N_17733,N_13153);
and U22882 (N_22882,N_16486,N_17339);
xor U22883 (N_22883,N_17763,N_13918);
and U22884 (N_22884,N_15322,N_12417);
and U22885 (N_22885,N_17139,N_12758);
and U22886 (N_22886,N_14523,N_14710);
xnor U22887 (N_22887,N_13718,N_17962);
nand U22888 (N_22888,N_15617,N_16635);
xnor U22889 (N_22889,N_14457,N_12231);
nand U22890 (N_22890,N_12363,N_13745);
xor U22891 (N_22891,N_16807,N_15263);
and U22892 (N_22892,N_14773,N_16454);
or U22893 (N_22893,N_13934,N_12629);
and U22894 (N_22894,N_14056,N_16562);
and U22895 (N_22895,N_14692,N_16547);
nor U22896 (N_22896,N_13721,N_12309);
or U22897 (N_22897,N_15239,N_16913);
nor U22898 (N_22898,N_16832,N_12573);
and U22899 (N_22899,N_16704,N_13642);
or U22900 (N_22900,N_14529,N_17541);
nor U22901 (N_22901,N_14523,N_12129);
nor U22902 (N_22902,N_15589,N_15213);
nand U22903 (N_22903,N_17036,N_15940);
xor U22904 (N_22904,N_14546,N_16574);
and U22905 (N_22905,N_17296,N_17839);
or U22906 (N_22906,N_13366,N_14552);
nand U22907 (N_22907,N_16446,N_13128);
xnor U22908 (N_22908,N_16630,N_17096);
or U22909 (N_22909,N_17248,N_17847);
xnor U22910 (N_22910,N_16587,N_13732);
nor U22911 (N_22911,N_14779,N_16567);
nand U22912 (N_22912,N_14715,N_15650);
nand U22913 (N_22913,N_16956,N_12369);
xor U22914 (N_22914,N_17205,N_14776);
nor U22915 (N_22915,N_16987,N_15547);
nor U22916 (N_22916,N_16695,N_16675);
nand U22917 (N_22917,N_12979,N_13607);
nor U22918 (N_22918,N_17960,N_14778);
nand U22919 (N_22919,N_12531,N_14950);
nand U22920 (N_22920,N_15936,N_14692);
nor U22921 (N_22921,N_14200,N_13997);
or U22922 (N_22922,N_14488,N_12885);
or U22923 (N_22923,N_17583,N_17999);
xor U22924 (N_22924,N_14570,N_14614);
and U22925 (N_22925,N_14316,N_17038);
xor U22926 (N_22926,N_16736,N_15602);
and U22927 (N_22927,N_13137,N_12606);
nand U22928 (N_22928,N_13934,N_15241);
and U22929 (N_22929,N_13751,N_14765);
or U22930 (N_22930,N_13013,N_16192);
xor U22931 (N_22931,N_15965,N_16978);
nand U22932 (N_22932,N_14525,N_14526);
and U22933 (N_22933,N_14679,N_16590);
nor U22934 (N_22934,N_14526,N_16073);
and U22935 (N_22935,N_13914,N_15312);
xor U22936 (N_22936,N_17201,N_16884);
nand U22937 (N_22937,N_12088,N_16851);
or U22938 (N_22938,N_17530,N_15122);
xnor U22939 (N_22939,N_12421,N_12288);
and U22940 (N_22940,N_15032,N_16461);
nand U22941 (N_22941,N_14286,N_15178);
nor U22942 (N_22942,N_12635,N_16445);
or U22943 (N_22943,N_13825,N_13740);
nor U22944 (N_22944,N_13858,N_13651);
nor U22945 (N_22945,N_17793,N_16697);
xor U22946 (N_22946,N_13919,N_12776);
or U22947 (N_22947,N_13015,N_16234);
nand U22948 (N_22948,N_15046,N_14068);
nor U22949 (N_22949,N_17114,N_14369);
xor U22950 (N_22950,N_15102,N_16071);
nand U22951 (N_22951,N_14410,N_17342);
nor U22952 (N_22952,N_12514,N_17696);
nand U22953 (N_22953,N_16808,N_17044);
xnor U22954 (N_22954,N_15322,N_14678);
nand U22955 (N_22955,N_17463,N_16755);
and U22956 (N_22956,N_17237,N_15646);
nand U22957 (N_22957,N_13893,N_16064);
xor U22958 (N_22958,N_17067,N_17863);
nand U22959 (N_22959,N_12067,N_13627);
and U22960 (N_22960,N_13906,N_13632);
or U22961 (N_22961,N_13964,N_15784);
and U22962 (N_22962,N_15537,N_17777);
nor U22963 (N_22963,N_13345,N_16571);
and U22964 (N_22964,N_13741,N_14922);
nor U22965 (N_22965,N_12465,N_15061);
or U22966 (N_22966,N_17411,N_17047);
xor U22967 (N_22967,N_17291,N_14280);
or U22968 (N_22968,N_15383,N_16073);
or U22969 (N_22969,N_16137,N_17114);
nand U22970 (N_22970,N_17971,N_15303);
and U22971 (N_22971,N_14973,N_14021);
nor U22972 (N_22972,N_17027,N_15668);
xor U22973 (N_22973,N_16677,N_16573);
and U22974 (N_22974,N_17998,N_17967);
xnor U22975 (N_22975,N_14555,N_15860);
and U22976 (N_22976,N_12215,N_16697);
or U22977 (N_22977,N_12686,N_13122);
and U22978 (N_22978,N_14523,N_16469);
or U22979 (N_22979,N_12033,N_15254);
nor U22980 (N_22980,N_16748,N_16117);
and U22981 (N_22981,N_13253,N_16543);
and U22982 (N_22982,N_15618,N_15871);
nor U22983 (N_22983,N_12737,N_12781);
or U22984 (N_22984,N_16603,N_14447);
or U22985 (N_22985,N_12982,N_13591);
or U22986 (N_22986,N_16944,N_12154);
nand U22987 (N_22987,N_16220,N_16518);
nor U22988 (N_22988,N_16656,N_13332);
and U22989 (N_22989,N_17086,N_17576);
nor U22990 (N_22990,N_15907,N_14979);
and U22991 (N_22991,N_13456,N_15960);
and U22992 (N_22992,N_17987,N_15507);
or U22993 (N_22993,N_14848,N_15135);
nand U22994 (N_22994,N_15205,N_15051);
xnor U22995 (N_22995,N_14079,N_17489);
xnor U22996 (N_22996,N_13460,N_13130);
and U22997 (N_22997,N_14924,N_13016);
and U22998 (N_22998,N_12346,N_15139);
or U22999 (N_22999,N_14628,N_14589);
xor U23000 (N_23000,N_14588,N_17078);
and U23001 (N_23001,N_13569,N_16231);
nor U23002 (N_23002,N_17775,N_13466);
or U23003 (N_23003,N_14583,N_17840);
xor U23004 (N_23004,N_14899,N_14781);
nor U23005 (N_23005,N_16063,N_13984);
nand U23006 (N_23006,N_12551,N_15564);
nor U23007 (N_23007,N_15325,N_17185);
and U23008 (N_23008,N_15785,N_16221);
and U23009 (N_23009,N_13893,N_15508);
or U23010 (N_23010,N_17731,N_17273);
nor U23011 (N_23011,N_15712,N_12534);
or U23012 (N_23012,N_15779,N_17771);
and U23013 (N_23013,N_16015,N_14236);
nand U23014 (N_23014,N_14078,N_16356);
xnor U23015 (N_23015,N_14323,N_17120);
and U23016 (N_23016,N_15852,N_16003);
nor U23017 (N_23017,N_16039,N_12476);
nand U23018 (N_23018,N_16947,N_14391);
or U23019 (N_23019,N_14561,N_13811);
nor U23020 (N_23020,N_12124,N_16922);
nand U23021 (N_23021,N_12599,N_16783);
and U23022 (N_23022,N_14490,N_15434);
nand U23023 (N_23023,N_15282,N_12310);
nand U23024 (N_23024,N_14485,N_16668);
nor U23025 (N_23025,N_13401,N_16027);
or U23026 (N_23026,N_16965,N_16499);
nor U23027 (N_23027,N_17557,N_16126);
nand U23028 (N_23028,N_13764,N_13165);
xnor U23029 (N_23029,N_17578,N_13227);
nand U23030 (N_23030,N_17859,N_17483);
nand U23031 (N_23031,N_12378,N_15228);
or U23032 (N_23032,N_15946,N_13824);
and U23033 (N_23033,N_13473,N_16963);
nand U23034 (N_23034,N_17287,N_14201);
xor U23035 (N_23035,N_12402,N_14317);
nand U23036 (N_23036,N_12690,N_13163);
and U23037 (N_23037,N_16832,N_16854);
xnor U23038 (N_23038,N_17311,N_17954);
nor U23039 (N_23039,N_12127,N_12632);
nand U23040 (N_23040,N_12438,N_17208);
nand U23041 (N_23041,N_15432,N_12768);
and U23042 (N_23042,N_12783,N_17438);
nand U23043 (N_23043,N_17099,N_12704);
xor U23044 (N_23044,N_12117,N_12156);
xor U23045 (N_23045,N_15358,N_16289);
nor U23046 (N_23046,N_13895,N_14048);
nor U23047 (N_23047,N_15741,N_12160);
nand U23048 (N_23048,N_15477,N_13546);
nand U23049 (N_23049,N_16856,N_16455);
nand U23050 (N_23050,N_13209,N_16854);
xor U23051 (N_23051,N_12327,N_16492);
nand U23052 (N_23052,N_17500,N_12290);
xnor U23053 (N_23053,N_12296,N_17212);
or U23054 (N_23054,N_17227,N_17506);
xor U23055 (N_23055,N_14494,N_12376);
or U23056 (N_23056,N_14520,N_14993);
or U23057 (N_23057,N_17212,N_15400);
nor U23058 (N_23058,N_17788,N_13892);
nor U23059 (N_23059,N_17272,N_17850);
xor U23060 (N_23060,N_17895,N_16883);
nor U23061 (N_23061,N_12064,N_15706);
nand U23062 (N_23062,N_16263,N_14099);
xnor U23063 (N_23063,N_16988,N_12591);
and U23064 (N_23064,N_16266,N_16232);
or U23065 (N_23065,N_15961,N_15786);
or U23066 (N_23066,N_17726,N_12695);
nor U23067 (N_23067,N_15819,N_13613);
nor U23068 (N_23068,N_17210,N_12762);
and U23069 (N_23069,N_13085,N_12261);
or U23070 (N_23070,N_12706,N_16449);
nand U23071 (N_23071,N_17022,N_16765);
nand U23072 (N_23072,N_16909,N_16136);
xnor U23073 (N_23073,N_12390,N_17487);
nand U23074 (N_23074,N_13925,N_14202);
nor U23075 (N_23075,N_16377,N_14086);
xnor U23076 (N_23076,N_15712,N_17195);
nand U23077 (N_23077,N_15147,N_15355);
nor U23078 (N_23078,N_15357,N_12972);
xnor U23079 (N_23079,N_12511,N_12456);
or U23080 (N_23080,N_17237,N_15723);
or U23081 (N_23081,N_13902,N_14815);
nor U23082 (N_23082,N_16108,N_16195);
xnor U23083 (N_23083,N_13780,N_13222);
nand U23084 (N_23084,N_17866,N_16727);
nor U23085 (N_23085,N_14671,N_14502);
or U23086 (N_23086,N_16164,N_15825);
xor U23087 (N_23087,N_14909,N_14269);
xor U23088 (N_23088,N_16742,N_16282);
or U23089 (N_23089,N_13548,N_13061);
xnor U23090 (N_23090,N_17754,N_16739);
xor U23091 (N_23091,N_16527,N_16570);
nor U23092 (N_23092,N_14527,N_13036);
or U23093 (N_23093,N_16001,N_12519);
and U23094 (N_23094,N_16706,N_14824);
xnor U23095 (N_23095,N_17366,N_17766);
nand U23096 (N_23096,N_14641,N_17419);
nand U23097 (N_23097,N_14057,N_17530);
and U23098 (N_23098,N_15687,N_17551);
xor U23099 (N_23099,N_12552,N_14428);
nand U23100 (N_23100,N_17194,N_17933);
or U23101 (N_23101,N_17666,N_14133);
or U23102 (N_23102,N_13621,N_12570);
nand U23103 (N_23103,N_13118,N_12102);
nor U23104 (N_23104,N_12975,N_17543);
nand U23105 (N_23105,N_17624,N_17497);
and U23106 (N_23106,N_14462,N_15099);
nor U23107 (N_23107,N_12479,N_17752);
nand U23108 (N_23108,N_15114,N_14902);
and U23109 (N_23109,N_15931,N_16611);
xor U23110 (N_23110,N_14607,N_13926);
nor U23111 (N_23111,N_13422,N_13054);
and U23112 (N_23112,N_16207,N_16013);
nand U23113 (N_23113,N_16020,N_12961);
and U23114 (N_23114,N_17128,N_15557);
and U23115 (N_23115,N_14531,N_13371);
or U23116 (N_23116,N_12150,N_14172);
and U23117 (N_23117,N_16449,N_14571);
and U23118 (N_23118,N_14421,N_15520);
and U23119 (N_23119,N_12965,N_16761);
and U23120 (N_23120,N_15994,N_12959);
nor U23121 (N_23121,N_17474,N_16002);
and U23122 (N_23122,N_14922,N_17617);
nand U23123 (N_23123,N_16422,N_12254);
or U23124 (N_23124,N_16870,N_16964);
or U23125 (N_23125,N_12651,N_16619);
nor U23126 (N_23126,N_14821,N_16600);
nor U23127 (N_23127,N_16651,N_13327);
or U23128 (N_23128,N_17482,N_15329);
or U23129 (N_23129,N_15623,N_16631);
nand U23130 (N_23130,N_16040,N_13410);
nand U23131 (N_23131,N_15598,N_15357);
nand U23132 (N_23132,N_17513,N_14506);
or U23133 (N_23133,N_16367,N_17714);
nand U23134 (N_23134,N_14749,N_13699);
nand U23135 (N_23135,N_17205,N_16690);
nand U23136 (N_23136,N_16452,N_17145);
nand U23137 (N_23137,N_13262,N_16010);
xor U23138 (N_23138,N_14744,N_12041);
or U23139 (N_23139,N_14568,N_17699);
nor U23140 (N_23140,N_15334,N_15498);
xnor U23141 (N_23141,N_15686,N_15629);
xor U23142 (N_23142,N_16805,N_15028);
nor U23143 (N_23143,N_16401,N_17522);
nand U23144 (N_23144,N_13341,N_15042);
or U23145 (N_23145,N_13750,N_13206);
and U23146 (N_23146,N_15832,N_15684);
nor U23147 (N_23147,N_13039,N_13457);
nor U23148 (N_23148,N_17247,N_13521);
xnor U23149 (N_23149,N_16937,N_12180);
xnor U23150 (N_23150,N_17858,N_12109);
xnor U23151 (N_23151,N_13745,N_13929);
nand U23152 (N_23152,N_17021,N_17137);
xnor U23153 (N_23153,N_15425,N_13866);
or U23154 (N_23154,N_12848,N_14938);
xor U23155 (N_23155,N_16854,N_16293);
and U23156 (N_23156,N_17433,N_14809);
xnor U23157 (N_23157,N_17331,N_12199);
or U23158 (N_23158,N_16811,N_12624);
nor U23159 (N_23159,N_17136,N_14795);
and U23160 (N_23160,N_12875,N_16402);
nand U23161 (N_23161,N_13391,N_16507);
or U23162 (N_23162,N_16464,N_15477);
or U23163 (N_23163,N_15065,N_17760);
and U23164 (N_23164,N_12066,N_16292);
or U23165 (N_23165,N_14060,N_14749);
or U23166 (N_23166,N_12779,N_12675);
xor U23167 (N_23167,N_14403,N_14402);
xnor U23168 (N_23168,N_15467,N_14877);
and U23169 (N_23169,N_15013,N_15536);
nor U23170 (N_23170,N_12765,N_13627);
nand U23171 (N_23171,N_16024,N_17468);
nand U23172 (N_23172,N_12871,N_16723);
nor U23173 (N_23173,N_17921,N_13545);
xnor U23174 (N_23174,N_17554,N_17537);
nor U23175 (N_23175,N_16686,N_17372);
xor U23176 (N_23176,N_17970,N_14443);
and U23177 (N_23177,N_16599,N_13930);
nor U23178 (N_23178,N_13477,N_17576);
or U23179 (N_23179,N_15321,N_15158);
or U23180 (N_23180,N_12554,N_16919);
xnor U23181 (N_23181,N_17684,N_16361);
or U23182 (N_23182,N_17233,N_15941);
nor U23183 (N_23183,N_13344,N_17699);
xor U23184 (N_23184,N_17960,N_13375);
nand U23185 (N_23185,N_14154,N_17594);
nor U23186 (N_23186,N_12794,N_17200);
or U23187 (N_23187,N_16323,N_16676);
and U23188 (N_23188,N_13287,N_16372);
or U23189 (N_23189,N_16659,N_16836);
xnor U23190 (N_23190,N_12929,N_16487);
xnor U23191 (N_23191,N_12941,N_12413);
and U23192 (N_23192,N_17518,N_15382);
and U23193 (N_23193,N_17098,N_13907);
xnor U23194 (N_23194,N_12286,N_17874);
and U23195 (N_23195,N_14820,N_15133);
and U23196 (N_23196,N_17956,N_17736);
and U23197 (N_23197,N_16081,N_17638);
nor U23198 (N_23198,N_16720,N_17606);
and U23199 (N_23199,N_16541,N_17573);
nand U23200 (N_23200,N_13709,N_14993);
nand U23201 (N_23201,N_16211,N_12311);
or U23202 (N_23202,N_17914,N_16561);
xor U23203 (N_23203,N_15004,N_16100);
or U23204 (N_23204,N_13202,N_16669);
nor U23205 (N_23205,N_14881,N_12365);
nor U23206 (N_23206,N_13248,N_16831);
xnor U23207 (N_23207,N_15595,N_17566);
or U23208 (N_23208,N_14557,N_13153);
or U23209 (N_23209,N_14264,N_17276);
xnor U23210 (N_23210,N_13335,N_14551);
and U23211 (N_23211,N_12921,N_17618);
nor U23212 (N_23212,N_12178,N_13497);
nand U23213 (N_23213,N_12432,N_16958);
and U23214 (N_23214,N_12387,N_12353);
xor U23215 (N_23215,N_15385,N_14880);
nand U23216 (N_23216,N_13731,N_14564);
and U23217 (N_23217,N_13707,N_12724);
nand U23218 (N_23218,N_17589,N_16132);
nand U23219 (N_23219,N_16038,N_14701);
or U23220 (N_23220,N_12218,N_12282);
xor U23221 (N_23221,N_12908,N_15703);
nand U23222 (N_23222,N_14705,N_13355);
and U23223 (N_23223,N_16246,N_14250);
or U23224 (N_23224,N_17200,N_15024);
nor U23225 (N_23225,N_13459,N_14897);
and U23226 (N_23226,N_13078,N_12376);
nand U23227 (N_23227,N_13118,N_14795);
xor U23228 (N_23228,N_15099,N_17885);
and U23229 (N_23229,N_17940,N_17887);
nor U23230 (N_23230,N_17027,N_16001);
nand U23231 (N_23231,N_13317,N_13768);
and U23232 (N_23232,N_14258,N_13362);
nor U23233 (N_23233,N_12949,N_12320);
or U23234 (N_23234,N_17875,N_17372);
xor U23235 (N_23235,N_14007,N_15823);
and U23236 (N_23236,N_15362,N_12902);
nand U23237 (N_23237,N_17456,N_14060);
or U23238 (N_23238,N_12470,N_16153);
xnor U23239 (N_23239,N_15751,N_14485);
or U23240 (N_23240,N_16306,N_16588);
nand U23241 (N_23241,N_14495,N_17577);
nor U23242 (N_23242,N_17026,N_13956);
nor U23243 (N_23243,N_15254,N_12983);
nand U23244 (N_23244,N_17579,N_13103);
nor U23245 (N_23245,N_16207,N_15191);
nand U23246 (N_23246,N_14959,N_17858);
xnor U23247 (N_23247,N_16540,N_15040);
nor U23248 (N_23248,N_13988,N_17888);
nor U23249 (N_23249,N_17867,N_14084);
and U23250 (N_23250,N_13918,N_15804);
nor U23251 (N_23251,N_16825,N_14105);
nand U23252 (N_23252,N_14513,N_16158);
xnor U23253 (N_23253,N_17101,N_14307);
or U23254 (N_23254,N_12974,N_14080);
nor U23255 (N_23255,N_13079,N_14563);
or U23256 (N_23256,N_14437,N_14842);
xor U23257 (N_23257,N_13332,N_17038);
nand U23258 (N_23258,N_16410,N_12723);
nor U23259 (N_23259,N_13627,N_12708);
xnor U23260 (N_23260,N_17532,N_17462);
xnor U23261 (N_23261,N_14717,N_13701);
nor U23262 (N_23262,N_13782,N_15452);
xor U23263 (N_23263,N_16325,N_13680);
nor U23264 (N_23264,N_15087,N_13142);
or U23265 (N_23265,N_12728,N_17878);
xnor U23266 (N_23266,N_14107,N_12568);
nor U23267 (N_23267,N_16261,N_12625);
xnor U23268 (N_23268,N_13341,N_17437);
and U23269 (N_23269,N_15136,N_12355);
and U23270 (N_23270,N_12754,N_14776);
or U23271 (N_23271,N_13262,N_13264);
or U23272 (N_23272,N_17626,N_13236);
xor U23273 (N_23273,N_16202,N_12085);
and U23274 (N_23274,N_13603,N_15257);
xnor U23275 (N_23275,N_17809,N_14865);
nor U23276 (N_23276,N_17127,N_14718);
xnor U23277 (N_23277,N_14406,N_15545);
and U23278 (N_23278,N_12651,N_15567);
nor U23279 (N_23279,N_13865,N_14398);
xnor U23280 (N_23280,N_13975,N_13657);
nand U23281 (N_23281,N_15364,N_12435);
nor U23282 (N_23282,N_15969,N_14930);
and U23283 (N_23283,N_13402,N_16242);
and U23284 (N_23284,N_17236,N_13046);
and U23285 (N_23285,N_14245,N_17638);
nand U23286 (N_23286,N_12501,N_14142);
or U23287 (N_23287,N_12204,N_13868);
xor U23288 (N_23288,N_12347,N_13089);
or U23289 (N_23289,N_17064,N_16221);
nand U23290 (N_23290,N_15863,N_15064);
and U23291 (N_23291,N_15215,N_15516);
xnor U23292 (N_23292,N_12822,N_12571);
nand U23293 (N_23293,N_14221,N_14352);
or U23294 (N_23294,N_13999,N_16544);
nand U23295 (N_23295,N_14056,N_16459);
or U23296 (N_23296,N_13770,N_14284);
nand U23297 (N_23297,N_14896,N_16508);
and U23298 (N_23298,N_17420,N_13558);
or U23299 (N_23299,N_15742,N_13489);
nand U23300 (N_23300,N_13054,N_17369);
or U23301 (N_23301,N_16063,N_14219);
nand U23302 (N_23302,N_17679,N_14422);
nand U23303 (N_23303,N_17606,N_12190);
xor U23304 (N_23304,N_12957,N_17142);
nand U23305 (N_23305,N_17027,N_13349);
nand U23306 (N_23306,N_13635,N_13667);
or U23307 (N_23307,N_15866,N_16190);
nor U23308 (N_23308,N_14193,N_17283);
nand U23309 (N_23309,N_12764,N_13593);
or U23310 (N_23310,N_14228,N_15419);
and U23311 (N_23311,N_13060,N_14061);
and U23312 (N_23312,N_13744,N_15478);
and U23313 (N_23313,N_15902,N_15035);
nor U23314 (N_23314,N_14755,N_15799);
and U23315 (N_23315,N_14766,N_14995);
xor U23316 (N_23316,N_12782,N_17091);
xor U23317 (N_23317,N_13163,N_17695);
xor U23318 (N_23318,N_17877,N_16296);
or U23319 (N_23319,N_14579,N_14710);
nor U23320 (N_23320,N_17575,N_17045);
or U23321 (N_23321,N_14953,N_14610);
nor U23322 (N_23322,N_16752,N_12257);
nor U23323 (N_23323,N_15406,N_13592);
and U23324 (N_23324,N_14239,N_16465);
and U23325 (N_23325,N_14727,N_16883);
or U23326 (N_23326,N_14650,N_17312);
or U23327 (N_23327,N_16924,N_16305);
nand U23328 (N_23328,N_13640,N_12199);
or U23329 (N_23329,N_14781,N_13829);
xor U23330 (N_23330,N_16480,N_17902);
and U23331 (N_23331,N_17537,N_14536);
nand U23332 (N_23332,N_12397,N_14562);
nor U23333 (N_23333,N_15172,N_16960);
nand U23334 (N_23334,N_12555,N_12492);
xor U23335 (N_23335,N_13578,N_14769);
nor U23336 (N_23336,N_15496,N_17506);
nand U23337 (N_23337,N_14227,N_16647);
nor U23338 (N_23338,N_17779,N_15618);
xnor U23339 (N_23339,N_14090,N_14022);
and U23340 (N_23340,N_16280,N_16300);
or U23341 (N_23341,N_15621,N_14142);
xnor U23342 (N_23342,N_15036,N_15505);
and U23343 (N_23343,N_17832,N_17049);
and U23344 (N_23344,N_13310,N_12644);
and U23345 (N_23345,N_12224,N_14613);
or U23346 (N_23346,N_17027,N_12489);
nand U23347 (N_23347,N_15324,N_17705);
or U23348 (N_23348,N_13554,N_17055);
xor U23349 (N_23349,N_15376,N_16966);
or U23350 (N_23350,N_17313,N_13204);
nand U23351 (N_23351,N_12754,N_15017);
xor U23352 (N_23352,N_16416,N_15347);
and U23353 (N_23353,N_15826,N_15246);
xnor U23354 (N_23354,N_12407,N_12782);
xnor U23355 (N_23355,N_17822,N_12865);
and U23356 (N_23356,N_14243,N_15594);
nor U23357 (N_23357,N_14236,N_14986);
or U23358 (N_23358,N_16006,N_12879);
nand U23359 (N_23359,N_13611,N_16404);
or U23360 (N_23360,N_17732,N_14149);
and U23361 (N_23361,N_17537,N_17425);
xor U23362 (N_23362,N_16558,N_15300);
xor U23363 (N_23363,N_13146,N_12686);
and U23364 (N_23364,N_15630,N_13098);
and U23365 (N_23365,N_13507,N_16032);
or U23366 (N_23366,N_17483,N_16257);
xor U23367 (N_23367,N_14176,N_12207);
nor U23368 (N_23368,N_12102,N_12538);
xor U23369 (N_23369,N_13451,N_17158);
nor U23370 (N_23370,N_16039,N_12340);
nor U23371 (N_23371,N_17520,N_14909);
or U23372 (N_23372,N_17789,N_13887);
and U23373 (N_23373,N_17167,N_16566);
and U23374 (N_23374,N_16016,N_14197);
and U23375 (N_23375,N_15002,N_17039);
nand U23376 (N_23376,N_12162,N_13610);
nor U23377 (N_23377,N_15045,N_16696);
and U23378 (N_23378,N_15430,N_12584);
xor U23379 (N_23379,N_15743,N_17890);
nor U23380 (N_23380,N_15862,N_12688);
xor U23381 (N_23381,N_14236,N_16425);
and U23382 (N_23382,N_15633,N_14924);
xnor U23383 (N_23383,N_13155,N_14785);
nand U23384 (N_23384,N_16187,N_14768);
and U23385 (N_23385,N_16841,N_12798);
or U23386 (N_23386,N_12967,N_14260);
nor U23387 (N_23387,N_13124,N_14057);
nor U23388 (N_23388,N_15667,N_12841);
and U23389 (N_23389,N_13605,N_15760);
nor U23390 (N_23390,N_12373,N_13289);
nand U23391 (N_23391,N_17899,N_13867);
and U23392 (N_23392,N_15739,N_12394);
xnor U23393 (N_23393,N_14036,N_15980);
nand U23394 (N_23394,N_15274,N_15038);
nor U23395 (N_23395,N_15193,N_13249);
nand U23396 (N_23396,N_13890,N_17119);
nand U23397 (N_23397,N_14348,N_17332);
nand U23398 (N_23398,N_13441,N_16870);
or U23399 (N_23399,N_15065,N_13372);
xor U23400 (N_23400,N_14934,N_16223);
xnor U23401 (N_23401,N_13458,N_12938);
xor U23402 (N_23402,N_14976,N_13017);
or U23403 (N_23403,N_14519,N_13358);
nand U23404 (N_23404,N_17097,N_17305);
and U23405 (N_23405,N_17421,N_12690);
nand U23406 (N_23406,N_15188,N_16163);
nand U23407 (N_23407,N_16867,N_13394);
and U23408 (N_23408,N_13680,N_17305);
and U23409 (N_23409,N_14908,N_16996);
nor U23410 (N_23410,N_13236,N_17730);
and U23411 (N_23411,N_15546,N_15993);
or U23412 (N_23412,N_16136,N_15203);
nor U23413 (N_23413,N_12195,N_13164);
and U23414 (N_23414,N_16302,N_13851);
xnor U23415 (N_23415,N_15290,N_13298);
xor U23416 (N_23416,N_17108,N_14859);
nor U23417 (N_23417,N_17386,N_15426);
nand U23418 (N_23418,N_15584,N_12711);
nor U23419 (N_23419,N_12244,N_12514);
xor U23420 (N_23420,N_13597,N_13733);
or U23421 (N_23421,N_15163,N_16447);
and U23422 (N_23422,N_14768,N_16623);
or U23423 (N_23423,N_14360,N_16158);
xnor U23424 (N_23424,N_12320,N_13250);
xor U23425 (N_23425,N_16073,N_17457);
or U23426 (N_23426,N_15250,N_14855);
and U23427 (N_23427,N_17810,N_15998);
nand U23428 (N_23428,N_17464,N_14758);
nand U23429 (N_23429,N_15752,N_13602);
or U23430 (N_23430,N_16440,N_12019);
nand U23431 (N_23431,N_17289,N_17356);
nor U23432 (N_23432,N_16245,N_16483);
or U23433 (N_23433,N_12340,N_17817);
nand U23434 (N_23434,N_13218,N_13559);
nor U23435 (N_23435,N_13595,N_16560);
nor U23436 (N_23436,N_16317,N_13270);
nor U23437 (N_23437,N_12287,N_14716);
xor U23438 (N_23438,N_16973,N_13044);
nand U23439 (N_23439,N_17413,N_14594);
or U23440 (N_23440,N_15131,N_14189);
nor U23441 (N_23441,N_15468,N_13177);
nor U23442 (N_23442,N_15763,N_15167);
or U23443 (N_23443,N_13081,N_14646);
and U23444 (N_23444,N_12595,N_12387);
xnor U23445 (N_23445,N_15104,N_17518);
nand U23446 (N_23446,N_17445,N_15955);
nand U23447 (N_23447,N_14574,N_12284);
and U23448 (N_23448,N_15739,N_15198);
nor U23449 (N_23449,N_17601,N_12906);
and U23450 (N_23450,N_14420,N_17158);
nand U23451 (N_23451,N_16814,N_17833);
or U23452 (N_23452,N_14122,N_13390);
or U23453 (N_23453,N_17134,N_17210);
or U23454 (N_23454,N_15990,N_13358);
nand U23455 (N_23455,N_13016,N_12908);
xnor U23456 (N_23456,N_17437,N_14521);
or U23457 (N_23457,N_17053,N_17947);
nand U23458 (N_23458,N_13245,N_13485);
nor U23459 (N_23459,N_14624,N_13406);
or U23460 (N_23460,N_12151,N_16059);
nand U23461 (N_23461,N_14155,N_13027);
and U23462 (N_23462,N_16996,N_17527);
and U23463 (N_23463,N_12602,N_15220);
nand U23464 (N_23464,N_12164,N_12333);
nor U23465 (N_23465,N_17802,N_13973);
nand U23466 (N_23466,N_14290,N_14771);
nand U23467 (N_23467,N_14651,N_15279);
and U23468 (N_23468,N_17049,N_14531);
and U23469 (N_23469,N_15900,N_14890);
nand U23470 (N_23470,N_12974,N_14022);
or U23471 (N_23471,N_15262,N_12744);
or U23472 (N_23472,N_14752,N_15675);
nand U23473 (N_23473,N_14797,N_17916);
xor U23474 (N_23474,N_13696,N_17020);
and U23475 (N_23475,N_16626,N_15971);
nand U23476 (N_23476,N_14640,N_16984);
nand U23477 (N_23477,N_13110,N_16835);
and U23478 (N_23478,N_14984,N_12082);
and U23479 (N_23479,N_17983,N_15768);
nand U23480 (N_23480,N_14591,N_16256);
nand U23481 (N_23481,N_16884,N_16748);
and U23482 (N_23482,N_13870,N_16836);
and U23483 (N_23483,N_14072,N_13287);
nand U23484 (N_23484,N_13668,N_14087);
nand U23485 (N_23485,N_16305,N_14800);
nor U23486 (N_23486,N_12805,N_15144);
and U23487 (N_23487,N_12449,N_15008);
nor U23488 (N_23488,N_13248,N_15854);
nor U23489 (N_23489,N_13806,N_12918);
nor U23490 (N_23490,N_17751,N_14899);
and U23491 (N_23491,N_16806,N_16314);
and U23492 (N_23492,N_13124,N_13756);
and U23493 (N_23493,N_17081,N_12295);
xnor U23494 (N_23494,N_12218,N_12509);
nor U23495 (N_23495,N_17746,N_17388);
nand U23496 (N_23496,N_13186,N_13334);
or U23497 (N_23497,N_12475,N_12979);
nor U23498 (N_23498,N_12323,N_16529);
or U23499 (N_23499,N_17575,N_16318);
xnor U23500 (N_23500,N_17798,N_15876);
and U23501 (N_23501,N_14486,N_13959);
xnor U23502 (N_23502,N_14924,N_17049);
and U23503 (N_23503,N_17720,N_17300);
and U23504 (N_23504,N_13633,N_13467);
nand U23505 (N_23505,N_13333,N_14794);
nand U23506 (N_23506,N_12759,N_14440);
or U23507 (N_23507,N_13801,N_12352);
and U23508 (N_23508,N_17447,N_17167);
nand U23509 (N_23509,N_17461,N_15850);
nor U23510 (N_23510,N_15198,N_13968);
or U23511 (N_23511,N_12707,N_12053);
nand U23512 (N_23512,N_16754,N_17833);
and U23513 (N_23513,N_16499,N_15981);
xor U23514 (N_23514,N_17189,N_14684);
nand U23515 (N_23515,N_13445,N_12110);
or U23516 (N_23516,N_14026,N_13096);
xnor U23517 (N_23517,N_16998,N_15292);
or U23518 (N_23518,N_17980,N_15187);
nor U23519 (N_23519,N_15520,N_14358);
nor U23520 (N_23520,N_17072,N_12594);
or U23521 (N_23521,N_15842,N_17048);
xnor U23522 (N_23522,N_17908,N_17035);
or U23523 (N_23523,N_17489,N_13594);
nand U23524 (N_23524,N_15247,N_16320);
nor U23525 (N_23525,N_17334,N_16220);
xor U23526 (N_23526,N_14290,N_14835);
xnor U23527 (N_23527,N_13960,N_17401);
or U23528 (N_23528,N_14576,N_16791);
xor U23529 (N_23529,N_14884,N_14883);
xnor U23530 (N_23530,N_17477,N_16893);
and U23531 (N_23531,N_12775,N_13361);
nand U23532 (N_23532,N_15182,N_17740);
xnor U23533 (N_23533,N_16840,N_16412);
nand U23534 (N_23534,N_14700,N_15198);
and U23535 (N_23535,N_14711,N_15398);
xnor U23536 (N_23536,N_16360,N_12368);
and U23537 (N_23537,N_14724,N_17050);
or U23538 (N_23538,N_12215,N_17796);
and U23539 (N_23539,N_15887,N_12871);
nor U23540 (N_23540,N_14316,N_12005);
or U23541 (N_23541,N_17484,N_13374);
or U23542 (N_23542,N_16155,N_17604);
or U23543 (N_23543,N_12200,N_14343);
and U23544 (N_23544,N_13361,N_15014);
nand U23545 (N_23545,N_17193,N_17254);
nor U23546 (N_23546,N_16267,N_13720);
nor U23547 (N_23547,N_12487,N_16185);
xor U23548 (N_23548,N_12933,N_15873);
nand U23549 (N_23549,N_13767,N_14678);
nand U23550 (N_23550,N_14391,N_17028);
nor U23551 (N_23551,N_16726,N_12234);
or U23552 (N_23552,N_16855,N_17646);
nand U23553 (N_23553,N_14305,N_15950);
xor U23554 (N_23554,N_16604,N_16584);
or U23555 (N_23555,N_13871,N_12666);
nand U23556 (N_23556,N_15990,N_12330);
nand U23557 (N_23557,N_13341,N_17509);
or U23558 (N_23558,N_15822,N_17328);
or U23559 (N_23559,N_14993,N_14158);
nor U23560 (N_23560,N_14725,N_17892);
and U23561 (N_23561,N_14732,N_14124);
nand U23562 (N_23562,N_12116,N_15881);
nor U23563 (N_23563,N_17105,N_13593);
nand U23564 (N_23564,N_16507,N_13758);
nand U23565 (N_23565,N_16576,N_16344);
nor U23566 (N_23566,N_14277,N_15880);
nand U23567 (N_23567,N_13050,N_16919);
nor U23568 (N_23568,N_17815,N_16752);
nand U23569 (N_23569,N_12783,N_13768);
xnor U23570 (N_23570,N_15536,N_12538);
or U23571 (N_23571,N_12733,N_14379);
and U23572 (N_23572,N_13236,N_15235);
and U23573 (N_23573,N_13931,N_16570);
or U23574 (N_23574,N_16320,N_12037);
and U23575 (N_23575,N_16210,N_13507);
and U23576 (N_23576,N_14496,N_12033);
nand U23577 (N_23577,N_17904,N_13458);
xnor U23578 (N_23578,N_12375,N_15903);
or U23579 (N_23579,N_13566,N_17060);
xnor U23580 (N_23580,N_17195,N_12621);
nand U23581 (N_23581,N_15493,N_14905);
and U23582 (N_23582,N_12603,N_17976);
nand U23583 (N_23583,N_13920,N_17313);
nand U23584 (N_23584,N_17842,N_13253);
nor U23585 (N_23585,N_15581,N_14101);
nand U23586 (N_23586,N_14637,N_14045);
nand U23587 (N_23587,N_13985,N_15602);
xor U23588 (N_23588,N_17042,N_12975);
xor U23589 (N_23589,N_13977,N_13006);
nand U23590 (N_23590,N_16710,N_13626);
xnor U23591 (N_23591,N_16230,N_15527);
and U23592 (N_23592,N_12199,N_16926);
nand U23593 (N_23593,N_13733,N_13388);
or U23594 (N_23594,N_14109,N_13894);
and U23595 (N_23595,N_14935,N_17084);
and U23596 (N_23596,N_12047,N_17026);
or U23597 (N_23597,N_16854,N_14437);
or U23598 (N_23598,N_16018,N_17133);
nor U23599 (N_23599,N_12878,N_14092);
nor U23600 (N_23600,N_13834,N_12744);
or U23601 (N_23601,N_13527,N_12758);
nand U23602 (N_23602,N_14449,N_13515);
and U23603 (N_23603,N_16083,N_14683);
xor U23604 (N_23604,N_12200,N_13525);
or U23605 (N_23605,N_15499,N_12655);
nand U23606 (N_23606,N_15288,N_17904);
nand U23607 (N_23607,N_16064,N_12845);
or U23608 (N_23608,N_14539,N_15161);
and U23609 (N_23609,N_12139,N_12355);
or U23610 (N_23610,N_14076,N_13875);
xnor U23611 (N_23611,N_12731,N_16890);
or U23612 (N_23612,N_12521,N_15341);
nor U23613 (N_23613,N_14810,N_17610);
xnor U23614 (N_23614,N_17907,N_17390);
or U23615 (N_23615,N_16261,N_12879);
nor U23616 (N_23616,N_15142,N_14258);
or U23617 (N_23617,N_12585,N_12959);
and U23618 (N_23618,N_17025,N_16861);
or U23619 (N_23619,N_17796,N_12196);
and U23620 (N_23620,N_16677,N_17537);
nor U23621 (N_23621,N_13587,N_17901);
or U23622 (N_23622,N_17085,N_13382);
nor U23623 (N_23623,N_12216,N_12222);
or U23624 (N_23624,N_16075,N_14030);
xor U23625 (N_23625,N_13307,N_16045);
nor U23626 (N_23626,N_17321,N_17638);
nor U23627 (N_23627,N_17394,N_13106);
nor U23628 (N_23628,N_15584,N_17564);
xor U23629 (N_23629,N_17553,N_13824);
xor U23630 (N_23630,N_14179,N_16796);
or U23631 (N_23631,N_12967,N_17789);
or U23632 (N_23632,N_16816,N_12582);
and U23633 (N_23633,N_13069,N_16705);
nand U23634 (N_23634,N_12912,N_12815);
and U23635 (N_23635,N_12771,N_16495);
and U23636 (N_23636,N_12921,N_16684);
nor U23637 (N_23637,N_15989,N_17132);
nand U23638 (N_23638,N_17026,N_13357);
nand U23639 (N_23639,N_16183,N_17540);
nor U23640 (N_23640,N_16629,N_13100);
or U23641 (N_23641,N_17081,N_13733);
xnor U23642 (N_23642,N_16083,N_17834);
xor U23643 (N_23643,N_12134,N_14396);
xor U23644 (N_23644,N_16866,N_17750);
or U23645 (N_23645,N_13598,N_16624);
nor U23646 (N_23646,N_15182,N_17508);
and U23647 (N_23647,N_15814,N_13262);
and U23648 (N_23648,N_13822,N_13451);
or U23649 (N_23649,N_12380,N_14816);
nand U23650 (N_23650,N_17349,N_14858);
or U23651 (N_23651,N_13295,N_17536);
or U23652 (N_23652,N_17582,N_17512);
xor U23653 (N_23653,N_16495,N_16438);
xnor U23654 (N_23654,N_17523,N_12131);
nor U23655 (N_23655,N_15509,N_13110);
and U23656 (N_23656,N_16908,N_17014);
nand U23657 (N_23657,N_15931,N_12685);
xor U23658 (N_23658,N_16334,N_12138);
or U23659 (N_23659,N_15183,N_14736);
xor U23660 (N_23660,N_17805,N_12688);
and U23661 (N_23661,N_13939,N_17817);
xor U23662 (N_23662,N_14339,N_16317);
or U23663 (N_23663,N_14468,N_12110);
xnor U23664 (N_23664,N_14931,N_15923);
nor U23665 (N_23665,N_12384,N_12095);
nor U23666 (N_23666,N_17741,N_17302);
and U23667 (N_23667,N_16418,N_14006);
xnor U23668 (N_23668,N_13537,N_15227);
nor U23669 (N_23669,N_15532,N_15572);
and U23670 (N_23670,N_17440,N_15419);
xor U23671 (N_23671,N_14808,N_14692);
nor U23672 (N_23672,N_15682,N_15075);
and U23673 (N_23673,N_13122,N_15673);
nor U23674 (N_23674,N_13144,N_17330);
nor U23675 (N_23675,N_13615,N_16028);
xnor U23676 (N_23676,N_13403,N_15757);
nand U23677 (N_23677,N_16801,N_13446);
and U23678 (N_23678,N_14772,N_16582);
or U23679 (N_23679,N_12059,N_14539);
and U23680 (N_23680,N_14395,N_12051);
and U23681 (N_23681,N_17220,N_14713);
xor U23682 (N_23682,N_12080,N_16459);
xnor U23683 (N_23683,N_16900,N_12363);
xor U23684 (N_23684,N_12154,N_13312);
nand U23685 (N_23685,N_15467,N_13834);
and U23686 (N_23686,N_12202,N_15465);
nor U23687 (N_23687,N_17000,N_12032);
nand U23688 (N_23688,N_14235,N_14016);
and U23689 (N_23689,N_14811,N_12412);
or U23690 (N_23690,N_17326,N_17426);
xor U23691 (N_23691,N_15644,N_15805);
nand U23692 (N_23692,N_12218,N_15096);
or U23693 (N_23693,N_14714,N_16672);
nand U23694 (N_23694,N_15512,N_15378);
xnor U23695 (N_23695,N_12650,N_14800);
nand U23696 (N_23696,N_14431,N_14638);
xor U23697 (N_23697,N_12236,N_16859);
or U23698 (N_23698,N_15015,N_16602);
nand U23699 (N_23699,N_16753,N_17878);
or U23700 (N_23700,N_16168,N_16206);
and U23701 (N_23701,N_12187,N_17562);
xor U23702 (N_23702,N_14222,N_16174);
and U23703 (N_23703,N_14873,N_17143);
nor U23704 (N_23704,N_12353,N_14056);
or U23705 (N_23705,N_15023,N_16478);
or U23706 (N_23706,N_15735,N_17353);
nand U23707 (N_23707,N_12647,N_15175);
xnor U23708 (N_23708,N_12157,N_16750);
nand U23709 (N_23709,N_13373,N_17549);
and U23710 (N_23710,N_15660,N_17952);
xor U23711 (N_23711,N_13556,N_17927);
nor U23712 (N_23712,N_15112,N_13131);
nand U23713 (N_23713,N_12812,N_13800);
xnor U23714 (N_23714,N_15026,N_13111);
or U23715 (N_23715,N_16570,N_14348);
xnor U23716 (N_23716,N_13362,N_17971);
nor U23717 (N_23717,N_17910,N_12204);
xor U23718 (N_23718,N_17301,N_13494);
or U23719 (N_23719,N_14682,N_16153);
xnor U23720 (N_23720,N_17285,N_17051);
nor U23721 (N_23721,N_12760,N_16288);
nand U23722 (N_23722,N_15414,N_15888);
xnor U23723 (N_23723,N_15410,N_14115);
or U23724 (N_23724,N_17824,N_14031);
or U23725 (N_23725,N_14767,N_12551);
and U23726 (N_23726,N_16402,N_16387);
xnor U23727 (N_23727,N_17469,N_14983);
nor U23728 (N_23728,N_15041,N_14294);
nand U23729 (N_23729,N_16123,N_12671);
and U23730 (N_23730,N_16385,N_16675);
xnor U23731 (N_23731,N_12729,N_12774);
xor U23732 (N_23732,N_12652,N_13565);
or U23733 (N_23733,N_15982,N_15761);
nor U23734 (N_23734,N_16996,N_14305);
and U23735 (N_23735,N_15693,N_17969);
xor U23736 (N_23736,N_17122,N_12005);
or U23737 (N_23737,N_15068,N_17803);
nand U23738 (N_23738,N_15586,N_15471);
or U23739 (N_23739,N_14565,N_12515);
nand U23740 (N_23740,N_17214,N_13182);
nor U23741 (N_23741,N_12275,N_17720);
nand U23742 (N_23742,N_14887,N_14584);
and U23743 (N_23743,N_12802,N_13067);
or U23744 (N_23744,N_15803,N_14526);
and U23745 (N_23745,N_17963,N_14306);
and U23746 (N_23746,N_16964,N_13362);
nor U23747 (N_23747,N_15373,N_13400);
nand U23748 (N_23748,N_16142,N_17993);
xor U23749 (N_23749,N_14623,N_17737);
or U23750 (N_23750,N_14917,N_16174);
xor U23751 (N_23751,N_14189,N_16057);
xnor U23752 (N_23752,N_17886,N_12809);
nor U23753 (N_23753,N_12824,N_13708);
xor U23754 (N_23754,N_14868,N_16526);
or U23755 (N_23755,N_12279,N_14556);
or U23756 (N_23756,N_16952,N_12510);
and U23757 (N_23757,N_13369,N_16914);
nand U23758 (N_23758,N_14253,N_12273);
nor U23759 (N_23759,N_17389,N_15029);
nor U23760 (N_23760,N_12461,N_12137);
or U23761 (N_23761,N_13262,N_12986);
nand U23762 (N_23762,N_13772,N_15950);
and U23763 (N_23763,N_12019,N_17152);
nand U23764 (N_23764,N_12184,N_14588);
or U23765 (N_23765,N_13303,N_16274);
or U23766 (N_23766,N_12133,N_16496);
and U23767 (N_23767,N_12245,N_12522);
and U23768 (N_23768,N_13637,N_17983);
nand U23769 (N_23769,N_13803,N_13450);
and U23770 (N_23770,N_16797,N_12243);
xnor U23771 (N_23771,N_15116,N_13048);
or U23772 (N_23772,N_15598,N_17907);
nor U23773 (N_23773,N_14766,N_13325);
xnor U23774 (N_23774,N_12434,N_12700);
or U23775 (N_23775,N_17861,N_15761);
and U23776 (N_23776,N_17929,N_12020);
nor U23777 (N_23777,N_16592,N_17941);
or U23778 (N_23778,N_12981,N_15872);
xnor U23779 (N_23779,N_14638,N_12098);
xor U23780 (N_23780,N_16900,N_16807);
or U23781 (N_23781,N_13562,N_15280);
xnor U23782 (N_23782,N_13349,N_16813);
nand U23783 (N_23783,N_16760,N_13192);
nor U23784 (N_23784,N_14123,N_16446);
nor U23785 (N_23785,N_12752,N_13918);
xnor U23786 (N_23786,N_15486,N_15323);
xor U23787 (N_23787,N_12502,N_16650);
nand U23788 (N_23788,N_15070,N_15542);
or U23789 (N_23789,N_13651,N_16205);
nand U23790 (N_23790,N_16899,N_14479);
and U23791 (N_23791,N_14418,N_17046);
or U23792 (N_23792,N_17570,N_16748);
and U23793 (N_23793,N_15336,N_17549);
and U23794 (N_23794,N_12946,N_12711);
and U23795 (N_23795,N_13072,N_12476);
xor U23796 (N_23796,N_12191,N_15657);
nand U23797 (N_23797,N_13269,N_15421);
or U23798 (N_23798,N_16010,N_16100);
nand U23799 (N_23799,N_14762,N_13056);
or U23800 (N_23800,N_16694,N_15593);
nor U23801 (N_23801,N_14702,N_12723);
and U23802 (N_23802,N_14884,N_13008);
nand U23803 (N_23803,N_12126,N_17383);
nor U23804 (N_23804,N_12356,N_12166);
nor U23805 (N_23805,N_16173,N_17497);
xor U23806 (N_23806,N_16863,N_13204);
xnor U23807 (N_23807,N_15263,N_12312);
nand U23808 (N_23808,N_12816,N_17260);
nor U23809 (N_23809,N_12974,N_16993);
nor U23810 (N_23810,N_16489,N_15202);
or U23811 (N_23811,N_16897,N_15392);
xnor U23812 (N_23812,N_17604,N_17652);
and U23813 (N_23813,N_13946,N_14181);
nand U23814 (N_23814,N_14238,N_15844);
and U23815 (N_23815,N_12915,N_17708);
and U23816 (N_23816,N_16948,N_15590);
or U23817 (N_23817,N_14919,N_15001);
or U23818 (N_23818,N_13850,N_16288);
nor U23819 (N_23819,N_16874,N_17472);
xor U23820 (N_23820,N_15351,N_14899);
nand U23821 (N_23821,N_13076,N_16150);
xor U23822 (N_23822,N_13954,N_17312);
nor U23823 (N_23823,N_13852,N_16463);
nand U23824 (N_23824,N_12302,N_14921);
or U23825 (N_23825,N_16115,N_14950);
nand U23826 (N_23826,N_16422,N_17304);
nor U23827 (N_23827,N_16777,N_15148);
and U23828 (N_23828,N_12241,N_15432);
nand U23829 (N_23829,N_14381,N_12324);
xnor U23830 (N_23830,N_17689,N_15919);
nand U23831 (N_23831,N_17912,N_15193);
nand U23832 (N_23832,N_12069,N_13315);
or U23833 (N_23833,N_15285,N_17383);
or U23834 (N_23834,N_13476,N_17180);
and U23835 (N_23835,N_14493,N_13894);
or U23836 (N_23836,N_17653,N_17287);
nor U23837 (N_23837,N_16271,N_16519);
nor U23838 (N_23838,N_13607,N_15933);
or U23839 (N_23839,N_12143,N_16139);
nor U23840 (N_23840,N_15931,N_12174);
or U23841 (N_23841,N_17149,N_17827);
or U23842 (N_23842,N_14826,N_14331);
nand U23843 (N_23843,N_16740,N_16403);
and U23844 (N_23844,N_15141,N_12332);
nand U23845 (N_23845,N_14670,N_16838);
and U23846 (N_23846,N_12065,N_17577);
xor U23847 (N_23847,N_17378,N_14343);
nand U23848 (N_23848,N_17660,N_16465);
nand U23849 (N_23849,N_12963,N_14711);
xnor U23850 (N_23850,N_16366,N_15687);
xnor U23851 (N_23851,N_12301,N_16614);
and U23852 (N_23852,N_12790,N_14101);
or U23853 (N_23853,N_17016,N_16348);
and U23854 (N_23854,N_17790,N_16454);
and U23855 (N_23855,N_14122,N_16673);
or U23856 (N_23856,N_17325,N_14638);
and U23857 (N_23857,N_15269,N_14263);
nor U23858 (N_23858,N_13806,N_16616);
nor U23859 (N_23859,N_14538,N_16474);
nand U23860 (N_23860,N_15161,N_12275);
xnor U23861 (N_23861,N_17025,N_14229);
nor U23862 (N_23862,N_16603,N_16277);
and U23863 (N_23863,N_13021,N_13544);
nor U23864 (N_23864,N_17403,N_13769);
nor U23865 (N_23865,N_14944,N_16746);
and U23866 (N_23866,N_13001,N_17028);
xor U23867 (N_23867,N_16657,N_12093);
and U23868 (N_23868,N_14915,N_14439);
or U23869 (N_23869,N_12171,N_15103);
nor U23870 (N_23870,N_17876,N_14480);
nand U23871 (N_23871,N_14471,N_13708);
or U23872 (N_23872,N_15115,N_14264);
and U23873 (N_23873,N_13515,N_17957);
xor U23874 (N_23874,N_16614,N_13561);
xor U23875 (N_23875,N_15676,N_15378);
xor U23876 (N_23876,N_16488,N_15201);
or U23877 (N_23877,N_17499,N_16353);
or U23878 (N_23878,N_16389,N_12070);
xnor U23879 (N_23879,N_13693,N_16436);
nor U23880 (N_23880,N_16908,N_15621);
nand U23881 (N_23881,N_16571,N_15834);
or U23882 (N_23882,N_14997,N_17170);
nor U23883 (N_23883,N_12654,N_15665);
nor U23884 (N_23884,N_15566,N_15854);
and U23885 (N_23885,N_15431,N_13056);
xor U23886 (N_23886,N_15326,N_16938);
nor U23887 (N_23887,N_17558,N_15212);
xor U23888 (N_23888,N_13480,N_16058);
nand U23889 (N_23889,N_17060,N_15489);
or U23890 (N_23890,N_17219,N_16094);
and U23891 (N_23891,N_12078,N_14157);
or U23892 (N_23892,N_14357,N_13419);
or U23893 (N_23893,N_15335,N_17068);
nor U23894 (N_23894,N_16709,N_15064);
nand U23895 (N_23895,N_12237,N_16177);
or U23896 (N_23896,N_16939,N_17018);
and U23897 (N_23897,N_12648,N_16864);
and U23898 (N_23898,N_16544,N_16220);
nor U23899 (N_23899,N_14558,N_15881);
nor U23900 (N_23900,N_16141,N_15996);
and U23901 (N_23901,N_16738,N_14345);
nor U23902 (N_23902,N_14225,N_13233);
nor U23903 (N_23903,N_13507,N_15468);
or U23904 (N_23904,N_12913,N_14785);
and U23905 (N_23905,N_17406,N_12485);
or U23906 (N_23906,N_12599,N_17092);
and U23907 (N_23907,N_13386,N_12500);
nand U23908 (N_23908,N_12265,N_17892);
nor U23909 (N_23909,N_15051,N_13509);
nand U23910 (N_23910,N_12354,N_17872);
nor U23911 (N_23911,N_12920,N_16639);
nor U23912 (N_23912,N_13503,N_16404);
and U23913 (N_23913,N_14665,N_15399);
and U23914 (N_23914,N_15196,N_14843);
xor U23915 (N_23915,N_16325,N_14138);
or U23916 (N_23916,N_12718,N_12109);
or U23917 (N_23917,N_16883,N_12198);
xor U23918 (N_23918,N_17612,N_17456);
nor U23919 (N_23919,N_13145,N_16051);
nand U23920 (N_23920,N_15998,N_14393);
xor U23921 (N_23921,N_12599,N_16486);
and U23922 (N_23922,N_12739,N_16487);
and U23923 (N_23923,N_13253,N_14549);
nand U23924 (N_23924,N_15092,N_17595);
and U23925 (N_23925,N_13196,N_15791);
nor U23926 (N_23926,N_12471,N_12748);
and U23927 (N_23927,N_14980,N_17407);
or U23928 (N_23928,N_16947,N_16259);
nor U23929 (N_23929,N_14491,N_17329);
and U23930 (N_23930,N_14047,N_14696);
nor U23931 (N_23931,N_15908,N_12765);
and U23932 (N_23932,N_16217,N_16399);
and U23933 (N_23933,N_16591,N_15551);
xor U23934 (N_23934,N_16666,N_16432);
nor U23935 (N_23935,N_16273,N_17080);
nand U23936 (N_23936,N_13080,N_14082);
xor U23937 (N_23937,N_15596,N_14433);
nor U23938 (N_23938,N_16231,N_16008);
or U23939 (N_23939,N_17056,N_14290);
nand U23940 (N_23940,N_14762,N_12499);
or U23941 (N_23941,N_17389,N_15917);
nand U23942 (N_23942,N_16432,N_13996);
xor U23943 (N_23943,N_12063,N_15287);
nand U23944 (N_23944,N_12615,N_17620);
and U23945 (N_23945,N_17166,N_16589);
nor U23946 (N_23946,N_17660,N_15765);
or U23947 (N_23947,N_17432,N_15275);
nand U23948 (N_23948,N_16534,N_13266);
nand U23949 (N_23949,N_12151,N_17540);
and U23950 (N_23950,N_12873,N_12675);
nor U23951 (N_23951,N_14393,N_17138);
nor U23952 (N_23952,N_12401,N_15416);
nand U23953 (N_23953,N_15042,N_17717);
or U23954 (N_23954,N_13355,N_15414);
nand U23955 (N_23955,N_15071,N_16568);
or U23956 (N_23956,N_13146,N_12059);
and U23957 (N_23957,N_17827,N_16484);
xor U23958 (N_23958,N_12941,N_12115);
nor U23959 (N_23959,N_14405,N_13030);
and U23960 (N_23960,N_17086,N_17392);
and U23961 (N_23961,N_17525,N_15187);
nand U23962 (N_23962,N_13016,N_16345);
nor U23963 (N_23963,N_17792,N_15435);
or U23964 (N_23964,N_16935,N_17481);
nand U23965 (N_23965,N_12730,N_14060);
or U23966 (N_23966,N_16092,N_12053);
xor U23967 (N_23967,N_16155,N_17801);
nor U23968 (N_23968,N_13085,N_13735);
nand U23969 (N_23969,N_12332,N_13231);
nand U23970 (N_23970,N_16788,N_17208);
nand U23971 (N_23971,N_12770,N_12132);
nand U23972 (N_23972,N_17749,N_13738);
and U23973 (N_23973,N_15893,N_17904);
xor U23974 (N_23974,N_15000,N_12124);
nand U23975 (N_23975,N_14740,N_14971);
xnor U23976 (N_23976,N_12312,N_14082);
nand U23977 (N_23977,N_12213,N_14785);
nand U23978 (N_23978,N_15840,N_17049);
or U23979 (N_23979,N_12034,N_14480);
xor U23980 (N_23980,N_12245,N_17619);
or U23981 (N_23981,N_16910,N_13683);
nor U23982 (N_23982,N_13420,N_12664);
nor U23983 (N_23983,N_15146,N_14298);
xnor U23984 (N_23984,N_13024,N_15246);
nand U23985 (N_23985,N_15676,N_12692);
xnor U23986 (N_23986,N_17571,N_14554);
or U23987 (N_23987,N_15837,N_13778);
xor U23988 (N_23988,N_16607,N_13025);
and U23989 (N_23989,N_16482,N_16071);
and U23990 (N_23990,N_13298,N_17812);
nor U23991 (N_23991,N_14069,N_15422);
xnor U23992 (N_23992,N_14080,N_17059);
nand U23993 (N_23993,N_16025,N_13844);
nand U23994 (N_23994,N_14327,N_14975);
or U23995 (N_23995,N_14281,N_14438);
nor U23996 (N_23996,N_15228,N_17231);
xnor U23997 (N_23997,N_13273,N_13651);
or U23998 (N_23998,N_14570,N_15549);
xor U23999 (N_23999,N_13579,N_15640);
or U24000 (N_24000,N_22350,N_19826);
nand U24001 (N_24001,N_19930,N_23222);
xnor U24002 (N_24002,N_20433,N_22346);
nor U24003 (N_24003,N_19424,N_22620);
nor U24004 (N_24004,N_19965,N_18279);
or U24005 (N_24005,N_20424,N_20191);
or U24006 (N_24006,N_18717,N_22038);
nor U24007 (N_24007,N_22923,N_20374);
or U24008 (N_24008,N_18673,N_21746);
and U24009 (N_24009,N_21541,N_20089);
and U24010 (N_24010,N_20227,N_19455);
xnor U24011 (N_24011,N_19548,N_18839);
nand U24012 (N_24012,N_23463,N_23601);
and U24013 (N_24013,N_23701,N_19083);
nand U24014 (N_24014,N_20345,N_20228);
nor U24015 (N_24015,N_20949,N_20455);
xnor U24016 (N_24016,N_22883,N_22843);
and U24017 (N_24017,N_22353,N_20229);
nand U24018 (N_24018,N_18502,N_22608);
nor U24019 (N_24019,N_19315,N_20784);
nand U24020 (N_24020,N_18406,N_19243);
nor U24021 (N_24021,N_22800,N_19231);
and U24022 (N_24022,N_19665,N_22977);
or U24023 (N_24023,N_20823,N_21635);
nand U24024 (N_24024,N_23148,N_21190);
or U24025 (N_24025,N_23248,N_20250);
or U24026 (N_24026,N_22590,N_18667);
and U24027 (N_24027,N_23696,N_20377);
nor U24028 (N_24028,N_22441,N_23312);
and U24029 (N_24029,N_21744,N_23615);
or U24030 (N_24030,N_18982,N_20830);
and U24031 (N_24031,N_18598,N_21538);
nor U24032 (N_24032,N_23414,N_18904);
and U24033 (N_24033,N_19606,N_23585);
and U24034 (N_24034,N_22339,N_23996);
or U24035 (N_24035,N_23018,N_23054);
nor U24036 (N_24036,N_23849,N_20308);
xnor U24037 (N_24037,N_22670,N_20033);
nand U24038 (N_24038,N_18046,N_18226);
and U24039 (N_24039,N_21971,N_22762);
and U24040 (N_24040,N_18072,N_20491);
xnor U24041 (N_24041,N_20218,N_22139);
nor U24042 (N_24042,N_22133,N_21355);
xor U24043 (N_24043,N_23706,N_20103);
and U24044 (N_24044,N_18298,N_18810);
and U24045 (N_24045,N_21842,N_21693);
nand U24046 (N_24046,N_21872,N_21247);
xnor U24047 (N_24047,N_23198,N_20220);
and U24048 (N_24048,N_18217,N_18802);
nand U24049 (N_24049,N_22284,N_22950);
and U24050 (N_24050,N_18396,N_18293);
nor U24051 (N_24051,N_18332,N_22953);
and U24052 (N_24052,N_19452,N_21051);
xor U24053 (N_24053,N_19471,N_20596);
nand U24054 (N_24054,N_18702,N_22786);
or U24055 (N_24055,N_19076,N_22974);
xor U24056 (N_24056,N_22048,N_19065);
and U24057 (N_24057,N_20853,N_19582);
nor U24058 (N_24058,N_22372,N_22510);
or U24059 (N_24059,N_18537,N_19211);
nor U24060 (N_24060,N_19882,N_23032);
xnor U24061 (N_24061,N_22111,N_23741);
xnor U24062 (N_24062,N_22261,N_20872);
or U24063 (N_24063,N_21453,N_20663);
or U24064 (N_24064,N_23598,N_23058);
nand U24065 (N_24065,N_19331,N_21040);
nand U24066 (N_24066,N_23718,N_23142);
or U24067 (N_24067,N_20039,N_21486);
nand U24068 (N_24068,N_18196,N_20054);
nor U24069 (N_24069,N_18912,N_22965);
nor U24070 (N_24070,N_20956,N_18594);
xor U24071 (N_24071,N_22719,N_19189);
and U24072 (N_24072,N_19728,N_19380);
nor U24073 (N_24073,N_19150,N_22035);
xnor U24074 (N_24074,N_22092,N_18112);
nor U24075 (N_24075,N_20756,N_21509);
xor U24076 (N_24076,N_22918,N_20165);
xor U24077 (N_24077,N_22498,N_21447);
and U24078 (N_24078,N_23606,N_19744);
and U24079 (N_24079,N_19311,N_22702);
nand U24080 (N_24080,N_20193,N_19916);
nor U24081 (N_24081,N_23124,N_22234);
nor U24082 (N_24082,N_19546,N_20800);
xnor U24083 (N_24083,N_18587,N_19614);
xnor U24084 (N_24084,N_21895,N_18765);
nor U24085 (N_24085,N_20870,N_19403);
xor U24086 (N_24086,N_22336,N_22575);
and U24087 (N_24087,N_18808,N_23812);
or U24088 (N_24088,N_19601,N_22129);
nor U24089 (N_24089,N_20877,N_20267);
or U24090 (N_24090,N_22070,N_20141);
and U24091 (N_24091,N_23294,N_19658);
or U24092 (N_24092,N_22016,N_22387);
xor U24093 (N_24093,N_20164,N_23587);
nor U24094 (N_24094,N_21537,N_20609);
or U24095 (N_24095,N_23302,N_21898);
xnor U24096 (N_24096,N_22089,N_20897);
or U24097 (N_24097,N_19472,N_20898);
xnor U24098 (N_24098,N_19956,N_21417);
xnor U24099 (N_24099,N_22807,N_18955);
nor U24100 (N_24100,N_22173,N_18249);
and U24101 (N_24101,N_19038,N_23260);
nor U24102 (N_24102,N_20874,N_23013);
or U24103 (N_24103,N_18187,N_19643);
or U24104 (N_24104,N_18116,N_21512);
and U24105 (N_24105,N_18843,N_21863);
and U24106 (N_24106,N_20614,N_18304);
xor U24107 (N_24107,N_21268,N_19531);
nor U24108 (N_24108,N_18377,N_23899);
or U24109 (N_24109,N_21146,N_20966);
or U24110 (N_24110,N_18254,N_18054);
nand U24111 (N_24111,N_23494,N_19099);
or U24112 (N_24112,N_22793,N_19904);
nor U24113 (N_24113,N_23255,N_20010);
nor U24114 (N_24114,N_18427,N_21603);
nor U24115 (N_24115,N_21937,N_20703);
xnor U24116 (N_24116,N_19763,N_18022);
and U24117 (N_24117,N_21779,N_21936);
and U24118 (N_24118,N_19864,N_19048);
and U24119 (N_24119,N_21911,N_20389);
nor U24120 (N_24120,N_20632,N_18593);
nand U24121 (N_24121,N_21217,N_18443);
xnor U24122 (N_24122,N_18696,N_20025);
and U24123 (N_24123,N_19079,N_20590);
nor U24124 (N_24124,N_20537,N_21564);
or U24125 (N_24125,N_23462,N_19990);
or U24126 (N_24126,N_22056,N_21934);
and U24127 (N_24127,N_23523,N_21701);
and U24128 (N_24128,N_21695,N_22219);
and U24129 (N_24129,N_18891,N_23898);
nor U24130 (N_24130,N_19256,N_19874);
xor U24131 (N_24131,N_19397,N_21715);
xnor U24132 (N_24132,N_22979,N_19418);
or U24133 (N_24133,N_19732,N_23945);
nand U24134 (N_24134,N_19829,N_23189);
nor U24135 (N_24135,N_18846,N_18523);
nand U24136 (N_24136,N_23573,N_19407);
or U24137 (N_24137,N_19707,N_19723);
nand U24138 (N_24138,N_18071,N_22235);
and U24139 (N_24139,N_21712,N_18481);
and U24140 (N_24140,N_21350,N_23197);
nand U24141 (N_24141,N_23663,N_21605);
or U24142 (N_24142,N_21063,N_18970);
or U24143 (N_24143,N_20148,N_19610);
nor U24144 (N_24144,N_20113,N_18687);
nand U24145 (N_24145,N_19368,N_21200);
xor U24146 (N_24146,N_23345,N_21590);
and U24147 (N_24147,N_21554,N_21865);
nand U24148 (N_24148,N_23402,N_18633);
nand U24149 (N_24149,N_20684,N_22078);
and U24150 (N_24150,N_23081,N_19290);
or U24151 (N_24151,N_22712,N_19837);
nor U24152 (N_24152,N_19174,N_21749);
and U24153 (N_24153,N_21826,N_23524);
nor U24154 (N_24154,N_23332,N_20402);
nand U24155 (N_24155,N_23121,N_23817);
and U24156 (N_24156,N_23661,N_18625);
nor U24157 (N_24157,N_22975,N_23906);
nand U24158 (N_24158,N_18563,N_23333);
xnor U24159 (N_24159,N_20231,N_22424);
nor U24160 (N_24160,N_20293,N_18206);
and U24161 (N_24161,N_18322,N_22373);
nand U24162 (N_24162,N_23570,N_23888);
or U24163 (N_24163,N_21873,N_18829);
nand U24164 (N_24164,N_20114,N_23976);
xnor U24165 (N_24165,N_23891,N_20503);
xnor U24166 (N_24166,N_20379,N_21242);
nand U24167 (N_24167,N_19487,N_21333);
and U24168 (N_24168,N_21346,N_21961);
and U24169 (N_24169,N_19267,N_19664);
nand U24170 (N_24170,N_19266,N_20811);
xnor U24171 (N_24171,N_18620,N_18547);
and U24172 (N_24172,N_20728,N_20393);
nor U24173 (N_24173,N_18452,N_21751);
nor U24174 (N_24174,N_21392,N_22463);
and U24175 (N_24175,N_20436,N_18714);
nor U24176 (N_24176,N_18162,N_20734);
nor U24177 (N_24177,N_22401,N_21144);
or U24178 (N_24178,N_22468,N_22383);
nand U24179 (N_24179,N_21794,N_20787);
nand U24180 (N_24180,N_23111,N_19302);
nand U24181 (N_24181,N_20333,N_23386);
or U24182 (N_24182,N_18818,N_18422);
nand U24183 (N_24183,N_22976,N_23153);
nor U24184 (N_24184,N_20901,N_22370);
nand U24185 (N_24185,N_22748,N_21648);
xnor U24186 (N_24186,N_22897,N_20076);
or U24187 (N_24187,N_18734,N_23832);
or U24188 (N_24188,N_22506,N_18343);
xor U24189 (N_24189,N_21815,N_18880);
or U24190 (N_24190,N_19627,N_23383);
or U24191 (N_24191,N_19633,N_21490);
xnor U24192 (N_24192,N_22471,N_21958);
and U24193 (N_24193,N_21782,N_20629);
xnor U24194 (N_24194,N_22710,N_23559);
or U24195 (N_24195,N_20413,N_21406);
nor U24196 (N_24196,N_20349,N_23688);
xnor U24197 (N_24197,N_22808,N_19694);
nor U24198 (N_24198,N_21639,N_19815);
xnor U24199 (N_24199,N_21774,N_20244);
nor U24200 (N_24200,N_22836,N_22671);
and U24201 (N_24201,N_20156,N_23025);
xor U24202 (N_24202,N_19514,N_19856);
xnor U24203 (N_24203,N_21353,N_20647);
nand U24204 (N_24204,N_19045,N_19399);
and U24205 (N_24205,N_21152,N_18713);
or U24206 (N_24206,N_18921,N_20137);
and U24207 (N_24207,N_18960,N_18104);
xor U24208 (N_24208,N_18291,N_21092);
nand U24209 (N_24209,N_18312,N_20304);
nor U24210 (N_24210,N_22533,N_21641);
nor U24211 (N_24211,N_19604,N_22992);
nor U24212 (N_24212,N_21822,N_20236);
nand U24213 (N_24213,N_18643,N_22202);
nand U24214 (N_24214,N_20206,N_19912);
or U24215 (N_24215,N_21844,N_18954);
nand U24216 (N_24216,N_19207,N_19233);
or U24217 (N_24217,N_18488,N_23893);
or U24218 (N_24218,N_20051,N_23131);
xnor U24219 (N_24219,N_18240,N_22701);
nor U24220 (N_24220,N_20525,N_23648);
xor U24221 (N_24221,N_20275,N_23053);
nor U24222 (N_24222,N_19940,N_22698);
nand U24223 (N_24223,N_23940,N_22999);
nand U24224 (N_24224,N_22410,N_20181);
and U24225 (N_24225,N_22771,N_22004);
nand U24226 (N_24226,N_21606,N_22480);
or U24227 (N_24227,N_21470,N_19634);
and U24228 (N_24228,N_21656,N_20200);
nand U24229 (N_24229,N_21279,N_23036);
nor U24230 (N_24230,N_23526,N_22729);
nand U24231 (N_24231,N_19495,N_21983);
nand U24232 (N_24232,N_20741,N_21228);
nor U24233 (N_24233,N_18911,N_23129);
or U24234 (N_24234,N_22587,N_19730);
xor U24235 (N_24235,N_23242,N_21617);
nand U24236 (N_24236,N_21282,N_18819);
nor U24237 (N_24237,N_22032,N_18387);
xnor U24238 (N_24238,N_23012,N_23481);
nand U24239 (N_24239,N_22272,N_20465);
xor U24240 (N_24240,N_21404,N_18163);
nor U24241 (N_24241,N_21445,N_23501);
and U24242 (N_24242,N_20794,N_20023);
nand U24243 (N_24243,N_20183,N_20550);
xor U24244 (N_24244,N_19536,N_18480);
xnor U24245 (N_24245,N_18825,N_22830);
and U24246 (N_24246,N_18169,N_22983);
nor U24247 (N_24247,N_20685,N_20927);
and U24248 (N_24248,N_19624,N_18616);
nand U24249 (N_24249,N_18002,N_18340);
xnor U24250 (N_24250,N_18948,N_19237);
and U24251 (N_24251,N_18416,N_20972);
and U24252 (N_24252,N_20392,N_19800);
and U24253 (N_24253,N_19499,N_23361);
nor U24254 (N_24254,N_21377,N_18335);
xor U24255 (N_24255,N_22937,N_23617);
nor U24256 (N_24256,N_18521,N_22083);
xnor U24257 (N_24257,N_22451,N_23313);
nand U24258 (N_24258,N_18498,N_18417);
nand U24259 (N_24259,N_21189,N_22128);
xnor U24260 (N_24260,N_19966,N_19303);
and U24261 (N_24261,N_23925,N_22728);
nand U24262 (N_24262,N_18067,N_23871);
or U24263 (N_24263,N_20930,N_19794);
or U24264 (N_24264,N_21487,N_22638);
nor U24265 (N_24265,N_21364,N_18872);
or U24266 (N_24266,N_20239,N_18401);
nor U24267 (N_24267,N_23584,N_22639);
xor U24268 (N_24268,N_18010,N_22209);
and U24269 (N_24269,N_20401,N_18231);
xnor U24270 (N_24270,N_23212,N_21325);
or U24271 (N_24271,N_23014,N_21597);
nor U24272 (N_24272,N_19326,N_20878);
nor U24273 (N_24273,N_18868,N_22804);
nor U24274 (N_24274,N_20423,N_18986);
xnor U24275 (N_24275,N_20835,N_23581);
nand U24276 (N_24276,N_19192,N_18993);
and U24277 (N_24277,N_23243,N_18391);
or U24278 (N_24278,N_19889,N_20223);
nor U24279 (N_24279,N_18739,N_20235);
nor U24280 (N_24280,N_23542,N_22791);
and U24281 (N_24281,N_22177,N_22612);
nand U24282 (N_24282,N_21477,N_20667);
nor U24283 (N_24283,N_21742,N_23767);
or U24284 (N_24284,N_23985,N_22947);
nand U24285 (N_24285,N_19466,N_22732);
xor U24286 (N_24286,N_19792,N_20668);
nand U24287 (N_24287,N_23049,N_22672);
nor U24288 (N_24288,N_23346,N_18573);
and U24289 (N_24289,N_18100,N_22708);
and U24290 (N_24290,N_19492,N_23075);
and U24291 (N_24291,N_18357,N_21616);
xnor U24292 (N_24292,N_18870,N_21059);
or U24293 (N_24293,N_20605,N_23983);
and U24294 (N_24294,N_21438,N_18320);
nand U24295 (N_24295,N_23751,N_18113);
nor U24296 (N_24296,N_23842,N_18828);
xnor U24297 (N_24297,N_18177,N_19274);
or U24298 (N_24298,N_22279,N_23577);
and U24299 (N_24299,N_19892,N_20857);
nor U24300 (N_24300,N_20264,N_23534);
nand U24301 (N_24301,N_18830,N_21772);
nand U24302 (N_24302,N_22314,N_21967);
and U24303 (N_24303,N_21941,N_19067);
nand U24304 (N_24304,N_19494,N_21460);
nand U24305 (N_24305,N_20542,N_19638);
or U24306 (N_24306,N_18185,N_18565);
nor U24307 (N_24307,N_21518,N_20234);
or U24308 (N_24308,N_22570,N_21568);
nand U24309 (N_24309,N_20572,N_23461);
nand U24310 (N_24310,N_19578,N_22379);
xnor U24311 (N_24311,N_23182,N_20026);
nand U24312 (N_24312,N_19597,N_23196);
or U24313 (N_24313,N_18555,N_22674);
or U24314 (N_24314,N_22206,N_21985);
xnor U24315 (N_24315,N_20101,N_19814);
xnor U24316 (N_24316,N_20924,N_20505);
nor U24317 (N_24317,N_20160,N_22020);
xnor U24318 (N_24318,N_18289,N_18174);
or U24319 (N_24319,N_21516,N_22442);
or U24320 (N_24320,N_20636,N_21707);
and U24321 (N_24321,N_21968,N_22170);
xnor U24322 (N_24322,N_18740,N_22029);
nand U24323 (N_24323,N_23082,N_20692);
or U24324 (N_24324,N_22690,N_22594);
or U24325 (N_24325,N_21640,N_23820);
nor U24326 (N_24326,N_21116,N_21332);
and U24327 (N_24327,N_18030,N_19100);
xor U24328 (N_24328,N_19996,N_23761);
xor U24329 (N_24329,N_19628,N_20736);
xnor U24330 (N_24330,N_23062,N_23855);
nand U24331 (N_24331,N_19972,N_22742);
and U24332 (N_24332,N_21811,N_18194);
nand U24333 (N_24333,N_23132,N_20129);
or U24334 (N_24334,N_23856,N_23530);
xnor U24335 (N_24335,N_23726,N_20052);
or U24336 (N_24336,N_21959,N_21072);
nor U24337 (N_24337,N_18974,N_19570);
xnor U24338 (N_24338,N_21182,N_18500);
or U24339 (N_24339,N_23739,N_19078);
or U24340 (N_24340,N_19084,N_23913);
and U24341 (N_24341,N_18944,N_20077);
or U24342 (N_24342,N_18630,N_18156);
xor U24343 (N_24343,N_20404,N_19574);
nor U24344 (N_24344,N_21814,N_18769);
xor U24345 (N_24345,N_19000,N_22665);
or U24346 (N_24346,N_20182,N_23057);
nor U24347 (N_24347,N_20405,N_20788);
or U24348 (N_24348,N_20318,N_20289);
or U24349 (N_24349,N_19253,N_23933);
nand U24350 (N_24350,N_18223,N_23391);
and U24351 (N_24351,N_23728,N_20694);
nand U24352 (N_24352,N_22778,N_22260);
nor U24353 (N_24353,N_19733,N_22425);
xnor U24354 (N_24354,N_23550,N_23787);
and U24355 (N_24355,N_19064,N_19544);
nand U24356 (N_24356,N_21970,N_18068);
or U24357 (N_24357,N_21101,N_19722);
and U24358 (N_24358,N_23490,N_21244);
nand U24359 (N_24359,N_22103,N_20184);
nand U24360 (N_24360,N_22136,N_20305);
xnor U24361 (N_24361,N_22535,N_21266);
and U24362 (N_24362,N_21055,N_20963);
nand U24363 (N_24363,N_23865,N_22359);
xor U24364 (N_24364,N_23145,N_18398);
nand U24365 (N_24365,N_21046,N_22585);
or U24366 (N_24366,N_22752,N_20407);
nor U24367 (N_24367,N_19112,N_23935);
nor U24368 (N_24368,N_18404,N_23972);
and U24369 (N_24369,N_20579,N_23815);
nor U24370 (N_24370,N_20824,N_18455);
nor U24371 (N_24371,N_20288,N_23677);
and U24372 (N_24372,N_20152,N_18018);
nor U24373 (N_24373,N_23791,N_20842);
or U24374 (N_24374,N_23716,N_20613);
nor U24375 (N_24375,N_22600,N_20648);
xor U24376 (N_24376,N_23349,N_20669);
nor U24377 (N_24377,N_18679,N_20773);
nand U24378 (N_24378,N_19491,N_21168);
or U24379 (N_24379,N_23154,N_21206);
or U24380 (N_24380,N_19206,N_22096);
nand U24381 (N_24381,N_18977,N_19660);
and U24382 (N_24382,N_21699,N_23747);
nand U24383 (N_24383,N_20678,N_19028);
or U24384 (N_24384,N_18812,N_19925);
nand U24385 (N_24385,N_22114,N_23758);
xor U24386 (N_24386,N_20154,N_22358);
nand U24387 (N_24387,N_19545,N_18049);
nor U24388 (N_24388,N_20472,N_20130);
and U24389 (N_24389,N_21618,N_20739);
nor U24390 (N_24390,N_21314,N_18755);
or U24391 (N_24391,N_20202,N_20271);
or U24392 (N_24392,N_23381,N_20671);
nand U24393 (N_24393,N_19310,N_18757);
nor U24394 (N_24394,N_21737,N_21812);
nor U24395 (N_24395,N_23202,N_21381);
nor U24396 (N_24396,N_19104,N_18848);
and U24397 (N_24397,N_18577,N_19054);
nor U24398 (N_24398,N_22908,N_19567);
nand U24399 (N_24399,N_20693,N_23457);
or U24400 (N_24400,N_18450,N_21057);
or U24401 (N_24401,N_21419,N_20290);
nand U24402 (N_24402,N_20845,N_20742);
nand U24403 (N_24403,N_18631,N_21535);
nand U24404 (N_24404,N_21067,N_23309);
and U24405 (N_24405,N_19980,N_18753);
or U24406 (N_24406,N_23502,N_18351);
and U24407 (N_24407,N_22138,N_18815);
or U24408 (N_24408,N_20351,N_18635);
or U24409 (N_24409,N_23233,N_21604);
xnor U24410 (N_24410,N_20820,N_23884);
nor U24411 (N_24411,N_19154,N_18016);
xnor U24412 (N_24412,N_19566,N_21321);
nor U24413 (N_24413,N_20551,N_19823);
or U24414 (N_24414,N_20494,N_22958);
or U24415 (N_24415,N_22795,N_18436);
nor U24416 (N_24416,N_23643,N_23757);
nor U24417 (N_24417,N_23164,N_18778);
and U24418 (N_24418,N_20048,N_22715);
nand U24419 (N_24419,N_19724,N_20925);
xor U24420 (N_24420,N_19085,N_22924);
nor U24421 (N_24421,N_18090,N_19106);
and U24422 (N_24422,N_19603,N_22101);
xnor U24423 (N_24423,N_18583,N_20448);
nand U24424 (N_24424,N_18556,N_21017);
nor U24425 (N_24425,N_22325,N_22640);
nor U24426 (N_24426,N_23498,N_20122);
or U24427 (N_24427,N_19308,N_23277);
xnor U24428 (N_24428,N_18814,N_22935);
xnor U24429 (N_24429,N_20630,N_21308);
nor U24430 (N_24430,N_19595,N_23022);
or U24431 (N_24431,N_23136,N_21035);
nor U24432 (N_24432,N_19373,N_21855);
and U24433 (N_24433,N_18119,N_21389);
nand U24434 (N_24434,N_19299,N_21192);
nor U24435 (N_24435,N_18373,N_21164);
nand U24436 (N_24436,N_19214,N_19511);
nand U24437 (N_24437,N_21663,N_18285);
and U24438 (N_24438,N_21093,N_20687);
or U24439 (N_24439,N_19002,N_18472);
or U24440 (N_24440,N_23557,N_18560);
nand U24441 (N_24441,N_18303,N_19391);
nor U24442 (N_24442,N_19777,N_23672);
or U24443 (N_24443,N_23566,N_21837);
nand U24444 (N_24444,N_21205,N_19314);
nor U24445 (N_24445,N_22432,N_22654);
and U24446 (N_24446,N_22073,N_19618);
xor U24447 (N_24447,N_22302,N_18719);
or U24448 (N_24448,N_21047,N_18766);
xor U24449 (N_24449,N_21303,N_18761);
or U24450 (N_24450,N_22782,N_18632);
or U24451 (N_24451,N_18967,N_20778);
xnor U24452 (N_24452,N_22155,N_18255);
or U24453 (N_24453,N_19212,N_20726);
or U24454 (N_24454,N_22881,N_18987);
or U24455 (N_24455,N_22684,N_23063);
xnor U24456 (N_24456,N_19528,N_22152);
and U24457 (N_24457,N_19900,N_21162);
xnor U24458 (N_24458,N_18862,N_22236);
nand U24459 (N_24459,N_21584,N_20725);
nor U24460 (N_24460,N_20654,N_21692);
xor U24461 (N_24461,N_21033,N_18997);
xnor U24462 (N_24462,N_20135,N_22525);
or U24463 (N_24463,N_20056,N_22760);
nand U24464 (N_24464,N_23947,N_18898);
or U24465 (N_24465,N_19917,N_22928);
xor U24466 (N_24466,N_21547,N_21241);
nand U24467 (N_24467,N_23844,N_18805);
nor U24468 (N_24468,N_20681,N_22581);
and U24469 (N_24469,N_22559,N_22223);
or U24470 (N_24470,N_21140,N_22829);
xnor U24471 (N_24471,N_22806,N_21995);
nand U24472 (N_24472,N_19767,N_20798);
and U24473 (N_24473,N_20149,N_23268);
nor U24474 (N_24474,N_19802,N_21850);
nor U24475 (N_24475,N_23476,N_21220);
and U24476 (N_24476,N_23705,N_19841);
nand U24477 (N_24477,N_18209,N_22650);
nor U24478 (N_24478,N_18886,N_23816);
and U24479 (N_24479,N_23365,N_22704);
nand U24480 (N_24480,N_19370,N_20804);
and U24481 (N_24481,N_20695,N_21974);
xnor U24482 (N_24482,N_21529,N_20109);
or U24483 (N_24483,N_18659,N_22632);
or U24484 (N_24484,N_21876,N_21714);
or U24485 (N_24485,N_22488,N_20699);
and U24486 (N_24486,N_19766,N_20997);
nand U24487 (N_24487,N_21560,N_21919);
and U24488 (N_24488,N_22435,N_20485);
or U24489 (N_24489,N_20514,N_22695);
or U24490 (N_24490,N_21566,N_20059);
nand U24491 (N_24491,N_19442,N_20520);
xnor U24492 (N_24492,N_22440,N_20241);
and U24493 (N_24493,N_22427,N_23017);
xor U24494 (N_24494,N_18208,N_22856);
nor U24495 (N_24495,N_18053,N_21634);
or U24496 (N_24496,N_18055,N_22232);
or U24497 (N_24497,N_21860,N_19131);
nor U24498 (N_24498,N_22069,N_22902);
or U24499 (N_24499,N_19714,N_18813);
and U24500 (N_24500,N_23533,N_23266);
xnor U24501 (N_24501,N_19286,N_21711);
nor U24502 (N_24502,N_22319,N_23575);
and U24503 (N_24503,N_18961,N_21444);
or U24504 (N_24504,N_22085,N_20753);
xnor U24505 (N_24505,N_21925,N_18690);
nand U24506 (N_24506,N_20513,N_20529);
or U24507 (N_24507,N_23679,N_22356);
xor U24508 (N_24508,N_23097,N_19727);
or U24509 (N_24509,N_20545,N_21909);
nor U24510 (N_24510,N_18314,N_21412);
and U24511 (N_24511,N_20608,N_23669);
nand U24512 (N_24512,N_19451,N_19888);
or U24513 (N_24513,N_21363,N_19832);
or U24514 (N_24514,N_21233,N_21643);
and U24515 (N_24515,N_19523,N_19655);
nor U24516 (N_24516,N_22838,N_19143);
nor U24517 (N_24517,N_19877,N_21478);
nand U24518 (N_24518,N_21757,N_22515);
nand U24519 (N_24519,N_20245,N_23885);
nor U24520 (N_24520,N_21395,N_20037);
and U24521 (N_24521,N_21178,N_20873);
nand U24522 (N_24522,N_20649,N_22502);
or U24523 (N_24523,N_18073,N_22584);
or U24524 (N_24524,N_23796,N_21249);
and U24525 (N_24525,N_23930,N_20658);
and U24526 (N_24526,N_19945,N_21288);
nor U24527 (N_24527,N_18423,N_21722);
and U24528 (N_24528,N_23558,N_19312);
nand U24529 (N_24529,N_19273,N_20475);
and U24530 (N_24530,N_19044,N_23919);
or U24531 (N_24531,N_23191,N_21300);
xor U24532 (N_24532,N_20087,N_20471);
nand U24533 (N_24533,N_19598,N_22090);
or U24534 (N_24534,N_21976,N_19879);
nor U24535 (N_24535,N_18330,N_19780);
xnor U24536 (N_24536,N_22814,N_20805);
nand U24537 (N_24537,N_21209,N_23924);
or U24538 (N_24538,N_18579,N_22796);
xnor U24539 (N_24539,N_18437,N_18964);
nand U24540 (N_24540,N_18897,N_20586);
xor U24541 (N_24541,N_21006,N_18321);
nor U24542 (N_24542,N_20958,N_20387);
nor U24543 (N_24543,N_18148,N_22662);
xor U24544 (N_24544,N_22968,N_19711);
nand U24545 (N_24545,N_20100,N_18852);
nor U24546 (N_24546,N_21548,N_22963);
or U24547 (N_24547,N_18259,N_20221);
nor U24548 (N_24548,N_23777,N_19489);
and U24549 (N_24549,N_18371,N_19751);
nor U24550 (N_24550,N_20783,N_19988);
xnor U24551 (N_24551,N_23046,N_23829);
and U24552 (N_24552,N_20534,N_21423);
and U24553 (N_24553,N_22895,N_23675);
xnor U24554 (N_24554,N_18166,N_19801);
xor U24555 (N_24555,N_22143,N_21810);
or U24556 (N_24556,N_18487,N_19352);
nor U24557 (N_24557,N_19366,N_22108);
nor U24558 (N_24558,N_19057,N_21612);
or U24559 (N_24559,N_22371,N_22316);
xnor U24560 (N_24560,N_18675,N_18790);
xnor U24561 (N_24561,N_22879,N_20325);
nor U24562 (N_24562,N_23213,N_20480);
xnor U24563 (N_24563,N_23611,N_20283);
xor U24564 (N_24564,N_20546,N_19998);
xnor U24565 (N_24565,N_18584,N_19560);
nor U24566 (N_24566,N_20560,N_22333);
nor U24567 (N_24567,N_18801,N_22252);
nor U24568 (N_24568,N_18385,N_22428);
and U24569 (N_24569,N_18783,N_18668);
xnor U24570 (N_24570,N_20419,N_21665);
nand U24571 (N_24571,N_20073,N_19319);
xor U24572 (N_24572,N_18832,N_18433);
nand U24573 (N_24573,N_23835,N_18354);
xnor U24574 (N_24574,N_23128,N_21235);
and U24575 (N_24575,N_18520,N_22242);
and U24576 (N_24576,N_21677,N_20967);
or U24577 (N_24577,N_23125,N_18244);
and U24578 (N_24578,N_20606,N_20098);
xnor U24579 (N_24579,N_23733,N_22966);
and U24580 (N_24580,N_22349,N_18172);
and U24581 (N_24581,N_21907,N_23691);
nor U24582 (N_24582,N_20683,N_18511);
nor U24583 (N_24583,N_21986,N_19016);
nor U24584 (N_24584,N_18754,N_19865);
or U24585 (N_24585,N_21005,N_23803);
and U24586 (N_24586,N_18492,N_22826);
nand U24587 (N_24587,N_23921,N_22874);
or U24588 (N_24588,N_22126,N_18833);
and U24589 (N_24589,N_20259,N_22912);
nand U24590 (N_24590,N_21087,N_21408);
xnor U24591 (N_24591,N_21576,N_20088);
nand U24592 (N_24592,N_23236,N_22331);
nand U24593 (N_24593,N_18227,N_21037);
or U24594 (N_24594,N_22859,N_18362);
xor U24595 (N_24595,N_23269,N_18251);
and U24596 (N_24596,N_18130,N_22591);
and U24597 (N_24597,N_22224,N_20620);
or U24598 (N_24598,N_19062,N_20121);
nand U24599 (N_24599,N_18144,N_19046);
or U24600 (N_24600,N_19677,N_22158);
or U24601 (N_24601,N_22773,N_20604);
and U24602 (N_24602,N_23169,N_20945);
nor U24603 (N_24603,N_21646,N_20134);
and U24604 (N_24604,N_21565,N_21688);
or U24605 (N_24605,N_18914,N_23955);
or U24606 (N_24606,N_23469,N_23127);
or U24607 (N_24607,N_23418,N_20395);
nor U24608 (N_24608,N_19898,N_19787);
nand U24609 (N_24609,N_21328,N_23172);
nand U24610 (N_24610,N_23003,N_23095);
xnor U24611 (N_24611,N_18193,N_18542);
and U24612 (N_24612,N_21933,N_21666);
nor U24613 (N_24613,N_20929,N_21915);
nor U24614 (N_24614,N_23166,N_21657);
and U24615 (N_24615,N_23084,N_19863);
and U24616 (N_24616,N_23564,N_20984);
nor U24617 (N_24617,N_20983,N_19709);
xor U24618 (N_24618,N_19440,N_19637);
xnor U24619 (N_24619,N_19338,N_18655);
or U24620 (N_24620,N_19383,N_19672);
xor U24621 (N_24621,N_18256,N_22119);
or U24622 (N_24622,N_23499,N_19306);
or U24623 (N_24623,N_20519,N_20094);
nor U24624 (N_24624,N_19759,N_22244);
nor U24625 (N_24625,N_22682,N_22899);
xnor U24626 (N_24626,N_21031,N_21223);
and U24627 (N_24627,N_21758,N_20947);
nor U24628 (N_24628,N_19375,N_20680);
or U24629 (N_24629,N_21179,N_19363);
nor U24630 (N_24630,N_23618,N_23473);
nor U24631 (N_24631,N_23158,N_23326);
xor U24632 (N_24632,N_20920,N_21586);
and U24633 (N_24633,N_23968,N_18180);
or U24634 (N_24634,N_20744,N_23092);
xor U24635 (N_24635,N_20479,N_22526);
xnor U24636 (N_24636,N_20440,N_22516);
or U24637 (N_24637,N_20074,N_19845);
or U24638 (N_24638,N_23563,N_20310);
or U24639 (N_24639,N_21466,N_23298);
xor U24640 (N_24640,N_20598,N_23303);
xor U24641 (N_24641,N_19128,N_22492);
nand U24642 (N_24642,N_18538,N_22294);
nor U24643 (N_24643,N_23207,N_23765);
or U24644 (N_24644,N_20571,N_19500);
or U24645 (N_24645,N_20660,N_19576);
xor U24646 (N_24646,N_20359,N_23235);
nand U24647 (N_24647,N_23102,N_23999);
xor U24648 (N_24648,N_23226,N_22189);
nor U24649 (N_24649,N_23224,N_22885);
xor U24650 (N_24650,N_20530,N_21106);
nor U24651 (N_24651,N_19448,N_22469);
nor U24652 (N_24652,N_19470,N_23941);
or U24653 (N_24653,N_19817,N_22001);
nand U24654 (N_24654,N_18031,N_23998);
xnor U24655 (N_24655,N_20554,N_18027);
and U24656 (N_24656,N_19747,N_22277);
or U24657 (N_24657,N_23264,N_20816);
and U24658 (N_24658,N_18099,N_23527);
nand U24659 (N_24659,N_21904,N_19241);
nand U24660 (N_24660,N_18315,N_23546);
xnor U24661 (N_24661,N_20350,N_19066);
nand U24662 (N_24662,N_22547,N_22347);
nor U24663 (N_24663,N_20626,N_18061);
xnor U24664 (N_24664,N_22837,N_19803);
nor U24665 (N_24665,N_21080,N_22757);
nor U24666 (N_24666,N_18896,N_22904);
nor U24667 (N_24667,N_20331,N_20863);
or U24668 (N_24668,N_23149,N_20083);
and U24669 (N_24669,N_19105,N_22113);
nor U24670 (N_24670,N_20577,N_23375);
and U24671 (N_24671,N_20538,N_19260);
or U24672 (N_24672,N_21906,N_18597);
or U24673 (N_24673,N_18900,N_19033);
and U24674 (N_24674,N_23279,N_19467);
xnor U24675 (N_24675,N_19248,N_19720);
and U24676 (N_24676,N_22082,N_19382);
xor U24677 (N_24677,N_19152,N_18973);
and U24678 (N_24678,N_22628,N_20197);
or U24679 (N_24679,N_21098,N_20498);
xnor U24680 (N_24680,N_23645,N_21027);
or U24681 (N_24681,N_23105,N_19195);
and U24682 (N_24682,N_22039,N_20020);
nand U24683 (N_24683,N_22213,N_20322);
or U24684 (N_24684,N_20677,N_20611);
or U24685 (N_24685,N_20822,N_20211);
nand U24686 (N_24686,N_18310,N_20936);
nand U24687 (N_24687,N_19753,N_21304);
nor U24688 (N_24688,N_21600,N_22543);
and U24689 (N_24689,N_22956,N_18626);
nand U24690 (N_24690,N_21232,N_21181);
nor U24691 (N_24691,N_19939,N_22207);
nand U24692 (N_24692,N_18701,N_18797);
and U24693 (N_24693,N_21595,N_22756);
and U24694 (N_24694,N_18378,N_18804);
nand U24695 (N_24695,N_18892,N_19043);
xnor U24696 (N_24696,N_22867,N_22238);
nand U24697 (N_24697,N_19852,N_18541);
or U24698 (N_24698,N_20429,N_21854);
or U24699 (N_24699,N_20222,N_22758);
and U24700 (N_24700,N_23449,N_23528);
or U24701 (N_24701,N_22147,N_23157);
nor U24702 (N_24702,N_18269,N_22178);
nor U24703 (N_24703,N_22634,N_21498);
xor U24704 (N_24704,N_18860,N_20361);
xnor U24705 (N_24705,N_18693,N_23171);
or U24706 (N_24706,N_20896,N_21756);
nand U24707 (N_24707,N_21649,N_18658);
nor U24708 (N_24708,N_23840,N_21382);
xnor U24709 (N_24709,N_22886,N_19977);
or U24710 (N_24710,N_20767,N_22450);
and U24711 (N_24711,N_18370,N_18247);
and U24712 (N_24712,N_20907,N_19405);
or U24713 (N_24713,N_20727,N_19263);
nor U24714 (N_24714,N_18528,N_22211);
and U24715 (N_24715,N_23702,N_22303);
and U24716 (N_24716,N_18548,N_19821);
or U24717 (N_24717,N_21973,N_18058);
nand U24718 (N_24718,N_20763,N_20721);
xor U24719 (N_24719,N_20569,N_19622);
or U24720 (N_24720,N_22626,N_20633);
nand U24721 (N_24721,N_21048,N_22042);
and U24722 (N_24722,N_23305,N_22249);
or U24723 (N_24723,N_22664,N_21615);
nor U24724 (N_24724,N_19625,N_20957);
or U24725 (N_24725,N_22614,N_23347);
or U24726 (N_24726,N_19641,N_20902);
and U24727 (N_24727,N_22573,N_19542);
nor U24728 (N_24728,N_20814,N_22205);
or U24729 (N_24729,N_18842,N_22014);
nor U24730 (N_24730,N_23413,N_20585);
and U24731 (N_24731,N_22493,N_21251);
or U24732 (N_24732,N_21238,N_19329);
nor U24733 (N_24733,N_23740,N_20939);
and U24734 (N_24734,N_19639,N_20138);
and U24735 (N_24735,N_23508,N_21397);
xor U24736 (N_24736,N_19245,N_22381);
and U24737 (N_24737,N_19739,N_19293);
nor U24738 (N_24738,N_19818,N_18389);
nand U24739 (N_24739,N_21173,N_19388);
or U24740 (N_24740,N_18770,N_23511);
and U24741 (N_24741,N_22818,N_22382);
nor U24742 (N_24742,N_20321,N_18108);
or U24743 (N_24743,N_21187,N_23446);
xnor U24744 (N_24744,N_23364,N_18313);
nand U24745 (N_24745,N_23795,N_19262);
and U24746 (N_24746,N_21329,N_22743);
xnor U24747 (N_24747,N_23109,N_18399);
xnor U24748 (N_24748,N_20474,N_21183);
nand U24749 (N_24749,N_23962,N_23792);
or U24750 (N_24750,N_23431,N_21579);
nor U24751 (N_24751,N_21823,N_19341);
xor U24752 (N_24752,N_18489,N_19731);
or U24753 (N_24753,N_21239,N_23569);
or U24754 (N_24754,N_21867,N_23868);
or U24755 (N_24755,N_21954,N_21274);
nand U24756 (N_24756,N_19454,N_23745);
xor U24757 (N_24757,N_21099,N_20399);
nor U24758 (N_24758,N_20045,N_20478);
xor U24759 (N_24759,N_21494,N_21171);
xor U24760 (N_24760,N_18025,N_19635);
nor U24761 (N_24761,N_19258,N_22299);
and U24762 (N_24762,N_19547,N_18086);
and U24763 (N_24763,N_23650,N_23633);
and U24764 (N_24764,N_23272,N_19236);
nand U24765 (N_24765,N_23295,N_22002);
nand U24766 (N_24766,N_22892,N_23192);
nor U24767 (N_24767,N_20847,N_19170);
and U24768 (N_24768,N_18909,N_19486);
nor U24769 (N_24769,N_20718,N_20323);
xnor U24770 (N_24770,N_23657,N_18381);
nand U24771 (N_24771,N_21211,N_18941);
nand U24772 (N_24772,N_22419,N_19296);
or U24773 (N_24773,N_22280,N_22598);
and U24774 (N_24774,N_22775,N_22669);
or U24775 (N_24775,N_22596,N_21736);
nand U24776 (N_24776,N_19527,N_18728);
or U24777 (N_24777,N_19776,N_23324);
nand U24778 (N_24778,N_23343,N_23857);
nand U24779 (N_24779,N_20672,N_20933);
nand U24780 (N_24780,N_20559,N_20209);
nor U24781 (N_24781,N_20230,N_19060);
and U24782 (N_24782,N_20339,N_18168);
and U24783 (N_24783,N_20123,N_22946);
nor U24784 (N_24784,N_19647,N_21253);
and U24785 (N_24785,N_21258,N_21156);
nor U24786 (N_24786,N_19913,N_18924);
xnor U24787 (N_24787,N_19737,N_19721);
or U24788 (N_24788,N_19537,N_19844);
nand U24789 (N_24789,N_19132,N_21243);
nor U24790 (N_24790,N_21111,N_23595);
xnor U24791 (N_24791,N_19501,N_20306);
nand U24792 (N_24792,N_18484,N_18382);
nor U24793 (N_24793,N_20373,N_23887);
nor U24794 (N_24794,N_18903,N_18338);
nor U24795 (N_24795,N_22564,N_18402);
or U24796 (N_24796,N_19113,N_19789);
nor U24797 (N_24797,N_18079,N_18198);
xor U24798 (N_24798,N_19893,N_18709);
nor U24799 (N_24799,N_22030,N_23709);
and U24800 (N_24800,N_21058,N_21326);
nand U24801 (N_24801,N_22926,N_18907);
or U24802 (N_24802,N_19847,N_21456);
or U24803 (N_24803,N_18902,N_19269);
nor U24804 (N_24804,N_21638,N_19602);
and U24805 (N_24805,N_22631,N_21729);
nand U24806 (N_24806,N_20797,N_18132);
nor U24807 (N_24807,N_23421,N_22195);
nand U24808 (N_24808,N_19657,N_21532);
or U24809 (N_24809,N_18653,N_20749);
and U24810 (N_24810,N_18773,N_20096);
or U24811 (N_24811,N_21365,N_20948);
nand U24812 (N_24812,N_21551,N_21322);
or U24813 (N_24813,N_20990,N_22854);
nor U24814 (N_24814,N_22338,N_22984);
nand U24815 (N_24815,N_23056,N_19081);
nor U24816 (N_24816,N_23138,N_20219);
xnor U24817 (N_24817,N_20273,N_20512);
or U24818 (N_24818,N_21960,N_19168);
nor U24819 (N_24819,N_20425,N_22027);
or U24820 (N_24820,N_21097,N_18586);
and U24821 (N_24821,N_19773,N_23605);
nand U24822 (N_24822,N_18239,N_19316);
or U24823 (N_24823,N_21150,N_23736);
or U24824 (N_24824,N_21483,N_19157);
nor U24825 (N_24825,N_18934,N_18956);
xnor U24826 (N_24826,N_23146,N_20257);
nand U24827 (N_24827,N_18115,N_19781);
or U24828 (N_24828,N_23800,N_20543);
or U24829 (N_24829,N_21060,N_21263);
nor U24830 (N_24830,N_23519,N_22803);
nor U24831 (N_24831,N_18596,N_19631);
or U24832 (N_24832,N_18463,N_19282);
nand U24833 (N_24833,N_20642,N_19662);
nor U24834 (N_24834,N_20688,N_19367);
and U24835 (N_24835,N_18540,N_19052);
nor U24836 (N_24836,N_19991,N_18847);
nand U24837 (N_24837,N_19431,N_23047);
nor U24838 (N_24838,N_22456,N_18601);
nand U24839 (N_24839,N_23237,N_20720);
nor U24840 (N_24840,N_21452,N_20029);
or U24841 (N_24841,N_22192,N_21449);
nand U24842 (N_24842,N_23427,N_23444);
and U24843 (N_24843,N_20834,N_23896);
and U24844 (N_24844,N_22930,N_23183);
and U24845 (N_24845,N_21433,N_18822);
and U24846 (N_24846,N_20187,N_23108);
or U24847 (N_24847,N_21170,N_19122);
and U24848 (N_24848,N_19164,N_23028);
or U24849 (N_24849,N_20000,N_22860);
nor U24850 (N_24850,N_19322,N_22907);
or U24851 (N_24851,N_23310,N_20855);
nor U24852 (N_24852,N_19409,N_22499);
nor U24853 (N_24853,N_20295,N_20263);
nor U24854 (N_24854,N_19649,N_20774);
nor U24855 (N_24855,N_23074,N_23750);
nor U24856 (N_24856,N_18933,N_22098);
or U24857 (N_24857,N_21358,N_18212);
or U24858 (N_24858,N_21016,N_19398);
nor U24859 (N_24859,N_18179,N_21216);
xnor U24860 (N_24860,N_23586,N_20021);
nor U24861 (N_24861,N_21686,N_18296);
nand U24862 (N_24862,N_21503,N_20337);
xnor U24863 (N_24863,N_20476,N_18513);
and U24864 (N_24864,N_22072,N_19441);
xnor U24865 (N_24865,N_21913,N_18794);
nor U24866 (N_24866,N_23926,N_22723);
nand U24867 (N_24867,N_19089,N_20204);
xnor U24868 (N_24868,N_20561,N_23249);
nand U24869 (N_24869,N_20501,N_23442);
or U24870 (N_24870,N_18849,N_18131);
nand U24871 (N_24871,N_20510,N_20836);
or U24872 (N_24872,N_20844,N_18527);
nor U24873 (N_24873,N_20496,N_20185);
or U24874 (N_24874,N_20999,N_21598);
or U24875 (N_24875,N_23420,N_23552);
xor U24876 (N_24876,N_18441,N_19309);
xnor U24877 (N_24877,N_20921,N_22985);
or U24878 (N_24878,N_21871,N_18942);
or U24879 (N_24879,N_21764,N_19173);
or U24880 (N_24880,N_20441,N_23509);
xnor U24881 (N_24881,N_18442,N_21479);
and U24882 (N_24882,N_22768,N_18035);
xnor U24883 (N_24883,N_18915,N_19799);
or U24884 (N_24884,N_23664,N_19116);
and U24885 (N_24885,N_20057,N_20813);
nand U24886 (N_24886,N_19468,N_23915);
nand U24887 (N_24887,N_18841,N_23045);
nor U24888 (N_24888,N_18602,N_21042);
nand U24889 (N_24889,N_22396,N_23798);
xor U24890 (N_24890,N_23231,N_20769);
nor U24891 (N_24891,N_21001,N_20740);
nor U24892 (N_24892,N_21999,N_19333);
nand U24893 (N_24893,N_22653,N_18920);
nor U24894 (N_24894,N_18462,N_19870);
xnor U24895 (N_24895,N_22150,N_22047);
nand U24896 (N_24896,N_19127,N_19469);
xnor U24897 (N_24897,N_19463,N_23000);
nand U24898 (N_24898,N_21188,N_19532);
nand U24899 (N_24899,N_22971,N_22380);
nor U24900 (N_24900,N_20004,N_21000);
and U24901 (N_24901,N_22051,N_23368);
nor U24902 (N_24902,N_18328,N_20544);
xor U24903 (N_24903,N_19321,N_18013);
xnor U24904 (N_24904,N_20635,N_21422);
and U24905 (N_24905,N_18699,N_23479);
nand U24906 (N_24906,N_23977,N_20738);
or U24907 (N_24907,N_18857,N_20105);
xnor U24908 (N_24908,N_19124,N_19073);
xnor U24909 (N_24909,N_20282,N_21862);
nand U24910 (N_24910,N_21738,N_21945);
and U24911 (N_24911,N_22037,N_23641);
nand U24912 (N_24912,N_19871,N_20118);
or U24913 (N_24913,N_18300,N_23610);
and U24914 (N_24914,N_21102,N_22774);
nor U24915 (N_24915,N_21327,N_18951);
xor U24916 (N_24916,N_19325,N_18855);
xor U24917 (N_24917,N_23300,N_19752);
xnor U24918 (N_24918,N_18543,N_18273);
or U24919 (N_24919,N_23419,N_20049);
and U24920 (N_24920,N_18535,N_19292);
nand U24921 (N_24921,N_21998,N_21052);
and U24922 (N_24922,N_21044,N_22005);
or U24923 (N_24923,N_18858,N_18093);
nand U24924 (N_24924,N_19861,N_20366);
or U24925 (N_24925,N_20704,N_21698);
nor U24926 (N_24926,N_20781,N_23720);
or U24927 (N_24927,N_21458,N_23635);
xnor U24928 (N_24928,N_20006,N_20296);
nand U24929 (N_24929,N_18106,N_19580);
or U24930 (N_24930,N_18574,N_20065);
and U24931 (N_24931,N_18557,N_18785);
and U24932 (N_24932,N_23497,N_21409);
and U24933 (N_24933,N_18262,N_18678);
nand U24934 (N_24934,N_18749,N_23532);
or U24935 (N_24935,N_21653,N_18499);
nor U24936 (N_24936,N_22239,N_20932);
nor U24937 (N_24937,N_22057,N_22788);
nor U24938 (N_24938,N_19213,N_19223);
nor U24939 (N_24939,N_21914,N_19678);
nor U24940 (N_24940,N_22700,N_21949);
and U24941 (N_24941,N_22423,N_22344);
and U24942 (N_24942,N_18919,N_21857);
nor U24943 (N_24943,N_23465,N_22167);
nor U24944 (N_24944,N_19689,N_23215);
xnor U24945 (N_24945,N_19612,N_18517);
and U24946 (N_24946,N_23069,N_21236);
nand U24947 (N_24947,N_20018,N_21791);
nand U24948 (N_24948,N_18200,N_20132);
nor U24949 (N_24949,N_18051,N_23088);
and U24950 (N_24950,N_22183,N_22571);
nor U24951 (N_24951,N_22267,N_18937);
xnor U24952 (N_24952,N_21026,N_20871);
nor U24953 (N_24953,N_19857,N_23673);
and U24954 (N_24954,N_21086,N_18261);
nor U24955 (N_24955,N_20414,N_23116);
xnor U24956 (N_24956,N_19096,N_22633);
or U24957 (N_24957,N_21225,N_23877);
xor U24958 (N_24958,N_21193,N_19246);
nand U24959 (N_24959,N_22727,N_20128);
and U24960 (N_24960,N_19906,N_22529);
or U24961 (N_24961,N_21520,N_19530);
nand U24962 (N_24962,N_21360,N_23342);
and U24963 (N_24963,N_22473,N_20427);
or U24964 (N_24964,N_20353,N_23799);
or U24965 (N_24965,N_20974,N_20917);
xor U24966 (N_24966,N_22697,N_20178);
nand U24967 (N_24967,N_19390,N_23174);
nor U24968 (N_24968,N_19023,N_18670);
and U24969 (N_24969,N_20445,N_23824);
or U24970 (N_24970,N_21932,N_18575);
nor U24971 (N_24971,N_23825,N_20801);
xor U24972 (N_24972,N_20987,N_18656);
and U24973 (N_24973,N_22334,N_23482);
xnor U24974 (N_24974,N_21912,N_23101);
nor U24975 (N_24975,N_22250,N_18165);
or U24976 (N_24976,N_19430,N_20679);
nand U24977 (N_24977,N_20411,N_20327);
nand U24978 (N_24978,N_20652,N_18292);
nand U24979 (N_24979,N_19754,N_18908);
and U24980 (N_24980,N_21219,N_23685);
nor U24981 (N_24981,N_19175,N_23009);
nand U24982 (N_24982,N_19102,N_22176);
nand U24983 (N_24983,N_23770,N_18697);
xor U24984 (N_24984,N_23341,N_21781);
nand U24985 (N_24985,N_19410,N_20002);
xor U24986 (N_24986,N_21096,N_22054);
or U24987 (N_24987,N_19701,N_23730);
nor U24988 (N_24988,N_23488,N_20281);
and U24989 (N_24989,N_19729,N_21210);
nor U24990 (N_24990,N_19072,N_18578);
nor U24991 (N_24991,N_21462,N_19667);
xnor U24992 (N_24992,N_20292,N_20640);
nor U24993 (N_24993,N_20362,N_20656);
and U24994 (N_24994,N_18913,N_19209);
nor U24995 (N_24995,N_23551,N_23785);
or U24996 (N_24996,N_20451,N_19503);
and U24997 (N_24997,N_21559,N_22273);
nor U24998 (N_24998,N_19762,N_19793);
or U24999 (N_24999,N_20682,N_20484);
or U25000 (N_25000,N_18705,N_23329);
xnor U25001 (N_25001,N_20370,N_21338);
xor U25002 (N_25002,N_21840,N_18834);
and U25003 (N_25003,N_19588,N_22805);
nor U25004 (N_25004,N_22080,N_21078);
and U25005 (N_25005,N_22652,N_19480);
nor U25006 (N_25006,N_23067,N_21296);
nand U25007 (N_25007,N_21918,N_20449);
xnor U25008 (N_25008,N_21687,N_23357);
and U25009 (N_25009,N_21683,N_23579);
nor U25010 (N_25010,N_19987,N_21105);
nand U25011 (N_25011,N_18220,N_21887);
xnor U25012 (N_25012,N_20751,N_20277);
xnor U25013 (N_25013,N_21290,N_21184);
nand U25014 (N_25014,N_22889,N_23029);
nor U25015 (N_25015,N_19760,N_18029);
or U25016 (N_25016,N_18515,N_21882);
and U25017 (N_25017,N_22615,N_19652);
and U25018 (N_25018,N_21024,N_19149);
and U25019 (N_25019,N_19007,N_21902);
nor U25020 (N_25020,N_22987,N_18742);
nor U25021 (N_25021,N_23201,N_20341);
xor U25022 (N_25022,N_19910,N_23299);
nand U25023 (N_25023,N_20390,N_18392);
and U25024 (N_25024,N_22220,N_21118);
nand U25025 (N_25025,N_20151,N_18235);
and U25026 (N_25026,N_22637,N_21492);
or U25027 (N_25027,N_19911,N_18605);
and U25028 (N_25028,N_21951,N_18276);
nor U25029 (N_25029,N_19656,N_22132);
nand U25030 (N_25030,N_20938,N_21416);
xnor U25031 (N_25031,N_21583,N_18722);
or U25032 (N_25032,N_21539,N_18608);
nor U25033 (N_25033,N_18612,N_18968);
nor U25034 (N_25034,N_19238,N_22389);
and U25035 (N_25035,N_23719,N_18380);
or U25036 (N_25036,N_21839,N_18665);
nor U25037 (N_25037,N_20382,N_20188);
nor U25038 (N_25038,N_20159,N_22969);
nor U25039 (N_25039,N_22255,N_18518);
and U25040 (N_25040,N_19187,N_21336);
nor U25041 (N_25041,N_18600,N_18865);
or U25042 (N_25042,N_23412,N_22180);
or U25043 (N_25043,N_20408,N_22241);
nand U25044 (N_25044,N_18210,N_18853);
nor U25045 (N_25045,N_20439,N_18379);
and U25046 (N_25046,N_20953,N_18248);
xor U25047 (N_25047,N_20131,N_22636);
nor U25048 (N_25048,N_19037,N_22593);
nor U25049 (N_25049,N_21437,N_20467);
xor U25050 (N_25050,N_23042,N_18571);
xnor U25051 (N_25051,N_18889,N_20216);
or U25052 (N_25052,N_19320,N_19854);
nand U25053 (N_25053,N_21070,N_23889);
or U25054 (N_25054,N_22945,N_18554);
or U25055 (N_25055,N_23048,N_22074);
nand U25056 (N_25056,N_23008,N_22352);
and U25057 (N_25057,N_20246,N_21762);
or U25058 (N_25058,N_20565,N_22508);
xor U25059 (N_25059,N_21817,N_19685);
xor U25060 (N_25060,N_19114,N_23861);
xnor U25061 (N_25061,N_18110,N_23037);
nor U25062 (N_25062,N_21769,N_19668);
nor U25063 (N_25063,N_22842,N_21259);
and U25064 (N_25064,N_20639,N_19082);
nor U25065 (N_25065,N_19412,N_19690);
nand U25066 (N_25066,N_18109,N_22767);
xnor U25067 (N_25067,N_20595,N_21878);
and U25068 (N_25068,N_18721,N_18514);
or U25069 (N_25069,N_23204,N_18439);
or U25070 (N_25070,N_21344,N_18103);
nand U25071 (N_25071,N_22509,N_18275);
or U25072 (N_25072,N_21905,N_23435);
nand U25073 (N_25073,N_22429,N_23397);
xor U25074 (N_25074,N_22656,N_23135);
nand U25075 (N_25075,N_21089,N_23181);
or U25076 (N_25076,N_18477,N_21527);
nor U25077 (N_25077,N_22214,N_19805);
nor U25078 (N_25078,N_18336,N_19097);
and U25079 (N_25079,N_22880,N_21533);
nor U25080 (N_25080,N_23317,N_23271);
nand U25081 (N_25081,N_20112,N_22925);
or U25082 (N_25082,N_20986,N_23206);
xor U25083 (N_25083,N_22448,N_23396);
nor U25084 (N_25084,N_23604,N_21809);
xor U25085 (N_25085,N_21730,N_18101);
nor U25086 (N_25086,N_18283,N_22233);
xnor U25087 (N_25087,N_21908,N_20796);
xnor U25088 (N_25088,N_21775,N_23763);
nand U25089 (N_25089,N_21599,N_23480);
nand U25090 (N_25090,N_22839,N_20591);
and U25091 (N_25091,N_18299,N_22328);
nor U25092 (N_25092,N_21343,N_22513);
and U25093 (N_25093,N_23781,N_22894);
xnor U25094 (N_25094,N_20417,N_20369);
and U25095 (N_25095,N_18887,N_21121);
nor U25096 (N_25096,N_19868,N_20962);
xnor U25097 (N_25097,N_19936,N_19359);
nor U25098 (N_25098,N_20592,N_22780);
xor U25099 (N_25099,N_23939,N_23094);
xnor U25100 (N_25100,N_18066,N_18835);
and U25101 (N_25101,N_20207,N_18720);
or U25102 (N_25102,N_22927,N_21966);
xor U25103 (N_25103,N_23443,N_22645);
and U25104 (N_25104,N_21208,N_21030);
xnor U25105 (N_25105,N_22556,N_19279);
and U25106 (N_25106,N_18776,N_22363);
and U25107 (N_25107,N_23995,N_22124);
nor U25108 (N_25108,N_18505,N_21578);
and U25109 (N_25109,N_21369,N_23848);
and U25110 (N_25110,N_21056,N_18768);
and U25111 (N_25111,N_20698,N_20117);
or U25112 (N_25112,N_22052,N_20007);
and U25113 (N_25113,N_18490,N_19541);
nand U25114 (N_25114,N_22149,N_18512);
or U25115 (N_25115,N_21981,N_18004);
and U25116 (N_25116,N_21414,N_21115);
nor U25117 (N_25117,N_20291,N_19406);
xnor U25118 (N_25118,N_20931,N_23952);
xor U25119 (N_25119,N_19849,N_21376);
xnor U25120 (N_25120,N_19459,N_19691);
xor U25121 (N_25121,N_20469,N_18927);
nor U25122 (N_25122,N_21675,N_21623);
or U25123 (N_25123,N_21461,N_19989);
nor U25124 (N_25124,N_23141,N_21700);
nand U25125 (N_25125,N_19812,N_18345);
or U25126 (N_25126,N_23362,N_21167);
xor U25127 (N_25127,N_23356,N_19981);
nand U25128 (N_25128,N_18339,N_20365);
xor U25129 (N_25129,N_23416,N_20069);
xnor U25130 (N_25130,N_20597,N_20747);
nand U25131 (N_25131,N_23562,N_23223);
nand U25132 (N_25132,N_19934,N_20459);
xor U25133 (N_25133,N_23087,N_19644);
nand U25134 (N_25134,N_18809,N_23280);
and U25135 (N_25135,N_20581,N_21910);
nor U25136 (N_25136,N_22900,N_23229);
or U25137 (N_25137,N_22820,N_20247);
and U25138 (N_25138,N_20717,N_21398);
and U25139 (N_25139,N_20758,N_22606);
or U25140 (N_25140,N_23544,N_18730);
xor U25141 (N_25141,N_19976,N_22411);
xnor U25142 (N_25142,N_20009,N_19867);
nor U25143 (N_25143,N_20653,N_23974);
xnor U25144 (N_25144,N_20759,N_19330);
and U25145 (N_25145,N_23430,N_23291);
xnor U25146 (N_25146,N_22166,N_20675);
nor U25147 (N_25147,N_19557,N_19270);
xnor U25148 (N_25148,N_21771,N_23366);
xor U25149 (N_25149,N_22313,N_23485);
or U25150 (N_25150,N_18958,N_23110);
or U25151 (N_25151,N_23327,N_19661);
nand U25152 (N_25152,N_20950,N_18376);
or U25153 (N_25153,N_23880,N_23335);
nor U25154 (N_25154,N_21127,N_20110);
nand U25155 (N_25155,N_23971,N_22812);
and U25156 (N_25156,N_22409,N_23348);
xor U25157 (N_25157,N_18599,N_22351);
nand U25158 (N_25158,N_23670,N_23674);
nor U25159 (N_25159,N_23699,N_22485);
and U25160 (N_25160,N_21283,N_20980);
nor U25161 (N_25161,N_22097,N_23549);
and U25162 (N_25162,N_19219,N_21755);
and U25163 (N_25163,N_23894,N_23071);
nor U25164 (N_25164,N_23031,N_19392);
xor U25165 (N_25165,N_18506,N_21890);
and U25166 (N_25166,N_19923,N_18098);
nor U25167 (N_25167,N_19839,N_18906);
nor U25168 (N_25168,N_20426,N_22616);
nor U25169 (N_25169,N_21783,N_23766);
nand U25170 (N_25170,N_22741,N_20771);
and U25171 (N_25171,N_21280,N_23241);
and U25172 (N_25172,N_22959,N_23314);
nand U25173 (N_25173,N_23631,N_20319);
or U25174 (N_25174,N_22305,N_18959);
and U25175 (N_25175,N_22317,N_23548);
and U25176 (N_25176,N_18947,N_23624);
and U25177 (N_25177,N_19983,N_22703);
nand U25178 (N_25178,N_23683,N_21457);
and U25179 (N_25179,N_22388,N_18183);
nand U25180 (N_25180,N_23290,N_18946);
and U25181 (N_25181,N_18225,N_22011);
xor U25182 (N_25182,N_23016,N_23156);
xnor U25183 (N_25183,N_20533,N_23866);
or U25184 (N_25184,N_22497,N_20097);
nand U25185 (N_25185,N_19464,N_23123);
nor U25186 (N_25186,N_21334,N_21827);
nand U25187 (N_25187,N_20916,N_21451);
or U25188 (N_25188,N_21018,N_22391);
nand U25189 (N_25189,N_19726,N_20340);
nor U25190 (N_25190,N_22607,N_18059);
xnor U25191 (N_25191,N_23823,N_22171);
nor U25192 (N_25192,N_23813,N_23567);
xor U25193 (N_25193,N_18744,N_20482);
xor U25194 (N_25194,N_18309,N_23515);
nand U25195 (N_25195,N_19944,N_21759);
and U25196 (N_25196,N_22000,N_18854);
nand U25197 (N_25197,N_23103,N_18867);
nand U25198 (N_25198,N_22589,N_18012);
and U25199 (N_25199,N_19437,N_21948);
nand U25200 (N_25200,N_19005,N_19518);
and U25201 (N_25201,N_18265,N_21947);
and U25202 (N_25202,N_21472,N_23693);
nand U25203 (N_25203,N_21130,N_20093);
and U25204 (N_25204,N_21293,N_19304);
nand U25205 (N_25205,N_19230,N_18409);
xor U25206 (N_25206,N_23004,N_22861);
nand U25207 (N_25207,N_18470,N_18694);
and U25208 (N_25208,N_19673,N_21880);
nor U25209 (N_25209,N_18806,N_21988);
and U25210 (N_25210,N_18032,N_22680);
and U25211 (N_25211,N_22491,N_22061);
and U25212 (N_25212,N_18257,N_20383);
nand U25213 (N_25213,N_22688,N_22901);
xor U25214 (N_25214,N_19351,N_23311);
nand U25215 (N_25215,N_22973,N_20865);
and U25216 (N_25216,N_18779,N_21264);
xor U25217 (N_25217,N_21703,N_19654);
nor U25218 (N_25218,N_23850,N_18751);
and U25219 (N_25219,N_19347,N_23780);
nand U25220 (N_25220,N_19788,N_21428);
xor U25221 (N_25221,N_19130,N_23398);
and U25222 (N_25222,N_19462,N_20375);
nand U25223 (N_25223,N_22873,N_21157);
nor U25224 (N_25224,N_23211,N_18795);
or U25225 (N_25225,N_18995,N_20899);
xor U25226 (N_25226,N_20086,N_21585);
nor U25227 (N_25227,N_18039,N_19275);
xnor U25228 (N_25228,N_19259,N_19985);
or U25229 (N_25229,N_21681,N_22063);
nor U25230 (N_25230,N_19555,N_21530);
nor U25231 (N_25231,N_20507,N_23560);
nand U25232 (N_25232,N_23472,N_20757);
or U25233 (N_25233,N_22376,N_22481);
and U25234 (N_25234,N_18155,N_19493);
or U25235 (N_25235,N_18475,N_19978);
nor U25236 (N_25236,N_18421,N_21816);
and U25237 (N_25237,N_19343,N_18182);
and U25238 (N_25238,N_19693,N_22320);
nand U25239 (N_25239,N_22553,N_18939);
nand U25240 (N_25240,N_21256,N_18882);
xor U25241 (N_25241,N_19895,N_21271);
xnor U25242 (N_25242,N_23403,N_20812);
xnor U25243 (N_25243,N_22210,N_23782);
nand U25244 (N_25244,N_21155,N_21861);
and U25245 (N_25245,N_18628,N_19387);
and U25246 (N_25246,N_21573,N_18069);
xnor U25247 (N_25247,N_18372,N_21609);
nand U25248 (N_25248,N_20497,N_21095);
or U25249 (N_25249,N_21117,N_19361);
nor U25250 (N_25250,N_18729,N_22345);
nand U25251 (N_25251,N_21797,N_19216);
nor U25252 (N_25252,N_21002,N_23646);
and U25253 (N_25253,N_23666,N_22263);
and U25254 (N_25254,N_22586,N_19198);
nor U25255 (N_25255,N_18627,N_22148);
xor U25256 (N_25256,N_18642,N_20420);
nand U25257 (N_25257,N_19563,N_20186);
nor U25258 (N_25258,N_20090,N_18237);
and U25259 (N_25259,N_20486,N_18861);
and U25260 (N_25260,N_22026,N_21351);
nand U25261 (N_25261,N_19474,N_23319);
or U25262 (N_25262,N_20017,N_20993);
and U25263 (N_25263,N_21450,N_22486);
xnor U25264 (N_25264,N_23859,N_18562);
and U25265 (N_25265,N_20053,N_23258);
and U25266 (N_25266,N_19186,N_22475);
xnor U25267 (N_25267,N_20418,N_19538);
or U25268 (N_25268,N_21465,N_22577);
nor U25269 (N_25269,N_22066,N_22464);
nor U25270 (N_25270,N_19420,N_19932);
or U25271 (N_25271,N_21523,N_20276);
nand U25272 (N_25272,N_21980,N_19419);
nor U25273 (N_25273,N_23964,N_21169);
nand U25274 (N_25274,N_18952,N_22449);
nand U25275 (N_25275,N_21785,N_21629);
xor U25276 (N_25276,N_21992,N_19619);
and U25277 (N_25277,N_23263,N_19565);
nor U25278 (N_25278,N_18792,N_23949);
or U25279 (N_25279,N_20969,N_23252);
or U25280 (N_25280,N_18050,N_22770);
nor U25281 (N_25281,N_18525,N_18504);
or U25282 (N_25282,N_21165,N_19808);
or U25283 (N_25283,N_22392,N_20111);
nor U25284 (N_25284,N_23315,N_21955);
xor U25285 (N_25285,N_22130,N_19257);
xnor U25286 (N_25286,N_22747,N_21021);
or U25287 (N_25287,N_23471,N_22731);
and U25288 (N_25288,N_20708,N_22141);
xor U25289 (N_25289,N_21410,N_23602);
and U25290 (N_25290,N_21952,N_22226);
nand U25291 (N_25291,N_18234,N_22191);
and U25292 (N_25292,N_20696,N_21830);
nor U25293 (N_25293,N_23918,N_18123);
nand U25294 (N_25294,N_20285,N_20828);
and U25295 (N_25295,N_21476,N_19429);
nand U25296 (N_25296,N_21153,N_20645);
and U25297 (N_25297,N_20511,N_20066);
and U25298 (N_25298,N_19004,N_22393);
and U25299 (N_25299,N_20242,N_20888);
nor U25300 (N_25300,N_18150,N_21834);
nand U25301 (N_25301,N_21443,N_21032);
nor U25302 (N_25302,N_20064,N_22869);
or U25303 (N_25303,N_22916,N_23656);
and U25304 (N_25304,N_21440,N_23614);
nand U25305 (N_25305,N_19671,N_18859);
xnor U25306 (N_25306,N_22046,N_22949);
xnor U25307 (N_25307,N_21869,N_19450);
and U25308 (N_25308,N_19551,N_22549);
xnor U25309 (N_25309,N_19345,N_18311);
nor U25310 (N_25310,N_18003,N_23545);
xor U25311 (N_25311,N_18364,N_22936);
and U25312 (N_25312,N_18318,N_18057);
and U25313 (N_25313,N_22840,N_18871);
xnor U25314 (N_25314,N_18782,N_23378);
nor U25315 (N_25315,N_20238,N_18692);
or U25316 (N_25316,N_18866,N_19901);
nand U25317 (N_25317,N_23711,N_19120);
and U25318 (N_25318,N_18446,N_20376);
or U25319 (N_25319,N_22157,N_22407);
nor U25320 (N_25320,N_23408,N_22845);
nand U25321 (N_25321,N_22691,N_23890);
nand U25322 (N_25322,N_19042,N_23320);
or U25323 (N_25323,N_19962,N_18001);
nor U25324 (N_25324,N_18820,N_21278);
nor U25325 (N_25325,N_21426,N_21588);
and U25326 (N_25326,N_22734,N_22501);
or U25327 (N_25327,N_23707,N_19999);
nor U25328 (N_25328,N_22962,N_22763);
and U25329 (N_25329,N_23023,N_21319);
nor U25330 (N_25330,N_23654,N_21571);
or U25331 (N_25331,N_23190,N_22321);
nand U25332 (N_25332,N_22995,N_23860);
and U25333 (N_25333,N_20737,N_21265);
and U25334 (N_25334,N_21191,N_19961);
or U25335 (N_25335,N_21459,N_19609);
and U25336 (N_25336,N_18905,N_18173);
nor U25337 (N_25337,N_23282,N_19769);
and U25338 (N_25338,N_20777,N_20989);
nor U25339 (N_25339,N_21022,N_19881);
and U25340 (N_25340,N_18622,N_20522);
and U25341 (N_25341,N_23424,N_21158);
or U25342 (N_25342,N_19669,N_21706);
xor U25343 (N_25343,N_21593,N_18102);
or U25344 (N_25344,N_19161,N_19651);
nor U25345 (N_25345,N_18359,N_20826);
and U25346 (N_25346,N_23879,N_19790);
nand U25347 (N_25347,N_22378,N_22721);
and U25348 (N_25348,N_21592,N_23450);
xor U25349 (N_25349,N_21135,N_19705);
xor U25350 (N_25350,N_20879,N_21112);
or U25351 (N_25351,N_20793,N_19183);
nor U25352 (N_25352,N_22545,N_19646);
and U25353 (N_25353,N_18228,N_22709);
and U25354 (N_25354,N_20817,N_18444);
xor U25355 (N_25355,N_21740,N_21316);
or U25356 (N_25356,N_20657,N_23113);
and U25357 (N_25357,N_21824,N_22248);
nor U25358 (N_25358,N_21805,N_19688);
and U25359 (N_25359,N_18358,N_18465);
or U25360 (N_25360,N_19931,N_18965);
or U25361 (N_25361,N_20409,N_21262);
xor U25362 (N_25362,N_19063,N_19648);
or U25363 (N_25363,N_20707,N_20628);
and U25364 (N_25364,N_19519,N_23738);
and U25365 (N_25365,N_19846,N_21991);
or U25366 (N_25366,N_19291,N_22915);
nor U25367 (N_25367,N_18963,N_22426);
nor U25368 (N_25368,N_20515,N_22182);
and U25369 (N_25369,N_19093,N_19355);
nand U25370 (N_25370,N_20299,N_18640);
xor U25371 (N_25371,N_23583,N_18149);
and U25372 (N_25372,N_22738,N_22222);
and U25373 (N_25373,N_21889,N_20885);
or U25374 (N_25374,N_20254,N_18415);
xor U25375 (N_25375,N_22618,N_23609);
nand U25376 (N_25376,N_19630,N_21631);
xor U25377 (N_25377,N_22404,N_18996);
nor U25378 (N_25378,N_23613,N_22264);
xor U25379 (N_25379,N_18671,N_18393);
nor U25380 (N_25380,N_20028,N_22726);
xor U25381 (N_25381,N_19146,N_23400);
nand U25382 (N_25382,N_19975,N_19109);
and U25383 (N_25383,N_19017,N_20904);
and U25384 (N_25384,N_21301,N_20493);
and U25385 (N_25385,N_21644,N_23292);
or U25386 (N_25386,N_21222,N_21025);
nor U25387 (N_25387,N_22489,N_18074);
and U25388 (N_25388,N_18431,N_21195);
nor U25389 (N_25389,N_23928,N_20578);
xnor U25390 (N_25390,N_21953,N_22022);
or U25391 (N_25391,N_23668,N_18945);
xor U25392 (N_25392,N_19700,N_20876);
and U25393 (N_25393,N_19475,N_21859);
and U25394 (N_25394,N_23159,N_19771);
nor U25395 (N_25395,N_23379,N_23072);
nor U25396 (N_25396,N_21347,N_23478);
xnor U25397 (N_25397,N_18669,N_23536);
and U25398 (N_25398,N_21201,N_21825);
and U25399 (N_25399,N_20203,N_20914);
and U25400 (N_25400,N_22477,N_23505);
and U25401 (N_25401,N_21275,N_22307);
nor U25402 (N_25402,N_23882,N_20745);
nand U25403 (N_25403,N_23228,N_20386);
xnor U25404 (N_25404,N_19825,N_18764);
nor U25405 (N_25405,N_22476,N_18350);
nor U25406 (N_25406,N_23682,N_21454);
or U25407 (N_25407,N_18122,N_23234);
nor U25408 (N_25408,N_21790,N_18716);
nand U25409 (N_25409,N_23665,N_20153);
nor U25410 (N_25410,N_22071,N_23984);
or U25411 (N_25411,N_19342,N_21147);
nand U25412 (N_25412,N_23458,N_22846);
or U25413 (N_25413,N_19422,N_19583);
nor U25414 (N_25414,N_20650,N_23034);
nor U25415 (N_25415,N_19670,N_20384);
xor U25416 (N_25416,N_19328,N_22312);
or U25417 (N_25417,N_21963,N_20047);
nor U25418 (N_25418,N_18735,N_18712);
and U25419 (N_25419,N_20760,N_22605);
and U25420 (N_25420,N_20166,N_19348);
or U25421 (N_25421,N_21302,N_23988);
and U25422 (N_25422,N_22981,N_23965);
nor U25423 (N_25423,N_21806,N_18595);
and U25424 (N_25424,N_18453,N_20061);
nor U25425 (N_25425,N_18726,N_20941);
nor U25426 (N_25426,N_20887,N_18826);
xnor U25427 (N_25427,N_18796,N_23376);
or U25428 (N_25428,N_23784,N_22629);
and U25429 (N_25429,N_22609,N_21521);
nor U25430 (N_25430,N_21434,N_19031);
and U25431 (N_25431,N_19107,N_22482);
nor U25432 (N_25432,N_18925,N_20723);
xnor U25433 (N_25433,N_21197,N_23619);
and U25434 (N_25434,N_23704,N_18733);
nor U25435 (N_25435,N_23895,N_22326);
nor U25436 (N_25436,N_21137,N_22458);
xor U25437 (N_25437,N_20344,N_23936);
nor U25438 (N_25438,N_19205,N_19561);
nand U25439 (N_25439,N_22237,N_18468);
and U25440 (N_25440,N_22792,N_21776);
xor U25441 (N_25441,N_18623,N_21464);
xor U25442 (N_25442,N_20913,N_23943);
and U25443 (N_25443,N_20470,N_22997);
and U25444 (N_25444,N_18197,N_22197);
nand U25445 (N_25445,N_22348,N_23967);
and U25446 (N_25446,N_21589,N_22567);
xor U25447 (N_25447,N_23500,N_22399);
nand U25448 (N_25448,N_18618,N_20506);
and U25449 (N_25449,N_19119,N_22619);
or U25450 (N_25450,N_20104,N_20851);
or U25451 (N_25451,N_21286,N_22500);
nor U25452 (N_25452,N_20856,N_20457);
and U25453 (N_25453,N_23452,N_22828);
nand U25454 (N_25454,N_22641,N_19620);
xnor U25455 (N_25455,N_18772,N_20489);
xnor U25456 (N_25456,N_19811,N_18184);
or U25457 (N_25457,N_23355,N_18430);
and U25458 (N_25458,N_18893,N_23155);
or U25459 (N_25459,N_19376,N_22276);
nor U25460 (N_25460,N_23632,N_21507);
and U25461 (N_25461,N_19334,N_23385);
nand U25462 (N_25462,N_22081,N_19745);
nand U25463 (N_25463,N_20593,N_23649);
and U25464 (N_25464,N_22127,N_18789);
and U25465 (N_25465,N_18660,N_18214);
or U25466 (N_25466,N_20960,N_19047);
xor U25467 (N_25467,N_22849,N_23678);
xnor U25468 (N_25468,N_19075,N_21708);
nand U25469 (N_25469,N_19575,N_18988);
nor U25470 (N_25470,N_19830,N_19719);
and U25471 (N_25471,N_18926,N_18449);
or U25472 (N_25472,N_23061,N_18246);
or U25473 (N_25473,N_19227,N_21310);
xnor U25474 (N_25474,N_18551,N_20233);
xnor U25475 (N_25475,N_21545,N_21561);
and U25476 (N_25476,N_22679,N_23161);
nand U25477 (N_25477,N_20785,N_18390);
and U25478 (N_25478,N_20055,N_23963);
nand U25479 (N_25479,N_19402,N_21977);
or U25480 (N_25480,N_19221,N_19427);
nand U25481 (N_25481,N_22582,N_21662);
nand U25482 (N_25482,N_23565,N_22102);
and U25483 (N_25483,N_19039,N_19873);
or U25484 (N_25484,N_20976,N_19088);
and U25485 (N_25485,N_21407,N_21544);
xor U25486 (N_25486,N_18491,N_20713);
xnor U25487 (N_25487,N_23959,N_20908);
or U25488 (N_25488,N_20095,N_23591);
xnor U25489 (N_25489,N_19973,N_23989);
and U25490 (N_25490,N_22948,N_18120);
and U25491 (N_25491,N_23468,N_22686);
or U25492 (N_25492,N_21784,N_21849);
xor U25493 (N_25493,N_20732,N_22931);
or U25494 (N_25494,N_18672,N_21674);
nor U25495 (N_25495,N_21929,N_19324);
or U25496 (N_25496,N_20661,N_19679);
nand U25497 (N_25497,N_23144,N_19169);
or U25498 (N_25498,N_20557,N_20862);
and U25499 (N_25499,N_20266,N_21754);
or U25500 (N_25500,N_23847,N_18281);
nand U25501 (N_25501,N_18774,N_18803);
or U25502 (N_25502,N_23304,N_21760);
nor U25503 (N_25503,N_23638,N_20670);
xnor U25504 (N_25504,N_21391,N_18546);
xnor U25505 (N_25505,N_23278,N_18145);
or U25506 (N_25506,N_22580,N_20286);
nand U25507 (N_25507,N_20631,N_19184);
nand U25508 (N_25508,N_20194,N_20145);
xor U25509 (N_25509,N_21594,N_21119);
or U25510 (N_25510,N_20008,N_22059);
nand U25511 (N_25511,N_21747,N_21655);
xnor U25512 (N_25512,N_20078,N_20212);
nand U25513 (N_25513,N_18056,N_22146);
and U25514 (N_25514,N_18873,N_22699);
nand U25515 (N_25515,N_22693,N_19585);
and U25516 (N_25516,N_22275,N_23743);
and U25517 (N_25517,N_23178,N_20555);
and U25518 (N_25518,N_20081,N_19680);
and U25519 (N_25519,N_23467,N_22043);
nand U25520 (N_25520,N_21553,N_18282);
nor U25521 (N_25521,N_20768,N_23246);
and U25522 (N_25522,N_18082,N_21379);
and U25523 (N_25523,N_19715,N_19820);
or U25524 (N_25524,N_20849,N_19742);
or U25525 (N_25525,N_22400,N_21331);
and U25526 (N_25526,N_19850,N_23932);
nand U25527 (N_25527,N_18935,N_18877);
xor U25528 (N_25528,N_18384,N_18950);
and U25529 (N_25529,N_19682,N_23437);
and U25530 (N_25530,N_23321,N_23744);
nor U25531 (N_25531,N_21023,N_22644);
nor U25532 (N_25532,N_18875,N_22324);
nor U25533 (N_25533,N_21129,N_23085);
nor U25534 (N_25534,N_18188,N_23185);
nor U25535 (N_25535,N_19738,N_23520);
nand U25536 (N_25536,N_23772,N_21574);
nand U25537 (N_25537,N_22896,N_18044);
xor U25538 (N_25538,N_19621,N_23944);
nand U25539 (N_25539,N_20893,N_23801);
xor U25540 (N_25540,N_23878,N_18317);
xnor U25541 (N_25541,N_21893,N_23703);
nor U25542 (N_25542,N_22623,N_21337);
and U25543 (N_25543,N_20549,N_21088);
xnor U25544 (N_25544,N_18037,N_23622);
nor U25545 (N_25545,N_18456,N_20780);
nand U25546 (N_25546,N_21077,N_23395);
nor U25547 (N_25547,N_23425,N_23340);
or U25548 (N_25548,N_23634,N_21800);
xor U25549 (N_25549,N_19921,N_22246);
and U25550 (N_25550,N_23753,N_23692);
and U25551 (N_25551,N_19014,N_21028);
and U25552 (N_25552,N_19432,N_19074);
nand U25553 (N_25553,N_18467,N_21345);
or U25554 (N_25554,N_19069,N_20458);
and U25555 (N_25555,N_22375,N_20582);
and U25556 (N_25556,N_19764,N_19022);
or U25557 (N_25557,N_18807,N_18591);
and U25558 (N_25558,N_19822,N_19416);
or U25559 (N_25559,N_19025,N_18533);
xor U25560 (N_25560,N_21292,N_20655);
nand U25561 (N_25561,N_22835,N_21761);
xnor U25562 (N_25562,N_19947,N_23238);
nor U25563 (N_25563,N_22844,N_21215);
xor U25564 (N_25564,N_22431,N_18645);
and U25565 (N_25565,N_20909,N_21103);
or U25566 (N_25566,N_18170,N_18295);
or U25567 (N_25567,N_23774,N_23539);
xor U25568 (N_25568,N_22494,N_18539);
nand U25569 (N_25569,N_19240,N_21832);
nand U25570 (N_25570,N_23411,N_22281);
and U25571 (N_25571,N_18647,N_21793);
nand U25572 (N_25572,N_22416,N_19577);
and U25573 (N_25573,N_22405,N_20001);
and U25574 (N_25574,N_22461,N_18096);
nand U25575 (N_25575,N_20601,N_21524);
or U25576 (N_25576,N_18856,N_20438);
and U25577 (N_25577,N_19997,N_19834);
nor U25578 (N_25578,N_21728,N_18901);
nor U25579 (N_25579,N_20301,N_21900);
xnor U25580 (N_25580,N_23265,N_22882);
nor U25581 (N_25581,N_21151,N_20412);
and U25582 (N_25582,N_20161,N_23874);
and U25583 (N_25583,N_22058,N_18268);
nor U25584 (N_25584,N_21843,N_18710);
or U25585 (N_25585,N_20155,N_18366);
nand U25586 (N_25586,N_21357,N_18532);
nor U25587 (N_25587,N_21196,N_22259);
or U25588 (N_25588,N_20919,N_21367);
nand U25589 (N_25589,N_22991,N_19220);
and U25590 (N_25590,N_21120,N_18676);
nor U25591 (N_25591,N_23510,N_19029);
xor U25592 (N_25592,N_22520,N_22323);
or U25593 (N_25593,N_22467,N_23281);
and U25594 (N_25594,N_22285,N_23099);
or U25595 (N_25595,N_18400,N_23066);
nor U25596 (N_25596,N_19860,N_22541);
xor U25597 (N_25597,N_19703,N_19226);
nor U25598 (N_25598,N_21642,N_20410);
xnor U25599 (N_25599,N_19133,N_23358);
and U25600 (N_25600,N_22452,N_20035);
or U25601 (N_25601,N_18140,N_21475);
xnor U25602 (N_25602,N_23020,N_19126);
xor U25603 (N_25603,N_22642,N_23232);
and U25604 (N_25604,N_18199,N_20416);
nand U25605 (N_25605,N_23599,N_21741);
nand U25606 (N_25606,N_20644,N_20251);
or U25607 (N_25607,N_21207,N_23875);
nand U25608 (N_25608,N_20875,N_20563);
nor U25609 (N_25609,N_20422,N_20583);
and U25610 (N_25610,N_22044,N_18238);
nand U25611 (N_25611,N_21012,N_18308);
nand U25612 (N_25612,N_22539,N_22779);
nand U25613 (N_25613,N_21015,N_20157);
or U25614 (N_25614,N_21309,N_19605);
nor U25615 (N_25615,N_23516,N_22799);
nor U25616 (N_25616,N_23759,N_21045);
and U25617 (N_25617,N_23818,N_19136);
nor U25618 (N_25618,N_22789,N_20623);
xnor U25619 (N_25619,N_22327,N_18581);
nor U25620 (N_25620,N_19623,N_21126);
or U25621 (N_25621,N_20584,N_22998);
and U25622 (N_25622,N_23821,N_20302);
nand U25623 (N_25623,N_18953,N_22444);
or U25624 (N_25624,N_22169,N_19782);
nor U25625 (N_25625,N_18360,N_20499);
nand U25626 (N_25626,N_21009,N_19156);
nand U25627 (N_25627,N_18981,N_21922);
nand U25628 (N_25628,N_22343,N_23115);
xor U25629 (N_25629,N_22511,N_22622);
xnor U25630 (N_25630,N_19774,N_19869);
and U25631 (N_25631,N_20526,N_22569);
nor U25632 (N_25632,N_22528,N_18569);
nor U25633 (N_25633,N_20935,N_21678);
or U25634 (N_25634,N_20943,N_20889);
nand U25635 (N_25635,N_21029,N_21994);
xnor U25636 (N_25636,N_20450,N_22831);
nor U25637 (N_25637,N_20225,N_22933);
nor U25638 (N_25638,N_22919,N_21836);
or U25639 (N_25639,N_22184,N_19683);
or U25640 (N_25640,N_22870,N_18651);
nor U25641 (N_25641,N_23239,N_20343);
nand U25642 (N_25642,N_19145,N_18636);
and U25643 (N_25643,N_19434,N_21141);
and U25644 (N_25644,N_19969,N_19859);
or U25645 (N_25645,N_21386,N_23389);
and U25646 (N_25646,N_18748,N_21705);
nor U25647 (N_25647,N_18280,N_20803);
nor U25648 (N_25648,N_21957,N_19748);
and U25649 (N_25649,N_23636,N_22957);
nand U25650 (N_25650,N_20839,N_21883);
or U25651 (N_25651,N_21499,N_19317);
xnor U25652 (N_25652,N_20463,N_22724);
xor U25653 (N_25653,N_21950,N_19858);
nand U25654 (N_25654,N_22445,N_23286);
nand U25655 (N_25655,N_23788,N_18028);
xnor U25656 (N_25656,N_21254,N_23043);
and U25657 (N_25657,N_21122,N_22174);
xor U25658 (N_25658,N_19049,N_22534);
and U25659 (N_25659,N_20955,N_18143);
or U25660 (N_25660,N_21489,N_20142);
nor U25661 (N_25661,N_22109,N_19327);
and U25662 (N_25662,N_22067,N_18615);
or U25663 (N_25663,N_23723,N_21469);
nor U25664 (N_25664,N_21942,N_23903);
nand U25665 (N_25665,N_23296,N_23176);
or U25666 (N_25666,N_18767,N_18250);
nand U25667 (N_25667,N_20547,N_19098);
or U25668 (N_25668,N_21938,N_23244);
and U25669 (N_25669,N_21163,N_22797);
xor U25670 (N_25670,N_20256,N_23760);
nor U25671 (N_25671,N_22862,N_19919);
nand U25672 (N_25672,N_19277,N_23802);
nor U25673 (N_25673,N_18363,N_20553);
and U25674 (N_25674,N_21145,N_21550);
xnor U25675 (N_25675,N_22716,N_23762);
nand U25676 (N_25676,N_23881,N_21833);
xnor U25677 (N_25677,N_19853,N_21467);
nand U25678 (N_25678,N_18419,N_22994);
xor U25679 (N_25679,N_20127,N_20456);
and U25680 (N_25680,N_19071,N_23667);
and U25681 (N_25681,N_22008,N_19021);
xor U25682 (N_25682,N_21393,N_19517);
and U25683 (N_25683,N_22123,N_22599);
or U25684 (N_25684,N_23044,N_21160);
xnor U25685 (N_25685,N_20108,N_22318);
or U25686 (N_25686,N_18972,N_20617);
nor U25687 (N_25687,N_19400,N_18682);
nor U25688 (N_25688,N_20348,N_19190);
or U25689 (N_25689,N_19885,N_18062);
and U25690 (N_25690,N_20536,N_23336);
or U25691 (N_25691,N_22655,N_20067);
nand U25692 (N_25692,N_19372,N_22660);
xnor U25693 (N_25693,N_23073,N_21198);
nor U25694 (N_25694,N_22621,N_18414);
or U25695 (N_25695,N_20014,N_23987);
nand U25696 (N_25696,N_21563,N_19393);
xor U25697 (N_25697,N_21176,N_23507);
or U25698 (N_25698,N_20838,N_23662);
xor U25699 (N_25699,N_19958,N_23007);
and U25700 (N_25700,N_22010,N_18014);
nand U25701 (N_25701,N_18270,N_23354);
xor U25702 (N_25702,N_22563,N_23351);
or U25703 (N_25703,N_19423,N_23051);
xnor U25704 (N_25704,N_18036,N_20080);
and U25705 (N_25705,N_18005,N_21069);
or U25706 (N_25706,N_23623,N_18154);
xor U25707 (N_25707,N_20144,N_22646);
or U25708 (N_25708,N_19783,N_19926);
nand U25709 (N_25709,N_22203,N_18750);
or U25710 (N_25710,N_19851,N_20397);
xnor U25711 (N_25711,N_19775,N_22077);
xnor U25712 (N_25712,N_22116,N_21484);
nand U25713 (N_25713,N_23826,N_18895);
xnor U25714 (N_25714,N_21956,N_23518);
xnor U25715 (N_25715,N_22560,N_18743);
xnor U25716 (N_25716,N_18916,N_18334);
nand U25717 (N_25717,N_23200,N_23433);
and U25718 (N_25718,N_22200,N_21356);
xor U25719 (N_25719,N_23811,N_19535);
or U25720 (N_25720,N_18649,N_21277);
and U25721 (N_25721,N_23872,N_21804);
or U25722 (N_25722,N_20735,N_21227);
or U25723 (N_25723,N_21996,N_21671);
nand U25724 (N_25724,N_22104,N_18711);
and U25725 (N_25725,N_19498,N_22624);
xor U25726 (N_25726,N_18171,N_23843);
xor U25727 (N_25727,N_21939,N_20637);
nor U25728 (N_25728,N_20702,N_20868);
or U25729 (N_25729,N_23690,N_21074);
nand U25730 (N_25730,N_22406,N_18940);
nor U25731 (N_25731,N_20195,N_19140);
and U25732 (N_25732,N_22053,N_22932);
or U25733 (N_25733,N_19791,N_22503);
and U25734 (N_25734,N_23456,N_23600);
nand U25735 (N_25735,N_22941,N_18146);
or U25736 (N_25736,N_18885,N_21853);
nand U25737 (N_25737,N_20071,N_23323);
nand U25738 (N_25738,N_21628,N_20300);
or U25739 (N_25739,N_23393,N_21128);
nand U25740 (N_25740,N_23911,N_23732);
xor U25741 (N_25741,N_18811,N_22145);
and U25742 (N_25742,N_19357,N_21384);
or U25743 (N_25743,N_21285,N_21852);
or U25744 (N_25744,N_20625,N_20965);
nor U25745 (N_25745,N_21768,N_21270);
and U25746 (N_25746,N_23417,N_18928);
nand U25747 (N_25747,N_22153,N_22076);
and U25748 (N_25748,N_20279,N_23892);
or U25749 (N_25749,N_23969,N_23616);
nand U25750 (N_25750,N_19203,N_19505);
xor U25751 (N_25751,N_23845,N_23293);
nand U25752 (N_25752,N_20403,N_19507);
or U25753 (N_25753,N_21491,N_23270);
xnor U25754 (N_25754,N_19957,N_21620);
nor U25755 (N_25755,N_21405,N_18365);
and U25756 (N_25756,N_19967,N_20043);
nand U25757 (N_25757,N_20180,N_22602);
or U25758 (N_25758,N_20415,N_22420);
xnor U25759 (N_25759,N_19757,N_21082);
nor U25760 (N_25760,N_23809,N_18840);
nand U25761 (N_25761,N_19172,N_21306);
and U25762 (N_25762,N_22019,N_23177);
and U25763 (N_25763,N_20531,N_20867);
nand U25764 (N_25764,N_21735,N_19840);
nor U25765 (N_25765,N_22604,N_21930);
and U25766 (N_25766,N_22337,N_18089);
nand U25767 (N_25767,N_22135,N_22088);
nor U25768 (N_25768,N_22301,N_18341);
xor U25769 (N_25769,N_19594,N_22772);
nand U25770 (N_25770,N_22517,N_18932);
or U25771 (N_25771,N_19836,N_22749);
nand U25772 (N_25772,N_18677,N_23180);
and U25773 (N_25773,N_19746,N_23089);
nor U25774 (N_25774,N_21798,N_18153);
xnor U25775 (N_25775,N_18432,N_21780);
xor U25776 (N_25776,N_19139,N_22368);
nor U25777 (N_25777,N_19323,N_23193);
and U25778 (N_25778,N_18429,N_20452);
nand U25779 (N_25779,N_22920,N_22544);
or U25780 (N_25780,N_23846,N_23359);
or U25781 (N_25781,N_22530,N_19928);
and U25782 (N_25782,N_21795,N_20915);
nand U25783 (N_25783,N_18752,N_21577);
nor U25784 (N_25784,N_21661,N_22759);
nor U25785 (N_25785,N_19891,N_23275);
and U25786 (N_25786,N_20265,N_22023);
and U25787 (N_25787,N_20619,N_18621);
or U25788 (N_25788,N_18095,N_23651);
and U25789 (N_25789,N_20460,N_23553);
or U25790 (N_25790,N_23117,N_19369);
nand U25791 (N_25791,N_21100,N_19349);
nor U25792 (N_25792,N_23808,N_21841);
nand U25793 (N_25793,N_23503,N_19596);
nand U25794 (N_25794,N_19953,N_21218);
or U25795 (N_25795,N_18580,N_21596);
and U25796 (N_25796,N_20324,N_21212);
or U25797 (N_25797,N_22115,N_20172);
nand U25798 (N_25798,N_18685,N_18176);
or U25799 (N_25799,N_18460,N_18876);
nand U25800 (N_25800,N_20748,N_19695);
nor U25801 (N_25801,N_21610,N_23466);
nor U25802 (N_25802,N_19785,N_18403);
and U25803 (N_25803,N_21424,N_19943);
and U25804 (N_25804,N_20435,N_20866);
or U25805 (N_25805,N_22970,N_20686);
or U25806 (N_25806,N_18723,N_19970);
nand U25807 (N_25807,N_19950,N_21068);
and U25808 (N_25808,N_23363,N_21531);
nand U25809 (N_25809,N_22733,N_18650);
xor U25810 (N_25810,N_18798,N_19215);
nor U25811 (N_25811,N_19297,N_21515);
nand U25812 (N_25812,N_22851,N_18686);
xnor U25813 (N_25813,N_23529,N_20287);
xnor U25814 (N_25814,N_19650,N_20903);
xor U25815 (N_25815,N_18516,N_18023);
and U25816 (N_25816,N_23934,N_20714);
nand U25817 (N_25817,N_18698,N_22034);
and U25818 (N_25818,N_22852,N_23914);
and U25819 (N_25819,N_19948,N_20346);
and U25820 (N_25820,N_20662,N_19356);
nor U25821 (N_25821,N_19831,N_18211);
and U25822 (N_25822,N_22413,N_20765);
xor U25823 (N_25823,N_20372,N_20923);
nand U25824 (N_25824,N_23250,N_20523);
nand U25825 (N_25825,N_20363,N_20729);
or U25826 (N_25826,N_23208,N_18222);
nor U25827 (N_25827,N_19540,N_19684);
and U25828 (N_25828,N_18126,N_21385);
and U25829 (N_25829,N_19167,N_22802);
and U25830 (N_25830,N_19191,N_23251);
nor U25831 (N_25831,N_23330,N_22266);
nor U25832 (N_25832,N_19010,N_22201);
xnor U25833 (N_25833,N_22265,N_21608);
xnor U25834 (N_25834,N_21549,N_18307);
nand U25835 (N_25835,N_20934,N_19697);
nor U25836 (N_25836,N_23779,N_20977);
or U25837 (N_25837,N_22367,N_21313);
nor U25838 (N_25838,N_20068,N_19414);
xnor U25839 (N_25839,N_23929,N_23775);
and U25840 (N_25840,N_21317,N_18164);
nor U25841 (N_25841,N_19481,N_20750);
nor U25842 (N_25842,N_22470,N_21341);
and U25843 (N_25843,N_23541,N_21773);
nor U25844 (N_25844,N_22355,N_21838);
nor U25845 (N_25845,N_21305,N_22761);
and U25846 (N_25846,N_21065,N_22574);
nor U25847 (N_25847,N_20162,N_21891);
and U25848 (N_25848,N_19138,N_21650);
nand U25849 (N_25849,N_19842,N_22472);
and U25850 (N_25850,N_19160,N_23556);
nor U25851 (N_25851,N_23727,N_21734);
nor U25852 (N_25852,N_18786,N_18695);
or U25853 (N_25853,N_22230,N_20806);
and U25854 (N_25854,N_23576,N_19196);
xnor U25855 (N_25855,N_20532,N_22647);
xnor U25856 (N_25856,N_19524,N_22247);
or U25857 (N_25857,N_22784,N_20795);
nand U25858 (N_25858,N_23055,N_18791);
or U25859 (N_25859,N_22360,N_18681);
and U25860 (N_25860,N_20453,N_22278);
nor U25861 (N_25861,N_18306,N_18831);
or U25862 (N_25862,N_21845,N_20019);
xor U25863 (N_25863,N_21696,N_23853);
nand U25864 (N_25864,N_23525,N_20754);
nand U25865 (N_25865,N_22868,N_18294);
nand U25866 (N_25866,N_22766,N_21388);
xnor U25867 (N_25867,N_18614,N_21787);
nor U25868 (N_25868,N_22055,N_18737);
and U25869 (N_25869,N_19813,N_22459);
nand U25870 (N_25870,N_19015,N_19533);
nor U25871 (N_25871,N_23038,N_22561);
nor U25872 (N_25872,N_19129,N_18519);
xnor U25873 (N_25873,N_18230,N_22254);
xor U25874 (N_25874,N_21511,N_18038);
xnor U25875 (N_25875,N_19295,N_18775);
xor U25876 (N_25876,N_21177,N_22362);
or U25877 (N_25877,N_21802,N_20032);
nor U25878 (N_25878,N_18175,N_19374);
or U25879 (N_25879,N_21621,N_23627);
nor U25880 (N_25880,N_23447,N_20766);
xor U25881 (N_25881,N_18638,N_18724);
or U25882 (N_25882,N_18590,N_18800);
xnor U25883 (N_25883,N_18624,N_19300);
and U25884 (N_25884,N_23540,N_23006);
xnor U25885 (N_25885,N_23065,N_21441);
and U25886 (N_25886,N_21368,N_19903);
and U25887 (N_25887,N_18994,N_20041);
nand U25888 (N_25888,N_21413,N_21246);
nand U25889 (N_25889,N_22875,N_19534);
and U25890 (N_25890,N_21580,N_21342);
xor U25891 (N_25891,N_21672,N_19586);
or U25892 (N_25892,N_19607,N_18461);
nand U25893 (N_25893,N_22519,N_20466);
nor U25894 (N_25894,N_20848,N_20709);
or U25895 (N_25895,N_19750,N_19280);
xor U25896 (N_25896,N_20827,N_23423);
nand U25897 (N_25897,N_20892,N_22617);
and U25898 (N_25898,N_19415,N_21493);
and U25899 (N_25899,N_23353,N_20988);
and U25900 (N_25900,N_18619,N_21054);
nand U25901 (N_25901,N_18824,N_19920);
and U25902 (N_25902,N_23283,N_20355);
and U25903 (N_25903,N_19035,N_18127);
nand U25904 (N_25904,N_21390,N_23710);
nor U25905 (N_25905,N_22164,N_20900);
nand U25906 (N_25906,N_20038,N_20859);
nand U25907 (N_25907,N_20755,N_20177);
or U25908 (N_25908,N_20701,N_19358);
nand U25909 (N_25909,N_18476,N_23474);
or U25910 (N_25910,N_23052,N_23689);
and U25911 (N_25911,N_19979,N_22745);
and U25912 (N_25912,N_20981,N_21528);
nor U25913 (N_25913,N_18413,N_22204);
nand U25914 (N_25914,N_20829,N_23070);
nand U25915 (N_25915,N_18552,N_19271);
xor U25916 (N_25916,N_18663,N_21969);
nand U25917 (N_25917,N_23997,N_18097);
xnor U25918 (N_25918,N_22430,N_19866);
nand U25919 (N_25919,N_20886,N_21685);
nand U25920 (N_25920,N_22433,N_21899);
xor U25921 (N_25921,N_22087,N_23230);
and U25922 (N_25922,N_21281,N_21557);
nor U25923 (N_25923,N_23050,N_21847);
and U25924 (N_25924,N_19379,N_18691);
nor U25925 (N_25925,N_18979,N_19401);
and U25926 (N_25926,N_22989,N_19003);
nor U25927 (N_25927,N_23162,N_21471);
or U25928 (N_25928,N_21691,N_21645);
nor U25929 (N_25929,N_22110,N_22730);
xor U25930 (N_25930,N_22270,N_21864);
nand U25931 (N_25931,N_22361,N_18922);
nand U25932 (N_25932,N_18408,N_22841);
nand U25933 (N_25933,N_18349,N_20196);
nor U25934 (N_25934,N_20858,N_23590);
and U25935 (N_25935,N_18083,N_19091);
nor U25936 (N_25936,N_20106,N_23873);
nand U25937 (N_25937,N_18424,N_20603);
xor U25938 (N_25938,N_18641,N_20883);
xnor U25939 (N_25939,N_22079,N_20860);
and U25940 (N_25940,N_20809,N_23179);
nand U25941 (N_25941,N_19875,N_20996);
and U25942 (N_25942,N_19556,N_23626);
nand U25943 (N_25943,N_21820,N_22890);
or U25944 (N_25944,N_23830,N_21435);
and U25945 (N_25945,N_22144,N_19984);
nand U25946 (N_25946,N_21020,N_21083);
nand U25947 (N_25947,N_21546,N_23140);
nor U25948 (N_25948,N_22685,N_23629);
nand U25949 (N_25949,N_21267,N_22711);
nand U25950 (N_25950,N_21307,N_20528);
and U25951 (N_25951,N_19756,N_22532);
nand U25952 (N_25952,N_22658,N_19553);
nor U25953 (N_25953,N_19488,N_18738);
nor U25954 (N_25954,N_19568,N_20461);
nor U25955 (N_25955,N_20580,N_20562);
nand U25956 (N_25956,N_19058,N_23822);
and U25957 (N_25957,N_20792,N_18917);
nor U25958 (N_25958,N_19479,N_21481);
and U25959 (N_25959,N_20733,N_21633);
and U25960 (N_25960,N_20819,N_20326);
or U25961 (N_25961,N_18042,N_23640);
or U25962 (N_25962,N_22592,N_18158);
or U25963 (N_25963,N_19696,N_18943);
xnor U25964 (N_25964,N_18816,N_19151);
nor U25965 (N_25965,N_22540,N_21556);
xnor U25966 (N_25966,N_23789,N_21813);
nor U25967 (N_25967,N_21131,N_21676);
and U25968 (N_25968,N_22384,N_18576);
xnor U25969 (N_25969,N_18962,N_19055);
and U25970 (N_25970,N_22783,N_22086);
nor U25971 (N_25971,N_21946,N_19283);
or U25972 (N_25972,N_23429,N_22465);
nor U25973 (N_25973,N_21104,N_21237);
and U25974 (N_25974,N_18290,N_19344);
or U25975 (N_25975,N_22283,N_23122);
xor U25976 (N_25976,N_23453,N_23676);
nand U25977 (N_25977,N_22864,N_23680);
xor U25978 (N_25978,N_20881,N_22479);
and U25979 (N_25979,N_19350,N_19051);
and U25980 (N_25980,N_21500,N_19543);
nand U25981 (N_25981,N_19706,N_19735);
xnor U25982 (N_25982,N_23068,N_20564);
nor U25983 (N_25983,N_18821,N_20147);
nor U25984 (N_25984,N_20854,N_23041);
or U25985 (N_25985,N_18167,N_19009);
nor U25986 (N_25986,N_20719,N_21935);
nor U25987 (N_25987,N_18780,N_21501);
xor U25988 (N_25988,N_18117,N_22340);
and U25989 (N_25989,N_18508,N_18024);
and U25990 (N_25990,N_21630,N_18142);
and U25991 (N_25991,N_22117,N_22787);
nor U25992 (N_25992,N_21421,N_23422);
and U25993 (N_25993,N_23637,N_22311);
or U25994 (N_25994,N_18355,N_22274);
nor U25995 (N_25995,N_21289,N_22913);
xor U25996 (N_25996,N_23905,N_18000);
and U25997 (N_25997,N_19166,N_23225);
nor U25998 (N_25998,N_22105,N_20005);
nand U25999 (N_25999,N_22978,N_20044);
nor U26000 (N_26000,N_20602,N_18486);
or U26001 (N_26001,N_22292,N_21652);
and U26002 (N_26002,N_18159,N_18684);
and U26003 (N_26003,N_21374,N_21323);
nand U26004 (N_26004,N_21071,N_21229);
and U26005 (N_26005,N_22049,N_20360);
xor U26006 (N_26006,N_19148,N_19185);
and U26007 (N_26007,N_20612,N_19473);
nor U26008 (N_26008,N_21607,N_18930);
xor U26009 (N_26009,N_23917,N_22160);
nor U26010 (N_26010,N_20040,N_19963);
nand U26011 (N_26011,N_21255,N_18567);
xor U26012 (N_26012,N_21348,N_18975);
xor U26013 (N_26013,N_21066,N_18864);
xnor U26014 (N_26014,N_18242,N_23492);
nand U26015 (N_26015,N_23694,N_22776);
or U26016 (N_26016,N_23404,N_23639);
xor U26017 (N_26017,N_18190,N_21697);
nand U26018 (N_26018,N_18233,N_23214);
nor U26019 (N_26019,N_23337,N_23956);
xor U26020 (N_26020,N_22891,N_22315);
or U26021 (N_26021,N_21109,N_21972);
or U26022 (N_26022,N_18076,N_23247);
and U26023 (N_26023,N_22555,N_23360);
and U26024 (N_26024,N_20705,N_22940);
and U26025 (N_26025,N_20978,N_19460);
nand U26026 (N_26026,N_18374,N_21821);
and U26027 (N_26027,N_23954,N_23186);
nand U26028 (N_26028,N_21884,N_19922);
nand U26029 (N_26029,N_20937,N_21276);
and U26030 (N_26030,N_23460,N_22821);
nor U26031 (N_26031,N_19439,N_21361);
xor U26032 (N_26032,N_23708,N_22193);
and U26033 (N_26033,N_21931,N_21770);
or U26034 (N_26034,N_23647,N_21920);
nand U26035 (N_26035,N_23080,N_22813);
or U26036 (N_26036,N_21495,N_20354);
xnor U26037 (N_26037,N_22536,N_23596);
nor U26038 (N_26038,N_21680,N_19456);
nor U26039 (N_26039,N_18324,N_19993);
xnor U26040 (N_26040,N_19117,N_18356);
nor U26041 (N_26041,N_23210,N_23831);
or U26042 (N_26042,N_20840,N_23836);
xnor U26043 (N_26043,N_21036,N_21819);
and U26044 (N_26044,N_18297,N_20761);
or U26045 (N_26045,N_22179,N_19182);
nand U26046 (N_26046,N_20003,N_22798);
nand U26047 (N_26047,N_22335,N_20998);
nor U26048 (N_26048,N_18181,N_22161);
or U26049 (N_26049,N_19384,N_20268);
xor U26050 (N_26050,N_20627,N_20352);
xor U26051 (N_26051,N_23287,N_23220);
nand U26052 (N_26052,N_23580,N_18092);
xnor U26053 (N_26053,N_22505,N_22015);
and U26054 (N_26054,N_18085,N_20119);
xor U26055 (N_26055,N_21731,N_23289);
or U26056 (N_26056,N_18568,N_22422);
and U26057 (N_26057,N_20964,N_20615);
or U26058 (N_26058,N_20762,N_22377);
xnor U26059 (N_26059,N_19204,N_22137);
nor U26060 (N_26060,N_18064,N_19843);
nor U26061 (N_26061,N_23010,N_18745);
and U26062 (N_26062,N_22282,N_23406);
nand U26063 (N_26063,N_18286,N_20070);
nor U26064 (N_26064,N_22888,N_21011);
nand U26065 (N_26065,N_21636,N_19115);
nand U26066 (N_26066,N_21562,N_23582);
or U26067 (N_26067,N_19502,N_21125);
nor U26068 (N_26068,N_23746,N_18047);
nor U26069 (N_26069,N_22403,N_22871);
xnor U26070 (N_26070,N_23352,N_18666);
or U26071 (N_26071,N_22017,N_21944);
nor U26072 (N_26072,N_20890,N_22228);
xor U26073 (N_26073,N_19147,N_18425);
nor U26074 (N_26074,N_19254,N_22354);
or U26075 (N_26075,N_19632,N_21041);
and U26076 (N_26076,N_21010,N_23970);
xnor U26077 (N_26077,N_19041,N_23862);
xnor U26078 (N_26078,N_19077,N_19636);
nand U26079 (N_26079,N_18938,N_21038);
nand U26080 (N_26080,N_20378,N_21378);
xor U26081 (N_26081,N_22988,N_18337);
nand U26082 (N_26082,N_19163,N_23980);
nand U26083 (N_26083,N_21442,N_22366);
and U26084 (N_26084,N_20262,N_20588);
nor U26085 (N_26085,N_23907,N_21614);
nor U26086 (N_26086,N_18178,N_21673);
or U26087 (N_26087,N_23854,N_20676);
nand U26088 (N_26088,N_23307,N_22934);
xnor U26089 (N_26089,N_19179,N_18496);
or U26090 (N_26090,N_21892,N_22857);
nand U26091 (N_26091,N_22706,N_20248);
nand U26092 (N_26092,N_23374,N_21558);
or U26093 (N_26093,N_22938,N_18457);
xnor U26094 (N_26094,N_23137,N_22676);
and U26095 (N_26095,N_20618,N_20743);
xor U26096 (N_26096,N_22218,N_21335);
nand U26097 (N_26097,N_22990,N_18689);
xnor U26098 (N_26098,N_22462,N_19386);
xnor U26099 (N_26099,N_19704,N_21540);
nor U26100 (N_26100,N_20518,N_23687);
and U26101 (N_26101,N_19526,N_23134);
or U26102 (N_26102,N_18048,N_21064);
or U26103 (N_26103,N_19702,N_22013);
or U26104 (N_26104,N_21359,N_21720);
and U26105 (N_26105,N_21311,N_23254);
xnor U26106 (N_26106,N_19918,N_21613);
and U26107 (N_26107,N_21888,N_18793);
or U26108 (N_26108,N_19008,N_22357);
nand U26109 (N_26109,N_19717,N_19234);
xnor U26110 (N_26110,N_19743,N_21185);
and U26111 (N_26111,N_22466,N_22765);
or U26112 (N_26112,N_20711,N_18160);
nor U26113 (N_26113,N_23077,N_21581);
xor U26114 (N_26114,N_18850,N_23173);
or U26115 (N_26115,N_21807,N_22084);
xor U26116 (N_26116,N_21375,N_23628);
nor U26117 (N_26117,N_19068,N_19894);
nand U26118 (N_26118,N_18736,N_20548);
nand U26119 (N_26119,N_23512,N_22887);
nand U26120 (N_26120,N_22986,N_18078);
and U26121 (N_26121,N_18478,N_20710);
or U26122 (N_26122,N_21076,N_20338);
nor U26123 (N_26123,N_19896,N_18021);
and U26124 (N_26124,N_22696,N_20973);
nor U26125 (N_26125,N_22478,N_21877);
nand U26126 (N_26126,N_21885,N_21133);
or U26127 (N_26127,N_20946,N_18207);
and U26128 (N_26128,N_19013,N_19425);
nor U26129 (N_26129,N_22740,N_20400);
nor U26130 (N_26130,N_23778,N_21777);
nand U26131 (N_26131,N_19197,N_23331);
and U26132 (N_26132,N_23076,N_19718);
nand U26133 (N_26133,N_19924,N_20706);
and U26134 (N_26134,N_22668,N_21879);
and U26135 (N_26135,N_22369,N_18272);
nor U26136 (N_26136,N_22961,N_19496);
xor U26137 (N_26137,N_22903,N_21923);
xnor U26138 (N_26138,N_19287,N_22855);
nor U26139 (N_26139,N_21993,N_18725);
or U26140 (N_26140,N_19927,N_20170);
or U26141 (N_26141,N_20810,N_18661);
nor U26142 (N_26142,N_19411,N_21132);
or U26143 (N_26143,N_20659,N_20143);
nand U26144 (N_26144,N_22790,N_18134);
xnor U26145 (N_26145,N_21399,N_23205);
and U26146 (N_26146,N_20979,N_19176);
nor U26147 (N_26147,N_23093,N_22437);
and U26148 (N_26148,N_23561,N_18918);
or U26149 (N_26149,N_19490,N_22256);
or U26150 (N_26150,N_21284,N_19027);
and U26151 (N_26151,N_23475,N_20031);
nor U26152 (N_26152,N_22094,N_19848);
and U26153 (N_26153,N_21504,N_19478);
and U26154 (N_26154,N_18863,N_21114);
and U26155 (N_26155,N_19971,N_18482);
and U26156 (N_26156,N_23262,N_23920);
nor U26157 (N_26157,N_22107,N_21315);
and U26158 (N_26158,N_22610,N_18983);
nand U26159 (N_26159,N_22216,N_21732);
or U26160 (N_26160,N_23897,N_23328);
and U26161 (N_26161,N_23725,N_19111);
and U26162 (N_26162,N_23495,N_22093);
nor U26163 (N_26163,N_21194,N_23011);
xnor U26164 (N_26164,N_19404,N_22106);
nand U26165 (N_26165,N_23734,N_22186);
nand U26166 (N_26166,N_20697,N_21997);
nor U26167 (N_26167,N_18838,N_22287);
nor U26168 (N_26168,N_18084,N_20799);
xor U26169 (N_26169,N_21049,N_23863);
nand U26170 (N_26170,N_21514,N_21401);
or U26171 (N_26171,N_21984,N_19135);
and U26172 (N_26172,N_20146,N_18788);
nor U26173 (N_26173,N_18991,N_23547);
nand U26174 (N_26174,N_18707,N_23749);
or U26175 (N_26175,N_20906,N_19445);
and U26176 (N_26176,N_20634,N_20942);
nand U26177 (N_26177,N_22447,N_22833);
nor U26178 (N_26178,N_21670,N_21519);
and U26179 (N_26179,N_22065,N_19110);
xor U26180 (N_26180,N_22603,N_22865);
or U26181 (N_26181,N_18329,N_18369);
nor U26182 (N_26182,N_21402,N_23660);
nor U26183 (N_26183,N_22215,N_23521);
or U26184 (N_26184,N_21894,N_18703);
nor U26185 (N_26185,N_20724,N_23030);
or U26186 (N_26186,N_19908,N_21799);
nor U26187 (N_26187,N_22329,N_20959);
or U26188 (N_26188,N_18375,N_18606);
nand U26189 (N_26189,N_23916,N_19611);
xor U26190 (N_26190,N_21654,N_22025);
or U26191 (N_26191,N_20314,N_21622);
nor U26192 (N_26192,N_19086,N_21455);
nand U26193 (N_26193,N_19030,N_20730);
and U26194 (N_26194,N_23975,N_22827);
xnor U26195 (N_26195,N_23621,N_22661);
xnor U26196 (N_26196,N_23957,N_21230);
or U26197 (N_26197,N_21668,N_19162);
and U26198 (N_26198,N_20368,N_20951);
nor U26199 (N_26199,N_23401,N_20213);
nand U26200 (N_26200,N_22746,N_20599);
or U26201 (N_26201,N_23297,N_19589);
or U26202 (N_26202,N_20843,N_22815);
or U26203 (N_26203,N_18147,N_21926);
and U26204 (N_26204,N_18302,N_23344);
and U26205 (N_26205,N_22576,N_20918);
or U26206 (N_26206,N_22769,N_19740);
xor U26207 (N_26207,N_19476,N_22196);
and U26208 (N_26208,N_21174,N_22720);
and U26209 (N_26209,N_22942,N_20487);
and U26210 (N_26210,N_23274,N_20243);
nand U26211 (N_26211,N_22832,N_19716);
or U26212 (N_26212,N_20789,N_18756);
nand U26213 (N_26213,N_20168,N_23722);
xor U26214 (N_26214,N_21637,N_18065);
xor U26215 (N_26215,N_19232,N_21166);
xnor U26216 (N_26216,N_20575,N_22134);
and U26217 (N_26217,N_22825,N_19974);
or U26218 (N_26218,N_22980,N_22496);
nor U26219 (N_26219,N_19515,N_20910);
xor U26220 (N_26220,N_20163,N_23489);
nand U26221 (N_26221,N_19982,N_21989);
and U26222 (N_26222,N_21921,N_18700);
nand U26223 (N_26223,N_19019,N_19952);
nand U26224 (N_26224,N_21354,N_18931);
and U26225 (N_26225,N_19177,N_20970);
or U26226 (N_26226,N_19681,N_19144);
or U26227 (N_26227,N_19674,N_21927);
and U26228 (N_26228,N_20120,N_21436);
and U26229 (N_26229,N_18277,N_18386);
nand U26230 (N_26230,N_23735,N_18545);
nor U26231 (N_26231,N_18218,N_21901);
nand U26232 (N_26232,N_22007,N_18784);
nor U26233 (N_26233,N_23773,N_22601);
nor U26234 (N_26234,N_23493,N_19960);
nand U26235 (N_26235,N_23439,N_21874);
and U26236 (N_26236,N_21572,N_18361);
nor U26237 (N_26237,N_19516,N_22611);
or U26238 (N_26238,N_18397,N_19712);
or U26239 (N_26239,N_20690,N_22527);
or U26240 (N_26240,N_22172,N_20210);
and U26241 (N_26241,N_23827,N_21175);
or U26242 (N_26242,N_22737,N_19509);
xor U26243 (N_26243,N_20775,N_22365);
and U26244 (N_26244,N_18274,N_21110);
or U26245 (N_26245,N_18607,N_19056);
nor U26246 (N_26246,N_22689,N_19559);
or U26247 (N_26247,N_18203,N_22165);
xor U26248 (N_26248,N_19615,N_21727);
and U26249 (N_26249,N_23686,N_22417);
and U26250 (N_26250,N_18473,N_20312);
nand U26251 (N_26251,N_19666,N_19725);
and U26252 (N_26252,N_21061,N_20689);
nor U26253 (N_26253,N_18708,N_21624);
nand U26254 (N_26254,N_20490,N_21848);
and U26255 (N_26255,N_23748,N_18344);
or U26256 (N_26256,N_19307,N_23496);
nor U26257 (N_26257,N_21371,N_19465);
xor U26258 (N_26258,N_19937,N_18124);
or U26259 (N_26259,N_20058,N_18949);
nand U26260 (N_26260,N_21373,N_23768);
and U26261 (N_26261,N_23776,N_19592);
or U26262 (N_26262,N_21480,N_22523);
xnor U26263 (N_26263,N_18558,N_19335);
and U26264 (N_26264,N_22507,N_18503);
nor U26265 (N_26265,N_23334,N_19435);
or U26266 (N_26266,N_22120,N_23064);
or U26267 (N_26267,N_20406,N_21684);
and U26268 (N_26268,N_22666,N_21575);
nor U26269 (N_26269,N_19180,N_19103);
xnor U26270 (N_26270,N_23714,N_23589);
or U26271 (N_26271,N_19708,N_20171);
nand U26272 (N_26272,N_19804,N_18549);
and U26273 (N_26273,N_21214,N_18447);
or U26274 (N_26274,N_22504,N_19012);
or U26275 (N_26275,N_20447,N_20576);
nor U26276 (N_26276,N_19318,N_18553);
nor U26277 (N_26277,N_21473,N_23992);
nor U26278 (N_26278,N_23203,N_18844);
xnor U26279 (N_26279,N_18236,N_21008);
nand U26280 (N_26280,N_23147,N_21765);
and U26281 (N_26281,N_18883,N_18570);
nand U26282 (N_26282,N_20566,N_19995);
nor U26283 (N_26283,N_19827,N_23902);
nand U26284 (N_26284,N_23107,N_23833);
nor U26285 (N_26285,N_21725,N_22952);
xnor U26286 (N_26286,N_20034,N_21003);
xnor U26287 (N_26287,N_23322,N_22295);
nor U26288 (N_26288,N_22163,N_20024);
xnor U26289 (N_26289,N_23612,N_23267);
or U26290 (N_26290,N_23986,N_19816);
nand U26291 (N_26291,N_19887,N_23285);
xor U26292 (N_26292,N_22245,N_23338);
nand U26293 (N_26293,N_20462,N_20764);
and U26294 (N_26294,N_22512,N_23841);
or U26295 (N_26295,N_20821,N_19252);
nand U26296 (N_26296,N_22018,N_19433);
nor U26297 (N_26297,N_23079,N_19101);
xor U26298 (N_26298,N_20790,N_22243);
or U26299 (N_26299,N_21917,N_23655);
xor U26300 (N_26300,N_18458,N_19281);
and U26301 (N_26301,N_18319,N_23737);
nand U26302 (N_26302,N_18326,N_23377);
xor U26303 (N_26303,N_22418,N_23371);
and U26304 (N_26304,N_19244,N_21502);
nor U26305 (N_26305,N_19593,N_18301);
nand U26306 (N_26306,N_19158,N_20610);
or U26307 (N_26307,N_18817,N_23035);
nand U26308 (N_26308,N_20381,N_20189);
nor U26309 (N_26309,N_20012,N_19510);
xnor U26310 (N_26310,N_19032,N_18136);
nand U26311 (N_26311,N_22474,N_22033);
nand U26312 (N_26312,N_18258,N_20060);
xnor U26313 (N_26313,N_23078,N_19986);
or U26314 (N_26314,N_18611,N_23163);
xor U26315 (N_26315,N_20116,N_23958);
or U26316 (N_26316,N_22050,N_22651);
nor U26317 (N_26317,N_21903,N_20199);
nor U26318 (N_26318,N_22554,N_18617);
nand U26319 (N_26319,N_19202,N_21979);
nor U26320 (N_26320,N_22390,N_20622);
nand U26321 (N_26321,N_21851,N_18213);
xor U26322 (N_26322,N_22578,N_18267);
and U26323 (N_26323,N_23199,N_20205);
or U26324 (N_26324,N_21221,N_19676);
xor U26325 (N_26325,N_20030,N_18589);
or U26326 (N_26326,N_19938,N_18732);
nand U26327 (N_26327,N_20311,N_18011);
nor U26328 (N_26328,N_23867,N_19828);
or U26329 (N_26329,N_19094,N_22568);
and U26330 (N_26330,N_22705,N_20782);
nand U26331 (N_26331,N_21039,N_21506);
nor U26332 (N_26332,N_23194,N_19264);
xor U26333 (N_26333,N_23219,N_20504);
or U26334 (N_26334,N_18704,N_22785);
and U26335 (N_26335,N_22878,N_22630);
nand U26336 (N_26336,N_18139,N_22181);
or U26337 (N_26337,N_21213,N_20869);
or U26338 (N_26338,N_18052,N_19692);
and U26339 (N_26339,N_21468,N_19591);
and U26340 (N_26340,N_22212,N_23981);
or U26341 (N_26341,N_23316,N_21602);
nor U26342 (N_26342,N_20837,N_23806);
or U26343 (N_26343,N_23588,N_21704);
nand U26344 (N_26344,N_23712,N_20574);
nand U26345 (N_26345,N_22060,N_19346);
and U26346 (N_26346,N_19155,N_23910);
nand U26347 (N_26347,N_20280,N_20079);
and U26348 (N_26348,N_18224,N_22739);
xnor U26349 (N_26349,N_22297,N_21370);
and U26350 (N_26350,N_22112,N_22675);
nor U26351 (N_26351,N_23388,N_19458);
nor U26352 (N_26352,N_23409,N_18888);
and U26353 (N_26353,N_18137,N_20252);
xnor U26354 (N_26354,N_19284,N_22414);
nand U26355 (N_26355,N_18435,N_20075);
and U26356 (N_26356,N_22484,N_18428);
and U26357 (N_26357,N_21107,N_23168);
nor U26358 (N_26358,N_23104,N_18559);
or U26359 (N_26359,N_22095,N_21320);
and U26360 (N_26360,N_19339,N_19686);
and U26361 (N_26361,N_22848,N_23951);
and U26362 (N_26362,N_22683,N_23372);
xor U26363 (N_26363,N_23184,N_21990);
nand U26364 (N_26364,N_20624,N_19819);
and U26365 (N_26365,N_18688,N_21004);
nor U26366 (N_26366,N_20940,N_23697);
or U26367 (N_26367,N_21943,N_23756);
and U26368 (N_26368,N_23717,N_22398);
nand U26369 (N_26369,N_21526,N_21138);
and U26370 (N_26370,N_22003,N_19090);
or U26371 (N_26371,N_20912,N_18664);
nor U26372 (N_26372,N_19562,N_22332);
or U26373 (N_26373,N_18652,N_21723);
nor U26374 (N_26374,N_20786,N_19807);
nand U26375 (N_26375,N_19564,N_18836);
and U26376 (N_26376,N_18129,N_20556);
xnor U26377 (N_26377,N_19360,N_22764);
nand U26378 (N_26378,N_19784,N_19092);
xnor U26379 (N_26379,N_23240,N_21273);
nand U26380 (N_26380,N_23731,N_23729);
nor U26381 (N_26381,N_21415,N_18759);
or U26382 (N_26382,N_18529,N_22298);
nor U26383 (N_26383,N_23851,N_18186);
and U26384 (N_26384,N_22673,N_19165);
xor U26385 (N_26385,N_19447,N_18992);
or U26386 (N_26386,N_22253,N_21829);
and U26387 (N_26387,N_23644,N_18881);
nor U26388 (N_26388,N_21372,N_21536);
nand U26389 (N_26389,N_19569,N_20802);
xor U26390 (N_26390,N_23814,N_22288);
xnor U26391 (N_26391,N_18474,N_22483);
nand U26392 (N_26392,N_23922,N_20861);
or U26393 (N_26393,N_23819,N_23308);
xnor U26394 (N_26394,N_21349,N_19810);
xor U26395 (N_26395,N_19251,N_19629);
xor U26396 (N_26396,N_18469,N_22659);
nor U26397 (N_26397,N_20607,N_19239);
or U26398 (N_26398,N_19872,N_22009);
xor U26399 (N_26399,N_22075,N_19453);
and U26400 (N_26400,N_23946,N_23876);
and U26401 (N_26401,N_21718,N_21318);
nor U26402 (N_26402,N_22217,N_18746);
nand U26403 (N_26403,N_19968,N_19613);
nor U26404 (N_26404,N_19087,N_23367);
or U26405 (N_26405,N_19779,N_19385);
nor U26406 (N_26406,N_18333,N_20022);
and U26407 (N_26407,N_21081,N_18327);
and U26408 (N_26408,N_22229,N_19929);
xor U26409 (N_26409,N_18410,N_21420);
nand U26410 (N_26410,N_22893,N_20587);
and U26411 (N_26411,N_21432,N_20124);
or U26412 (N_26412,N_19954,N_18845);
xnor U26413 (N_26413,N_20176,N_22291);
nor U26414 (N_26414,N_19200,N_19770);
nand U26415 (N_26415,N_23399,N_22777);
or U26416 (N_26416,N_19353,N_22175);
nor U26417 (N_26417,N_22960,N_22040);
xnor U26418 (N_26418,N_22538,N_18191);
nor U26419 (N_26419,N_22819,N_19395);
nand U26420 (N_26420,N_22955,N_18479);
and U26421 (N_26421,N_19444,N_22707);
and U26422 (N_26422,N_21569,N_23114);
or U26423 (N_26423,N_23953,N_20217);
xor U26424 (N_26424,N_20015,N_18216);
and U26425 (N_26425,N_18451,N_21928);
or U26426 (N_26426,N_23459,N_18604);
nand U26427 (N_26427,N_22162,N_22397);
and U26428 (N_26428,N_18278,N_23428);
and U26429 (N_26429,N_18989,N_21108);
xnor U26430 (N_26430,N_23771,N_23392);
nor U26431 (N_26431,N_19855,N_23950);
nor U26432 (N_26432,N_21079,N_20464);
or U26433 (N_26433,N_21295,N_21073);
nor U26434 (N_26434,N_18990,N_22364);
and U26435 (N_26435,N_22140,N_21448);
nor U26436 (N_26436,N_20944,N_18762);
or U26437 (N_26437,N_19268,N_22722);
or U26438 (N_26438,N_19761,N_20169);
xnor U26439 (N_26439,N_20477,N_22187);
nor U26440 (N_26440,N_20297,N_23090);
xor U26441 (N_26441,N_18325,N_18367);
xor U26442 (N_26442,N_22823,N_21019);
nor U26443 (N_26443,N_18459,N_19443);
nor U26444 (N_26444,N_19438,N_20508);
or U26445 (N_26445,N_18507,N_23143);
or U26446 (N_26446,N_20260,N_20483);
xor U26447 (N_26447,N_23455,N_19835);
or U26448 (N_26448,N_23982,N_21570);
and U26449 (N_26449,N_19778,N_19880);
xnor U26450 (N_26450,N_21664,N_22374);
or U26451 (N_26451,N_22542,N_21134);
or U26452 (N_26452,N_20589,N_18483);
nor U26453 (N_26453,N_23904,N_21870);
or U26454 (N_26454,N_21159,N_18264);
or U26455 (N_26455,N_21234,N_20294);
nand U26456 (N_26456,N_20791,N_23086);
nand U26457 (N_26457,N_19018,N_23477);
nor U26458 (N_26458,N_23769,N_22386);
nand U26459 (N_26459,N_18288,N_18524);
nor U26460 (N_26460,N_20568,N_22911);
xor U26461 (N_26461,N_20646,N_21591);
xnor U26462 (N_26462,N_23410,N_22884);
xnor U26463 (N_26463,N_20952,N_22583);
nand U26464 (N_26464,N_20831,N_19396);
nand U26465 (N_26465,N_22816,N_20674);
or U26466 (N_26466,N_19020,N_22131);
nor U26467 (N_26467,N_20158,N_18135);
nand U26468 (N_26468,N_18731,N_20398);
and U26469 (N_26469,N_20825,N_19289);
nand U26470 (N_26470,N_23961,N_18758);
and U26471 (N_26471,N_21136,N_18747);
and U26472 (N_26472,N_20891,N_18985);
nor U26473 (N_26473,N_23288,N_22330);
nand U26474 (N_26474,N_23170,N_20594);
nand U26475 (N_26475,N_20335,N_19428);
xor U26476 (N_26476,N_21294,N_20278);
xor U26477 (N_26477,N_19255,N_20336);
nor U26478 (N_26478,N_23387,N_22194);
and U26479 (N_26479,N_19734,N_18572);
nand U26480 (N_26480,N_23217,N_23218);
xor U26481 (N_26481,N_23653,N_20226);
nand U26482 (N_26482,N_19959,N_18760);
nand U26483 (N_26483,N_22490,N_23942);
xor U26484 (N_26484,N_20516,N_23572);
or U26485 (N_26485,N_21043,N_21050);
nor U26486 (N_26486,N_23948,N_22091);
nand U26487 (N_26487,N_18107,N_20926);
nand U26488 (N_26488,N_20249,N_23938);
nor U26489 (N_26489,N_23221,N_19645);
nand U26490 (N_26490,N_20852,N_21186);
or U26491 (N_26491,N_21660,N_19171);
and U26492 (N_26492,N_20968,N_20046);
nand U26493 (N_26493,N_19484,N_18936);
and U26494 (N_26494,N_22657,N_23432);
nand U26495 (N_26495,N_18741,N_19914);
and U26496 (N_26496,N_19034,N_20443);
nand U26497 (N_26497,N_20270,N_22286);
nor U26498 (N_26498,N_20342,N_18674);
and U26499 (N_26499,N_22495,N_21763);
or U26500 (N_26500,N_20535,N_22122);
nor U26501 (N_26501,N_22227,N_22118);
and U26502 (N_26502,N_18411,N_20994);
and U26503 (N_26503,N_19786,N_22755);
and U26504 (N_26504,N_19749,N_22455);
nand U26505 (N_26505,N_22943,N_21446);
nor U26506 (N_26506,N_18629,N_18426);
or U26507 (N_26507,N_23979,N_20673);
nor U26508 (N_26508,N_18133,N_23130);
or U26509 (N_26509,N_20502,N_23658);
nand U26510 (N_26510,N_20975,N_20570);
xnor U26511 (N_26511,N_22717,N_21766);
or U26512 (N_26512,N_22558,N_19394);
xor U26513 (N_26513,N_18466,N_18395);
xor U26514 (N_26514,N_18128,N_19525);
and U26515 (N_26515,N_20332,N_23671);
xnor U26516 (N_26516,N_20253,N_21964);
and U26517 (N_26517,N_22954,N_23339);
or U26518 (N_26518,N_22794,N_23535);
or U26519 (N_26519,N_22045,N_18536);
and U26520 (N_26520,N_19572,N_20016);
nand U26521 (N_26521,N_21261,N_20175);
or U26522 (N_26522,N_19485,N_23927);
and U26523 (N_26523,N_19590,N_22308);
nand U26524 (N_26524,N_23373,N_19617);
nand U26525 (N_26525,N_20091,N_21627);
nand U26526 (N_26526,N_19224,N_20552);
nor U26527 (N_26527,N_22817,N_23506);
and U26528 (N_26528,N_21260,N_23445);
or U26529 (N_26529,N_18464,N_21916);
and U26530 (N_26530,N_18727,N_21161);
nor U26531 (N_26531,N_19504,N_20214);
or U26532 (N_26532,N_18353,N_19194);
nor U26533 (N_26533,N_23684,N_22906);
and U26534 (N_26534,N_19600,N_22342);
or U26535 (N_26535,N_22692,N_20638);
xnor U26536 (N_26536,N_22627,N_20643);
or U26537 (N_26537,N_19134,N_22914);
nand U26538 (N_26538,N_19935,N_23165);
nand U26539 (N_26539,N_22190,N_20072);
or U26540 (N_26540,N_23380,N_21778);
nand U26541 (N_26541,N_22185,N_18405);
and U26542 (N_26542,N_18219,N_18485);
or U26543 (N_26543,N_21257,N_22667);
nand U26544 (N_26544,N_21525,N_21231);
or U26545 (N_26545,N_19809,N_18394);
xor U26546 (N_26546,N_23039,N_20173);
and U26547 (N_26547,N_21702,N_18438);
nand U26548 (N_26548,N_18510,N_19949);
nand U26549 (N_26549,N_21139,N_18879);
nor U26550 (N_26550,N_19378,N_21767);
and U26551 (N_26551,N_20731,N_20391);
xnor U26552 (N_26552,N_18561,N_23713);
nor U26553 (N_26553,N_18347,N_22310);
xor U26554 (N_26554,N_20521,N_18654);
or U26555 (N_26555,N_21803,N_20431);
nand U26556 (N_26556,N_21690,N_23160);
nor U26557 (N_26557,N_23886,N_21709);
xor U26558 (N_26558,N_21743,N_18125);
nand U26559 (N_26559,N_22522,N_18978);
or U26560 (N_26560,N_21084,N_19354);
xnor U26561 (N_26561,N_19153,N_23119);
nand U26562 (N_26562,N_19941,N_21324);
or U26563 (N_26563,N_19108,N_22811);
and U26564 (N_26564,N_18787,N_22412);
xnor U26565 (N_26565,N_21204,N_23538);
nor U26566 (N_26566,N_22457,N_22905);
and U26567 (N_26567,N_22909,N_21250);
nor U26568 (N_26568,N_19421,N_21748);
nand U26569 (N_26569,N_18138,N_20167);
nor U26570 (N_26570,N_20991,N_19512);
or U26571 (N_26571,N_22006,N_20125);
nor U26572 (N_26572,N_21856,N_21587);
xor U26573 (N_26573,N_23438,N_20995);
nor U26574 (N_26574,N_22100,N_23724);
and U26575 (N_26575,N_22824,N_18493);
nand U26576 (N_26576,N_21142,N_21123);
nor U26577 (N_26577,N_19951,N_18019);
xnor U26578 (N_26578,N_20437,N_23091);
nand U26579 (N_26579,N_22750,N_19653);
nor U26580 (N_26580,N_19201,N_22834);
xor U26581 (N_26581,N_19713,N_21387);
or U26582 (N_26582,N_23607,N_21224);
nor U26583 (N_26583,N_23106,N_21203);
nand U26584 (N_26584,N_22064,N_22262);
xnor U26585 (N_26585,N_23245,N_22068);
nand U26586 (N_26586,N_23555,N_19508);
xor U26587 (N_26587,N_18094,N_18342);
nand U26588 (N_26588,N_21679,N_22847);
nor U26589 (N_26589,N_19272,N_19159);
nor U26590 (N_26590,N_23537,N_20313);
and U26591 (N_26591,N_18331,N_21567);
nor U26592 (N_26592,N_19659,N_22877);
or U26593 (N_26593,N_22917,N_22643);
and U26594 (N_26594,N_20567,N_23369);
xor U26595 (N_26595,N_23253,N_21724);
and U26596 (N_26596,N_18874,N_21522);
nor U26597 (N_26597,N_18368,N_19758);
nor U26598 (N_26598,N_23257,N_20126);
or U26599 (N_26599,N_20454,N_18522);
xor U26600 (N_26600,N_23024,N_23259);
xnor U26601 (N_26601,N_22736,N_22487);
nor U26602 (N_26602,N_22898,N_19336);
nor U26603 (N_26603,N_21053,N_21669);
nand U26604 (N_26604,N_18683,N_19608);
and U26605 (N_26605,N_18564,N_19024);
and U26606 (N_26606,N_19741,N_21202);
nand U26607 (N_26607,N_23597,N_19902);
nand U26608 (N_26608,N_18305,N_22548);
or U26609 (N_26609,N_22951,N_23838);
or U26610 (N_26610,N_21366,N_20922);
nor U26611 (N_26611,N_18440,N_23440);
nand U26612 (N_26612,N_22514,N_18243);
or U26613 (N_26613,N_20818,N_21975);
nor U26614 (N_26614,N_23931,N_23574);
xor U26615 (N_26615,N_22735,N_23908);
nor U26616 (N_26616,N_23195,N_19768);
or U26617 (N_26617,N_19878,N_18715);
nor U26618 (N_26618,N_20421,N_22293);
nand U26619 (N_26619,N_18471,N_22649);
nor U26620 (N_26620,N_23869,N_21510);
nor U26621 (N_26621,N_22402,N_18009);
nor U26622 (N_26622,N_18020,N_21534);
nor U26623 (N_26623,N_19584,N_23937);
xor U26624 (N_26624,N_21632,N_21789);
xnor U26625 (N_26625,N_19554,N_23306);
nand U26626 (N_26626,N_22921,N_19520);
or U26627 (N_26627,N_23098,N_20272);
xnor U26628 (N_26628,N_23764,N_18899);
and U26629 (N_26629,N_21143,N_19579);
or U26630 (N_26630,N_23167,N_21497);
xnor U26631 (N_26631,N_22613,N_21682);
xor U26632 (N_26632,N_23810,N_22858);
and U26633 (N_26633,N_20261,N_22625);
nor U26634 (N_26634,N_23120,N_19529);
nand U26635 (N_26635,N_21380,N_18017);
nor U26636 (N_26636,N_18420,N_18501);
or U26637 (N_26637,N_20315,N_22415);
nand U26638 (N_26638,N_18229,N_23721);
nand U26639 (N_26639,N_19884,N_23592);
or U26640 (N_26640,N_21180,N_20880);
nor U26641 (N_26641,N_20320,N_21896);
xnor U26642 (N_26642,N_21710,N_21075);
nand U26643 (N_26643,N_19276,N_21014);
nor U26644 (N_26644,N_18550,N_23504);
nor U26645 (N_26645,N_18221,N_22385);
or U26646 (N_26646,N_21801,N_22062);
or U26647 (N_26647,N_23514,N_23021);
nand U26648 (N_26648,N_19059,N_21007);
and U26649 (N_26649,N_21978,N_23805);
or U26650 (N_26650,N_23384,N_19408);
or U26651 (N_26651,N_19210,N_21245);
or U26652 (N_26652,N_18494,N_23990);
nand U26653 (N_26653,N_19141,N_22290);
and U26654 (N_26654,N_18316,N_23642);
xor U26655 (N_26655,N_23256,N_21226);
xnor U26656 (N_26656,N_23407,N_22251);
and U26657 (N_26657,N_22341,N_20905);
nor U26658 (N_26658,N_18105,N_18192);
nand U26659 (N_26659,N_23426,N_23864);
xnor U26660 (N_26660,N_20527,N_18646);
and U26661 (N_26661,N_20954,N_19907);
and U26662 (N_26662,N_23828,N_18495);
xnor U26663 (N_26663,N_18412,N_23797);
nor U26664 (N_26664,N_23216,N_20600);
nor U26665 (N_26665,N_18497,N_21619);
nor U26666 (N_26666,N_19332,N_19933);
and U26667 (N_26667,N_21987,N_18837);
and U26668 (N_26668,N_20224,N_19616);
and U26669 (N_26669,N_22588,N_18648);
nor U26670 (N_26670,N_23804,N_22289);
xor U26671 (N_26671,N_20107,N_18976);
xnor U26672 (N_26672,N_20309,N_18544);
xor U26673 (N_26673,N_18827,N_19208);
nor U26674 (N_26674,N_21482,N_22257);
nand U26675 (N_26675,N_22151,N_21403);
and U26676 (N_26676,N_19288,N_23909);
nand U26677 (N_26677,N_19698,N_22531);
and U26678 (N_26678,N_19250,N_23015);
and U26679 (N_26679,N_22304,N_22681);
or U26680 (N_26680,N_23227,N_20776);
xnor U26681 (N_26681,N_19482,N_21463);
or U26682 (N_26682,N_22694,N_18008);
nand U26683 (N_26683,N_22648,N_21252);
and U26684 (N_26684,N_21485,N_18201);
nor U26685 (N_26685,N_19340,N_21154);
nand U26686 (N_26686,N_19417,N_19550);
nand U26687 (N_26687,N_22929,N_21034);
nor U26688 (N_26688,N_18610,N_21552);
nor U26689 (N_26689,N_18118,N_20488);
nor U26690 (N_26690,N_19225,N_18075);
or U26691 (N_26691,N_22876,N_21733);
xnor U26692 (N_26692,N_23483,N_22460);
nand U26693 (N_26693,N_21752,N_22300);
or U26694 (N_26694,N_19552,N_23261);
xor U26695 (N_26695,N_21013,N_23454);
nand U26696 (N_26696,N_23839,N_19371);
nand U26697 (N_26697,N_23470,N_21753);
nand U26698 (N_26698,N_22521,N_22678);
nand U26699 (N_26699,N_19337,N_22781);
and U26700 (N_26700,N_18869,N_19457);
nor U26701 (N_26701,N_22394,N_20430);
and U26702 (N_26702,N_19897,N_20716);
xor U26703 (N_26703,N_20473,N_23276);
xnor U26704 (N_26704,N_20232,N_19193);
and U26705 (N_26705,N_18045,N_21396);
and U26706 (N_26706,N_23755,N_20027);
xnor U26707 (N_26707,N_21124,N_19876);
and U26708 (N_26708,N_20330,N_22663);
and U26709 (N_26709,N_22967,N_21940);
or U26710 (N_26710,N_21611,N_23100);
or U26711 (N_26711,N_23382,N_19121);
nand U26712 (N_26712,N_21505,N_18060);
and U26713 (N_26713,N_21745,N_19955);
or U26714 (N_26714,N_21694,N_18006);
and U26715 (N_26715,N_23002,N_23973);
nor U26716 (N_26716,N_20329,N_20492);
nor U26717 (N_26717,N_22199,N_20084);
xnor U26718 (N_26718,N_18613,N_18530);
xor U26719 (N_26719,N_18260,N_18007);
xor U26720 (N_26720,N_19497,N_18189);
xor U26721 (N_26721,N_22635,N_19558);
nor U26722 (N_26722,N_22718,N_22939);
xor U26723 (N_26723,N_19278,N_18531);
and U26724 (N_26724,N_19364,N_18271);
nand U26725 (N_26725,N_20715,N_18644);
xnor U26726 (N_26726,N_22964,N_19413);
and U26727 (N_26727,N_22714,N_23681);
or U26728 (N_26728,N_18763,N_21866);
and U26729 (N_26729,N_20201,N_19137);
and U26730 (N_26730,N_22296,N_19381);
and U26731 (N_26731,N_23284,N_21474);
nor U26732 (N_26732,N_21542,N_20841);
or U26733 (N_26733,N_21750,N_18966);
xnor U26734 (N_26734,N_18448,N_23794);
xnor U26735 (N_26735,N_21582,N_20444);
or U26736 (N_26736,N_22972,N_22552);
and U26737 (N_26737,N_18111,N_20442);
nand U26738 (N_26738,N_20770,N_21149);
nand U26739 (N_26739,N_22268,N_19229);
nor U26740 (N_26740,N_20192,N_19899);
or U26741 (N_26741,N_20558,N_18894);
nor U26742 (N_26742,N_18969,N_18706);
nand U26743 (N_26743,N_23301,N_23390);
or U26744 (N_26744,N_22810,N_23486);
nor U26745 (N_26745,N_21298,N_20102);
nand U26746 (N_26746,N_21272,N_19824);
nand U26747 (N_26747,N_18609,N_21339);
nor U26748 (N_26748,N_23112,N_19797);
nand U26749 (N_26749,N_18781,N_23448);
or U26750 (N_26750,N_20691,N_20500);
nor U26751 (N_26751,N_22309,N_20894);
nand U26752 (N_26752,N_18910,N_18195);
and U26753 (N_26753,N_23484,N_20434);
and U26754 (N_26754,N_23152,N_20428);
xor U26755 (N_26755,N_20621,N_20371);
xnor U26756 (N_26756,N_21831,N_19178);
and U26757 (N_26757,N_23060,N_21717);
or U26758 (N_26758,N_19436,N_18929);
or U26759 (N_26759,N_22099,N_20380);
or U26760 (N_26760,N_23603,N_20307);
or U26761 (N_26761,N_23209,N_18070);
and U26762 (N_26762,N_23040,N_21427);
or U26763 (N_26763,N_23659,N_20334);
and U26764 (N_26764,N_19217,N_18015);
nand U26765 (N_26765,N_21430,N_18033);
and U26766 (N_26766,N_18971,N_22572);
xnor U26767 (N_26767,N_18534,N_22306);
nor U26768 (N_26768,N_21858,N_23858);
and U26769 (N_26769,N_22271,N_23273);
xor U26770 (N_26770,N_19301,N_20328);
nand U26771 (N_26771,N_19006,N_19070);
nand U26772 (N_26772,N_22225,N_19389);
and U26773 (N_26773,N_19181,N_22546);
and U26774 (N_26774,N_22910,N_19909);
or U26775 (N_26775,N_20895,N_21091);
nand U26776 (N_26776,N_20712,N_20772);
nor U26777 (N_26777,N_18152,N_22322);
and U26778 (N_26778,N_21248,N_20616);
and U26779 (N_26779,N_21726,N_23027);
xnor U26780 (N_26780,N_20198,N_21299);
xnor U26781 (N_26781,N_19249,N_19992);
or U26782 (N_26782,N_18418,N_19581);
xor U26783 (N_26783,N_20394,N_20357);
and U26784 (N_26784,N_19755,N_23698);
and U26785 (N_26785,N_21647,N_20240);
xnor U26786 (N_26786,N_21808,N_19506);
and U26787 (N_26787,N_21658,N_22677);
or U26788 (N_26788,N_21340,N_23993);
nor U26789 (N_26789,N_22562,N_21240);
xor U26790 (N_26790,N_19218,N_19377);
or U26791 (N_26791,N_19061,N_23900);
xnor U26792 (N_26792,N_19862,N_21425);
nor U26793 (N_26793,N_23834,N_23991);
and U26794 (N_26794,N_20208,N_20850);
or U26795 (N_26795,N_23434,N_21513);
nand U26796 (N_26796,N_19796,N_21625);
nor U26797 (N_26797,N_21786,N_21792);
or U26798 (N_26798,N_19521,N_20540);
nand U26799 (N_26799,N_18232,N_18718);
or U26800 (N_26800,N_23187,N_22801);
xnor U26801 (N_26801,N_18603,N_23033);
nor U26802 (N_26802,N_23625,N_23790);
and U26803 (N_26803,N_18063,N_18984);
and U26804 (N_26804,N_22922,N_18080);
or U26805 (N_26805,N_23133,N_22168);
and U26806 (N_26806,N_20651,N_18204);
and U26807 (N_26807,N_21788,N_18454);
nand U26808 (N_26808,N_22142,N_23188);
xnor U26809 (N_26809,N_23571,N_23464);
or U26810 (N_26810,N_19833,N_22438);
nand U26811 (N_26811,N_21886,N_22439);
and U26812 (N_26812,N_18266,N_22744);
nand U26813 (N_26813,N_20985,N_21897);
nor U26814 (N_26814,N_19626,N_23978);
xnor U26815 (N_26815,N_20573,N_23912);
nand U26816 (N_26816,N_20139,N_18823);
xnor U26817 (N_26817,N_21090,N_22240);
nand U26818 (N_26818,N_22866,N_18923);
and U26819 (N_26819,N_18215,N_19798);
nand U26820 (N_26820,N_18141,N_23370);
nand U26821 (N_26821,N_20174,N_18157);
xnor U26822 (N_26822,N_19477,N_18287);
or U26823 (N_26823,N_21269,N_20539);
or U26824 (N_26824,N_19365,N_21846);
xor U26825 (N_26825,N_19886,N_21362);
nand U26826 (N_26826,N_21667,N_23487);
xnor U26827 (N_26827,N_20884,N_19772);
nand U26828 (N_26828,N_18639,N_21601);
xor U26829 (N_26829,N_23325,N_23350);
xnor U26830 (N_26830,N_22258,N_20042);
and U26831 (N_26831,N_18884,N_18998);
and U26832 (N_26832,N_18777,N_18121);
or U26833 (N_26833,N_18043,N_22518);
or U26834 (N_26834,N_19011,N_22853);
or U26835 (N_26835,N_20284,N_21062);
nand U26836 (N_26836,N_23175,N_22753);
nor U26837 (N_26837,N_20269,N_22154);
or U26838 (N_26838,N_20140,N_20115);
nor U26839 (N_26839,N_23001,N_21488);
nand U26840 (N_26840,N_20982,N_20752);
and U26841 (N_26841,N_23568,N_22443);
and U26842 (N_26842,N_18252,N_19915);
xor U26843 (N_26843,N_22231,N_21818);
or U26844 (N_26844,N_23318,N_18348);
and U26845 (N_26845,N_19446,N_22198);
nor U26846 (N_26846,N_21312,N_19905);
xor U26847 (N_26847,N_19675,N_20396);
nor U26848 (N_26848,N_19235,N_18878);
nor U26849 (N_26849,N_23752,N_19305);
xnor U26850 (N_26850,N_18151,N_21626);
and U26851 (N_26851,N_22408,N_22809);
or U26852 (N_26852,N_19142,N_18662);
nand U26853 (N_26853,N_19461,N_22188);
nor U26854 (N_26854,N_18034,N_20524);
nand U26855 (N_26855,N_19483,N_20495);
or U26856 (N_26856,N_22595,N_23451);
nand U26857 (N_26857,N_23754,N_23608);
xor U26858 (N_26858,N_21828,N_20779);
and U26859 (N_26859,N_19765,N_20303);
and U26860 (N_26860,N_20992,N_19362);
or U26861 (N_26861,N_23436,N_18205);
or U26862 (N_26862,N_22159,N_21394);
and U26863 (N_26863,N_19994,N_20468);
nand U26864 (N_26864,N_22579,N_19426);
xor U26865 (N_26865,N_21496,N_20298);
and U26866 (N_26866,N_18657,N_20832);
nor U26867 (N_26867,N_23715,N_20215);
and U26868 (N_26868,N_21199,N_23630);
xnor U26869 (N_26869,N_18091,N_22121);
xor U26870 (N_26870,N_19188,N_18588);
nand U26871 (N_26871,N_19222,N_18407);
nor U26872 (N_26872,N_20317,N_23441);
xor U26873 (N_26873,N_19573,N_21431);
xor U26874 (N_26874,N_19242,N_23578);
nor U26875 (N_26875,N_21962,N_23901);
nor U26876 (N_26876,N_22028,N_23005);
nand U26877 (N_26877,N_19946,N_21352);
or U26878 (N_26878,N_23531,N_20258);
nand U26879 (N_26879,N_23793,N_20179);
or U26880 (N_26880,N_19883,N_19964);
nand U26881 (N_26881,N_23096,N_18088);
or U26882 (N_26882,N_23652,N_23543);
and U26883 (N_26883,N_20517,N_19838);
xnor U26884 (N_26884,N_19806,N_20911);
and U26885 (N_26885,N_19795,N_20509);
or U26886 (N_26886,N_19095,N_20846);
nand U26887 (N_26887,N_19294,N_21651);
and U26888 (N_26888,N_20063,N_20722);
nor U26889 (N_26889,N_20133,N_18114);
and U26890 (N_26890,N_21287,N_19890);
and U26891 (N_26891,N_21429,N_21659);
nand U26892 (N_26892,N_18077,N_22537);
nor U26893 (N_26893,N_19036,N_18040);
nand U26894 (N_26894,N_19261,N_22446);
nor U26895 (N_26895,N_19026,N_21330);
and U26896 (N_26896,N_23700,N_23960);
nor U26897 (N_26897,N_21400,N_22395);
and U26898 (N_26898,N_20664,N_19942);
xnor U26899 (N_26899,N_18999,N_20666);
and U26900 (N_26900,N_22944,N_23742);
xor U26901 (N_26901,N_21716,N_23026);
nor U26902 (N_26902,N_20665,N_19050);
nand U26903 (N_26903,N_23783,N_22434);
or U26904 (N_26904,N_21418,N_20237);
nand U26905 (N_26905,N_19118,N_23852);
nor U26906 (N_26906,N_19513,N_20961);
or U26907 (N_26907,N_20432,N_22454);
and U26908 (N_26908,N_20446,N_22850);
xor U26909 (N_26909,N_22725,N_18087);
xor U26910 (N_26910,N_19699,N_23059);
or U26911 (N_26911,N_23620,N_22557);
and U26912 (N_26912,N_18041,N_23966);
nor U26913 (N_26913,N_18890,N_22863);
nand U26914 (N_26914,N_18245,N_22421);
or U26915 (N_26915,N_23994,N_23126);
xnor U26916 (N_26916,N_23593,N_18585);
and U26917 (N_26917,N_23807,N_21965);
nor U26918 (N_26918,N_22208,N_21875);
or U26919 (N_26919,N_20388,N_21172);
or U26920 (N_26920,N_20050,N_21439);
nor U26921 (N_26921,N_23415,N_20190);
nor U26922 (N_26922,N_23695,N_21796);
and U26923 (N_26923,N_18634,N_19599);
nand U26924 (N_26924,N_23837,N_21113);
and U26925 (N_26925,N_22751,N_22125);
nand U26926 (N_26926,N_18434,N_22822);
nand U26927 (N_26927,N_18509,N_23517);
xor U26928 (N_26928,N_19080,N_22024);
or U26929 (N_26929,N_18957,N_23151);
and U26930 (N_26930,N_18637,N_19053);
xnor U26931 (N_26931,N_19549,N_21291);
xnor U26932 (N_26932,N_19001,N_19298);
or U26933 (N_26933,N_23491,N_19587);
or U26934 (N_26934,N_20808,N_20062);
xor U26935 (N_26935,N_20746,N_22551);
xor U26936 (N_26936,N_23522,N_18445);
nand U26937 (N_26937,N_20011,N_18346);
nand U26938 (N_26938,N_18592,N_21555);
xnor U26939 (N_26939,N_20036,N_20807);
and U26940 (N_26940,N_19687,N_22524);
xor U26941 (N_26941,N_22436,N_18161);
nand U26942 (N_26942,N_20347,N_23786);
and U26943 (N_26943,N_19539,N_21297);
and U26944 (N_26944,N_22687,N_21148);
xnor U26945 (N_26945,N_21835,N_21383);
nor U26946 (N_26946,N_20815,N_18352);
nand U26947 (N_26947,N_21094,N_18566);
and U26948 (N_26948,N_21982,N_23554);
and U26949 (N_26949,N_20541,N_23594);
xor U26950 (N_26950,N_21924,N_21721);
or U26951 (N_26951,N_18526,N_22597);
and U26952 (N_26952,N_22993,N_20882);
nand U26953 (N_26953,N_23083,N_19040);
xnor U26954 (N_26954,N_19571,N_19199);
nor U26955 (N_26955,N_20971,N_19449);
nor U26956 (N_26956,N_21508,N_22036);
and U26957 (N_26957,N_20082,N_19123);
and U26958 (N_26958,N_21719,N_19125);
xnor U26959 (N_26959,N_22996,N_22156);
and U26960 (N_26960,N_22021,N_21517);
nor U26961 (N_26961,N_23139,N_23513);
xnor U26962 (N_26962,N_21881,N_18026);
xnor U26963 (N_26963,N_19736,N_23923);
nand U26964 (N_26964,N_20641,N_22012);
or U26965 (N_26965,N_22754,N_22041);
nand U26966 (N_26966,N_20385,N_21713);
nand U26967 (N_26967,N_19228,N_20316);
xnor U26968 (N_26968,N_18253,N_23150);
xnor U26969 (N_26969,N_18851,N_18980);
nand U26970 (N_26970,N_21689,N_23883);
and U26971 (N_26971,N_22872,N_18771);
xor U26972 (N_26972,N_20481,N_20833);
or U26973 (N_26973,N_19663,N_20928);
nor U26974 (N_26974,N_20136,N_19265);
nand U26975 (N_26975,N_20367,N_22031);
and U26976 (N_26976,N_18582,N_18383);
xnor U26977 (N_26977,N_18081,N_23870);
xnor U26978 (N_26978,N_18323,N_21543);
or U26979 (N_26979,N_20364,N_22550);
nand U26980 (N_26980,N_21411,N_21868);
or U26981 (N_26981,N_20274,N_18202);
and U26982 (N_26982,N_22269,N_19640);
nand U26983 (N_26983,N_19642,N_20013);
nor U26984 (N_26984,N_20085,N_21739);
xor U26985 (N_26985,N_19285,N_22713);
nand U26986 (N_26986,N_19710,N_22221);
nand U26987 (N_26987,N_18263,N_19247);
and U26988 (N_26988,N_23019,N_20150);
nand U26989 (N_26989,N_19313,N_23394);
and U26990 (N_26990,N_22566,N_18388);
xor U26991 (N_26991,N_19522,N_20358);
nor U26992 (N_26992,N_18284,N_20356);
or U26993 (N_26993,N_22453,N_22565);
nor U26994 (N_26994,N_20255,N_20864);
nor U26995 (N_26995,N_18799,N_20092);
xnor U26996 (N_26996,N_23118,N_18680);
nand U26997 (N_26997,N_22982,N_20700);
and U26998 (N_26998,N_21085,N_23405);
nor U26999 (N_26999,N_18241,N_20099);
and U27000 (N_27000,N_21189,N_23555);
and U27001 (N_27001,N_22398,N_23809);
xor U27002 (N_27002,N_22683,N_23909);
nor U27003 (N_27003,N_21809,N_20525);
nor U27004 (N_27004,N_19940,N_23973);
xnor U27005 (N_27005,N_20356,N_20021);
nor U27006 (N_27006,N_19916,N_18258);
nand U27007 (N_27007,N_20924,N_20531);
or U27008 (N_27008,N_19784,N_22982);
and U27009 (N_27009,N_20045,N_21807);
and U27010 (N_27010,N_19145,N_18464);
xnor U27011 (N_27011,N_19377,N_20408);
nand U27012 (N_27012,N_21117,N_23207);
and U27013 (N_27013,N_21781,N_21416);
nor U27014 (N_27014,N_21438,N_21864);
and U27015 (N_27015,N_20960,N_23316);
xor U27016 (N_27016,N_19954,N_19732);
xor U27017 (N_27017,N_19559,N_23068);
nor U27018 (N_27018,N_22260,N_20862);
or U27019 (N_27019,N_23126,N_20321);
nand U27020 (N_27020,N_23164,N_20444);
nor U27021 (N_27021,N_21165,N_18169);
nand U27022 (N_27022,N_19938,N_19857);
and U27023 (N_27023,N_18192,N_21029);
nand U27024 (N_27024,N_23913,N_19617);
or U27025 (N_27025,N_21927,N_19533);
and U27026 (N_27026,N_19228,N_20567);
and U27027 (N_27027,N_20608,N_18835);
nor U27028 (N_27028,N_23577,N_19353);
and U27029 (N_27029,N_20147,N_21467);
xor U27030 (N_27030,N_18120,N_19936);
nor U27031 (N_27031,N_23223,N_23108);
xnor U27032 (N_27032,N_23460,N_18394);
xnor U27033 (N_27033,N_20837,N_18226);
xor U27034 (N_27034,N_20270,N_20774);
xor U27035 (N_27035,N_22757,N_19328);
nor U27036 (N_27036,N_21493,N_20828);
and U27037 (N_27037,N_18383,N_19714);
nand U27038 (N_27038,N_21183,N_19315);
nor U27039 (N_27039,N_21500,N_18814);
and U27040 (N_27040,N_19194,N_20426);
xor U27041 (N_27041,N_21659,N_19429);
nor U27042 (N_27042,N_23799,N_22084);
nor U27043 (N_27043,N_22174,N_21807);
or U27044 (N_27044,N_21731,N_18805);
and U27045 (N_27045,N_23173,N_23730);
nand U27046 (N_27046,N_21879,N_19744);
xor U27047 (N_27047,N_19676,N_23659);
and U27048 (N_27048,N_20338,N_18314);
xnor U27049 (N_27049,N_22090,N_23727);
and U27050 (N_27050,N_23912,N_23792);
nor U27051 (N_27051,N_20113,N_23133);
xor U27052 (N_27052,N_19767,N_21412);
or U27053 (N_27053,N_20171,N_23715);
and U27054 (N_27054,N_21703,N_19637);
nor U27055 (N_27055,N_22609,N_21124);
or U27056 (N_27056,N_23639,N_18620);
and U27057 (N_27057,N_19219,N_18483);
xor U27058 (N_27058,N_21213,N_22780);
and U27059 (N_27059,N_19789,N_19401);
nand U27060 (N_27060,N_22143,N_18140);
nor U27061 (N_27061,N_23348,N_19667);
nor U27062 (N_27062,N_20026,N_23999);
nand U27063 (N_27063,N_20339,N_22859);
or U27064 (N_27064,N_22686,N_20267);
nand U27065 (N_27065,N_19368,N_18923);
nor U27066 (N_27066,N_22035,N_18246);
nor U27067 (N_27067,N_21819,N_23187);
or U27068 (N_27068,N_23957,N_20990);
nor U27069 (N_27069,N_18264,N_23498);
xnor U27070 (N_27070,N_18832,N_22476);
nand U27071 (N_27071,N_23603,N_19760);
nand U27072 (N_27072,N_23587,N_19851);
and U27073 (N_27073,N_22339,N_23673);
nand U27074 (N_27074,N_23384,N_21144);
nor U27075 (N_27075,N_21884,N_19207);
or U27076 (N_27076,N_19609,N_23739);
or U27077 (N_27077,N_22810,N_19934);
and U27078 (N_27078,N_19395,N_21689);
nand U27079 (N_27079,N_18469,N_20595);
nor U27080 (N_27080,N_19831,N_20540);
or U27081 (N_27081,N_18377,N_20202);
nor U27082 (N_27082,N_18128,N_18964);
nand U27083 (N_27083,N_22897,N_21697);
nor U27084 (N_27084,N_23181,N_20308);
nor U27085 (N_27085,N_18248,N_22944);
xnor U27086 (N_27086,N_18687,N_22426);
xor U27087 (N_27087,N_19931,N_22083);
xnor U27088 (N_27088,N_20948,N_23740);
and U27089 (N_27089,N_23338,N_18878);
and U27090 (N_27090,N_23919,N_22150);
nor U27091 (N_27091,N_23559,N_19143);
or U27092 (N_27092,N_23367,N_22374);
and U27093 (N_27093,N_19018,N_18916);
or U27094 (N_27094,N_23842,N_21992);
nor U27095 (N_27095,N_21363,N_18364);
nor U27096 (N_27096,N_19690,N_21811);
or U27097 (N_27097,N_22491,N_19402);
nand U27098 (N_27098,N_23077,N_19442);
nor U27099 (N_27099,N_23703,N_23687);
nor U27100 (N_27100,N_19095,N_19939);
xor U27101 (N_27101,N_22048,N_22906);
and U27102 (N_27102,N_23441,N_22426);
nand U27103 (N_27103,N_18301,N_20946);
nand U27104 (N_27104,N_19982,N_21197);
xnor U27105 (N_27105,N_20871,N_20747);
nor U27106 (N_27106,N_21007,N_18451);
and U27107 (N_27107,N_21247,N_22693);
nor U27108 (N_27108,N_22136,N_23575);
nand U27109 (N_27109,N_18367,N_18970);
nand U27110 (N_27110,N_18720,N_18736);
nor U27111 (N_27111,N_20076,N_21616);
xor U27112 (N_27112,N_20679,N_21612);
nor U27113 (N_27113,N_23509,N_21817);
xor U27114 (N_27114,N_21629,N_23924);
xnor U27115 (N_27115,N_23816,N_23774);
nand U27116 (N_27116,N_18348,N_22077);
or U27117 (N_27117,N_22860,N_21974);
nand U27118 (N_27118,N_22510,N_21030);
or U27119 (N_27119,N_21492,N_18942);
nand U27120 (N_27120,N_18151,N_19199);
nor U27121 (N_27121,N_21749,N_19810);
and U27122 (N_27122,N_21948,N_23274);
or U27123 (N_27123,N_21833,N_23517);
nand U27124 (N_27124,N_22563,N_18096);
nor U27125 (N_27125,N_18340,N_23485);
and U27126 (N_27126,N_19608,N_20090);
nand U27127 (N_27127,N_22699,N_21951);
nor U27128 (N_27128,N_22361,N_23938);
or U27129 (N_27129,N_21097,N_20397);
nor U27130 (N_27130,N_19068,N_22407);
nor U27131 (N_27131,N_18917,N_18904);
and U27132 (N_27132,N_20217,N_18836);
nor U27133 (N_27133,N_22126,N_20129);
nand U27134 (N_27134,N_19712,N_18387);
and U27135 (N_27135,N_21531,N_18399);
nand U27136 (N_27136,N_19397,N_21072);
nor U27137 (N_27137,N_21211,N_20646);
xor U27138 (N_27138,N_20610,N_18222);
and U27139 (N_27139,N_21597,N_23972);
xnor U27140 (N_27140,N_21291,N_21020);
nand U27141 (N_27141,N_22484,N_18018);
nand U27142 (N_27142,N_22252,N_20464);
and U27143 (N_27143,N_21451,N_19063);
and U27144 (N_27144,N_18809,N_18052);
xor U27145 (N_27145,N_21755,N_20045);
nand U27146 (N_27146,N_21773,N_18877);
xnor U27147 (N_27147,N_22133,N_19188);
and U27148 (N_27148,N_23785,N_18718);
nor U27149 (N_27149,N_20630,N_22731);
xnor U27150 (N_27150,N_21190,N_20183);
xor U27151 (N_27151,N_20504,N_20935);
nor U27152 (N_27152,N_22553,N_20011);
nor U27153 (N_27153,N_21638,N_19231);
nor U27154 (N_27154,N_19923,N_21086);
or U27155 (N_27155,N_19583,N_22616);
nand U27156 (N_27156,N_18046,N_23778);
and U27157 (N_27157,N_20595,N_21962);
nor U27158 (N_27158,N_19939,N_19292);
or U27159 (N_27159,N_20066,N_18642);
nand U27160 (N_27160,N_22610,N_23856);
nand U27161 (N_27161,N_19277,N_18881);
and U27162 (N_27162,N_23878,N_21496);
and U27163 (N_27163,N_22579,N_20568);
xnor U27164 (N_27164,N_22662,N_18606);
xnor U27165 (N_27165,N_19405,N_21746);
and U27166 (N_27166,N_20889,N_19921);
and U27167 (N_27167,N_18590,N_21081);
and U27168 (N_27168,N_23525,N_22900);
nor U27169 (N_27169,N_23241,N_22888);
xor U27170 (N_27170,N_23937,N_18138);
or U27171 (N_27171,N_20307,N_20219);
or U27172 (N_27172,N_18071,N_18097);
and U27173 (N_27173,N_22234,N_20998);
nand U27174 (N_27174,N_18783,N_19131);
xor U27175 (N_27175,N_19921,N_19193);
nand U27176 (N_27176,N_22426,N_23185);
nor U27177 (N_27177,N_19407,N_19212);
or U27178 (N_27178,N_20451,N_20637);
nor U27179 (N_27179,N_19662,N_19794);
xor U27180 (N_27180,N_22830,N_21984);
and U27181 (N_27181,N_20345,N_21355);
and U27182 (N_27182,N_19509,N_22158);
nand U27183 (N_27183,N_22619,N_18584);
nand U27184 (N_27184,N_20059,N_22801);
and U27185 (N_27185,N_23235,N_20557);
xor U27186 (N_27186,N_23852,N_18814);
nand U27187 (N_27187,N_22271,N_23610);
nand U27188 (N_27188,N_20286,N_23952);
xor U27189 (N_27189,N_22859,N_20797);
nand U27190 (N_27190,N_22769,N_21725);
and U27191 (N_27191,N_21684,N_18404);
or U27192 (N_27192,N_19554,N_18884);
xor U27193 (N_27193,N_22228,N_18230);
xnor U27194 (N_27194,N_23997,N_19684);
nor U27195 (N_27195,N_19931,N_22654);
and U27196 (N_27196,N_21256,N_19788);
xnor U27197 (N_27197,N_23418,N_20666);
and U27198 (N_27198,N_19042,N_21212);
xor U27199 (N_27199,N_23378,N_18258);
xor U27200 (N_27200,N_21193,N_21035);
xnor U27201 (N_27201,N_18941,N_21429);
xnor U27202 (N_27202,N_21325,N_19617);
nand U27203 (N_27203,N_20375,N_21563);
xor U27204 (N_27204,N_20174,N_23136);
nand U27205 (N_27205,N_20699,N_21242);
xor U27206 (N_27206,N_19795,N_23996);
nor U27207 (N_27207,N_23117,N_23674);
xnor U27208 (N_27208,N_23931,N_21743);
nor U27209 (N_27209,N_22648,N_22230);
xor U27210 (N_27210,N_21810,N_18225);
nand U27211 (N_27211,N_19180,N_20919);
xnor U27212 (N_27212,N_23622,N_22770);
and U27213 (N_27213,N_20229,N_22432);
xnor U27214 (N_27214,N_19348,N_21250);
and U27215 (N_27215,N_22675,N_22965);
and U27216 (N_27216,N_23595,N_18313);
xor U27217 (N_27217,N_19750,N_21359);
nor U27218 (N_27218,N_20525,N_18882);
nor U27219 (N_27219,N_21072,N_18434);
nand U27220 (N_27220,N_22604,N_18787);
and U27221 (N_27221,N_20644,N_21840);
nor U27222 (N_27222,N_18463,N_21249);
or U27223 (N_27223,N_22424,N_19991);
or U27224 (N_27224,N_22747,N_20425);
or U27225 (N_27225,N_23780,N_19458);
or U27226 (N_27226,N_18009,N_22552);
nand U27227 (N_27227,N_20399,N_21568);
and U27228 (N_27228,N_18627,N_20551);
and U27229 (N_27229,N_18470,N_19723);
or U27230 (N_27230,N_21146,N_22046);
or U27231 (N_27231,N_20222,N_21882);
nor U27232 (N_27232,N_20268,N_20058);
nand U27233 (N_27233,N_19510,N_20279);
nand U27234 (N_27234,N_18220,N_19971);
nor U27235 (N_27235,N_19657,N_22206);
or U27236 (N_27236,N_18519,N_23278);
nor U27237 (N_27237,N_22477,N_22634);
nor U27238 (N_27238,N_19985,N_21829);
or U27239 (N_27239,N_23743,N_22251);
nor U27240 (N_27240,N_22872,N_18192);
or U27241 (N_27241,N_21503,N_18816);
nand U27242 (N_27242,N_20144,N_20264);
nor U27243 (N_27243,N_18334,N_21706);
nor U27244 (N_27244,N_22608,N_20777);
or U27245 (N_27245,N_19067,N_22934);
or U27246 (N_27246,N_18347,N_22426);
nor U27247 (N_27247,N_22110,N_22233);
xor U27248 (N_27248,N_22636,N_23381);
or U27249 (N_27249,N_22931,N_21179);
nand U27250 (N_27250,N_23117,N_18868);
nand U27251 (N_27251,N_23228,N_22989);
xor U27252 (N_27252,N_21960,N_22922);
xnor U27253 (N_27253,N_19259,N_18163);
nor U27254 (N_27254,N_20631,N_23076);
and U27255 (N_27255,N_19299,N_21964);
nand U27256 (N_27256,N_19168,N_23417);
or U27257 (N_27257,N_21520,N_19236);
and U27258 (N_27258,N_19785,N_23808);
nor U27259 (N_27259,N_22401,N_22231);
and U27260 (N_27260,N_18024,N_23932);
nand U27261 (N_27261,N_21755,N_18394);
or U27262 (N_27262,N_19234,N_18057);
nor U27263 (N_27263,N_21868,N_22384);
and U27264 (N_27264,N_18030,N_20145);
nor U27265 (N_27265,N_20189,N_22981);
nor U27266 (N_27266,N_19058,N_21766);
nand U27267 (N_27267,N_23260,N_18588);
nor U27268 (N_27268,N_19169,N_20565);
xor U27269 (N_27269,N_21923,N_20417);
or U27270 (N_27270,N_20898,N_23858);
nor U27271 (N_27271,N_20148,N_21105);
nor U27272 (N_27272,N_23724,N_23347);
and U27273 (N_27273,N_23925,N_21109);
nor U27274 (N_27274,N_20360,N_20230);
and U27275 (N_27275,N_20582,N_21987);
nor U27276 (N_27276,N_20348,N_21586);
nand U27277 (N_27277,N_18808,N_21464);
or U27278 (N_27278,N_22069,N_18405);
xnor U27279 (N_27279,N_20993,N_20086);
nor U27280 (N_27280,N_18431,N_21423);
or U27281 (N_27281,N_18531,N_22011);
nand U27282 (N_27282,N_19962,N_18861);
nand U27283 (N_27283,N_23808,N_18795);
nand U27284 (N_27284,N_19336,N_21316);
xor U27285 (N_27285,N_18937,N_23348);
xnor U27286 (N_27286,N_21540,N_22932);
nand U27287 (N_27287,N_22832,N_20965);
nor U27288 (N_27288,N_19778,N_23469);
xor U27289 (N_27289,N_20243,N_23849);
xnor U27290 (N_27290,N_20452,N_18039);
nor U27291 (N_27291,N_23657,N_22097);
nor U27292 (N_27292,N_21722,N_23664);
or U27293 (N_27293,N_21799,N_20698);
and U27294 (N_27294,N_19901,N_23039);
and U27295 (N_27295,N_18792,N_23144);
xnor U27296 (N_27296,N_23524,N_19482);
nor U27297 (N_27297,N_18541,N_18954);
nand U27298 (N_27298,N_18505,N_19781);
nand U27299 (N_27299,N_23666,N_22566);
nor U27300 (N_27300,N_19600,N_19506);
or U27301 (N_27301,N_19125,N_23520);
xor U27302 (N_27302,N_22421,N_21662);
nor U27303 (N_27303,N_23395,N_23342);
nor U27304 (N_27304,N_22869,N_19349);
xnor U27305 (N_27305,N_23230,N_22558);
or U27306 (N_27306,N_20063,N_21883);
and U27307 (N_27307,N_23474,N_20660);
and U27308 (N_27308,N_20773,N_20946);
nand U27309 (N_27309,N_22888,N_19289);
nor U27310 (N_27310,N_19491,N_20775);
xor U27311 (N_27311,N_19815,N_23170);
nand U27312 (N_27312,N_19298,N_19373);
or U27313 (N_27313,N_19821,N_21658);
or U27314 (N_27314,N_22187,N_21324);
nor U27315 (N_27315,N_21124,N_23452);
xnor U27316 (N_27316,N_23440,N_19140);
nand U27317 (N_27317,N_22474,N_18639);
and U27318 (N_27318,N_19093,N_21186);
and U27319 (N_27319,N_23679,N_22618);
and U27320 (N_27320,N_20742,N_18051);
and U27321 (N_27321,N_22171,N_23241);
and U27322 (N_27322,N_22417,N_21821);
xnor U27323 (N_27323,N_18916,N_18532);
xnor U27324 (N_27324,N_19334,N_19734);
nor U27325 (N_27325,N_19340,N_19316);
nor U27326 (N_27326,N_22990,N_22605);
xor U27327 (N_27327,N_20151,N_20503);
nor U27328 (N_27328,N_18471,N_21630);
and U27329 (N_27329,N_22750,N_19029);
xnor U27330 (N_27330,N_20934,N_22627);
nor U27331 (N_27331,N_18385,N_20345);
or U27332 (N_27332,N_23985,N_18600);
or U27333 (N_27333,N_23922,N_18489);
nor U27334 (N_27334,N_19409,N_21474);
nand U27335 (N_27335,N_22354,N_20427);
and U27336 (N_27336,N_22880,N_23004);
or U27337 (N_27337,N_20875,N_21957);
and U27338 (N_27338,N_22263,N_23017);
xnor U27339 (N_27339,N_19122,N_20705);
nor U27340 (N_27340,N_21375,N_21728);
xor U27341 (N_27341,N_18417,N_22867);
nand U27342 (N_27342,N_18927,N_19591);
nand U27343 (N_27343,N_22513,N_18728);
and U27344 (N_27344,N_22614,N_18372);
or U27345 (N_27345,N_21983,N_22825);
or U27346 (N_27346,N_21132,N_20636);
and U27347 (N_27347,N_22761,N_22031);
or U27348 (N_27348,N_20007,N_21174);
or U27349 (N_27349,N_18429,N_22515);
and U27350 (N_27350,N_19178,N_20144);
nor U27351 (N_27351,N_22687,N_23119);
and U27352 (N_27352,N_23233,N_19960);
nor U27353 (N_27353,N_19442,N_21221);
nor U27354 (N_27354,N_21329,N_19583);
nor U27355 (N_27355,N_23291,N_20340);
xnor U27356 (N_27356,N_23781,N_22099);
nand U27357 (N_27357,N_18114,N_21761);
nor U27358 (N_27358,N_18927,N_23195);
nor U27359 (N_27359,N_21159,N_21351);
and U27360 (N_27360,N_20228,N_19806);
xor U27361 (N_27361,N_23972,N_20894);
or U27362 (N_27362,N_22844,N_20347);
xnor U27363 (N_27363,N_20125,N_20544);
nor U27364 (N_27364,N_18719,N_21038);
xnor U27365 (N_27365,N_22444,N_23173);
nor U27366 (N_27366,N_23541,N_23860);
nand U27367 (N_27367,N_19122,N_22288);
or U27368 (N_27368,N_19452,N_22481);
xor U27369 (N_27369,N_22052,N_19123);
xor U27370 (N_27370,N_19230,N_18886);
nand U27371 (N_27371,N_22949,N_19998);
nand U27372 (N_27372,N_18515,N_23097);
or U27373 (N_27373,N_19144,N_23830);
nand U27374 (N_27374,N_21069,N_23442);
nor U27375 (N_27375,N_19428,N_21065);
nor U27376 (N_27376,N_22430,N_22747);
or U27377 (N_27377,N_23499,N_18259);
and U27378 (N_27378,N_23183,N_23685);
nand U27379 (N_27379,N_21262,N_18574);
nor U27380 (N_27380,N_20720,N_23351);
and U27381 (N_27381,N_21214,N_20345);
and U27382 (N_27382,N_21261,N_20009);
and U27383 (N_27383,N_22452,N_20529);
nand U27384 (N_27384,N_18374,N_21891);
and U27385 (N_27385,N_18060,N_18817);
nand U27386 (N_27386,N_21039,N_19023);
and U27387 (N_27387,N_18735,N_21964);
nor U27388 (N_27388,N_23838,N_21333);
xnor U27389 (N_27389,N_22607,N_19692);
or U27390 (N_27390,N_21444,N_22692);
nor U27391 (N_27391,N_18944,N_18873);
and U27392 (N_27392,N_18462,N_22417);
nand U27393 (N_27393,N_20235,N_18714);
nand U27394 (N_27394,N_18033,N_19561);
or U27395 (N_27395,N_23447,N_23137);
nand U27396 (N_27396,N_20289,N_21782);
nor U27397 (N_27397,N_19614,N_23599);
nor U27398 (N_27398,N_18396,N_20080);
nand U27399 (N_27399,N_22297,N_20592);
or U27400 (N_27400,N_19598,N_20114);
nor U27401 (N_27401,N_23207,N_18335);
nand U27402 (N_27402,N_22614,N_21697);
and U27403 (N_27403,N_18738,N_18876);
or U27404 (N_27404,N_21619,N_22223);
nor U27405 (N_27405,N_21459,N_18287);
or U27406 (N_27406,N_23268,N_20637);
nand U27407 (N_27407,N_21228,N_20114);
nand U27408 (N_27408,N_21583,N_22590);
xor U27409 (N_27409,N_23528,N_23958);
nor U27410 (N_27410,N_22577,N_21533);
or U27411 (N_27411,N_21547,N_20292);
and U27412 (N_27412,N_18527,N_19174);
nor U27413 (N_27413,N_23242,N_22732);
nand U27414 (N_27414,N_18666,N_21158);
nor U27415 (N_27415,N_22612,N_22803);
xor U27416 (N_27416,N_23258,N_19298);
nor U27417 (N_27417,N_21501,N_22218);
or U27418 (N_27418,N_19905,N_22885);
nor U27419 (N_27419,N_18026,N_18736);
nand U27420 (N_27420,N_23476,N_23465);
nor U27421 (N_27421,N_19944,N_23511);
nand U27422 (N_27422,N_21948,N_18349);
nor U27423 (N_27423,N_20380,N_20230);
nand U27424 (N_27424,N_18862,N_19747);
xor U27425 (N_27425,N_19522,N_19806);
xnor U27426 (N_27426,N_21063,N_21111);
xor U27427 (N_27427,N_18496,N_19347);
nand U27428 (N_27428,N_23936,N_21137);
and U27429 (N_27429,N_20140,N_19920);
or U27430 (N_27430,N_21342,N_19560);
nor U27431 (N_27431,N_19219,N_23174);
xor U27432 (N_27432,N_20739,N_20337);
nor U27433 (N_27433,N_18282,N_22398);
nor U27434 (N_27434,N_23310,N_23594);
nand U27435 (N_27435,N_22777,N_18027);
and U27436 (N_27436,N_23396,N_19906);
nor U27437 (N_27437,N_19202,N_22281);
xor U27438 (N_27438,N_23539,N_18135);
xor U27439 (N_27439,N_22134,N_20139);
or U27440 (N_27440,N_22518,N_19925);
nor U27441 (N_27441,N_23234,N_18769);
xnor U27442 (N_27442,N_19050,N_18728);
xnor U27443 (N_27443,N_21363,N_18150);
nand U27444 (N_27444,N_23081,N_18449);
nand U27445 (N_27445,N_20903,N_20635);
nor U27446 (N_27446,N_20413,N_19414);
nor U27447 (N_27447,N_20598,N_21411);
xor U27448 (N_27448,N_20171,N_22034);
nand U27449 (N_27449,N_21073,N_23031);
nand U27450 (N_27450,N_18300,N_19046);
nor U27451 (N_27451,N_20564,N_20712);
nor U27452 (N_27452,N_22654,N_23099);
xnor U27453 (N_27453,N_18305,N_19950);
xnor U27454 (N_27454,N_20755,N_23333);
or U27455 (N_27455,N_20899,N_21410);
nor U27456 (N_27456,N_21018,N_21948);
and U27457 (N_27457,N_23432,N_19936);
xor U27458 (N_27458,N_19442,N_21772);
nor U27459 (N_27459,N_23604,N_18563);
nand U27460 (N_27460,N_21249,N_19506);
or U27461 (N_27461,N_23706,N_20663);
and U27462 (N_27462,N_22699,N_21590);
nor U27463 (N_27463,N_18857,N_18159);
xnor U27464 (N_27464,N_19069,N_19413);
and U27465 (N_27465,N_19218,N_23830);
and U27466 (N_27466,N_20985,N_19510);
and U27467 (N_27467,N_22149,N_22592);
xnor U27468 (N_27468,N_21673,N_20959);
xor U27469 (N_27469,N_20568,N_20326);
or U27470 (N_27470,N_18897,N_19672);
or U27471 (N_27471,N_19397,N_21346);
xor U27472 (N_27472,N_18890,N_22931);
nor U27473 (N_27473,N_23999,N_20659);
nor U27474 (N_27474,N_19269,N_22176);
xor U27475 (N_27475,N_23970,N_23132);
or U27476 (N_27476,N_19677,N_22571);
or U27477 (N_27477,N_18325,N_19092);
or U27478 (N_27478,N_22121,N_22040);
or U27479 (N_27479,N_22743,N_18174);
or U27480 (N_27480,N_20695,N_20148);
xnor U27481 (N_27481,N_18990,N_22598);
xor U27482 (N_27482,N_22594,N_20719);
xnor U27483 (N_27483,N_19357,N_21753);
nand U27484 (N_27484,N_21243,N_22935);
and U27485 (N_27485,N_19849,N_23388);
and U27486 (N_27486,N_19833,N_19188);
nand U27487 (N_27487,N_21986,N_23731);
or U27488 (N_27488,N_20772,N_21175);
nand U27489 (N_27489,N_23977,N_21006);
nor U27490 (N_27490,N_21118,N_19315);
nor U27491 (N_27491,N_21853,N_22651);
or U27492 (N_27492,N_20975,N_20889);
or U27493 (N_27493,N_23411,N_20316);
xnor U27494 (N_27494,N_21788,N_23185);
nand U27495 (N_27495,N_21297,N_19369);
or U27496 (N_27496,N_18508,N_21713);
xnor U27497 (N_27497,N_23450,N_18418);
xnor U27498 (N_27498,N_20502,N_22635);
and U27499 (N_27499,N_19347,N_21215);
and U27500 (N_27500,N_22062,N_23424);
or U27501 (N_27501,N_23907,N_23891);
or U27502 (N_27502,N_18566,N_22534);
xor U27503 (N_27503,N_18599,N_19592);
nand U27504 (N_27504,N_22117,N_19387);
or U27505 (N_27505,N_23702,N_21162);
nand U27506 (N_27506,N_22754,N_23050);
nor U27507 (N_27507,N_19865,N_20638);
nor U27508 (N_27508,N_20531,N_23891);
and U27509 (N_27509,N_18128,N_22429);
nor U27510 (N_27510,N_23116,N_23211);
nand U27511 (N_27511,N_22123,N_23477);
xnor U27512 (N_27512,N_22264,N_21584);
or U27513 (N_27513,N_19226,N_18215);
nand U27514 (N_27514,N_23495,N_20555);
and U27515 (N_27515,N_22559,N_19570);
or U27516 (N_27516,N_21064,N_18596);
or U27517 (N_27517,N_19757,N_22924);
xnor U27518 (N_27518,N_21440,N_20809);
nand U27519 (N_27519,N_20274,N_21852);
or U27520 (N_27520,N_18013,N_23027);
and U27521 (N_27521,N_22218,N_23666);
nand U27522 (N_27522,N_18186,N_22701);
nor U27523 (N_27523,N_20567,N_23441);
xor U27524 (N_27524,N_22498,N_20171);
xnor U27525 (N_27525,N_19287,N_22710);
and U27526 (N_27526,N_18397,N_22075);
and U27527 (N_27527,N_23605,N_23934);
and U27528 (N_27528,N_18150,N_18608);
nor U27529 (N_27529,N_21718,N_18830);
or U27530 (N_27530,N_22950,N_21301);
nand U27531 (N_27531,N_22955,N_23563);
nor U27532 (N_27532,N_22860,N_18954);
and U27533 (N_27533,N_21529,N_18072);
xnor U27534 (N_27534,N_23076,N_18661);
nor U27535 (N_27535,N_23517,N_21333);
or U27536 (N_27536,N_18234,N_18836);
nor U27537 (N_27537,N_22591,N_22184);
nand U27538 (N_27538,N_20602,N_23120);
xor U27539 (N_27539,N_19881,N_22917);
nand U27540 (N_27540,N_19707,N_22880);
xnor U27541 (N_27541,N_20051,N_18580);
nor U27542 (N_27542,N_20053,N_19594);
or U27543 (N_27543,N_19718,N_19619);
nand U27544 (N_27544,N_23947,N_23468);
xor U27545 (N_27545,N_21195,N_23539);
xnor U27546 (N_27546,N_20083,N_20405);
nand U27547 (N_27547,N_22943,N_18040);
xor U27548 (N_27548,N_18346,N_23540);
nor U27549 (N_27549,N_19585,N_20817);
nand U27550 (N_27550,N_20963,N_22377);
and U27551 (N_27551,N_22507,N_22222);
and U27552 (N_27552,N_20037,N_21495);
and U27553 (N_27553,N_18062,N_19066);
xnor U27554 (N_27554,N_22994,N_23132);
or U27555 (N_27555,N_23274,N_22163);
or U27556 (N_27556,N_21795,N_18687);
nand U27557 (N_27557,N_22363,N_20249);
or U27558 (N_27558,N_20101,N_23268);
xnor U27559 (N_27559,N_19679,N_21152);
and U27560 (N_27560,N_23346,N_23157);
or U27561 (N_27561,N_19745,N_19427);
nor U27562 (N_27562,N_20509,N_20961);
xor U27563 (N_27563,N_21877,N_21287);
xor U27564 (N_27564,N_19683,N_22248);
nor U27565 (N_27565,N_19963,N_20684);
xor U27566 (N_27566,N_19301,N_18100);
nand U27567 (N_27567,N_21015,N_22559);
xor U27568 (N_27568,N_21396,N_18064);
nor U27569 (N_27569,N_23543,N_20556);
or U27570 (N_27570,N_20366,N_18511);
and U27571 (N_27571,N_21479,N_23763);
or U27572 (N_27572,N_21753,N_21703);
nor U27573 (N_27573,N_19265,N_23516);
nand U27574 (N_27574,N_20001,N_22349);
nand U27575 (N_27575,N_18735,N_22159);
and U27576 (N_27576,N_18915,N_21517);
and U27577 (N_27577,N_19700,N_21646);
or U27578 (N_27578,N_20465,N_20350);
nor U27579 (N_27579,N_23780,N_19331);
and U27580 (N_27580,N_21894,N_21738);
xnor U27581 (N_27581,N_22792,N_22030);
and U27582 (N_27582,N_19600,N_20164);
or U27583 (N_27583,N_20660,N_18282);
nand U27584 (N_27584,N_18205,N_21339);
or U27585 (N_27585,N_20555,N_19729);
and U27586 (N_27586,N_19839,N_19441);
and U27587 (N_27587,N_21557,N_19608);
or U27588 (N_27588,N_18903,N_20659);
and U27589 (N_27589,N_22396,N_19755);
or U27590 (N_27590,N_23921,N_23694);
nor U27591 (N_27591,N_21992,N_20039);
or U27592 (N_27592,N_20991,N_19724);
nand U27593 (N_27593,N_22172,N_18476);
xor U27594 (N_27594,N_21414,N_22989);
nand U27595 (N_27595,N_18194,N_20494);
and U27596 (N_27596,N_22106,N_19408);
xor U27597 (N_27597,N_19607,N_21476);
nor U27598 (N_27598,N_18718,N_21343);
nor U27599 (N_27599,N_20837,N_22438);
or U27600 (N_27600,N_18207,N_21530);
nand U27601 (N_27601,N_20216,N_21566);
nand U27602 (N_27602,N_20588,N_22036);
or U27603 (N_27603,N_20194,N_21068);
nor U27604 (N_27604,N_20859,N_23528);
and U27605 (N_27605,N_20173,N_20131);
nor U27606 (N_27606,N_19318,N_19997);
and U27607 (N_27607,N_21587,N_19336);
or U27608 (N_27608,N_18870,N_18373);
nand U27609 (N_27609,N_22335,N_21357);
or U27610 (N_27610,N_19975,N_20907);
nor U27611 (N_27611,N_22055,N_23384);
nor U27612 (N_27612,N_23466,N_19822);
nor U27613 (N_27613,N_23056,N_19802);
nand U27614 (N_27614,N_19512,N_20753);
nor U27615 (N_27615,N_20232,N_21519);
and U27616 (N_27616,N_18384,N_22757);
nand U27617 (N_27617,N_22218,N_19163);
or U27618 (N_27618,N_20345,N_20191);
nor U27619 (N_27619,N_19451,N_23846);
or U27620 (N_27620,N_23219,N_18262);
nor U27621 (N_27621,N_18487,N_19369);
nand U27622 (N_27622,N_23258,N_22330);
and U27623 (N_27623,N_20923,N_21688);
or U27624 (N_27624,N_21157,N_20541);
and U27625 (N_27625,N_23462,N_18219);
or U27626 (N_27626,N_19132,N_21982);
or U27627 (N_27627,N_19813,N_18471);
nand U27628 (N_27628,N_19739,N_20239);
or U27629 (N_27629,N_19613,N_18522);
xnor U27630 (N_27630,N_19970,N_22302);
xor U27631 (N_27631,N_21470,N_18166);
xor U27632 (N_27632,N_21043,N_20974);
and U27633 (N_27633,N_19619,N_18022);
or U27634 (N_27634,N_19781,N_18579);
or U27635 (N_27635,N_19077,N_19417);
or U27636 (N_27636,N_21033,N_18124);
nand U27637 (N_27637,N_19466,N_19661);
or U27638 (N_27638,N_20038,N_19195);
and U27639 (N_27639,N_19953,N_22104);
nand U27640 (N_27640,N_22357,N_23590);
nor U27641 (N_27641,N_23352,N_22333);
and U27642 (N_27642,N_18103,N_23632);
nand U27643 (N_27643,N_18871,N_18373);
nand U27644 (N_27644,N_22512,N_19879);
nor U27645 (N_27645,N_20402,N_19098);
nor U27646 (N_27646,N_19128,N_23140);
or U27647 (N_27647,N_21164,N_21512);
or U27648 (N_27648,N_22548,N_22426);
nor U27649 (N_27649,N_21761,N_18979);
xnor U27650 (N_27650,N_23813,N_20661);
and U27651 (N_27651,N_22421,N_18810);
and U27652 (N_27652,N_21268,N_20820);
or U27653 (N_27653,N_20299,N_21793);
and U27654 (N_27654,N_19794,N_20423);
xnor U27655 (N_27655,N_20871,N_21039);
xor U27656 (N_27656,N_20752,N_22554);
and U27657 (N_27657,N_19610,N_21904);
nand U27658 (N_27658,N_22285,N_23448);
nor U27659 (N_27659,N_19451,N_19779);
and U27660 (N_27660,N_19343,N_23371);
nor U27661 (N_27661,N_18629,N_23283);
or U27662 (N_27662,N_19755,N_18786);
nor U27663 (N_27663,N_21038,N_20649);
and U27664 (N_27664,N_22395,N_22549);
nand U27665 (N_27665,N_18652,N_20362);
and U27666 (N_27666,N_21510,N_22120);
or U27667 (N_27667,N_23676,N_22874);
nand U27668 (N_27668,N_23233,N_21116);
or U27669 (N_27669,N_19779,N_20970);
nand U27670 (N_27670,N_23724,N_20553);
and U27671 (N_27671,N_19792,N_18899);
nand U27672 (N_27672,N_22751,N_21922);
xnor U27673 (N_27673,N_20036,N_21724);
nor U27674 (N_27674,N_20040,N_19301);
nand U27675 (N_27675,N_19869,N_21108);
xor U27676 (N_27676,N_21138,N_21272);
and U27677 (N_27677,N_21175,N_22080);
or U27678 (N_27678,N_23956,N_22956);
nor U27679 (N_27679,N_21051,N_19450);
and U27680 (N_27680,N_19808,N_20503);
nand U27681 (N_27681,N_20572,N_18235);
and U27682 (N_27682,N_21113,N_23342);
nand U27683 (N_27683,N_23118,N_20915);
and U27684 (N_27684,N_22247,N_23132);
nor U27685 (N_27685,N_19674,N_23311);
and U27686 (N_27686,N_20274,N_18265);
or U27687 (N_27687,N_18469,N_19474);
nor U27688 (N_27688,N_18994,N_21554);
nor U27689 (N_27689,N_18005,N_23766);
nor U27690 (N_27690,N_18481,N_19684);
nor U27691 (N_27691,N_19015,N_22107);
or U27692 (N_27692,N_19212,N_21878);
and U27693 (N_27693,N_22608,N_19315);
and U27694 (N_27694,N_20950,N_19947);
and U27695 (N_27695,N_19188,N_23378);
or U27696 (N_27696,N_23083,N_22943);
nor U27697 (N_27697,N_21365,N_22409);
and U27698 (N_27698,N_18610,N_23269);
and U27699 (N_27699,N_22442,N_23101);
or U27700 (N_27700,N_20449,N_23105);
nor U27701 (N_27701,N_19453,N_21874);
or U27702 (N_27702,N_21191,N_19744);
xnor U27703 (N_27703,N_18475,N_19717);
and U27704 (N_27704,N_20751,N_19615);
and U27705 (N_27705,N_21782,N_23674);
xor U27706 (N_27706,N_19577,N_18808);
xnor U27707 (N_27707,N_23345,N_20947);
or U27708 (N_27708,N_19950,N_19208);
or U27709 (N_27709,N_23899,N_18957);
xor U27710 (N_27710,N_20831,N_19089);
and U27711 (N_27711,N_21106,N_20299);
or U27712 (N_27712,N_20980,N_18370);
and U27713 (N_27713,N_18765,N_22871);
nor U27714 (N_27714,N_20934,N_21612);
or U27715 (N_27715,N_20460,N_23283);
or U27716 (N_27716,N_19491,N_21736);
and U27717 (N_27717,N_23466,N_20390);
nand U27718 (N_27718,N_22756,N_21361);
nand U27719 (N_27719,N_20424,N_18175);
or U27720 (N_27720,N_20535,N_19954);
and U27721 (N_27721,N_18731,N_18542);
xnor U27722 (N_27722,N_19063,N_21915);
and U27723 (N_27723,N_21988,N_19320);
or U27724 (N_27724,N_20384,N_21904);
or U27725 (N_27725,N_19037,N_23525);
or U27726 (N_27726,N_18890,N_22272);
nor U27727 (N_27727,N_18662,N_20075);
or U27728 (N_27728,N_20004,N_21712);
nand U27729 (N_27729,N_22100,N_23955);
nor U27730 (N_27730,N_21079,N_20375);
nand U27731 (N_27731,N_22467,N_21932);
xnor U27732 (N_27732,N_20181,N_18311);
xnor U27733 (N_27733,N_21676,N_21627);
and U27734 (N_27734,N_22775,N_22628);
xnor U27735 (N_27735,N_18243,N_21823);
xnor U27736 (N_27736,N_21982,N_23048);
or U27737 (N_27737,N_20382,N_19999);
nor U27738 (N_27738,N_19215,N_19977);
xnor U27739 (N_27739,N_20665,N_20425);
or U27740 (N_27740,N_23321,N_19883);
xor U27741 (N_27741,N_22439,N_20524);
or U27742 (N_27742,N_18308,N_22486);
nor U27743 (N_27743,N_22838,N_20974);
or U27744 (N_27744,N_23320,N_21421);
xnor U27745 (N_27745,N_23615,N_19172);
nand U27746 (N_27746,N_20789,N_18225);
and U27747 (N_27747,N_22105,N_20996);
nand U27748 (N_27748,N_23028,N_19595);
or U27749 (N_27749,N_19177,N_22020);
and U27750 (N_27750,N_18620,N_23776);
nor U27751 (N_27751,N_18289,N_23404);
and U27752 (N_27752,N_21054,N_20069);
nor U27753 (N_27753,N_21292,N_21590);
nand U27754 (N_27754,N_19892,N_20201);
and U27755 (N_27755,N_20095,N_23946);
nand U27756 (N_27756,N_22363,N_23583);
or U27757 (N_27757,N_23128,N_21903);
nor U27758 (N_27758,N_23537,N_18329);
nand U27759 (N_27759,N_19289,N_18203);
or U27760 (N_27760,N_19287,N_18380);
nor U27761 (N_27761,N_19812,N_18050);
nand U27762 (N_27762,N_22687,N_23825);
xor U27763 (N_27763,N_21749,N_22683);
nand U27764 (N_27764,N_18202,N_22779);
or U27765 (N_27765,N_21630,N_18840);
nand U27766 (N_27766,N_21183,N_21230);
or U27767 (N_27767,N_21852,N_22926);
nand U27768 (N_27768,N_22858,N_22161);
nor U27769 (N_27769,N_23661,N_23269);
or U27770 (N_27770,N_18215,N_18655);
and U27771 (N_27771,N_22067,N_18105);
or U27772 (N_27772,N_21209,N_22582);
or U27773 (N_27773,N_20568,N_18480);
or U27774 (N_27774,N_21422,N_23535);
xor U27775 (N_27775,N_21466,N_19170);
or U27776 (N_27776,N_21778,N_20302);
or U27777 (N_27777,N_19336,N_19440);
or U27778 (N_27778,N_23713,N_23021);
xnor U27779 (N_27779,N_20810,N_19329);
or U27780 (N_27780,N_22155,N_20074);
nor U27781 (N_27781,N_19549,N_20249);
nand U27782 (N_27782,N_23496,N_18596);
nor U27783 (N_27783,N_19470,N_20026);
nor U27784 (N_27784,N_18250,N_22444);
nand U27785 (N_27785,N_20652,N_23904);
or U27786 (N_27786,N_20654,N_20989);
xnor U27787 (N_27787,N_22129,N_21638);
and U27788 (N_27788,N_19201,N_22175);
or U27789 (N_27789,N_21263,N_23242);
nand U27790 (N_27790,N_20268,N_20319);
nand U27791 (N_27791,N_21782,N_23734);
or U27792 (N_27792,N_22557,N_20256);
nand U27793 (N_27793,N_23235,N_19262);
or U27794 (N_27794,N_18338,N_22966);
nand U27795 (N_27795,N_23675,N_23446);
xnor U27796 (N_27796,N_21901,N_19362);
and U27797 (N_27797,N_21309,N_21154);
or U27798 (N_27798,N_23287,N_21675);
or U27799 (N_27799,N_22095,N_20177);
or U27800 (N_27800,N_21351,N_20491);
and U27801 (N_27801,N_21269,N_20135);
nand U27802 (N_27802,N_21380,N_18806);
and U27803 (N_27803,N_20859,N_19450);
or U27804 (N_27804,N_23121,N_18531);
nand U27805 (N_27805,N_23873,N_22829);
xnor U27806 (N_27806,N_18332,N_18006);
or U27807 (N_27807,N_22778,N_23235);
and U27808 (N_27808,N_18409,N_19103);
nor U27809 (N_27809,N_23408,N_18332);
nor U27810 (N_27810,N_22975,N_21334);
nand U27811 (N_27811,N_22516,N_23314);
or U27812 (N_27812,N_23091,N_21211);
xnor U27813 (N_27813,N_23961,N_18326);
nor U27814 (N_27814,N_19431,N_19974);
xnor U27815 (N_27815,N_20855,N_23628);
or U27816 (N_27816,N_21215,N_20546);
and U27817 (N_27817,N_22111,N_22113);
or U27818 (N_27818,N_23471,N_23132);
or U27819 (N_27819,N_21725,N_22365);
and U27820 (N_27820,N_19388,N_20962);
and U27821 (N_27821,N_20324,N_23277);
xor U27822 (N_27822,N_23254,N_20932);
or U27823 (N_27823,N_18140,N_18231);
nand U27824 (N_27824,N_18672,N_21039);
or U27825 (N_27825,N_19324,N_18658);
and U27826 (N_27826,N_20228,N_19324);
nand U27827 (N_27827,N_18963,N_23919);
and U27828 (N_27828,N_20261,N_20460);
and U27829 (N_27829,N_22781,N_22834);
or U27830 (N_27830,N_22878,N_18511);
xor U27831 (N_27831,N_22216,N_19243);
and U27832 (N_27832,N_21478,N_18117);
or U27833 (N_27833,N_21953,N_21966);
or U27834 (N_27834,N_19780,N_18536);
or U27835 (N_27835,N_23410,N_20231);
nand U27836 (N_27836,N_23533,N_21231);
and U27837 (N_27837,N_18606,N_22749);
nand U27838 (N_27838,N_21142,N_20571);
nand U27839 (N_27839,N_23058,N_20617);
xor U27840 (N_27840,N_19629,N_23714);
nor U27841 (N_27841,N_21309,N_20594);
nand U27842 (N_27842,N_23578,N_22572);
nand U27843 (N_27843,N_22705,N_19369);
or U27844 (N_27844,N_21746,N_20322);
nand U27845 (N_27845,N_23678,N_21339);
and U27846 (N_27846,N_18598,N_18433);
nor U27847 (N_27847,N_22005,N_23234);
or U27848 (N_27848,N_20417,N_23176);
nand U27849 (N_27849,N_23107,N_18705);
nor U27850 (N_27850,N_23420,N_20490);
nand U27851 (N_27851,N_20035,N_20437);
nand U27852 (N_27852,N_21870,N_20847);
xor U27853 (N_27853,N_21535,N_23437);
nor U27854 (N_27854,N_20158,N_23416);
nand U27855 (N_27855,N_22928,N_22582);
nand U27856 (N_27856,N_23744,N_19638);
or U27857 (N_27857,N_21099,N_21962);
xnor U27858 (N_27858,N_22493,N_19524);
nor U27859 (N_27859,N_22098,N_21216);
and U27860 (N_27860,N_21676,N_18529);
and U27861 (N_27861,N_22953,N_21303);
and U27862 (N_27862,N_18722,N_18252);
nor U27863 (N_27863,N_22310,N_21919);
xor U27864 (N_27864,N_22672,N_18896);
and U27865 (N_27865,N_23542,N_22897);
or U27866 (N_27866,N_19311,N_23443);
or U27867 (N_27867,N_23470,N_21873);
nor U27868 (N_27868,N_23556,N_18123);
nor U27869 (N_27869,N_18126,N_23677);
nor U27870 (N_27870,N_20771,N_19427);
xnor U27871 (N_27871,N_18385,N_20737);
nand U27872 (N_27872,N_21338,N_23308);
or U27873 (N_27873,N_21973,N_20640);
or U27874 (N_27874,N_21668,N_21790);
nand U27875 (N_27875,N_19671,N_21828);
nor U27876 (N_27876,N_19950,N_20329);
nor U27877 (N_27877,N_19756,N_22299);
nand U27878 (N_27878,N_20221,N_18462);
xnor U27879 (N_27879,N_23383,N_21669);
or U27880 (N_27880,N_20135,N_21416);
nand U27881 (N_27881,N_23152,N_19577);
xnor U27882 (N_27882,N_19500,N_18101);
or U27883 (N_27883,N_19317,N_20387);
nor U27884 (N_27884,N_21339,N_22579);
or U27885 (N_27885,N_18125,N_22530);
nor U27886 (N_27886,N_21839,N_21268);
nor U27887 (N_27887,N_23413,N_22576);
xnor U27888 (N_27888,N_21559,N_21245);
nand U27889 (N_27889,N_21098,N_20122);
or U27890 (N_27890,N_19307,N_21708);
nor U27891 (N_27891,N_21592,N_20780);
or U27892 (N_27892,N_21403,N_22700);
xnor U27893 (N_27893,N_22214,N_19821);
or U27894 (N_27894,N_21206,N_23330);
nand U27895 (N_27895,N_23881,N_21927);
and U27896 (N_27896,N_19800,N_18025);
nor U27897 (N_27897,N_22456,N_21899);
and U27898 (N_27898,N_22771,N_19556);
or U27899 (N_27899,N_19598,N_18898);
or U27900 (N_27900,N_18070,N_23778);
or U27901 (N_27901,N_22283,N_22346);
and U27902 (N_27902,N_23935,N_23320);
and U27903 (N_27903,N_22271,N_21039);
nor U27904 (N_27904,N_19203,N_20671);
nand U27905 (N_27905,N_20832,N_19377);
xor U27906 (N_27906,N_22830,N_19006);
xor U27907 (N_27907,N_20760,N_18704);
nor U27908 (N_27908,N_18249,N_22859);
nand U27909 (N_27909,N_21828,N_23546);
nand U27910 (N_27910,N_19675,N_21385);
or U27911 (N_27911,N_23952,N_23756);
nand U27912 (N_27912,N_23631,N_22793);
nor U27913 (N_27913,N_18151,N_23836);
or U27914 (N_27914,N_19712,N_19119);
xor U27915 (N_27915,N_21748,N_21657);
nand U27916 (N_27916,N_19672,N_22629);
nand U27917 (N_27917,N_23863,N_18487);
and U27918 (N_27918,N_21512,N_18216);
or U27919 (N_27919,N_19634,N_20005);
nand U27920 (N_27920,N_19621,N_20705);
or U27921 (N_27921,N_22209,N_23078);
xor U27922 (N_27922,N_18846,N_23327);
xnor U27923 (N_27923,N_19209,N_18420);
or U27924 (N_27924,N_18589,N_18311);
xor U27925 (N_27925,N_20692,N_18248);
or U27926 (N_27926,N_23907,N_20513);
xnor U27927 (N_27927,N_21256,N_23940);
nand U27928 (N_27928,N_23258,N_23180);
nand U27929 (N_27929,N_22018,N_21325);
or U27930 (N_27930,N_18712,N_18112);
nand U27931 (N_27931,N_20381,N_23737);
or U27932 (N_27932,N_21495,N_21000);
xnor U27933 (N_27933,N_19798,N_22714);
nand U27934 (N_27934,N_18832,N_21931);
and U27935 (N_27935,N_21360,N_22120);
and U27936 (N_27936,N_19195,N_19966);
nand U27937 (N_27937,N_20162,N_22333);
xnor U27938 (N_27938,N_18443,N_23204);
or U27939 (N_27939,N_20680,N_20565);
or U27940 (N_27940,N_22056,N_19640);
and U27941 (N_27941,N_22452,N_21843);
nor U27942 (N_27942,N_18834,N_21777);
nor U27943 (N_27943,N_19622,N_22734);
nand U27944 (N_27944,N_20007,N_21265);
xnor U27945 (N_27945,N_18407,N_20324);
and U27946 (N_27946,N_21152,N_20160);
and U27947 (N_27947,N_20841,N_21803);
or U27948 (N_27948,N_21656,N_20982);
or U27949 (N_27949,N_20231,N_18094);
nor U27950 (N_27950,N_19112,N_18528);
or U27951 (N_27951,N_19971,N_23811);
and U27952 (N_27952,N_22717,N_18643);
nand U27953 (N_27953,N_20432,N_21222);
or U27954 (N_27954,N_19621,N_19371);
nand U27955 (N_27955,N_22143,N_22195);
or U27956 (N_27956,N_20566,N_23516);
and U27957 (N_27957,N_23979,N_19951);
nand U27958 (N_27958,N_19883,N_21332);
and U27959 (N_27959,N_23888,N_22208);
xnor U27960 (N_27960,N_19644,N_23161);
nand U27961 (N_27961,N_21915,N_18540);
xnor U27962 (N_27962,N_19104,N_22092);
and U27963 (N_27963,N_23390,N_22057);
nor U27964 (N_27964,N_23941,N_18791);
nor U27965 (N_27965,N_21929,N_23273);
and U27966 (N_27966,N_21515,N_21222);
or U27967 (N_27967,N_18703,N_22436);
or U27968 (N_27968,N_18250,N_22518);
and U27969 (N_27969,N_22321,N_18717);
nand U27970 (N_27970,N_20203,N_22388);
xnor U27971 (N_27971,N_21777,N_21553);
xor U27972 (N_27972,N_19787,N_22515);
nand U27973 (N_27973,N_21889,N_19848);
or U27974 (N_27974,N_20498,N_23301);
and U27975 (N_27975,N_23501,N_22753);
and U27976 (N_27976,N_23434,N_18853);
or U27977 (N_27977,N_21190,N_19035);
nand U27978 (N_27978,N_21799,N_19834);
nand U27979 (N_27979,N_18949,N_19415);
nor U27980 (N_27980,N_23676,N_23307);
nand U27981 (N_27981,N_18830,N_18992);
nor U27982 (N_27982,N_22744,N_20917);
nand U27983 (N_27983,N_23122,N_19087);
and U27984 (N_27984,N_19175,N_20275);
and U27985 (N_27985,N_18818,N_21372);
nor U27986 (N_27986,N_23981,N_19696);
nand U27987 (N_27987,N_19426,N_23110);
or U27988 (N_27988,N_20170,N_21573);
xor U27989 (N_27989,N_20315,N_20690);
and U27990 (N_27990,N_18796,N_19583);
xor U27991 (N_27991,N_22808,N_21196);
or U27992 (N_27992,N_20173,N_21353);
nor U27993 (N_27993,N_20976,N_23311);
nor U27994 (N_27994,N_19953,N_21332);
nand U27995 (N_27995,N_19793,N_20035);
xor U27996 (N_27996,N_22961,N_18359);
nand U27997 (N_27997,N_18313,N_20882);
nor U27998 (N_27998,N_20849,N_22571);
xnor U27999 (N_27999,N_20319,N_22667);
and U28000 (N_28000,N_19780,N_19967);
xor U28001 (N_28001,N_19668,N_21855);
nor U28002 (N_28002,N_23737,N_21493);
xor U28003 (N_28003,N_23736,N_23676);
or U28004 (N_28004,N_22494,N_22290);
nor U28005 (N_28005,N_23844,N_19264);
or U28006 (N_28006,N_19827,N_21926);
xor U28007 (N_28007,N_18961,N_21182);
xnor U28008 (N_28008,N_18537,N_18396);
xor U28009 (N_28009,N_21039,N_22913);
and U28010 (N_28010,N_21576,N_21632);
and U28011 (N_28011,N_22859,N_22805);
and U28012 (N_28012,N_22932,N_19071);
nand U28013 (N_28013,N_23745,N_19949);
nor U28014 (N_28014,N_21800,N_23990);
xnor U28015 (N_28015,N_23009,N_19759);
or U28016 (N_28016,N_18213,N_22859);
nand U28017 (N_28017,N_21728,N_21819);
nand U28018 (N_28018,N_23128,N_18146);
nand U28019 (N_28019,N_18945,N_23411);
nor U28020 (N_28020,N_19960,N_21526);
or U28021 (N_28021,N_18525,N_19961);
nand U28022 (N_28022,N_23044,N_20278);
nand U28023 (N_28023,N_23658,N_20065);
xor U28024 (N_28024,N_23711,N_23006);
or U28025 (N_28025,N_19244,N_19764);
xor U28026 (N_28026,N_21272,N_21581);
and U28027 (N_28027,N_21780,N_19436);
xnor U28028 (N_28028,N_19453,N_18218);
or U28029 (N_28029,N_19270,N_18526);
xnor U28030 (N_28030,N_21661,N_18191);
nor U28031 (N_28031,N_19995,N_20521);
or U28032 (N_28032,N_20344,N_23788);
nor U28033 (N_28033,N_22219,N_19144);
or U28034 (N_28034,N_19793,N_23684);
or U28035 (N_28035,N_21578,N_20762);
and U28036 (N_28036,N_20081,N_21940);
or U28037 (N_28037,N_23667,N_21885);
xor U28038 (N_28038,N_19859,N_18521);
xor U28039 (N_28039,N_22310,N_21700);
xnor U28040 (N_28040,N_18332,N_19202);
xnor U28041 (N_28041,N_18301,N_20739);
nor U28042 (N_28042,N_18481,N_23337);
and U28043 (N_28043,N_21124,N_23630);
nand U28044 (N_28044,N_18495,N_20401);
or U28045 (N_28045,N_23757,N_19148);
nand U28046 (N_28046,N_20521,N_23624);
xnor U28047 (N_28047,N_22126,N_20853);
or U28048 (N_28048,N_21345,N_23493);
nor U28049 (N_28049,N_18094,N_21642);
or U28050 (N_28050,N_21980,N_20931);
or U28051 (N_28051,N_21880,N_22531);
xor U28052 (N_28052,N_22238,N_19731);
or U28053 (N_28053,N_20685,N_22999);
and U28054 (N_28054,N_22418,N_22515);
or U28055 (N_28055,N_18173,N_18416);
nand U28056 (N_28056,N_20598,N_21198);
or U28057 (N_28057,N_22011,N_22061);
nor U28058 (N_28058,N_23300,N_22331);
and U28059 (N_28059,N_21450,N_23454);
and U28060 (N_28060,N_19463,N_23395);
nor U28061 (N_28061,N_18533,N_20501);
nor U28062 (N_28062,N_23989,N_21006);
or U28063 (N_28063,N_18165,N_20300);
and U28064 (N_28064,N_22859,N_18248);
or U28065 (N_28065,N_19188,N_23924);
and U28066 (N_28066,N_18029,N_19515);
nand U28067 (N_28067,N_22866,N_19688);
nand U28068 (N_28068,N_22812,N_23306);
nor U28069 (N_28069,N_19242,N_23342);
or U28070 (N_28070,N_19736,N_22807);
xnor U28071 (N_28071,N_19459,N_18129);
nor U28072 (N_28072,N_19571,N_22131);
and U28073 (N_28073,N_18515,N_22957);
xor U28074 (N_28074,N_22548,N_20416);
or U28075 (N_28075,N_23991,N_19626);
and U28076 (N_28076,N_23439,N_18043);
nand U28077 (N_28077,N_20783,N_23296);
and U28078 (N_28078,N_18053,N_22882);
nor U28079 (N_28079,N_19789,N_20781);
nand U28080 (N_28080,N_19116,N_21239);
nand U28081 (N_28081,N_23167,N_19372);
xnor U28082 (N_28082,N_19007,N_21632);
nor U28083 (N_28083,N_23573,N_19032);
and U28084 (N_28084,N_23183,N_21482);
nand U28085 (N_28085,N_20257,N_18675);
xor U28086 (N_28086,N_23212,N_18462);
nor U28087 (N_28087,N_22983,N_23938);
nand U28088 (N_28088,N_21582,N_20819);
nor U28089 (N_28089,N_18519,N_18897);
nor U28090 (N_28090,N_23606,N_19602);
nand U28091 (N_28091,N_19557,N_18690);
nand U28092 (N_28092,N_18263,N_23345);
xnor U28093 (N_28093,N_23384,N_23547);
xnor U28094 (N_28094,N_20428,N_18935);
or U28095 (N_28095,N_20500,N_18154);
xnor U28096 (N_28096,N_22831,N_21659);
nor U28097 (N_28097,N_18141,N_18432);
or U28098 (N_28098,N_22995,N_22852);
xor U28099 (N_28099,N_20655,N_22432);
nand U28100 (N_28100,N_18327,N_18306);
and U28101 (N_28101,N_22971,N_20844);
nand U28102 (N_28102,N_18139,N_21232);
nor U28103 (N_28103,N_20104,N_19243);
nor U28104 (N_28104,N_19340,N_18598);
nor U28105 (N_28105,N_18371,N_19370);
nand U28106 (N_28106,N_21620,N_19828);
nand U28107 (N_28107,N_22906,N_18451);
nand U28108 (N_28108,N_20846,N_21150);
or U28109 (N_28109,N_23289,N_18873);
or U28110 (N_28110,N_18230,N_19431);
nand U28111 (N_28111,N_18104,N_19420);
nand U28112 (N_28112,N_21683,N_22640);
nor U28113 (N_28113,N_20223,N_18926);
nand U28114 (N_28114,N_23538,N_21688);
xnor U28115 (N_28115,N_20822,N_20390);
and U28116 (N_28116,N_20377,N_20542);
and U28117 (N_28117,N_23017,N_20174);
xor U28118 (N_28118,N_20207,N_21083);
and U28119 (N_28119,N_18832,N_18149);
nand U28120 (N_28120,N_20698,N_20609);
xnor U28121 (N_28121,N_23666,N_21039);
nand U28122 (N_28122,N_18786,N_23403);
or U28123 (N_28123,N_23272,N_21959);
nand U28124 (N_28124,N_19526,N_19236);
and U28125 (N_28125,N_20700,N_20753);
and U28126 (N_28126,N_22561,N_22636);
nor U28127 (N_28127,N_19025,N_19801);
nand U28128 (N_28128,N_23547,N_20675);
and U28129 (N_28129,N_23267,N_22924);
or U28130 (N_28130,N_19269,N_21753);
and U28131 (N_28131,N_21219,N_23398);
or U28132 (N_28132,N_21548,N_20803);
nand U28133 (N_28133,N_18973,N_19211);
nand U28134 (N_28134,N_23276,N_22295);
and U28135 (N_28135,N_18094,N_22346);
or U28136 (N_28136,N_21842,N_23910);
xnor U28137 (N_28137,N_21188,N_21479);
xnor U28138 (N_28138,N_19801,N_22986);
nand U28139 (N_28139,N_19907,N_23606);
nor U28140 (N_28140,N_19956,N_22641);
or U28141 (N_28141,N_19831,N_19502);
or U28142 (N_28142,N_22255,N_23048);
nor U28143 (N_28143,N_22940,N_19850);
and U28144 (N_28144,N_21634,N_19179);
nand U28145 (N_28145,N_22708,N_20512);
nand U28146 (N_28146,N_23244,N_18884);
and U28147 (N_28147,N_20378,N_18391);
nand U28148 (N_28148,N_18584,N_20484);
and U28149 (N_28149,N_22822,N_20345);
or U28150 (N_28150,N_23847,N_23673);
or U28151 (N_28151,N_22153,N_22353);
or U28152 (N_28152,N_21691,N_18221);
nand U28153 (N_28153,N_23756,N_19333);
or U28154 (N_28154,N_18714,N_18522);
nand U28155 (N_28155,N_21870,N_21433);
xnor U28156 (N_28156,N_23944,N_19457);
or U28157 (N_28157,N_22634,N_21398);
nand U28158 (N_28158,N_23506,N_23883);
or U28159 (N_28159,N_18118,N_18025);
or U28160 (N_28160,N_20309,N_19181);
and U28161 (N_28161,N_22965,N_22585);
or U28162 (N_28162,N_18405,N_22809);
and U28163 (N_28163,N_23808,N_18229);
and U28164 (N_28164,N_21727,N_20757);
xor U28165 (N_28165,N_23545,N_23933);
or U28166 (N_28166,N_22856,N_23833);
nand U28167 (N_28167,N_21824,N_20384);
xnor U28168 (N_28168,N_20858,N_18216);
or U28169 (N_28169,N_18958,N_18159);
and U28170 (N_28170,N_21882,N_22934);
nor U28171 (N_28171,N_20248,N_22425);
nor U28172 (N_28172,N_18722,N_23083);
nor U28173 (N_28173,N_18978,N_22032);
and U28174 (N_28174,N_23159,N_23789);
or U28175 (N_28175,N_22074,N_18767);
nor U28176 (N_28176,N_23935,N_21342);
nand U28177 (N_28177,N_18908,N_20715);
xor U28178 (N_28178,N_23969,N_19810);
or U28179 (N_28179,N_19146,N_21913);
xor U28180 (N_28180,N_18009,N_23883);
nor U28181 (N_28181,N_23129,N_23173);
and U28182 (N_28182,N_18910,N_20634);
xor U28183 (N_28183,N_22188,N_22234);
nand U28184 (N_28184,N_21345,N_21965);
or U28185 (N_28185,N_18246,N_18490);
nand U28186 (N_28186,N_20026,N_20619);
or U28187 (N_28187,N_18061,N_21269);
nor U28188 (N_28188,N_22355,N_21686);
xnor U28189 (N_28189,N_19253,N_20265);
and U28190 (N_28190,N_22084,N_18179);
nor U28191 (N_28191,N_20656,N_19670);
nand U28192 (N_28192,N_22325,N_23187);
and U28193 (N_28193,N_20594,N_21930);
nor U28194 (N_28194,N_19745,N_21781);
and U28195 (N_28195,N_18582,N_19952);
nor U28196 (N_28196,N_18900,N_23787);
xnor U28197 (N_28197,N_23886,N_19145);
or U28198 (N_28198,N_20544,N_21053);
nand U28199 (N_28199,N_21918,N_20909);
nand U28200 (N_28200,N_23549,N_23008);
and U28201 (N_28201,N_18125,N_19711);
nor U28202 (N_28202,N_19688,N_20253);
or U28203 (N_28203,N_19971,N_23031);
or U28204 (N_28204,N_21330,N_18169);
and U28205 (N_28205,N_18600,N_21395);
nand U28206 (N_28206,N_18774,N_22692);
and U28207 (N_28207,N_23872,N_18149);
xor U28208 (N_28208,N_23527,N_18804);
nand U28209 (N_28209,N_23223,N_18514);
or U28210 (N_28210,N_21529,N_20102);
xnor U28211 (N_28211,N_18748,N_18073);
xor U28212 (N_28212,N_18315,N_20214);
nor U28213 (N_28213,N_19586,N_18819);
or U28214 (N_28214,N_21514,N_19682);
or U28215 (N_28215,N_20891,N_18384);
nand U28216 (N_28216,N_22960,N_22492);
xor U28217 (N_28217,N_19243,N_19633);
nor U28218 (N_28218,N_22371,N_21580);
or U28219 (N_28219,N_20246,N_18835);
nor U28220 (N_28220,N_21681,N_22215);
and U28221 (N_28221,N_23688,N_20086);
nor U28222 (N_28222,N_21102,N_23521);
or U28223 (N_28223,N_23611,N_20150);
nor U28224 (N_28224,N_23258,N_21367);
and U28225 (N_28225,N_22861,N_23903);
nor U28226 (N_28226,N_20908,N_21623);
nor U28227 (N_28227,N_22449,N_21853);
or U28228 (N_28228,N_18435,N_21975);
nand U28229 (N_28229,N_22248,N_20461);
or U28230 (N_28230,N_18540,N_20410);
nand U28231 (N_28231,N_21313,N_18606);
xor U28232 (N_28232,N_19395,N_19578);
nor U28233 (N_28233,N_18528,N_23798);
xnor U28234 (N_28234,N_23948,N_20878);
or U28235 (N_28235,N_20318,N_19100);
and U28236 (N_28236,N_20938,N_22623);
nand U28237 (N_28237,N_23946,N_19328);
nand U28238 (N_28238,N_21092,N_19877);
xnor U28239 (N_28239,N_18327,N_21385);
and U28240 (N_28240,N_20436,N_19379);
xor U28241 (N_28241,N_18896,N_18518);
nor U28242 (N_28242,N_18429,N_23777);
and U28243 (N_28243,N_18419,N_19246);
nand U28244 (N_28244,N_20228,N_20588);
nor U28245 (N_28245,N_18482,N_18595);
and U28246 (N_28246,N_22618,N_22974);
and U28247 (N_28247,N_19655,N_19040);
or U28248 (N_28248,N_19646,N_21951);
xnor U28249 (N_28249,N_21536,N_20063);
nor U28250 (N_28250,N_23189,N_18540);
nand U28251 (N_28251,N_21404,N_22424);
and U28252 (N_28252,N_21923,N_21303);
and U28253 (N_28253,N_18718,N_23606);
nand U28254 (N_28254,N_23747,N_22075);
nor U28255 (N_28255,N_21314,N_19926);
or U28256 (N_28256,N_23978,N_18173);
nor U28257 (N_28257,N_20095,N_21036);
nor U28258 (N_28258,N_18036,N_20194);
nand U28259 (N_28259,N_22491,N_22926);
and U28260 (N_28260,N_19499,N_22333);
nor U28261 (N_28261,N_22954,N_18260);
nor U28262 (N_28262,N_18530,N_21920);
and U28263 (N_28263,N_23883,N_21592);
xor U28264 (N_28264,N_19446,N_23082);
and U28265 (N_28265,N_18697,N_22728);
nand U28266 (N_28266,N_21752,N_19845);
or U28267 (N_28267,N_20219,N_19888);
nor U28268 (N_28268,N_19609,N_20270);
nand U28269 (N_28269,N_20353,N_21766);
or U28270 (N_28270,N_19313,N_18795);
xor U28271 (N_28271,N_23241,N_22944);
or U28272 (N_28272,N_18834,N_18099);
xnor U28273 (N_28273,N_22784,N_18142);
nand U28274 (N_28274,N_18526,N_21751);
nor U28275 (N_28275,N_21479,N_19905);
and U28276 (N_28276,N_22482,N_19148);
or U28277 (N_28277,N_23399,N_23437);
xnor U28278 (N_28278,N_22458,N_20926);
nand U28279 (N_28279,N_21189,N_18862);
nand U28280 (N_28280,N_22377,N_20997);
and U28281 (N_28281,N_22491,N_19721);
xnor U28282 (N_28282,N_23015,N_18965);
nor U28283 (N_28283,N_18020,N_21965);
xor U28284 (N_28284,N_22340,N_20250);
and U28285 (N_28285,N_21678,N_19236);
nand U28286 (N_28286,N_19344,N_22758);
nor U28287 (N_28287,N_19133,N_18890);
and U28288 (N_28288,N_18511,N_19905);
and U28289 (N_28289,N_21780,N_20184);
nor U28290 (N_28290,N_20462,N_22467);
or U28291 (N_28291,N_20736,N_21666);
or U28292 (N_28292,N_19578,N_19655);
nor U28293 (N_28293,N_23535,N_18350);
and U28294 (N_28294,N_20981,N_19508);
nand U28295 (N_28295,N_23698,N_23228);
and U28296 (N_28296,N_22223,N_19152);
nand U28297 (N_28297,N_22807,N_20955);
nand U28298 (N_28298,N_20872,N_19032);
nor U28299 (N_28299,N_23152,N_18081);
xor U28300 (N_28300,N_21706,N_19759);
or U28301 (N_28301,N_23646,N_23357);
and U28302 (N_28302,N_18172,N_22371);
or U28303 (N_28303,N_20341,N_19849);
nand U28304 (N_28304,N_20713,N_22871);
nand U28305 (N_28305,N_18217,N_19829);
nor U28306 (N_28306,N_21443,N_20243);
and U28307 (N_28307,N_19220,N_22391);
nand U28308 (N_28308,N_19686,N_22824);
nand U28309 (N_28309,N_23154,N_18034);
xnor U28310 (N_28310,N_23616,N_23937);
nor U28311 (N_28311,N_19672,N_22601);
nand U28312 (N_28312,N_22701,N_18377);
nor U28313 (N_28313,N_20772,N_19029);
nor U28314 (N_28314,N_19808,N_21368);
and U28315 (N_28315,N_22071,N_19123);
or U28316 (N_28316,N_22040,N_23643);
nand U28317 (N_28317,N_21217,N_20414);
xnor U28318 (N_28318,N_23329,N_23026);
nand U28319 (N_28319,N_19056,N_19895);
xnor U28320 (N_28320,N_20339,N_23145);
or U28321 (N_28321,N_23730,N_18859);
nand U28322 (N_28322,N_23714,N_21150);
xnor U28323 (N_28323,N_18335,N_20292);
nand U28324 (N_28324,N_23932,N_19050);
or U28325 (N_28325,N_21204,N_23910);
or U28326 (N_28326,N_23847,N_19358);
xnor U28327 (N_28327,N_18663,N_20171);
nor U28328 (N_28328,N_19223,N_19361);
nor U28329 (N_28329,N_21183,N_19820);
nand U28330 (N_28330,N_18611,N_19382);
or U28331 (N_28331,N_20884,N_18820);
xnor U28332 (N_28332,N_21169,N_19033);
nor U28333 (N_28333,N_20120,N_21957);
nand U28334 (N_28334,N_18231,N_20664);
nand U28335 (N_28335,N_21961,N_21419);
nor U28336 (N_28336,N_22186,N_19455);
nor U28337 (N_28337,N_22127,N_20705);
xnor U28338 (N_28338,N_21503,N_19263);
xor U28339 (N_28339,N_23055,N_19319);
xnor U28340 (N_28340,N_19190,N_19182);
nor U28341 (N_28341,N_19853,N_20167);
and U28342 (N_28342,N_22242,N_20530);
nor U28343 (N_28343,N_21032,N_20774);
nand U28344 (N_28344,N_22350,N_20835);
nand U28345 (N_28345,N_22798,N_22389);
and U28346 (N_28346,N_23312,N_23243);
and U28347 (N_28347,N_22057,N_23543);
or U28348 (N_28348,N_20238,N_21078);
nand U28349 (N_28349,N_19630,N_22940);
and U28350 (N_28350,N_21836,N_21755);
or U28351 (N_28351,N_21032,N_23323);
nand U28352 (N_28352,N_21375,N_19121);
xor U28353 (N_28353,N_22175,N_19942);
nand U28354 (N_28354,N_19220,N_20388);
xor U28355 (N_28355,N_21672,N_22012);
and U28356 (N_28356,N_19988,N_21648);
xor U28357 (N_28357,N_21057,N_22694);
and U28358 (N_28358,N_19988,N_18708);
and U28359 (N_28359,N_18876,N_19289);
xor U28360 (N_28360,N_18623,N_22532);
and U28361 (N_28361,N_19849,N_18898);
nor U28362 (N_28362,N_23279,N_21999);
and U28363 (N_28363,N_19864,N_20743);
xnor U28364 (N_28364,N_20353,N_21110);
or U28365 (N_28365,N_22534,N_18783);
or U28366 (N_28366,N_21790,N_21087);
or U28367 (N_28367,N_20551,N_23323);
and U28368 (N_28368,N_19967,N_18032);
nor U28369 (N_28369,N_21894,N_22735);
or U28370 (N_28370,N_23270,N_20630);
nand U28371 (N_28371,N_19744,N_21149);
or U28372 (N_28372,N_18451,N_18389);
nor U28373 (N_28373,N_19187,N_18033);
nand U28374 (N_28374,N_19840,N_22417);
or U28375 (N_28375,N_19190,N_19640);
and U28376 (N_28376,N_23108,N_20300);
nor U28377 (N_28377,N_18015,N_23610);
and U28378 (N_28378,N_19332,N_21153);
xor U28379 (N_28379,N_22973,N_22460);
xor U28380 (N_28380,N_21383,N_22211);
nor U28381 (N_28381,N_22878,N_21283);
or U28382 (N_28382,N_18653,N_21358);
xnor U28383 (N_28383,N_20263,N_23921);
nand U28384 (N_28384,N_21043,N_19090);
xor U28385 (N_28385,N_18826,N_18116);
nor U28386 (N_28386,N_23740,N_22573);
nor U28387 (N_28387,N_18400,N_21991);
xnor U28388 (N_28388,N_23477,N_22068);
xnor U28389 (N_28389,N_19082,N_19357);
or U28390 (N_28390,N_23851,N_20809);
nand U28391 (N_28391,N_20796,N_18598);
nand U28392 (N_28392,N_22721,N_23199);
xor U28393 (N_28393,N_21228,N_21749);
and U28394 (N_28394,N_19855,N_19226);
or U28395 (N_28395,N_23395,N_22935);
or U28396 (N_28396,N_21758,N_23403);
nor U28397 (N_28397,N_20820,N_22242);
xnor U28398 (N_28398,N_19967,N_23978);
nor U28399 (N_28399,N_20236,N_22018);
nand U28400 (N_28400,N_18192,N_23163);
and U28401 (N_28401,N_18726,N_22591);
nor U28402 (N_28402,N_23931,N_21711);
xor U28403 (N_28403,N_23670,N_21230);
nor U28404 (N_28404,N_23350,N_21396);
xnor U28405 (N_28405,N_23639,N_18573);
nor U28406 (N_28406,N_23648,N_19926);
nor U28407 (N_28407,N_23524,N_21774);
xor U28408 (N_28408,N_20817,N_20686);
or U28409 (N_28409,N_23952,N_22971);
xnor U28410 (N_28410,N_19141,N_19389);
xor U28411 (N_28411,N_23089,N_23027);
nand U28412 (N_28412,N_18997,N_19051);
or U28413 (N_28413,N_19690,N_20605);
nand U28414 (N_28414,N_20096,N_22871);
xnor U28415 (N_28415,N_23504,N_20478);
xor U28416 (N_28416,N_20959,N_18120);
nand U28417 (N_28417,N_23884,N_22718);
nand U28418 (N_28418,N_18681,N_20395);
xor U28419 (N_28419,N_18011,N_23011);
nand U28420 (N_28420,N_21094,N_20660);
nor U28421 (N_28421,N_18364,N_23091);
xnor U28422 (N_28422,N_21697,N_22843);
and U28423 (N_28423,N_23925,N_22143);
xor U28424 (N_28424,N_19286,N_23832);
xor U28425 (N_28425,N_18591,N_18636);
and U28426 (N_28426,N_23511,N_23650);
or U28427 (N_28427,N_18595,N_22240);
nand U28428 (N_28428,N_20290,N_19713);
xor U28429 (N_28429,N_20609,N_20165);
and U28430 (N_28430,N_23409,N_22358);
nor U28431 (N_28431,N_23160,N_21373);
and U28432 (N_28432,N_20775,N_19240);
nand U28433 (N_28433,N_22341,N_19078);
xnor U28434 (N_28434,N_18815,N_21731);
nand U28435 (N_28435,N_18052,N_22718);
or U28436 (N_28436,N_20104,N_20456);
xor U28437 (N_28437,N_23952,N_21450);
or U28438 (N_28438,N_19533,N_21435);
and U28439 (N_28439,N_18323,N_20199);
or U28440 (N_28440,N_22422,N_20935);
nand U28441 (N_28441,N_19389,N_18515);
and U28442 (N_28442,N_21043,N_23038);
or U28443 (N_28443,N_23732,N_23893);
nand U28444 (N_28444,N_22186,N_23907);
nand U28445 (N_28445,N_19041,N_21158);
xnor U28446 (N_28446,N_20200,N_20542);
nor U28447 (N_28447,N_20055,N_19104);
nor U28448 (N_28448,N_23950,N_23785);
and U28449 (N_28449,N_22097,N_19898);
xnor U28450 (N_28450,N_18750,N_19113);
xnor U28451 (N_28451,N_21106,N_20762);
nor U28452 (N_28452,N_22588,N_20786);
nor U28453 (N_28453,N_19714,N_20384);
nand U28454 (N_28454,N_21122,N_19705);
and U28455 (N_28455,N_18565,N_21909);
xnor U28456 (N_28456,N_21760,N_21963);
xor U28457 (N_28457,N_21393,N_19301);
nor U28458 (N_28458,N_18102,N_23659);
xor U28459 (N_28459,N_19779,N_20512);
and U28460 (N_28460,N_18010,N_22945);
xnor U28461 (N_28461,N_19166,N_19177);
or U28462 (N_28462,N_18159,N_21862);
or U28463 (N_28463,N_21668,N_21292);
nor U28464 (N_28464,N_20000,N_21350);
nand U28465 (N_28465,N_20083,N_22822);
nor U28466 (N_28466,N_22527,N_19852);
nand U28467 (N_28467,N_23317,N_19571);
nand U28468 (N_28468,N_18721,N_19641);
nor U28469 (N_28469,N_21879,N_18713);
nor U28470 (N_28470,N_22771,N_18999);
xnor U28471 (N_28471,N_22845,N_22789);
xnor U28472 (N_28472,N_19927,N_19239);
xor U28473 (N_28473,N_21257,N_20268);
and U28474 (N_28474,N_20463,N_19452);
nand U28475 (N_28475,N_23130,N_21701);
nand U28476 (N_28476,N_19603,N_23835);
and U28477 (N_28477,N_22453,N_23914);
or U28478 (N_28478,N_18960,N_20007);
nand U28479 (N_28479,N_20448,N_23873);
and U28480 (N_28480,N_18546,N_22325);
xor U28481 (N_28481,N_22464,N_22638);
or U28482 (N_28482,N_20059,N_18670);
nor U28483 (N_28483,N_22287,N_20106);
or U28484 (N_28484,N_22599,N_18109);
xor U28485 (N_28485,N_20148,N_22822);
or U28486 (N_28486,N_22482,N_22986);
and U28487 (N_28487,N_18295,N_23862);
xor U28488 (N_28488,N_22873,N_22519);
xnor U28489 (N_28489,N_23773,N_19543);
nor U28490 (N_28490,N_20321,N_19826);
or U28491 (N_28491,N_18584,N_19533);
and U28492 (N_28492,N_21607,N_23378);
nor U28493 (N_28493,N_18650,N_18027);
or U28494 (N_28494,N_20777,N_18571);
or U28495 (N_28495,N_22758,N_23743);
nor U28496 (N_28496,N_21341,N_22294);
nor U28497 (N_28497,N_18305,N_19243);
or U28498 (N_28498,N_20429,N_20168);
nor U28499 (N_28499,N_23438,N_21464);
and U28500 (N_28500,N_21207,N_23666);
nand U28501 (N_28501,N_21862,N_20310);
or U28502 (N_28502,N_21501,N_23571);
nand U28503 (N_28503,N_22291,N_21359);
nand U28504 (N_28504,N_19883,N_21468);
xnor U28505 (N_28505,N_22481,N_22868);
or U28506 (N_28506,N_23447,N_20848);
nor U28507 (N_28507,N_18434,N_21750);
xnor U28508 (N_28508,N_22193,N_21134);
nand U28509 (N_28509,N_19182,N_22013);
nor U28510 (N_28510,N_22861,N_23549);
or U28511 (N_28511,N_23633,N_20488);
and U28512 (N_28512,N_21675,N_23881);
nand U28513 (N_28513,N_22591,N_21055);
and U28514 (N_28514,N_19630,N_20278);
xnor U28515 (N_28515,N_19013,N_18174);
or U28516 (N_28516,N_19703,N_23766);
xnor U28517 (N_28517,N_18998,N_20058);
xnor U28518 (N_28518,N_22776,N_20105);
nor U28519 (N_28519,N_20312,N_19232);
nand U28520 (N_28520,N_20143,N_22745);
and U28521 (N_28521,N_20178,N_20340);
nor U28522 (N_28522,N_22676,N_20237);
nor U28523 (N_28523,N_20301,N_22571);
nand U28524 (N_28524,N_21063,N_20153);
nor U28525 (N_28525,N_20180,N_21176);
nor U28526 (N_28526,N_23852,N_20277);
and U28527 (N_28527,N_20185,N_21467);
nand U28528 (N_28528,N_23258,N_23655);
and U28529 (N_28529,N_22658,N_18277);
or U28530 (N_28530,N_22286,N_23625);
nor U28531 (N_28531,N_19348,N_19917);
or U28532 (N_28532,N_21765,N_20249);
nand U28533 (N_28533,N_23517,N_18071);
xor U28534 (N_28534,N_21912,N_18620);
nand U28535 (N_28535,N_21730,N_23243);
nand U28536 (N_28536,N_21529,N_21194);
nor U28537 (N_28537,N_22290,N_21211);
and U28538 (N_28538,N_22157,N_22822);
xnor U28539 (N_28539,N_20194,N_22711);
nand U28540 (N_28540,N_21749,N_19334);
nand U28541 (N_28541,N_21916,N_23320);
nand U28542 (N_28542,N_20638,N_18117);
nand U28543 (N_28543,N_18741,N_19627);
and U28544 (N_28544,N_23368,N_18399);
nand U28545 (N_28545,N_22813,N_18715);
or U28546 (N_28546,N_18175,N_21187);
xor U28547 (N_28547,N_19410,N_22000);
or U28548 (N_28548,N_20493,N_20500);
xnor U28549 (N_28549,N_18971,N_22165);
nand U28550 (N_28550,N_18504,N_19999);
or U28551 (N_28551,N_19494,N_23821);
and U28552 (N_28552,N_23487,N_22314);
or U28553 (N_28553,N_21833,N_21122);
nand U28554 (N_28554,N_19282,N_23107);
xnor U28555 (N_28555,N_20504,N_20939);
nand U28556 (N_28556,N_22079,N_18339);
xnor U28557 (N_28557,N_20137,N_23973);
and U28558 (N_28558,N_19179,N_20782);
and U28559 (N_28559,N_20874,N_19669);
xor U28560 (N_28560,N_21191,N_18748);
nand U28561 (N_28561,N_21431,N_20421);
and U28562 (N_28562,N_23284,N_18643);
nor U28563 (N_28563,N_21924,N_22769);
nand U28564 (N_28564,N_22637,N_21852);
and U28565 (N_28565,N_19917,N_18316);
nor U28566 (N_28566,N_18303,N_21629);
xnor U28567 (N_28567,N_19160,N_22800);
nand U28568 (N_28568,N_23937,N_20554);
nor U28569 (N_28569,N_20061,N_20610);
or U28570 (N_28570,N_23617,N_20877);
and U28571 (N_28571,N_18141,N_19021);
or U28572 (N_28572,N_18353,N_21766);
or U28573 (N_28573,N_20646,N_21963);
and U28574 (N_28574,N_18251,N_22250);
or U28575 (N_28575,N_22548,N_19781);
xnor U28576 (N_28576,N_22929,N_22569);
nand U28577 (N_28577,N_20129,N_21566);
xor U28578 (N_28578,N_23208,N_22997);
xnor U28579 (N_28579,N_23876,N_23713);
xnor U28580 (N_28580,N_21954,N_19393);
xor U28581 (N_28581,N_20263,N_23796);
or U28582 (N_28582,N_19720,N_22624);
nand U28583 (N_28583,N_20512,N_20854);
xnor U28584 (N_28584,N_19857,N_18081);
or U28585 (N_28585,N_22568,N_20900);
xor U28586 (N_28586,N_20168,N_20484);
nand U28587 (N_28587,N_22018,N_22282);
nand U28588 (N_28588,N_20627,N_18481);
nor U28589 (N_28589,N_20036,N_19889);
nand U28590 (N_28590,N_23794,N_18857);
nor U28591 (N_28591,N_19528,N_22191);
nand U28592 (N_28592,N_20499,N_19075);
xor U28593 (N_28593,N_21711,N_18884);
nor U28594 (N_28594,N_20532,N_22361);
nand U28595 (N_28595,N_22982,N_21889);
nand U28596 (N_28596,N_23957,N_21239);
nor U28597 (N_28597,N_23976,N_18573);
nor U28598 (N_28598,N_23288,N_20079);
or U28599 (N_28599,N_18093,N_22582);
or U28600 (N_28600,N_19158,N_19519);
nand U28601 (N_28601,N_21803,N_20027);
and U28602 (N_28602,N_20208,N_21768);
nor U28603 (N_28603,N_19459,N_20533);
nand U28604 (N_28604,N_18766,N_19076);
or U28605 (N_28605,N_22644,N_23152);
nor U28606 (N_28606,N_23976,N_20500);
xor U28607 (N_28607,N_20542,N_23029);
xor U28608 (N_28608,N_21147,N_23732);
xor U28609 (N_28609,N_23972,N_22985);
and U28610 (N_28610,N_18989,N_22099);
or U28611 (N_28611,N_21970,N_22847);
nand U28612 (N_28612,N_20641,N_20031);
xor U28613 (N_28613,N_21218,N_21949);
and U28614 (N_28614,N_18843,N_19990);
or U28615 (N_28615,N_19979,N_18474);
nor U28616 (N_28616,N_20749,N_23053);
nor U28617 (N_28617,N_22338,N_20305);
xnor U28618 (N_28618,N_23985,N_20380);
nor U28619 (N_28619,N_19432,N_23630);
or U28620 (N_28620,N_23767,N_21845);
xnor U28621 (N_28621,N_20394,N_20758);
nor U28622 (N_28622,N_22339,N_22331);
or U28623 (N_28623,N_19973,N_23577);
nand U28624 (N_28624,N_20089,N_19045);
nor U28625 (N_28625,N_19792,N_19871);
and U28626 (N_28626,N_19813,N_19889);
xnor U28627 (N_28627,N_18848,N_21691);
nand U28628 (N_28628,N_23714,N_19045);
or U28629 (N_28629,N_19138,N_22476);
or U28630 (N_28630,N_21423,N_18261);
xor U28631 (N_28631,N_18075,N_20232);
and U28632 (N_28632,N_22635,N_21160);
xnor U28633 (N_28633,N_21070,N_18208);
nand U28634 (N_28634,N_21516,N_23554);
and U28635 (N_28635,N_18160,N_21131);
nor U28636 (N_28636,N_22371,N_21555);
and U28637 (N_28637,N_19767,N_18035);
xnor U28638 (N_28638,N_20655,N_22546);
nand U28639 (N_28639,N_18619,N_21893);
xnor U28640 (N_28640,N_19021,N_20354);
xor U28641 (N_28641,N_20155,N_23098);
nor U28642 (N_28642,N_18978,N_18240);
and U28643 (N_28643,N_23948,N_22410);
or U28644 (N_28644,N_20836,N_21258);
nand U28645 (N_28645,N_19447,N_18788);
and U28646 (N_28646,N_21786,N_19952);
nand U28647 (N_28647,N_22874,N_22280);
nor U28648 (N_28648,N_22589,N_20635);
or U28649 (N_28649,N_22194,N_19287);
or U28650 (N_28650,N_20791,N_23440);
xor U28651 (N_28651,N_21511,N_21172);
and U28652 (N_28652,N_19411,N_20394);
nor U28653 (N_28653,N_23107,N_20218);
or U28654 (N_28654,N_20872,N_22189);
or U28655 (N_28655,N_21445,N_22242);
or U28656 (N_28656,N_23650,N_19953);
and U28657 (N_28657,N_21965,N_18540);
nand U28658 (N_28658,N_21734,N_19526);
xnor U28659 (N_28659,N_23217,N_18022);
xor U28660 (N_28660,N_19803,N_18551);
nor U28661 (N_28661,N_22129,N_23071);
or U28662 (N_28662,N_23856,N_22455);
and U28663 (N_28663,N_23114,N_20640);
or U28664 (N_28664,N_18638,N_23403);
and U28665 (N_28665,N_21987,N_22209);
or U28666 (N_28666,N_23802,N_22413);
xnor U28667 (N_28667,N_23315,N_19952);
and U28668 (N_28668,N_21162,N_20397);
nand U28669 (N_28669,N_21532,N_22977);
xor U28670 (N_28670,N_23915,N_22436);
and U28671 (N_28671,N_22314,N_18243);
xor U28672 (N_28672,N_19410,N_22052);
nand U28673 (N_28673,N_19255,N_21856);
and U28674 (N_28674,N_21637,N_20855);
or U28675 (N_28675,N_19111,N_20097);
nand U28676 (N_28676,N_18939,N_22491);
nor U28677 (N_28677,N_19785,N_22472);
or U28678 (N_28678,N_22694,N_18851);
xor U28679 (N_28679,N_18524,N_18208);
nor U28680 (N_28680,N_22657,N_18399);
nand U28681 (N_28681,N_19665,N_22442);
nand U28682 (N_28682,N_19021,N_22431);
xor U28683 (N_28683,N_23547,N_20621);
nand U28684 (N_28684,N_21066,N_22950);
nor U28685 (N_28685,N_23013,N_19187);
nor U28686 (N_28686,N_22220,N_19610);
xor U28687 (N_28687,N_19327,N_21508);
nand U28688 (N_28688,N_23553,N_18520);
or U28689 (N_28689,N_19373,N_21252);
or U28690 (N_28690,N_20515,N_19698);
nor U28691 (N_28691,N_23776,N_22553);
or U28692 (N_28692,N_23524,N_20645);
xnor U28693 (N_28693,N_23105,N_22035);
or U28694 (N_28694,N_22780,N_22059);
or U28695 (N_28695,N_18875,N_19697);
nor U28696 (N_28696,N_18136,N_18884);
and U28697 (N_28697,N_21335,N_22933);
nand U28698 (N_28698,N_22088,N_20652);
xnor U28699 (N_28699,N_19448,N_23082);
nand U28700 (N_28700,N_23165,N_23153);
nand U28701 (N_28701,N_21791,N_23138);
nor U28702 (N_28702,N_22829,N_20842);
and U28703 (N_28703,N_22935,N_22224);
nand U28704 (N_28704,N_19232,N_20582);
nand U28705 (N_28705,N_19165,N_19097);
or U28706 (N_28706,N_21559,N_23020);
nor U28707 (N_28707,N_23770,N_23830);
and U28708 (N_28708,N_23233,N_21053);
nand U28709 (N_28709,N_22611,N_20776);
xor U28710 (N_28710,N_18760,N_19275);
and U28711 (N_28711,N_18651,N_18472);
nand U28712 (N_28712,N_20828,N_18745);
xnor U28713 (N_28713,N_18316,N_20390);
or U28714 (N_28714,N_20212,N_18520);
nor U28715 (N_28715,N_19293,N_23904);
nand U28716 (N_28716,N_18573,N_19307);
xor U28717 (N_28717,N_23256,N_21809);
nor U28718 (N_28718,N_21838,N_21553);
or U28719 (N_28719,N_23665,N_22406);
or U28720 (N_28720,N_22180,N_22061);
xor U28721 (N_28721,N_23041,N_23721);
xor U28722 (N_28722,N_21493,N_22597);
xor U28723 (N_28723,N_21660,N_19331);
nand U28724 (N_28724,N_23661,N_20251);
xor U28725 (N_28725,N_22268,N_23461);
or U28726 (N_28726,N_21862,N_18595);
or U28727 (N_28727,N_20422,N_23548);
or U28728 (N_28728,N_23007,N_23474);
nor U28729 (N_28729,N_22141,N_18965);
and U28730 (N_28730,N_22475,N_20960);
xnor U28731 (N_28731,N_22246,N_20348);
nand U28732 (N_28732,N_22068,N_23721);
xor U28733 (N_28733,N_23889,N_21317);
nor U28734 (N_28734,N_23229,N_18007);
nor U28735 (N_28735,N_21284,N_23823);
or U28736 (N_28736,N_20266,N_18745);
xor U28737 (N_28737,N_23838,N_23048);
or U28738 (N_28738,N_22590,N_19131);
or U28739 (N_28739,N_22796,N_20462);
and U28740 (N_28740,N_20357,N_18167);
nor U28741 (N_28741,N_22604,N_22636);
and U28742 (N_28742,N_23041,N_21005);
nor U28743 (N_28743,N_21742,N_19369);
and U28744 (N_28744,N_20480,N_22874);
xor U28745 (N_28745,N_21919,N_19378);
or U28746 (N_28746,N_20163,N_21295);
and U28747 (N_28747,N_23485,N_20651);
xor U28748 (N_28748,N_20387,N_19372);
or U28749 (N_28749,N_19076,N_21784);
nand U28750 (N_28750,N_22548,N_19784);
nand U28751 (N_28751,N_21359,N_22249);
nor U28752 (N_28752,N_18765,N_23071);
nand U28753 (N_28753,N_23735,N_23161);
and U28754 (N_28754,N_20733,N_22306);
nor U28755 (N_28755,N_22496,N_22073);
or U28756 (N_28756,N_21504,N_18820);
and U28757 (N_28757,N_18984,N_22105);
nor U28758 (N_28758,N_18475,N_18828);
and U28759 (N_28759,N_19002,N_21656);
and U28760 (N_28760,N_19374,N_19749);
and U28761 (N_28761,N_21170,N_20411);
and U28762 (N_28762,N_19378,N_21865);
nand U28763 (N_28763,N_21156,N_23523);
or U28764 (N_28764,N_21454,N_19500);
and U28765 (N_28765,N_22532,N_18717);
xnor U28766 (N_28766,N_19356,N_18114);
or U28767 (N_28767,N_19783,N_19405);
or U28768 (N_28768,N_23786,N_23151);
nor U28769 (N_28769,N_18200,N_18761);
xnor U28770 (N_28770,N_23809,N_22658);
xnor U28771 (N_28771,N_23556,N_18768);
nand U28772 (N_28772,N_23551,N_23200);
nand U28773 (N_28773,N_19439,N_19369);
nor U28774 (N_28774,N_19708,N_23425);
nand U28775 (N_28775,N_23703,N_21497);
nand U28776 (N_28776,N_20843,N_20019);
and U28777 (N_28777,N_23847,N_23465);
xnor U28778 (N_28778,N_23609,N_22044);
or U28779 (N_28779,N_19539,N_19389);
and U28780 (N_28780,N_22719,N_19327);
and U28781 (N_28781,N_19728,N_22929);
xor U28782 (N_28782,N_23203,N_20630);
xnor U28783 (N_28783,N_22871,N_21597);
nor U28784 (N_28784,N_22751,N_23754);
xor U28785 (N_28785,N_23777,N_18929);
nand U28786 (N_28786,N_18127,N_22893);
and U28787 (N_28787,N_19258,N_19745);
and U28788 (N_28788,N_19686,N_22495);
nand U28789 (N_28789,N_23033,N_23622);
nand U28790 (N_28790,N_18005,N_19540);
and U28791 (N_28791,N_18095,N_20527);
nand U28792 (N_28792,N_22784,N_18264);
or U28793 (N_28793,N_23833,N_23894);
and U28794 (N_28794,N_22689,N_20267);
nand U28795 (N_28795,N_23613,N_21259);
xnor U28796 (N_28796,N_21800,N_22814);
nand U28797 (N_28797,N_18327,N_22974);
xnor U28798 (N_28798,N_23563,N_22428);
nor U28799 (N_28799,N_22259,N_20507);
nor U28800 (N_28800,N_21941,N_20639);
nor U28801 (N_28801,N_18303,N_19154);
and U28802 (N_28802,N_23214,N_23196);
xnor U28803 (N_28803,N_19639,N_21535);
and U28804 (N_28804,N_19006,N_19090);
xor U28805 (N_28805,N_19151,N_19105);
nand U28806 (N_28806,N_19718,N_21274);
and U28807 (N_28807,N_19933,N_20213);
nand U28808 (N_28808,N_18014,N_18855);
and U28809 (N_28809,N_22928,N_22638);
and U28810 (N_28810,N_20369,N_22329);
nand U28811 (N_28811,N_23289,N_23342);
nand U28812 (N_28812,N_21442,N_21308);
nand U28813 (N_28813,N_23425,N_19601);
xnor U28814 (N_28814,N_22624,N_21479);
and U28815 (N_28815,N_21316,N_22726);
nor U28816 (N_28816,N_19200,N_20701);
nand U28817 (N_28817,N_19401,N_23265);
nand U28818 (N_28818,N_21339,N_23906);
xnor U28819 (N_28819,N_20643,N_23201);
nor U28820 (N_28820,N_22066,N_18641);
nor U28821 (N_28821,N_22027,N_22882);
or U28822 (N_28822,N_23275,N_22199);
nor U28823 (N_28823,N_18001,N_20163);
or U28824 (N_28824,N_23924,N_19418);
and U28825 (N_28825,N_23198,N_21990);
xnor U28826 (N_28826,N_21752,N_23726);
nand U28827 (N_28827,N_20173,N_21813);
nand U28828 (N_28828,N_18457,N_20960);
xor U28829 (N_28829,N_21577,N_22800);
xor U28830 (N_28830,N_19556,N_18760);
xnor U28831 (N_28831,N_22944,N_21474);
and U28832 (N_28832,N_21412,N_22731);
or U28833 (N_28833,N_18017,N_23032);
nor U28834 (N_28834,N_22253,N_23102);
nor U28835 (N_28835,N_21825,N_22126);
and U28836 (N_28836,N_19961,N_18404);
nor U28837 (N_28837,N_20472,N_22563);
nand U28838 (N_28838,N_20820,N_23897);
xor U28839 (N_28839,N_23773,N_21415);
or U28840 (N_28840,N_18250,N_21613);
xnor U28841 (N_28841,N_19629,N_21595);
xor U28842 (N_28842,N_22353,N_18010);
and U28843 (N_28843,N_18714,N_21205);
nor U28844 (N_28844,N_19627,N_18883);
or U28845 (N_28845,N_21816,N_23663);
xor U28846 (N_28846,N_22116,N_20186);
xor U28847 (N_28847,N_22958,N_19170);
and U28848 (N_28848,N_20691,N_23360);
nand U28849 (N_28849,N_22428,N_18204);
or U28850 (N_28850,N_18910,N_23651);
or U28851 (N_28851,N_19151,N_21005);
xor U28852 (N_28852,N_22333,N_20943);
and U28853 (N_28853,N_23645,N_18560);
and U28854 (N_28854,N_23957,N_21285);
nand U28855 (N_28855,N_19988,N_22440);
nor U28856 (N_28856,N_23351,N_23541);
xor U28857 (N_28857,N_20988,N_20167);
nand U28858 (N_28858,N_23766,N_19681);
or U28859 (N_28859,N_20094,N_23888);
xor U28860 (N_28860,N_22904,N_19775);
or U28861 (N_28861,N_18505,N_20047);
xnor U28862 (N_28862,N_20654,N_22097);
xnor U28863 (N_28863,N_21647,N_21640);
nand U28864 (N_28864,N_23157,N_20209);
nor U28865 (N_28865,N_20203,N_20622);
and U28866 (N_28866,N_23355,N_21696);
nor U28867 (N_28867,N_23002,N_22176);
and U28868 (N_28868,N_20619,N_20097);
and U28869 (N_28869,N_21657,N_18299);
or U28870 (N_28870,N_19628,N_22965);
or U28871 (N_28871,N_22858,N_18478);
nor U28872 (N_28872,N_22877,N_23050);
nand U28873 (N_28873,N_22206,N_19716);
or U28874 (N_28874,N_20247,N_21211);
nand U28875 (N_28875,N_18068,N_21474);
nor U28876 (N_28876,N_21067,N_22004);
and U28877 (N_28877,N_22604,N_18652);
xor U28878 (N_28878,N_19958,N_23879);
nand U28879 (N_28879,N_22881,N_20326);
nand U28880 (N_28880,N_21156,N_22989);
nand U28881 (N_28881,N_22110,N_20593);
and U28882 (N_28882,N_19209,N_19274);
or U28883 (N_28883,N_23922,N_21449);
and U28884 (N_28884,N_22720,N_20047);
xor U28885 (N_28885,N_18025,N_21779);
nor U28886 (N_28886,N_23887,N_23480);
xnor U28887 (N_28887,N_18993,N_19253);
nor U28888 (N_28888,N_22236,N_22412);
nand U28889 (N_28889,N_23982,N_21495);
xor U28890 (N_28890,N_19911,N_20534);
or U28891 (N_28891,N_20400,N_19548);
nor U28892 (N_28892,N_22707,N_23140);
and U28893 (N_28893,N_23352,N_19484);
or U28894 (N_28894,N_22096,N_19213);
nor U28895 (N_28895,N_22364,N_23292);
and U28896 (N_28896,N_23644,N_19682);
nor U28897 (N_28897,N_21780,N_23591);
xnor U28898 (N_28898,N_18927,N_19189);
or U28899 (N_28899,N_23499,N_23636);
or U28900 (N_28900,N_21378,N_21794);
or U28901 (N_28901,N_23033,N_18856);
nand U28902 (N_28902,N_20553,N_20305);
nand U28903 (N_28903,N_20528,N_18808);
xor U28904 (N_28904,N_18861,N_23986);
xor U28905 (N_28905,N_18007,N_20052);
nand U28906 (N_28906,N_18847,N_18444);
and U28907 (N_28907,N_20385,N_22389);
or U28908 (N_28908,N_18745,N_23592);
and U28909 (N_28909,N_23710,N_19264);
xor U28910 (N_28910,N_20773,N_22065);
xor U28911 (N_28911,N_22317,N_20551);
nand U28912 (N_28912,N_23345,N_19952);
nand U28913 (N_28913,N_18195,N_20889);
xnor U28914 (N_28914,N_21108,N_22191);
and U28915 (N_28915,N_23592,N_18800);
nor U28916 (N_28916,N_22287,N_19218);
or U28917 (N_28917,N_18250,N_23810);
nand U28918 (N_28918,N_20969,N_19557);
nand U28919 (N_28919,N_23546,N_19470);
and U28920 (N_28920,N_22962,N_20159);
nand U28921 (N_28921,N_23326,N_19582);
nor U28922 (N_28922,N_18313,N_18607);
or U28923 (N_28923,N_21268,N_23990);
nor U28924 (N_28924,N_21995,N_20074);
nor U28925 (N_28925,N_18172,N_21222);
xnor U28926 (N_28926,N_19528,N_20098);
and U28927 (N_28927,N_21148,N_22441);
xor U28928 (N_28928,N_21193,N_19991);
nand U28929 (N_28929,N_18504,N_23631);
nand U28930 (N_28930,N_23386,N_22936);
xor U28931 (N_28931,N_20635,N_23692);
nor U28932 (N_28932,N_22222,N_23790);
and U28933 (N_28933,N_23414,N_21425);
and U28934 (N_28934,N_23284,N_23382);
nor U28935 (N_28935,N_20344,N_22988);
or U28936 (N_28936,N_19670,N_19996);
nor U28937 (N_28937,N_19850,N_23543);
or U28938 (N_28938,N_18084,N_18011);
nand U28939 (N_28939,N_22225,N_23899);
xor U28940 (N_28940,N_22652,N_21958);
nand U28941 (N_28941,N_20495,N_18207);
nor U28942 (N_28942,N_22774,N_21299);
nand U28943 (N_28943,N_23070,N_23554);
xor U28944 (N_28944,N_23692,N_23351);
and U28945 (N_28945,N_19695,N_18941);
and U28946 (N_28946,N_22466,N_18512);
xnor U28947 (N_28947,N_21518,N_21271);
or U28948 (N_28948,N_19664,N_19548);
xnor U28949 (N_28949,N_18009,N_21349);
nor U28950 (N_28950,N_19703,N_23496);
nor U28951 (N_28951,N_22978,N_21142);
nand U28952 (N_28952,N_23867,N_18326);
nor U28953 (N_28953,N_20505,N_22321);
nor U28954 (N_28954,N_19011,N_19427);
and U28955 (N_28955,N_20013,N_20234);
nand U28956 (N_28956,N_23879,N_21913);
nand U28957 (N_28957,N_18573,N_18142);
and U28958 (N_28958,N_22404,N_19069);
xnor U28959 (N_28959,N_22115,N_18904);
and U28960 (N_28960,N_18594,N_21158);
nand U28961 (N_28961,N_19636,N_20460);
nand U28962 (N_28962,N_18995,N_22033);
xor U28963 (N_28963,N_23597,N_22378);
nor U28964 (N_28964,N_18250,N_18723);
nor U28965 (N_28965,N_19152,N_21272);
xnor U28966 (N_28966,N_18639,N_21075);
or U28967 (N_28967,N_23886,N_23026);
and U28968 (N_28968,N_23215,N_22069);
or U28969 (N_28969,N_20742,N_19336);
or U28970 (N_28970,N_19498,N_21515);
xnor U28971 (N_28971,N_22352,N_18259);
nand U28972 (N_28972,N_18606,N_18042);
xor U28973 (N_28973,N_18469,N_19045);
and U28974 (N_28974,N_18264,N_19504);
or U28975 (N_28975,N_23059,N_22606);
and U28976 (N_28976,N_23160,N_23869);
and U28977 (N_28977,N_22441,N_23177);
nand U28978 (N_28978,N_20128,N_23736);
nand U28979 (N_28979,N_23843,N_21180);
nand U28980 (N_28980,N_21157,N_22968);
nor U28981 (N_28981,N_20126,N_23033);
and U28982 (N_28982,N_23263,N_23897);
nor U28983 (N_28983,N_22262,N_20963);
nor U28984 (N_28984,N_21660,N_19856);
xnor U28985 (N_28985,N_22758,N_20744);
or U28986 (N_28986,N_21564,N_21656);
xor U28987 (N_28987,N_20568,N_20629);
nor U28988 (N_28988,N_18853,N_18965);
xor U28989 (N_28989,N_19091,N_21684);
nor U28990 (N_28990,N_21452,N_18506);
nor U28991 (N_28991,N_23364,N_21053);
or U28992 (N_28992,N_23752,N_20858);
nor U28993 (N_28993,N_20967,N_22238);
xor U28994 (N_28994,N_21831,N_19736);
nor U28995 (N_28995,N_21918,N_23410);
xnor U28996 (N_28996,N_23616,N_21685);
and U28997 (N_28997,N_23044,N_22631);
or U28998 (N_28998,N_22558,N_20810);
nand U28999 (N_28999,N_23909,N_19528);
and U29000 (N_29000,N_22815,N_18442);
nand U29001 (N_29001,N_22686,N_21429);
nand U29002 (N_29002,N_21199,N_18424);
or U29003 (N_29003,N_19710,N_18444);
xnor U29004 (N_29004,N_21887,N_22225);
xor U29005 (N_29005,N_18481,N_21062);
xnor U29006 (N_29006,N_22708,N_20441);
nand U29007 (N_29007,N_19579,N_23044);
xor U29008 (N_29008,N_20000,N_22498);
nor U29009 (N_29009,N_23627,N_22536);
nor U29010 (N_29010,N_23437,N_18031);
or U29011 (N_29011,N_23166,N_23794);
nand U29012 (N_29012,N_21846,N_22785);
xor U29013 (N_29013,N_18005,N_21124);
nor U29014 (N_29014,N_21166,N_22998);
nand U29015 (N_29015,N_21511,N_18996);
or U29016 (N_29016,N_18590,N_22330);
and U29017 (N_29017,N_18202,N_19195);
nand U29018 (N_29018,N_22136,N_23781);
nand U29019 (N_29019,N_23881,N_18411);
and U29020 (N_29020,N_19688,N_19181);
or U29021 (N_29021,N_22905,N_18755);
or U29022 (N_29022,N_18352,N_19721);
or U29023 (N_29023,N_18558,N_23899);
nor U29024 (N_29024,N_23196,N_19007);
and U29025 (N_29025,N_18642,N_23226);
nand U29026 (N_29026,N_18198,N_21600);
nor U29027 (N_29027,N_23838,N_22828);
xnor U29028 (N_29028,N_21591,N_22342);
nand U29029 (N_29029,N_20358,N_18716);
nand U29030 (N_29030,N_22964,N_20518);
and U29031 (N_29031,N_23741,N_19962);
or U29032 (N_29032,N_18516,N_21612);
xnor U29033 (N_29033,N_21070,N_19581);
xnor U29034 (N_29034,N_20196,N_18416);
xor U29035 (N_29035,N_23232,N_18619);
or U29036 (N_29036,N_22506,N_23032);
nand U29037 (N_29037,N_21595,N_19427);
xnor U29038 (N_29038,N_22027,N_20915);
and U29039 (N_29039,N_20791,N_20186);
xor U29040 (N_29040,N_21347,N_18986);
xor U29041 (N_29041,N_19638,N_21555);
xor U29042 (N_29042,N_20810,N_18361);
nand U29043 (N_29043,N_19053,N_21091);
and U29044 (N_29044,N_21907,N_18765);
xnor U29045 (N_29045,N_21956,N_21292);
xor U29046 (N_29046,N_19261,N_19972);
xnor U29047 (N_29047,N_20942,N_19684);
and U29048 (N_29048,N_20755,N_19962);
nand U29049 (N_29049,N_23648,N_19692);
nor U29050 (N_29050,N_18143,N_18896);
or U29051 (N_29051,N_23934,N_22499);
and U29052 (N_29052,N_20511,N_23163);
nor U29053 (N_29053,N_22320,N_23190);
and U29054 (N_29054,N_18642,N_23784);
and U29055 (N_29055,N_20815,N_18338);
and U29056 (N_29056,N_20314,N_23218);
nor U29057 (N_29057,N_21694,N_22333);
and U29058 (N_29058,N_23753,N_19749);
and U29059 (N_29059,N_21755,N_23322);
or U29060 (N_29060,N_23576,N_20454);
nor U29061 (N_29061,N_23871,N_22236);
and U29062 (N_29062,N_22004,N_19030);
xnor U29063 (N_29063,N_22842,N_18800);
nand U29064 (N_29064,N_21698,N_20334);
nor U29065 (N_29065,N_19608,N_22463);
nor U29066 (N_29066,N_22103,N_21687);
xnor U29067 (N_29067,N_19437,N_18061);
or U29068 (N_29068,N_18124,N_23702);
nand U29069 (N_29069,N_23222,N_20187);
nand U29070 (N_29070,N_19515,N_21127);
nor U29071 (N_29071,N_18846,N_22992);
xor U29072 (N_29072,N_20871,N_23079);
and U29073 (N_29073,N_21274,N_18668);
xnor U29074 (N_29074,N_22938,N_20074);
and U29075 (N_29075,N_23267,N_23228);
and U29076 (N_29076,N_18173,N_21230);
nor U29077 (N_29077,N_22881,N_20167);
or U29078 (N_29078,N_21248,N_20709);
and U29079 (N_29079,N_22502,N_21972);
nand U29080 (N_29080,N_18241,N_22604);
nand U29081 (N_29081,N_20149,N_23202);
nor U29082 (N_29082,N_23094,N_19794);
nor U29083 (N_29083,N_18738,N_18512);
nor U29084 (N_29084,N_19278,N_21317);
xor U29085 (N_29085,N_21497,N_18120);
nor U29086 (N_29086,N_18038,N_22389);
or U29087 (N_29087,N_22671,N_18717);
xor U29088 (N_29088,N_20840,N_20884);
or U29089 (N_29089,N_18269,N_22053);
and U29090 (N_29090,N_20893,N_23738);
and U29091 (N_29091,N_22073,N_20734);
and U29092 (N_29092,N_21544,N_23026);
xor U29093 (N_29093,N_18275,N_23410);
and U29094 (N_29094,N_22647,N_21461);
nor U29095 (N_29095,N_19079,N_23563);
and U29096 (N_29096,N_21207,N_19491);
xnor U29097 (N_29097,N_19993,N_23882);
or U29098 (N_29098,N_21127,N_23823);
nor U29099 (N_29099,N_19624,N_20430);
or U29100 (N_29100,N_19803,N_20070);
or U29101 (N_29101,N_18688,N_23226);
xnor U29102 (N_29102,N_23115,N_18026);
or U29103 (N_29103,N_20133,N_23974);
or U29104 (N_29104,N_23622,N_21202);
nand U29105 (N_29105,N_23587,N_22372);
nand U29106 (N_29106,N_18016,N_19554);
nor U29107 (N_29107,N_22622,N_23409);
nand U29108 (N_29108,N_22464,N_20223);
or U29109 (N_29109,N_23816,N_22280);
and U29110 (N_29110,N_20632,N_19475);
and U29111 (N_29111,N_20407,N_18368);
nor U29112 (N_29112,N_23074,N_22593);
nand U29113 (N_29113,N_18398,N_18655);
nand U29114 (N_29114,N_18408,N_19798);
or U29115 (N_29115,N_20304,N_18038);
nor U29116 (N_29116,N_22008,N_23107);
or U29117 (N_29117,N_22559,N_19475);
nor U29118 (N_29118,N_18821,N_20075);
nor U29119 (N_29119,N_22822,N_20223);
xnor U29120 (N_29120,N_20320,N_19210);
nand U29121 (N_29121,N_20428,N_23503);
nor U29122 (N_29122,N_20239,N_23737);
nor U29123 (N_29123,N_22955,N_22639);
and U29124 (N_29124,N_22474,N_22011);
xnor U29125 (N_29125,N_18698,N_20169);
nor U29126 (N_29126,N_20501,N_21465);
and U29127 (N_29127,N_20595,N_23507);
xor U29128 (N_29128,N_22743,N_22830);
and U29129 (N_29129,N_22479,N_21201);
or U29130 (N_29130,N_22904,N_20018);
or U29131 (N_29131,N_22370,N_21283);
nand U29132 (N_29132,N_22998,N_18406);
nand U29133 (N_29133,N_21129,N_18548);
xnor U29134 (N_29134,N_21235,N_21006);
nor U29135 (N_29135,N_19035,N_22145);
nand U29136 (N_29136,N_20662,N_22607);
nor U29137 (N_29137,N_21959,N_22264);
nor U29138 (N_29138,N_20422,N_23239);
and U29139 (N_29139,N_22961,N_23949);
and U29140 (N_29140,N_21536,N_23609);
or U29141 (N_29141,N_22354,N_20606);
nor U29142 (N_29142,N_20733,N_18004);
and U29143 (N_29143,N_21879,N_22070);
xnor U29144 (N_29144,N_21942,N_21748);
nand U29145 (N_29145,N_20284,N_20639);
xor U29146 (N_29146,N_22261,N_18504);
or U29147 (N_29147,N_22089,N_23890);
xnor U29148 (N_29148,N_20850,N_20553);
xnor U29149 (N_29149,N_20994,N_21373);
nand U29150 (N_29150,N_19148,N_20088);
or U29151 (N_29151,N_18909,N_21809);
and U29152 (N_29152,N_22494,N_22510);
nor U29153 (N_29153,N_20375,N_20915);
nand U29154 (N_29154,N_20607,N_19251);
xor U29155 (N_29155,N_19942,N_18539);
and U29156 (N_29156,N_18124,N_23689);
or U29157 (N_29157,N_22855,N_20710);
or U29158 (N_29158,N_18564,N_18569);
nand U29159 (N_29159,N_23499,N_21731);
or U29160 (N_29160,N_22306,N_23515);
nand U29161 (N_29161,N_22692,N_19288);
or U29162 (N_29162,N_19582,N_20448);
and U29163 (N_29163,N_21467,N_23335);
or U29164 (N_29164,N_21808,N_23183);
nor U29165 (N_29165,N_21948,N_21351);
nor U29166 (N_29166,N_20237,N_21085);
nand U29167 (N_29167,N_18872,N_21408);
xor U29168 (N_29168,N_23809,N_19917);
nand U29169 (N_29169,N_19817,N_19231);
xnor U29170 (N_29170,N_23322,N_22333);
and U29171 (N_29171,N_20326,N_23455);
and U29172 (N_29172,N_22648,N_23719);
nor U29173 (N_29173,N_23153,N_19285);
nand U29174 (N_29174,N_20851,N_23968);
xnor U29175 (N_29175,N_22332,N_20061);
or U29176 (N_29176,N_20198,N_21663);
or U29177 (N_29177,N_21424,N_20134);
and U29178 (N_29178,N_22244,N_19947);
nor U29179 (N_29179,N_18030,N_18848);
nor U29180 (N_29180,N_19366,N_19231);
nor U29181 (N_29181,N_19278,N_19990);
nor U29182 (N_29182,N_22116,N_20535);
nor U29183 (N_29183,N_18827,N_20013);
nand U29184 (N_29184,N_23676,N_22751);
or U29185 (N_29185,N_19118,N_18884);
xor U29186 (N_29186,N_20858,N_23522);
nor U29187 (N_29187,N_19610,N_20049);
xor U29188 (N_29188,N_20585,N_21110);
nor U29189 (N_29189,N_21375,N_23225);
and U29190 (N_29190,N_19828,N_19366);
or U29191 (N_29191,N_19234,N_18390);
or U29192 (N_29192,N_22249,N_21570);
nand U29193 (N_29193,N_20709,N_20317);
nand U29194 (N_29194,N_23518,N_18621);
or U29195 (N_29195,N_21242,N_21492);
xnor U29196 (N_29196,N_19756,N_21670);
nor U29197 (N_29197,N_21944,N_19507);
or U29198 (N_29198,N_18629,N_20733);
or U29199 (N_29199,N_21223,N_20068);
and U29200 (N_29200,N_23560,N_21880);
nor U29201 (N_29201,N_23964,N_19616);
nand U29202 (N_29202,N_20158,N_21679);
and U29203 (N_29203,N_19483,N_23545);
and U29204 (N_29204,N_19769,N_23392);
xor U29205 (N_29205,N_22270,N_20463);
or U29206 (N_29206,N_23905,N_23867);
or U29207 (N_29207,N_21923,N_22802);
nor U29208 (N_29208,N_23146,N_20124);
and U29209 (N_29209,N_21554,N_19093);
xnor U29210 (N_29210,N_23931,N_22089);
nand U29211 (N_29211,N_19997,N_19398);
nor U29212 (N_29212,N_21789,N_19448);
xnor U29213 (N_29213,N_20738,N_20478);
or U29214 (N_29214,N_22498,N_18120);
nand U29215 (N_29215,N_23331,N_22950);
nand U29216 (N_29216,N_23738,N_20209);
and U29217 (N_29217,N_21372,N_20867);
nor U29218 (N_29218,N_19444,N_21051);
or U29219 (N_29219,N_22757,N_19885);
xnor U29220 (N_29220,N_23105,N_22437);
or U29221 (N_29221,N_22302,N_20931);
xor U29222 (N_29222,N_19136,N_22056);
xnor U29223 (N_29223,N_23997,N_21531);
xor U29224 (N_29224,N_18527,N_21663);
nor U29225 (N_29225,N_20386,N_22287);
or U29226 (N_29226,N_19866,N_19691);
nand U29227 (N_29227,N_20354,N_19271);
and U29228 (N_29228,N_20754,N_23562);
nand U29229 (N_29229,N_22212,N_21384);
nand U29230 (N_29230,N_20337,N_23220);
or U29231 (N_29231,N_23941,N_22523);
nor U29232 (N_29232,N_20108,N_21042);
or U29233 (N_29233,N_22334,N_21777);
nand U29234 (N_29234,N_22703,N_22743);
and U29235 (N_29235,N_18075,N_18858);
xor U29236 (N_29236,N_19338,N_19607);
or U29237 (N_29237,N_22851,N_18950);
xnor U29238 (N_29238,N_19156,N_19040);
and U29239 (N_29239,N_20728,N_22056);
nor U29240 (N_29240,N_20375,N_18079);
nor U29241 (N_29241,N_23944,N_19995);
nor U29242 (N_29242,N_18021,N_23224);
nor U29243 (N_29243,N_22331,N_20364);
or U29244 (N_29244,N_23000,N_22256);
nor U29245 (N_29245,N_23999,N_18950);
nor U29246 (N_29246,N_19919,N_22054);
nor U29247 (N_29247,N_19045,N_19964);
nand U29248 (N_29248,N_19783,N_21640);
nor U29249 (N_29249,N_21054,N_19546);
nor U29250 (N_29250,N_18676,N_22598);
nor U29251 (N_29251,N_21689,N_22351);
and U29252 (N_29252,N_19222,N_23099);
xor U29253 (N_29253,N_22376,N_23173);
nor U29254 (N_29254,N_20386,N_18878);
nand U29255 (N_29255,N_21571,N_20723);
or U29256 (N_29256,N_20749,N_21812);
xnor U29257 (N_29257,N_20672,N_21985);
or U29258 (N_29258,N_19721,N_22828);
nand U29259 (N_29259,N_18476,N_19663);
nand U29260 (N_29260,N_19089,N_21375);
or U29261 (N_29261,N_18436,N_20100);
and U29262 (N_29262,N_18875,N_21810);
or U29263 (N_29263,N_19806,N_22737);
and U29264 (N_29264,N_23751,N_22778);
nand U29265 (N_29265,N_19321,N_23205);
nand U29266 (N_29266,N_19807,N_23630);
nor U29267 (N_29267,N_21593,N_21465);
and U29268 (N_29268,N_21468,N_22309);
nand U29269 (N_29269,N_22083,N_18069);
nor U29270 (N_29270,N_18208,N_20838);
or U29271 (N_29271,N_19336,N_23450);
and U29272 (N_29272,N_21049,N_21337);
or U29273 (N_29273,N_21854,N_18455);
or U29274 (N_29274,N_18456,N_23611);
or U29275 (N_29275,N_22838,N_23756);
nor U29276 (N_29276,N_23344,N_21376);
or U29277 (N_29277,N_20513,N_18980);
xor U29278 (N_29278,N_20204,N_18016);
xnor U29279 (N_29279,N_21900,N_18723);
xnor U29280 (N_29280,N_18505,N_21481);
xor U29281 (N_29281,N_21565,N_20045);
or U29282 (N_29282,N_18375,N_19818);
and U29283 (N_29283,N_21381,N_22356);
and U29284 (N_29284,N_20159,N_20609);
nor U29285 (N_29285,N_21957,N_23266);
xor U29286 (N_29286,N_21839,N_22528);
or U29287 (N_29287,N_18748,N_18999);
nor U29288 (N_29288,N_18250,N_22119);
xor U29289 (N_29289,N_21388,N_18042);
and U29290 (N_29290,N_20791,N_22201);
nand U29291 (N_29291,N_22205,N_20773);
xor U29292 (N_29292,N_18999,N_19576);
or U29293 (N_29293,N_22419,N_20368);
xnor U29294 (N_29294,N_20317,N_20179);
nand U29295 (N_29295,N_20588,N_19947);
xor U29296 (N_29296,N_18357,N_20040);
or U29297 (N_29297,N_20212,N_18996);
xnor U29298 (N_29298,N_23042,N_19226);
or U29299 (N_29299,N_23972,N_23084);
nand U29300 (N_29300,N_20854,N_20618);
nand U29301 (N_29301,N_18287,N_22216);
nor U29302 (N_29302,N_19312,N_20726);
and U29303 (N_29303,N_23172,N_23129);
and U29304 (N_29304,N_21677,N_18507);
nand U29305 (N_29305,N_19801,N_18210);
nor U29306 (N_29306,N_21326,N_18158);
nor U29307 (N_29307,N_20581,N_19392);
xnor U29308 (N_29308,N_23517,N_20671);
nand U29309 (N_29309,N_22213,N_20369);
and U29310 (N_29310,N_23452,N_23905);
nand U29311 (N_29311,N_18275,N_18118);
or U29312 (N_29312,N_21044,N_19093);
xor U29313 (N_29313,N_22560,N_21351);
and U29314 (N_29314,N_20110,N_23245);
or U29315 (N_29315,N_21575,N_21456);
nor U29316 (N_29316,N_18604,N_21920);
nor U29317 (N_29317,N_19025,N_18896);
xnor U29318 (N_29318,N_18368,N_19702);
or U29319 (N_29319,N_22803,N_18198);
xnor U29320 (N_29320,N_19389,N_21070);
and U29321 (N_29321,N_18596,N_23851);
nand U29322 (N_29322,N_22057,N_22110);
xnor U29323 (N_29323,N_21888,N_19289);
nand U29324 (N_29324,N_20268,N_21169);
nand U29325 (N_29325,N_22085,N_23260);
nor U29326 (N_29326,N_19955,N_18767);
and U29327 (N_29327,N_21953,N_20516);
nand U29328 (N_29328,N_18668,N_23415);
and U29329 (N_29329,N_20961,N_22131);
nand U29330 (N_29330,N_21791,N_18173);
xnor U29331 (N_29331,N_22707,N_23101);
nor U29332 (N_29332,N_19941,N_19083);
nand U29333 (N_29333,N_23001,N_20908);
or U29334 (N_29334,N_23679,N_18619);
nand U29335 (N_29335,N_22192,N_19308);
nand U29336 (N_29336,N_22662,N_20733);
and U29337 (N_29337,N_20067,N_19637);
or U29338 (N_29338,N_19249,N_22157);
nor U29339 (N_29339,N_22840,N_22658);
nor U29340 (N_29340,N_20397,N_19461);
xnor U29341 (N_29341,N_23735,N_20259);
and U29342 (N_29342,N_21618,N_19832);
nand U29343 (N_29343,N_18336,N_18007);
or U29344 (N_29344,N_22286,N_22788);
nor U29345 (N_29345,N_18294,N_23021);
or U29346 (N_29346,N_23922,N_23238);
nor U29347 (N_29347,N_19094,N_20066);
xor U29348 (N_29348,N_23860,N_23596);
nor U29349 (N_29349,N_21547,N_22555);
xnor U29350 (N_29350,N_18629,N_19286);
and U29351 (N_29351,N_20566,N_18019);
or U29352 (N_29352,N_19268,N_23318);
or U29353 (N_29353,N_20739,N_18876);
xor U29354 (N_29354,N_18581,N_21838);
xnor U29355 (N_29355,N_22503,N_19825);
xor U29356 (N_29356,N_19440,N_19225);
nor U29357 (N_29357,N_19663,N_20969);
or U29358 (N_29358,N_20473,N_22479);
xor U29359 (N_29359,N_20883,N_21046);
nand U29360 (N_29360,N_20242,N_18589);
or U29361 (N_29361,N_21220,N_18354);
or U29362 (N_29362,N_23736,N_18573);
and U29363 (N_29363,N_23388,N_19290);
or U29364 (N_29364,N_21543,N_19007);
nor U29365 (N_29365,N_22306,N_23563);
nand U29366 (N_29366,N_23644,N_19386);
and U29367 (N_29367,N_20214,N_21002);
xor U29368 (N_29368,N_23398,N_23238);
and U29369 (N_29369,N_22568,N_19000);
nand U29370 (N_29370,N_18926,N_23098);
nand U29371 (N_29371,N_18446,N_23931);
xor U29372 (N_29372,N_18682,N_21408);
and U29373 (N_29373,N_21087,N_20836);
xnor U29374 (N_29374,N_22749,N_18807);
nor U29375 (N_29375,N_21177,N_22011);
or U29376 (N_29376,N_20582,N_23514);
xnor U29377 (N_29377,N_19664,N_19244);
or U29378 (N_29378,N_18653,N_22121);
nand U29379 (N_29379,N_21480,N_20749);
and U29380 (N_29380,N_20456,N_22898);
nand U29381 (N_29381,N_23587,N_18427);
nand U29382 (N_29382,N_23336,N_21965);
or U29383 (N_29383,N_19360,N_19255);
xnor U29384 (N_29384,N_19774,N_23918);
and U29385 (N_29385,N_23238,N_18574);
and U29386 (N_29386,N_20962,N_18696);
nor U29387 (N_29387,N_20992,N_20723);
nor U29388 (N_29388,N_19070,N_23917);
or U29389 (N_29389,N_23751,N_18155);
nor U29390 (N_29390,N_23376,N_18699);
and U29391 (N_29391,N_21592,N_18878);
or U29392 (N_29392,N_22593,N_19152);
or U29393 (N_29393,N_20881,N_23326);
or U29394 (N_29394,N_19006,N_20667);
or U29395 (N_29395,N_18505,N_22305);
xnor U29396 (N_29396,N_19358,N_20786);
xor U29397 (N_29397,N_18337,N_18886);
xor U29398 (N_29398,N_20026,N_23713);
nand U29399 (N_29399,N_23310,N_20476);
and U29400 (N_29400,N_19299,N_19860);
and U29401 (N_29401,N_21368,N_18552);
or U29402 (N_29402,N_19172,N_20229);
and U29403 (N_29403,N_20730,N_18866);
nor U29404 (N_29404,N_22388,N_19734);
or U29405 (N_29405,N_21991,N_23800);
nor U29406 (N_29406,N_20102,N_18978);
nand U29407 (N_29407,N_18590,N_19779);
nor U29408 (N_29408,N_18166,N_23063);
and U29409 (N_29409,N_23457,N_22502);
nand U29410 (N_29410,N_19705,N_18866);
nor U29411 (N_29411,N_18817,N_19547);
xnor U29412 (N_29412,N_21653,N_19254);
xor U29413 (N_29413,N_18146,N_19436);
xnor U29414 (N_29414,N_21396,N_20762);
xnor U29415 (N_29415,N_18200,N_19790);
or U29416 (N_29416,N_23514,N_21526);
and U29417 (N_29417,N_22758,N_22505);
nor U29418 (N_29418,N_23411,N_19947);
xor U29419 (N_29419,N_18004,N_21796);
nand U29420 (N_29420,N_22065,N_21977);
and U29421 (N_29421,N_19873,N_21256);
and U29422 (N_29422,N_18668,N_20931);
or U29423 (N_29423,N_23632,N_19389);
and U29424 (N_29424,N_21460,N_22500);
or U29425 (N_29425,N_18274,N_18567);
nand U29426 (N_29426,N_18665,N_20426);
nor U29427 (N_29427,N_22591,N_21419);
and U29428 (N_29428,N_19655,N_23602);
and U29429 (N_29429,N_22340,N_23856);
and U29430 (N_29430,N_19132,N_19647);
and U29431 (N_29431,N_23543,N_18547);
nand U29432 (N_29432,N_23102,N_23549);
and U29433 (N_29433,N_19560,N_20372);
or U29434 (N_29434,N_19493,N_20579);
nor U29435 (N_29435,N_18328,N_23254);
nand U29436 (N_29436,N_22749,N_20858);
nor U29437 (N_29437,N_22136,N_19176);
and U29438 (N_29438,N_22418,N_23505);
xor U29439 (N_29439,N_21178,N_21490);
or U29440 (N_29440,N_20273,N_22948);
nor U29441 (N_29441,N_23689,N_22726);
nor U29442 (N_29442,N_20959,N_22564);
nand U29443 (N_29443,N_20116,N_20631);
nor U29444 (N_29444,N_19983,N_22778);
nand U29445 (N_29445,N_18984,N_23608);
xnor U29446 (N_29446,N_22881,N_20235);
xor U29447 (N_29447,N_20377,N_22735);
or U29448 (N_29448,N_22439,N_21450);
nor U29449 (N_29449,N_21396,N_18622);
nor U29450 (N_29450,N_18137,N_23373);
xnor U29451 (N_29451,N_23029,N_21334);
nand U29452 (N_29452,N_23328,N_18344);
and U29453 (N_29453,N_20130,N_22814);
or U29454 (N_29454,N_21666,N_18015);
xnor U29455 (N_29455,N_23950,N_19875);
xor U29456 (N_29456,N_20451,N_23576);
and U29457 (N_29457,N_18275,N_21300);
and U29458 (N_29458,N_20821,N_22319);
or U29459 (N_29459,N_18480,N_21577);
nor U29460 (N_29460,N_21266,N_19090);
nor U29461 (N_29461,N_18567,N_18135);
nor U29462 (N_29462,N_20695,N_20477);
nor U29463 (N_29463,N_23954,N_18683);
xnor U29464 (N_29464,N_20440,N_19343);
or U29465 (N_29465,N_23370,N_20322);
xnor U29466 (N_29466,N_22897,N_18617);
nor U29467 (N_29467,N_20064,N_23350);
xor U29468 (N_29468,N_22226,N_18965);
nor U29469 (N_29469,N_23279,N_20176);
nand U29470 (N_29470,N_18995,N_22630);
or U29471 (N_29471,N_21446,N_20958);
nor U29472 (N_29472,N_23562,N_18028);
nand U29473 (N_29473,N_19719,N_23979);
and U29474 (N_29474,N_19532,N_20886);
and U29475 (N_29475,N_20255,N_22388);
and U29476 (N_29476,N_21617,N_23227);
nand U29477 (N_29477,N_23161,N_20405);
or U29478 (N_29478,N_21927,N_21111);
nor U29479 (N_29479,N_19916,N_23949);
nand U29480 (N_29480,N_23816,N_20913);
nor U29481 (N_29481,N_19224,N_22027);
nor U29482 (N_29482,N_23831,N_19805);
xnor U29483 (N_29483,N_19255,N_23091);
nor U29484 (N_29484,N_18832,N_19245);
nor U29485 (N_29485,N_21732,N_23688);
nor U29486 (N_29486,N_19041,N_22469);
xnor U29487 (N_29487,N_19693,N_21886);
nor U29488 (N_29488,N_21698,N_22168);
nor U29489 (N_29489,N_22366,N_18225);
and U29490 (N_29490,N_20860,N_21102);
xnor U29491 (N_29491,N_23955,N_18476);
or U29492 (N_29492,N_20389,N_22528);
xnor U29493 (N_29493,N_23153,N_19735);
and U29494 (N_29494,N_22292,N_18673);
and U29495 (N_29495,N_18166,N_23310);
and U29496 (N_29496,N_19908,N_23872);
nand U29497 (N_29497,N_21300,N_20587);
and U29498 (N_29498,N_19781,N_18274);
nand U29499 (N_29499,N_21825,N_22615);
and U29500 (N_29500,N_19590,N_20681);
nand U29501 (N_29501,N_20455,N_19530);
or U29502 (N_29502,N_19127,N_23945);
or U29503 (N_29503,N_22032,N_23770);
and U29504 (N_29504,N_21713,N_19384);
xnor U29505 (N_29505,N_22503,N_21702);
xor U29506 (N_29506,N_22940,N_18001);
or U29507 (N_29507,N_20642,N_23223);
or U29508 (N_29508,N_19432,N_19933);
nand U29509 (N_29509,N_23959,N_18669);
nor U29510 (N_29510,N_20116,N_20212);
or U29511 (N_29511,N_22395,N_23522);
nand U29512 (N_29512,N_20857,N_23835);
or U29513 (N_29513,N_19477,N_21179);
or U29514 (N_29514,N_19604,N_21674);
or U29515 (N_29515,N_22210,N_23620);
or U29516 (N_29516,N_19971,N_21225);
nand U29517 (N_29517,N_20262,N_23438);
nor U29518 (N_29518,N_19927,N_21211);
and U29519 (N_29519,N_20365,N_22863);
and U29520 (N_29520,N_18868,N_23084);
and U29521 (N_29521,N_21829,N_23152);
or U29522 (N_29522,N_19114,N_22757);
nand U29523 (N_29523,N_19759,N_18236);
nor U29524 (N_29524,N_22479,N_21767);
or U29525 (N_29525,N_18785,N_20878);
xor U29526 (N_29526,N_19349,N_20583);
xor U29527 (N_29527,N_18872,N_18186);
or U29528 (N_29528,N_18087,N_22728);
xnor U29529 (N_29529,N_18194,N_22204);
nor U29530 (N_29530,N_21158,N_21117);
nor U29531 (N_29531,N_18793,N_23993);
or U29532 (N_29532,N_18531,N_18366);
and U29533 (N_29533,N_19080,N_22727);
or U29534 (N_29534,N_23100,N_20062);
xnor U29535 (N_29535,N_21248,N_21272);
nand U29536 (N_29536,N_21825,N_20875);
xnor U29537 (N_29537,N_19352,N_19219);
and U29538 (N_29538,N_22280,N_19598);
xnor U29539 (N_29539,N_23910,N_22685);
nor U29540 (N_29540,N_21805,N_22049);
xnor U29541 (N_29541,N_18882,N_21651);
nor U29542 (N_29542,N_22028,N_18125);
nand U29543 (N_29543,N_18835,N_20923);
and U29544 (N_29544,N_19662,N_22943);
and U29545 (N_29545,N_22934,N_18179);
xnor U29546 (N_29546,N_21004,N_20278);
or U29547 (N_29547,N_22115,N_21035);
nand U29548 (N_29548,N_23950,N_21829);
nor U29549 (N_29549,N_18901,N_22337);
and U29550 (N_29550,N_19849,N_21063);
nor U29551 (N_29551,N_20988,N_23050);
or U29552 (N_29552,N_22300,N_19174);
nand U29553 (N_29553,N_18784,N_18380);
nor U29554 (N_29554,N_20187,N_19355);
and U29555 (N_29555,N_20070,N_22089);
nor U29556 (N_29556,N_20431,N_20444);
nor U29557 (N_29557,N_18438,N_18047);
and U29558 (N_29558,N_18761,N_21945);
and U29559 (N_29559,N_22514,N_20388);
nor U29560 (N_29560,N_23157,N_21282);
nand U29561 (N_29561,N_21895,N_22697);
xor U29562 (N_29562,N_23186,N_19632);
and U29563 (N_29563,N_18636,N_19591);
nand U29564 (N_29564,N_22060,N_20037);
nand U29565 (N_29565,N_20348,N_21940);
nand U29566 (N_29566,N_22861,N_19312);
or U29567 (N_29567,N_22236,N_19418);
and U29568 (N_29568,N_18034,N_19452);
nor U29569 (N_29569,N_21246,N_21195);
and U29570 (N_29570,N_18600,N_18791);
xnor U29571 (N_29571,N_21287,N_22724);
or U29572 (N_29572,N_18456,N_19598);
nand U29573 (N_29573,N_22169,N_21290);
and U29574 (N_29574,N_20495,N_21437);
and U29575 (N_29575,N_23368,N_19573);
xor U29576 (N_29576,N_22240,N_21054);
nor U29577 (N_29577,N_19003,N_21118);
xor U29578 (N_29578,N_21391,N_20432);
or U29579 (N_29579,N_19660,N_21338);
xor U29580 (N_29580,N_20648,N_21476);
and U29581 (N_29581,N_18879,N_21370);
and U29582 (N_29582,N_18430,N_18811);
or U29583 (N_29583,N_19165,N_18774);
xor U29584 (N_29584,N_22623,N_23907);
xnor U29585 (N_29585,N_22373,N_18341);
nand U29586 (N_29586,N_20917,N_22690);
nor U29587 (N_29587,N_23932,N_22645);
nor U29588 (N_29588,N_22008,N_22414);
and U29589 (N_29589,N_18738,N_23037);
or U29590 (N_29590,N_18715,N_18830);
xor U29591 (N_29591,N_21487,N_23833);
nand U29592 (N_29592,N_18455,N_22265);
nand U29593 (N_29593,N_18362,N_21130);
and U29594 (N_29594,N_20949,N_19205);
nor U29595 (N_29595,N_23201,N_22914);
and U29596 (N_29596,N_21398,N_23204);
nand U29597 (N_29597,N_19234,N_23764);
and U29598 (N_29598,N_20100,N_23005);
or U29599 (N_29599,N_20519,N_22167);
and U29600 (N_29600,N_22402,N_20145);
and U29601 (N_29601,N_19368,N_19401);
or U29602 (N_29602,N_19907,N_21986);
nand U29603 (N_29603,N_23562,N_23510);
or U29604 (N_29604,N_21368,N_21650);
nor U29605 (N_29605,N_19265,N_20814);
or U29606 (N_29606,N_18512,N_21049);
nor U29607 (N_29607,N_20334,N_23205);
nor U29608 (N_29608,N_20100,N_21558);
xnor U29609 (N_29609,N_22066,N_23854);
nor U29610 (N_29610,N_23407,N_19396);
nand U29611 (N_29611,N_23569,N_21584);
nand U29612 (N_29612,N_22514,N_20473);
and U29613 (N_29613,N_20791,N_20587);
xor U29614 (N_29614,N_19580,N_18196);
nor U29615 (N_29615,N_21763,N_20982);
xor U29616 (N_29616,N_20328,N_18894);
and U29617 (N_29617,N_20629,N_22664);
nand U29618 (N_29618,N_18460,N_21468);
nor U29619 (N_29619,N_18978,N_23092);
xor U29620 (N_29620,N_22058,N_22893);
xnor U29621 (N_29621,N_22652,N_19784);
or U29622 (N_29622,N_20564,N_18916);
xor U29623 (N_29623,N_21364,N_20188);
nor U29624 (N_29624,N_21133,N_18994);
nand U29625 (N_29625,N_20341,N_21739);
and U29626 (N_29626,N_21189,N_18872);
nor U29627 (N_29627,N_18651,N_22466);
nor U29628 (N_29628,N_20884,N_20410);
nor U29629 (N_29629,N_21426,N_21473);
nand U29630 (N_29630,N_22186,N_21765);
nand U29631 (N_29631,N_19286,N_21507);
nor U29632 (N_29632,N_21406,N_23980);
xnor U29633 (N_29633,N_20400,N_18732);
or U29634 (N_29634,N_21937,N_21845);
xor U29635 (N_29635,N_22245,N_20189);
xor U29636 (N_29636,N_20814,N_20200);
xor U29637 (N_29637,N_21296,N_19937);
xnor U29638 (N_29638,N_19428,N_20896);
nor U29639 (N_29639,N_21369,N_22317);
xor U29640 (N_29640,N_19293,N_22112);
xor U29641 (N_29641,N_20466,N_21508);
nor U29642 (N_29642,N_18217,N_21090);
nand U29643 (N_29643,N_21546,N_22791);
xor U29644 (N_29644,N_22326,N_18778);
or U29645 (N_29645,N_18154,N_22737);
nand U29646 (N_29646,N_20536,N_21692);
xnor U29647 (N_29647,N_19172,N_22735);
and U29648 (N_29648,N_23429,N_19121);
or U29649 (N_29649,N_18538,N_22296);
or U29650 (N_29650,N_20331,N_22315);
and U29651 (N_29651,N_21655,N_22569);
or U29652 (N_29652,N_21416,N_23946);
xnor U29653 (N_29653,N_19040,N_21535);
nand U29654 (N_29654,N_22302,N_21268);
or U29655 (N_29655,N_23986,N_23067);
nor U29656 (N_29656,N_21578,N_19916);
and U29657 (N_29657,N_19647,N_19558);
xnor U29658 (N_29658,N_21745,N_18615);
or U29659 (N_29659,N_21198,N_23607);
xor U29660 (N_29660,N_21030,N_21440);
xnor U29661 (N_29661,N_18465,N_22578);
nor U29662 (N_29662,N_22290,N_22100);
nand U29663 (N_29663,N_19405,N_19248);
nor U29664 (N_29664,N_19907,N_19040);
nor U29665 (N_29665,N_20195,N_23805);
nand U29666 (N_29666,N_22910,N_18407);
xor U29667 (N_29667,N_23081,N_21730);
xor U29668 (N_29668,N_22188,N_18754);
nor U29669 (N_29669,N_21056,N_18566);
and U29670 (N_29670,N_23483,N_23373);
and U29671 (N_29671,N_23103,N_23261);
xor U29672 (N_29672,N_19871,N_22104);
and U29673 (N_29673,N_21521,N_21427);
and U29674 (N_29674,N_20599,N_18118);
xor U29675 (N_29675,N_21174,N_21729);
and U29676 (N_29676,N_20555,N_18159);
xnor U29677 (N_29677,N_23622,N_22494);
xnor U29678 (N_29678,N_19240,N_21128);
xnor U29679 (N_29679,N_19029,N_22719);
or U29680 (N_29680,N_18937,N_19233);
xnor U29681 (N_29681,N_19539,N_18362);
and U29682 (N_29682,N_20158,N_20755);
or U29683 (N_29683,N_19970,N_21967);
and U29684 (N_29684,N_22379,N_22219);
and U29685 (N_29685,N_22209,N_21978);
or U29686 (N_29686,N_23414,N_23609);
xor U29687 (N_29687,N_19875,N_19090);
or U29688 (N_29688,N_21622,N_23888);
nor U29689 (N_29689,N_22717,N_19975);
and U29690 (N_29690,N_20742,N_22183);
nor U29691 (N_29691,N_21197,N_22461);
and U29692 (N_29692,N_20754,N_21803);
and U29693 (N_29693,N_22215,N_20725);
or U29694 (N_29694,N_20906,N_22557);
nor U29695 (N_29695,N_19172,N_19415);
nor U29696 (N_29696,N_23618,N_23296);
nand U29697 (N_29697,N_19254,N_23988);
or U29698 (N_29698,N_20063,N_20212);
nor U29699 (N_29699,N_23827,N_18031);
nor U29700 (N_29700,N_22006,N_22851);
nand U29701 (N_29701,N_20822,N_22632);
nand U29702 (N_29702,N_18221,N_18624);
xnor U29703 (N_29703,N_20029,N_20084);
or U29704 (N_29704,N_21809,N_18639);
and U29705 (N_29705,N_22532,N_18113);
nor U29706 (N_29706,N_23330,N_23078);
nand U29707 (N_29707,N_22149,N_22540);
nand U29708 (N_29708,N_21860,N_22595);
xnor U29709 (N_29709,N_22840,N_21475);
or U29710 (N_29710,N_20111,N_18620);
and U29711 (N_29711,N_21474,N_21837);
and U29712 (N_29712,N_18281,N_20178);
xnor U29713 (N_29713,N_23204,N_21910);
or U29714 (N_29714,N_21562,N_22509);
or U29715 (N_29715,N_19251,N_22778);
and U29716 (N_29716,N_22954,N_18672);
nor U29717 (N_29717,N_20224,N_21551);
nor U29718 (N_29718,N_23654,N_19299);
xnor U29719 (N_29719,N_22945,N_18348);
nand U29720 (N_29720,N_22619,N_18111);
nor U29721 (N_29721,N_23509,N_23245);
or U29722 (N_29722,N_23591,N_18767);
nor U29723 (N_29723,N_22873,N_19110);
and U29724 (N_29724,N_18228,N_21423);
or U29725 (N_29725,N_20724,N_21193);
or U29726 (N_29726,N_23695,N_23656);
xor U29727 (N_29727,N_23718,N_22318);
and U29728 (N_29728,N_21958,N_19398);
xnor U29729 (N_29729,N_22788,N_19681);
nand U29730 (N_29730,N_21688,N_20682);
xor U29731 (N_29731,N_19342,N_18127);
nor U29732 (N_29732,N_18550,N_22026);
or U29733 (N_29733,N_20119,N_23248);
xor U29734 (N_29734,N_20741,N_20646);
nand U29735 (N_29735,N_22107,N_23170);
and U29736 (N_29736,N_18111,N_18956);
nand U29737 (N_29737,N_23617,N_18719);
or U29738 (N_29738,N_21260,N_19739);
and U29739 (N_29739,N_18332,N_23612);
xor U29740 (N_29740,N_18155,N_21278);
nor U29741 (N_29741,N_23285,N_21226);
or U29742 (N_29742,N_23776,N_21304);
xor U29743 (N_29743,N_18281,N_22835);
or U29744 (N_29744,N_18483,N_22971);
nor U29745 (N_29745,N_22587,N_18480);
or U29746 (N_29746,N_20255,N_18364);
or U29747 (N_29747,N_20748,N_20645);
xnor U29748 (N_29748,N_23707,N_22719);
and U29749 (N_29749,N_18522,N_22145);
xnor U29750 (N_29750,N_20076,N_19328);
or U29751 (N_29751,N_19142,N_18499);
and U29752 (N_29752,N_20030,N_21173);
or U29753 (N_29753,N_21059,N_20876);
xor U29754 (N_29754,N_21050,N_19080);
xor U29755 (N_29755,N_20289,N_23738);
xnor U29756 (N_29756,N_22779,N_19368);
nor U29757 (N_29757,N_20979,N_23692);
or U29758 (N_29758,N_18760,N_22641);
or U29759 (N_29759,N_22017,N_19531);
nand U29760 (N_29760,N_20310,N_21129);
nand U29761 (N_29761,N_18397,N_19310);
xor U29762 (N_29762,N_21918,N_22324);
or U29763 (N_29763,N_23400,N_22317);
nor U29764 (N_29764,N_21475,N_21096);
nand U29765 (N_29765,N_18859,N_22381);
and U29766 (N_29766,N_22464,N_18652);
nor U29767 (N_29767,N_20523,N_21826);
and U29768 (N_29768,N_19238,N_18572);
and U29769 (N_29769,N_18600,N_19403);
nand U29770 (N_29770,N_18790,N_18146);
nand U29771 (N_29771,N_20851,N_20301);
nand U29772 (N_29772,N_18460,N_22747);
and U29773 (N_29773,N_21708,N_23998);
nand U29774 (N_29774,N_20706,N_20817);
or U29775 (N_29775,N_21895,N_23147);
and U29776 (N_29776,N_23813,N_18925);
nand U29777 (N_29777,N_23782,N_21699);
or U29778 (N_29778,N_18717,N_19924);
nand U29779 (N_29779,N_21192,N_19514);
nor U29780 (N_29780,N_21522,N_23300);
nand U29781 (N_29781,N_22661,N_22715);
nor U29782 (N_29782,N_18128,N_23295);
nand U29783 (N_29783,N_21442,N_21772);
and U29784 (N_29784,N_19981,N_22615);
nand U29785 (N_29785,N_23799,N_18773);
xor U29786 (N_29786,N_22484,N_18723);
and U29787 (N_29787,N_21659,N_18784);
nor U29788 (N_29788,N_22239,N_20598);
nand U29789 (N_29789,N_23182,N_18233);
or U29790 (N_29790,N_18864,N_22944);
nand U29791 (N_29791,N_23764,N_21888);
nand U29792 (N_29792,N_21260,N_18360);
or U29793 (N_29793,N_19822,N_19656);
nor U29794 (N_29794,N_19565,N_22139);
nand U29795 (N_29795,N_23225,N_18290);
nor U29796 (N_29796,N_23280,N_21727);
nor U29797 (N_29797,N_23597,N_18713);
nor U29798 (N_29798,N_20581,N_19454);
nand U29799 (N_29799,N_19603,N_23634);
nor U29800 (N_29800,N_20295,N_22683);
xnor U29801 (N_29801,N_22258,N_22923);
xnor U29802 (N_29802,N_20279,N_18199);
xor U29803 (N_29803,N_20468,N_22110);
nand U29804 (N_29804,N_22119,N_18302);
and U29805 (N_29805,N_18643,N_21255);
or U29806 (N_29806,N_23577,N_21790);
nand U29807 (N_29807,N_20157,N_20855);
or U29808 (N_29808,N_22181,N_22946);
and U29809 (N_29809,N_21111,N_18381);
xor U29810 (N_29810,N_23875,N_23909);
and U29811 (N_29811,N_21967,N_23464);
or U29812 (N_29812,N_19916,N_19541);
nand U29813 (N_29813,N_19223,N_22487);
nor U29814 (N_29814,N_23585,N_23297);
and U29815 (N_29815,N_20552,N_19033);
xor U29816 (N_29816,N_19419,N_19502);
or U29817 (N_29817,N_19872,N_21437);
xnor U29818 (N_29818,N_18836,N_19469);
nand U29819 (N_29819,N_20938,N_23391);
nand U29820 (N_29820,N_19106,N_21220);
or U29821 (N_29821,N_23743,N_22356);
or U29822 (N_29822,N_18606,N_18888);
nand U29823 (N_29823,N_21509,N_21026);
xnor U29824 (N_29824,N_21549,N_20605);
and U29825 (N_29825,N_23933,N_21615);
nand U29826 (N_29826,N_20807,N_21080);
xnor U29827 (N_29827,N_22670,N_19305);
nor U29828 (N_29828,N_20454,N_18870);
xnor U29829 (N_29829,N_21649,N_23607);
nand U29830 (N_29830,N_18040,N_21631);
and U29831 (N_29831,N_22059,N_20743);
nand U29832 (N_29832,N_18241,N_18878);
nor U29833 (N_29833,N_23083,N_19013);
or U29834 (N_29834,N_23076,N_22239);
xnor U29835 (N_29835,N_23554,N_23191);
nor U29836 (N_29836,N_20439,N_22646);
xor U29837 (N_29837,N_18669,N_20414);
nor U29838 (N_29838,N_20846,N_18420);
and U29839 (N_29839,N_23685,N_18319);
nand U29840 (N_29840,N_23195,N_21426);
nor U29841 (N_29841,N_18822,N_22247);
nor U29842 (N_29842,N_23168,N_22469);
nor U29843 (N_29843,N_18938,N_20362);
or U29844 (N_29844,N_20298,N_20636);
nor U29845 (N_29845,N_21121,N_19092);
nand U29846 (N_29846,N_19279,N_20551);
or U29847 (N_29847,N_18426,N_20916);
nand U29848 (N_29848,N_20055,N_20606);
or U29849 (N_29849,N_19507,N_22879);
nand U29850 (N_29850,N_22503,N_22756);
or U29851 (N_29851,N_22289,N_19215);
or U29852 (N_29852,N_22276,N_18833);
or U29853 (N_29853,N_19110,N_19291);
nor U29854 (N_29854,N_21787,N_21244);
nor U29855 (N_29855,N_21873,N_19525);
nor U29856 (N_29856,N_20457,N_22828);
nand U29857 (N_29857,N_23660,N_19534);
or U29858 (N_29858,N_18797,N_21617);
nor U29859 (N_29859,N_22696,N_18415);
or U29860 (N_29860,N_18396,N_22725);
nor U29861 (N_29861,N_18318,N_19924);
nor U29862 (N_29862,N_18182,N_20204);
nand U29863 (N_29863,N_19183,N_20776);
nor U29864 (N_29864,N_21939,N_23919);
or U29865 (N_29865,N_22401,N_22576);
nor U29866 (N_29866,N_21781,N_19065);
nor U29867 (N_29867,N_23412,N_22920);
or U29868 (N_29868,N_19078,N_23266);
or U29869 (N_29869,N_23419,N_20846);
xor U29870 (N_29870,N_22716,N_22701);
nand U29871 (N_29871,N_22687,N_19383);
or U29872 (N_29872,N_21475,N_21572);
and U29873 (N_29873,N_20901,N_18604);
and U29874 (N_29874,N_19100,N_23711);
xor U29875 (N_29875,N_23676,N_21193);
nor U29876 (N_29876,N_19694,N_18721);
and U29877 (N_29877,N_23540,N_23928);
xnor U29878 (N_29878,N_18352,N_23402);
or U29879 (N_29879,N_18665,N_20226);
nand U29880 (N_29880,N_18875,N_22053);
nand U29881 (N_29881,N_18395,N_23011);
nor U29882 (N_29882,N_22228,N_19332);
or U29883 (N_29883,N_18021,N_18613);
and U29884 (N_29884,N_22237,N_19263);
nor U29885 (N_29885,N_19939,N_23874);
or U29886 (N_29886,N_21832,N_21721);
or U29887 (N_29887,N_18691,N_23460);
nor U29888 (N_29888,N_22954,N_22798);
or U29889 (N_29889,N_18583,N_22691);
or U29890 (N_29890,N_21878,N_21406);
nand U29891 (N_29891,N_19109,N_19521);
and U29892 (N_29892,N_18258,N_23148);
and U29893 (N_29893,N_19900,N_19367);
nand U29894 (N_29894,N_21234,N_21986);
nand U29895 (N_29895,N_19510,N_21496);
and U29896 (N_29896,N_20418,N_19663);
or U29897 (N_29897,N_23712,N_22226);
or U29898 (N_29898,N_23264,N_22285);
nor U29899 (N_29899,N_20190,N_19073);
or U29900 (N_29900,N_22160,N_22988);
or U29901 (N_29901,N_19566,N_22359);
nor U29902 (N_29902,N_21715,N_21821);
and U29903 (N_29903,N_23847,N_19748);
xnor U29904 (N_29904,N_21138,N_19125);
nand U29905 (N_29905,N_20309,N_20030);
nor U29906 (N_29906,N_18129,N_18352);
or U29907 (N_29907,N_22320,N_22559);
or U29908 (N_29908,N_18982,N_23691);
nand U29909 (N_29909,N_23684,N_23852);
xor U29910 (N_29910,N_20732,N_21555);
or U29911 (N_29911,N_20826,N_22175);
nand U29912 (N_29912,N_22078,N_22261);
and U29913 (N_29913,N_19867,N_22578);
xor U29914 (N_29914,N_18070,N_23280);
nor U29915 (N_29915,N_22477,N_19417);
and U29916 (N_29916,N_20081,N_23971);
nand U29917 (N_29917,N_18759,N_21916);
or U29918 (N_29918,N_20962,N_23283);
xnor U29919 (N_29919,N_22183,N_23820);
nand U29920 (N_29920,N_18069,N_21321);
xnor U29921 (N_29921,N_23771,N_20307);
and U29922 (N_29922,N_18181,N_23983);
or U29923 (N_29923,N_20355,N_19099);
and U29924 (N_29924,N_20809,N_20929);
or U29925 (N_29925,N_18664,N_20865);
xor U29926 (N_29926,N_20576,N_19824);
nor U29927 (N_29927,N_21650,N_21287);
and U29928 (N_29928,N_23148,N_20914);
nand U29929 (N_29929,N_18782,N_21797);
and U29930 (N_29930,N_22891,N_20240);
and U29931 (N_29931,N_19146,N_22163);
or U29932 (N_29932,N_19485,N_21169);
or U29933 (N_29933,N_23170,N_18970);
or U29934 (N_29934,N_22347,N_18698);
or U29935 (N_29935,N_18444,N_19495);
nand U29936 (N_29936,N_22038,N_20994);
or U29937 (N_29937,N_20734,N_20590);
xor U29938 (N_29938,N_23463,N_18377);
nand U29939 (N_29939,N_18611,N_19168);
or U29940 (N_29940,N_20473,N_20817);
nor U29941 (N_29941,N_21349,N_18459);
or U29942 (N_29942,N_20178,N_18633);
xor U29943 (N_29943,N_22794,N_21205);
nor U29944 (N_29944,N_19165,N_18107);
nand U29945 (N_29945,N_21816,N_20345);
nand U29946 (N_29946,N_18983,N_21330);
xor U29947 (N_29947,N_22050,N_19889);
xor U29948 (N_29948,N_19070,N_18600);
nand U29949 (N_29949,N_22999,N_19540);
nor U29950 (N_29950,N_23947,N_18846);
xnor U29951 (N_29951,N_18946,N_23348);
nor U29952 (N_29952,N_19109,N_22629);
xor U29953 (N_29953,N_22920,N_20773);
nor U29954 (N_29954,N_22523,N_20543);
xor U29955 (N_29955,N_22738,N_23070);
and U29956 (N_29956,N_23744,N_22785);
and U29957 (N_29957,N_19101,N_19331);
and U29958 (N_29958,N_21348,N_22762);
xnor U29959 (N_29959,N_21390,N_23238);
nand U29960 (N_29960,N_23563,N_20419);
nand U29961 (N_29961,N_18562,N_18159);
and U29962 (N_29962,N_22013,N_21364);
xnor U29963 (N_29963,N_21234,N_18821);
nand U29964 (N_29964,N_23251,N_19445);
nand U29965 (N_29965,N_20116,N_21197);
nor U29966 (N_29966,N_19163,N_18967);
nand U29967 (N_29967,N_22775,N_21130);
xnor U29968 (N_29968,N_22505,N_20403);
xnor U29969 (N_29969,N_23496,N_18000);
and U29970 (N_29970,N_21220,N_23382);
or U29971 (N_29971,N_19919,N_18347);
and U29972 (N_29972,N_21885,N_21198);
or U29973 (N_29973,N_22111,N_18511);
and U29974 (N_29974,N_23483,N_20212);
and U29975 (N_29975,N_18196,N_18262);
nor U29976 (N_29976,N_21182,N_18098);
nand U29977 (N_29977,N_20390,N_22550);
nand U29978 (N_29978,N_22152,N_21194);
and U29979 (N_29979,N_18676,N_18070);
nor U29980 (N_29980,N_20918,N_22212);
xor U29981 (N_29981,N_20464,N_23082);
xor U29982 (N_29982,N_18542,N_18462);
xnor U29983 (N_29983,N_18541,N_18933);
xnor U29984 (N_29984,N_22116,N_20174);
xor U29985 (N_29985,N_23290,N_18334);
nand U29986 (N_29986,N_20397,N_23765);
xor U29987 (N_29987,N_20182,N_19651);
nand U29988 (N_29988,N_18586,N_21774);
xor U29989 (N_29989,N_23629,N_22850);
or U29990 (N_29990,N_23939,N_19682);
xnor U29991 (N_29991,N_23105,N_22006);
nor U29992 (N_29992,N_18953,N_22864);
xor U29993 (N_29993,N_19367,N_22923);
nor U29994 (N_29994,N_22664,N_18289);
nor U29995 (N_29995,N_23385,N_23650);
or U29996 (N_29996,N_22563,N_19817);
nand U29997 (N_29997,N_18801,N_21447);
or U29998 (N_29998,N_21710,N_21925);
or U29999 (N_29999,N_22076,N_18717);
and UO_0 (O_0,N_25281,N_29961);
and UO_1 (O_1,N_28511,N_24657);
nand UO_2 (O_2,N_27466,N_26607);
nor UO_3 (O_3,N_24938,N_26047);
nand UO_4 (O_4,N_27085,N_27922);
or UO_5 (O_5,N_25630,N_29099);
nand UO_6 (O_6,N_27733,N_25979);
and UO_7 (O_7,N_29692,N_25320);
or UO_8 (O_8,N_26615,N_29309);
nand UO_9 (O_9,N_27462,N_26221);
or UO_10 (O_10,N_29997,N_28243);
nor UO_11 (O_11,N_24733,N_29451);
and UO_12 (O_12,N_25670,N_25330);
and UO_13 (O_13,N_24168,N_25438);
nand UO_14 (O_14,N_27881,N_27442);
or UO_15 (O_15,N_25987,N_28573);
nand UO_16 (O_16,N_24174,N_27164);
nor UO_17 (O_17,N_26336,N_27293);
and UO_18 (O_18,N_27183,N_26954);
or UO_19 (O_19,N_24526,N_28223);
nor UO_20 (O_20,N_29085,N_25268);
nand UO_21 (O_21,N_27334,N_25805);
nor UO_22 (O_22,N_28280,N_28784);
nor UO_23 (O_23,N_25389,N_28208);
nor UO_24 (O_24,N_26125,N_27326);
xnor UO_25 (O_25,N_26229,N_29206);
nor UO_26 (O_26,N_29069,N_28173);
and UO_27 (O_27,N_26650,N_28268);
and UO_28 (O_28,N_26814,N_28982);
and UO_29 (O_29,N_26981,N_27540);
nor UO_30 (O_30,N_28883,N_26794);
nor UO_31 (O_31,N_25218,N_26302);
xor UO_32 (O_32,N_25624,N_26265);
and UO_33 (O_33,N_27910,N_28427);
and UO_34 (O_34,N_24661,N_27701);
nor UO_35 (O_35,N_24267,N_27628);
or UO_36 (O_36,N_25398,N_27286);
nand UO_37 (O_37,N_25322,N_29237);
nand UO_38 (O_38,N_28150,N_24787);
nor UO_39 (O_39,N_26807,N_25215);
and UO_40 (O_40,N_29732,N_27460);
and UO_41 (O_41,N_24291,N_26094);
and UO_42 (O_42,N_26044,N_29635);
nor UO_43 (O_43,N_25549,N_25460);
nor UO_44 (O_44,N_27974,N_27985);
nor UO_45 (O_45,N_26550,N_25459);
and UO_46 (O_46,N_29136,N_28136);
or UO_47 (O_47,N_28458,N_25074);
xor UO_48 (O_48,N_29531,N_24510);
nor UO_49 (O_49,N_29789,N_27621);
nor UO_50 (O_50,N_25850,N_25232);
nand UO_51 (O_51,N_24914,N_28611);
nand UO_52 (O_52,N_27674,N_25939);
and UO_53 (O_53,N_27122,N_29037);
xor UO_54 (O_54,N_27088,N_29221);
and UO_55 (O_55,N_26142,N_25350);
and UO_56 (O_56,N_29190,N_27015);
nand UO_57 (O_57,N_28507,N_25575);
and UO_58 (O_58,N_29046,N_28297);
nand UO_59 (O_59,N_25697,N_25636);
and UO_60 (O_60,N_28559,N_26874);
xor UO_61 (O_61,N_28501,N_25253);
and UO_62 (O_62,N_26519,N_25981);
nor UO_63 (O_63,N_29222,N_28586);
xnor UO_64 (O_64,N_28951,N_26668);
nor UO_65 (O_65,N_29124,N_24975);
nor UO_66 (O_66,N_26710,N_27981);
or UO_67 (O_67,N_24829,N_24410);
xnor UO_68 (O_68,N_27377,N_25401);
or UO_69 (O_69,N_26080,N_29935);
xnor UO_70 (O_70,N_29538,N_24557);
xor UO_71 (O_71,N_25024,N_24537);
and UO_72 (O_72,N_28454,N_24558);
and UO_73 (O_73,N_24808,N_29627);
nand UO_74 (O_74,N_24889,N_24732);
xor UO_75 (O_75,N_26452,N_27480);
and UO_76 (O_76,N_29024,N_25968);
nand UO_77 (O_77,N_24461,N_24005);
or UO_78 (O_78,N_27408,N_29158);
nor UO_79 (O_79,N_29054,N_25442);
nor UO_80 (O_80,N_26701,N_26252);
nand UO_81 (O_81,N_29161,N_26511);
nor UO_82 (O_82,N_27801,N_27118);
or UO_83 (O_83,N_27786,N_27129);
nand UO_84 (O_84,N_28017,N_27723);
and UO_85 (O_85,N_27053,N_29980);
nor UO_86 (O_86,N_26068,N_25952);
or UO_87 (O_87,N_26597,N_28546);
nand UO_88 (O_88,N_26778,N_29077);
xnor UO_89 (O_89,N_25525,N_26030);
or UO_90 (O_90,N_27211,N_29100);
and UO_91 (O_91,N_28051,N_24752);
xor UO_92 (O_92,N_27142,N_26632);
nor UO_93 (O_93,N_27648,N_29553);
nor UO_94 (O_94,N_24129,N_28814);
or UO_95 (O_95,N_25715,N_24762);
xor UO_96 (O_96,N_26061,N_28588);
or UO_97 (O_97,N_27896,N_27359);
xnor UO_98 (O_98,N_28340,N_28610);
and UO_99 (O_99,N_27045,N_25731);
and UO_100 (O_100,N_26903,N_27979);
nor UO_101 (O_101,N_25794,N_27320);
and UO_102 (O_102,N_26174,N_26277);
nor UO_103 (O_103,N_28683,N_24313);
nand UO_104 (O_104,N_28253,N_29003);
or UO_105 (O_105,N_26666,N_29757);
or UO_106 (O_106,N_24239,N_24446);
xnor UO_107 (O_107,N_24241,N_24498);
and UO_108 (O_108,N_27920,N_26189);
or UO_109 (O_109,N_25693,N_28531);
xor UO_110 (O_110,N_29341,N_24877);
nor UO_111 (O_111,N_26023,N_27439);
and UO_112 (O_112,N_24896,N_25373);
xor UO_113 (O_113,N_29671,N_26885);
and UO_114 (O_114,N_29532,N_29141);
and UO_115 (O_115,N_25434,N_28566);
or UO_116 (O_116,N_24660,N_26284);
nand UO_117 (O_117,N_24918,N_27303);
nand UO_118 (O_118,N_29042,N_28276);
xnor UO_119 (O_119,N_25814,N_27630);
or UO_120 (O_120,N_26799,N_27178);
nor UO_121 (O_121,N_26951,N_27806);
nor UO_122 (O_122,N_26259,N_28486);
nor UO_123 (O_123,N_27274,N_27880);
nor UO_124 (O_124,N_24268,N_24160);
or UO_125 (O_125,N_28889,N_29408);
nor UO_126 (O_126,N_29007,N_28134);
or UO_127 (O_127,N_27642,N_25907);
and UO_128 (O_128,N_29375,N_25280);
xnor UO_129 (O_129,N_28129,N_28707);
nor UO_130 (O_130,N_29474,N_28795);
or UO_131 (O_131,N_25708,N_28016);
and UO_132 (O_132,N_25722,N_27421);
nand UO_133 (O_133,N_26627,N_28605);
nor UO_134 (O_134,N_28740,N_28483);
nor UO_135 (O_135,N_28895,N_29092);
nor UO_136 (O_136,N_28663,N_27073);
xnor UO_137 (O_137,N_26845,N_29536);
nor UO_138 (O_138,N_27483,N_29514);
and UO_139 (O_139,N_28023,N_24468);
nor UO_140 (O_140,N_29949,N_26427);
nor UO_141 (O_141,N_29027,N_24491);
nor UO_142 (O_142,N_24587,N_25931);
or UO_143 (O_143,N_28639,N_24915);
or UO_144 (O_144,N_28272,N_27339);
or UO_145 (O_145,N_24588,N_27782);
xor UO_146 (O_146,N_24081,N_26722);
nor UO_147 (O_147,N_28445,N_28823);
nand UO_148 (O_148,N_27301,N_29972);
nand UO_149 (O_149,N_24130,N_24951);
or UO_150 (O_150,N_26934,N_27354);
nand UO_151 (O_151,N_29038,N_29296);
xnor UO_152 (O_152,N_29860,N_24770);
and UO_153 (O_153,N_29633,N_27969);
xnor UO_154 (O_154,N_28443,N_26060);
xnor UO_155 (O_155,N_27162,N_24109);
and UO_156 (O_156,N_25552,N_26456);
nor UO_157 (O_157,N_27472,N_26609);
or UO_158 (O_158,N_24012,N_26151);
nand UO_159 (O_159,N_25516,N_27493);
nor UO_160 (O_160,N_29624,N_27874);
xor UO_161 (O_161,N_28909,N_25256);
or UO_162 (O_162,N_25088,N_26931);
xor UO_163 (O_163,N_25823,N_25245);
and UO_164 (O_164,N_26897,N_26398);
nand UO_165 (O_165,N_28396,N_27983);
nor UO_166 (O_166,N_26725,N_25784);
and UO_167 (O_167,N_24105,N_24325);
or UO_168 (O_168,N_28420,N_26949);
or UO_169 (O_169,N_27090,N_28167);
and UO_170 (O_170,N_25341,N_28222);
nand UO_171 (O_171,N_29189,N_24441);
xor UO_172 (O_172,N_25340,N_27269);
or UO_173 (O_173,N_25622,N_28689);
and UO_174 (O_174,N_27524,N_28447);
nor UO_175 (O_175,N_27279,N_26136);
nand UO_176 (O_176,N_27464,N_29788);
and UO_177 (O_177,N_26143,N_29978);
and UO_178 (O_178,N_26875,N_29062);
xor UO_179 (O_179,N_29043,N_27858);
nand UO_180 (O_180,N_24155,N_24036);
nand UO_181 (O_181,N_27202,N_28470);
nor UO_182 (O_182,N_24845,N_28660);
xor UO_183 (O_183,N_24977,N_27878);
nor UO_184 (O_184,N_25573,N_24224);
nand UO_185 (O_185,N_24063,N_24691);
xor UO_186 (O_186,N_24935,N_25277);
xnor UO_187 (O_187,N_24380,N_28065);
nor UO_188 (O_188,N_27672,N_29744);
and UO_189 (O_189,N_25743,N_24764);
or UO_190 (O_190,N_28186,N_28868);
and UO_191 (O_191,N_26117,N_28440);
nand UO_192 (O_192,N_29772,N_27867);
and UO_193 (O_193,N_24144,N_27823);
or UO_194 (O_194,N_26973,N_25514);
nor UO_195 (O_195,N_24574,N_24804);
or UO_196 (O_196,N_29599,N_28950);
xor UO_197 (O_197,N_28344,N_25977);
nand UO_198 (O_198,N_27932,N_28166);
and UO_199 (O_199,N_28721,N_24102);
xor UO_200 (O_200,N_25651,N_29241);
nor UO_201 (O_201,N_29262,N_24706);
or UO_202 (O_202,N_25596,N_26870);
xnor UO_203 (O_203,N_24548,N_26665);
or UO_204 (O_204,N_26629,N_26112);
and UO_205 (O_205,N_25701,N_25423);
nand UO_206 (O_206,N_27516,N_28783);
nor UO_207 (O_207,N_24353,N_28928);
nor UO_208 (O_208,N_24016,N_29689);
or UO_209 (O_209,N_28158,N_27347);
and UO_210 (O_210,N_25358,N_28037);
nor UO_211 (O_211,N_24058,N_29750);
nor UO_212 (O_212,N_24791,N_29397);
and UO_213 (O_213,N_25139,N_28917);
xor UO_214 (O_214,N_27297,N_25916);
and UO_215 (O_215,N_26707,N_26362);
xor UO_216 (O_216,N_28845,N_26618);
nor UO_217 (O_217,N_26860,N_28727);
xnor UO_218 (O_218,N_25451,N_24112);
nand UO_219 (O_219,N_24522,N_28782);
nor UO_220 (O_220,N_28007,N_28006);
and UO_221 (O_221,N_25095,N_24354);
or UO_222 (O_222,N_27533,N_27125);
and UO_223 (O_223,N_26434,N_25956);
nand UO_224 (O_224,N_24810,N_26408);
and UO_225 (O_225,N_29389,N_25485);
and UO_226 (O_226,N_28499,N_28698);
xor UO_227 (O_227,N_25383,N_24482);
nor UO_228 (O_228,N_27554,N_26965);
nor UO_229 (O_229,N_29798,N_26738);
xnor UO_230 (O_230,N_24653,N_25849);
nand UO_231 (O_231,N_26758,N_27222);
nor UO_232 (O_232,N_26461,N_24844);
or UO_233 (O_233,N_24251,N_24848);
or UO_234 (O_234,N_24438,N_24542);
xor UO_235 (O_235,N_27188,N_27384);
or UO_236 (O_236,N_29172,N_28637);
nand UO_237 (O_237,N_26246,N_28953);
or UO_238 (O_238,N_27050,N_28640);
nor UO_239 (O_239,N_27266,N_27098);
nor UO_240 (O_240,N_27115,N_26032);
nor UO_241 (O_241,N_26782,N_29709);
and UO_242 (O_242,N_26990,N_26438);
and UO_243 (O_243,N_24705,N_26101);
or UO_244 (O_244,N_29785,N_26800);
nor UO_245 (O_245,N_26655,N_26342);
nand UO_246 (O_246,N_25209,N_26601);
xnor UO_247 (O_247,N_25255,N_27608);
xnor UO_248 (O_248,N_27909,N_26848);
and UO_249 (O_249,N_27004,N_26058);
xnor UO_250 (O_250,N_25528,N_29706);
xnor UO_251 (O_251,N_25983,N_27190);
nor UO_252 (O_252,N_27433,N_26017);
xor UO_253 (O_253,N_27119,N_25774);
nor UO_254 (O_254,N_29891,N_26553);
nor UO_255 (O_255,N_25188,N_25479);
or UO_256 (O_256,N_28043,N_28720);
or UO_257 (O_257,N_28418,N_26436);
or UO_258 (O_258,N_25821,N_29110);
nand UO_259 (O_259,N_26829,N_29613);
nand UO_260 (O_260,N_27371,N_26444);
or UO_261 (O_261,N_26187,N_28085);
xor UO_262 (O_262,N_26639,N_29210);
nand UO_263 (O_263,N_25854,N_24989);
nor UO_264 (O_264,N_29121,N_28931);
nand UO_265 (O_265,N_28314,N_24901);
or UO_266 (O_266,N_29930,N_24755);
nor UO_267 (O_267,N_25906,N_24383);
or UO_268 (O_268,N_29500,N_29347);
nor UO_269 (O_269,N_24959,N_28350);
or UO_270 (O_270,N_29990,N_29999);
xnor UO_271 (O_271,N_27411,N_25580);
or UO_272 (O_272,N_24275,N_26357);
and UO_273 (O_273,N_28380,N_26881);
nand UO_274 (O_274,N_27020,N_28487);
nor UO_275 (O_275,N_25577,N_29729);
nand UO_276 (O_276,N_27657,N_28729);
or UO_277 (O_277,N_29376,N_27394);
nor UO_278 (O_278,N_27268,N_24176);
xnor UO_279 (O_279,N_28662,N_24134);
xor UO_280 (O_280,N_28147,N_29877);
nand UO_281 (O_281,N_27089,N_28351);
nor UO_282 (O_282,N_27406,N_27459);
and UO_283 (O_283,N_26106,N_26442);
or UO_284 (O_284,N_28188,N_25740);
and UO_285 (O_285,N_24198,N_26380);
and UO_286 (O_286,N_24186,N_28291);
xnor UO_287 (O_287,N_24912,N_26279);
nand UO_288 (O_288,N_26126,N_29944);
and UO_289 (O_289,N_28579,N_26703);
nor UO_290 (O_290,N_25683,N_28735);
nand UO_291 (O_291,N_26584,N_24925);
and UO_292 (O_292,N_26880,N_26008);
or UO_293 (O_293,N_28210,N_29734);
or UO_294 (O_294,N_26388,N_28769);
or UO_295 (O_295,N_26209,N_24610);
nand UO_296 (O_296,N_26547,N_24017);
xnor UO_297 (O_297,N_25863,N_26285);
or UO_298 (O_298,N_28091,N_26761);
and UO_299 (O_299,N_24142,N_29898);
and UO_300 (O_300,N_29508,N_27236);
nor UO_301 (O_301,N_25160,N_25117);
and UO_302 (O_302,N_26077,N_26218);
xnor UO_303 (O_303,N_25879,N_24259);
xor UO_304 (O_304,N_29597,N_25834);
or UO_305 (O_305,N_24776,N_27912);
nand UO_306 (O_306,N_28890,N_29286);
nor UO_307 (O_307,N_24760,N_29236);
and UO_308 (O_308,N_24431,N_26081);
nand UO_309 (O_309,N_29078,N_29321);
and UO_310 (O_310,N_28189,N_24919);
or UO_311 (O_311,N_26788,N_29466);
xnor UO_312 (O_312,N_27248,N_29014);
and UO_313 (O_313,N_26536,N_28927);
nor UO_314 (O_314,N_29114,N_28386);
and UO_315 (O_315,N_25703,N_25410);
nand UO_316 (O_316,N_25015,N_27237);
xnor UO_317 (O_317,N_25217,N_28666);
nor UO_318 (O_318,N_26206,N_27124);
nand UO_319 (O_319,N_29628,N_28765);
xnor UO_320 (O_320,N_28533,N_24612);
nand UO_321 (O_321,N_28383,N_26103);
nor UO_322 (O_322,N_28817,N_28366);
xnor UO_323 (O_323,N_28970,N_29256);
xor UO_324 (O_324,N_27150,N_28847);
nor UO_325 (O_325,N_27663,N_25537);
nor UO_326 (O_326,N_24107,N_27604);
nand UO_327 (O_327,N_25282,N_28233);
nand UO_328 (O_328,N_27742,N_24903);
nor UO_329 (O_329,N_27963,N_28432);
xor UO_330 (O_330,N_25785,N_29383);
xnor UO_331 (O_331,N_29993,N_27949);
nand UO_332 (O_332,N_24674,N_27926);
nor UO_333 (O_333,N_27416,N_25586);
and UO_334 (O_334,N_25084,N_27677);
xnor UO_335 (O_335,N_25421,N_24249);
nand UO_336 (O_336,N_27927,N_24227);
and UO_337 (O_337,N_26670,N_26836);
and UO_338 (O_338,N_27513,N_26680);
nand UO_339 (O_339,N_25853,N_29398);
nor UO_340 (O_340,N_29368,N_24245);
nor UO_341 (O_341,N_25621,N_24265);
or UO_342 (O_342,N_25140,N_26440);
nor UO_343 (O_343,N_25418,N_29079);
nand UO_344 (O_344,N_24080,N_28771);
or UO_345 (O_345,N_27361,N_25929);
nor UO_346 (O_346,N_24866,N_29609);
nand UO_347 (O_347,N_24262,N_28613);
or UO_348 (O_348,N_24690,N_27114);
or UO_349 (O_349,N_28625,N_27403);
and UO_350 (O_350,N_25530,N_25543);
nand UO_351 (O_351,N_24456,N_24496);
or UO_352 (O_352,N_26825,N_25632);
xnor UO_353 (O_353,N_26123,N_24604);
nor UO_354 (O_354,N_29677,N_27560);
nor UO_355 (O_355,N_25331,N_29984);
nor UO_356 (O_356,N_28263,N_28382);
and UO_357 (O_357,N_24511,N_24763);
xor UO_358 (O_358,N_25590,N_28372);
xnor UO_359 (O_359,N_27620,N_29979);
and UO_360 (O_360,N_24432,N_29143);
or UO_361 (O_361,N_25993,N_28265);
nand UO_362 (O_362,N_27842,N_24440);
nand UO_363 (O_363,N_28554,N_24695);
nand UO_364 (O_364,N_27948,N_29872);
nand UO_365 (O_365,N_28529,N_28976);
xor UO_366 (O_366,N_24230,N_27631);
xnor UO_367 (O_367,N_25037,N_24933);
or UO_368 (O_368,N_28844,N_27117);
or UO_369 (O_369,N_24566,N_26334);
nor UO_370 (O_370,N_27214,N_26478);
nor UO_371 (O_371,N_27532,N_29819);
xor UO_372 (O_372,N_27961,N_27288);
and UO_373 (O_373,N_24614,N_25976);
nand UO_374 (O_374,N_29138,N_29716);
or UO_375 (O_375,N_24985,N_25546);
nor UO_376 (O_376,N_24435,N_26378);
nand UO_377 (O_377,N_29995,N_25749);
or UO_378 (O_378,N_24549,N_24226);
and UO_379 (O_379,N_24639,N_29847);
nor UO_380 (O_380,N_24351,N_27105);
and UO_381 (O_381,N_27684,N_26010);
and UO_382 (O_382,N_28852,N_27841);
and UO_383 (O_383,N_26222,N_24971);
and UO_384 (O_384,N_27369,N_28884);
nor UO_385 (O_385,N_29491,N_27103);
and UO_386 (O_386,N_26720,N_29820);
xnor UO_387 (O_387,N_28552,N_28671);
nor UO_388 (O_388,N_26531,N_27319);
and UO_389 (O_389,N_24932,N_29968);
nand UO_390 (O_390,N_27750,N_25947);
nand UO_391 (O_391,N_24937,N_27893);
and UO_392 (O_392,N_27399,N_26678);
and UO_393 (O_393,N_27883,N_26643);
xnor UO_394 (O_394,N_25387,N_29093);
nand UO_395 (O_395,N_28240,N_25704);
and UO_396 (O_396,N_28563,N_24960);
nand UO_397 (O_397,N_25603,N_28273);
nand UO_398 (O_398,N_24712,N_28336);
and UO_399 (O_399,N_24961,N_29087);
and UO_400 (O_400,N_25150,N_29595);
or UO_401 (O_401,N_25604,N_25732);
or UO_402 (O_402,N_26619,N_25538);
nand UO_403 (O_403,N_29173,N_27541);
nand UO_404 (O_404,N_26429,N_26122);
nand UO_405 (O_405,N_26626,N_25382);
xor UO_406 (O_406,N_27312,N_24970);
xnor UO_407 (O_407,N_26503,N_25121);
or UO_408 (O_408,N_27653,N_25036);
xor UO_409 (O_409,N_24309,N_26353);
and UO_410 (O_410,N_25922,N_25089);
nor UO_411 (O_411,N_29645,N_27804);
nor UO_412 (O_412,N_24768,N_28622);
xor UO_413 (O_413,N_25143,N_27915);
nand UO_414 (O_414,N_25103,N_29289);
xnor UO_415 (O_415,N_27925,N_29539);
xnor UO_416 (O_416,N_26268,N_25100);
and UO_417 (O_417,N_26056,N_26631);
xor UO_418 (O_418,N_24713,N_27768);
xor UO_419 (O_419,N_26613,N_29184);
nand UO_420 (O_420,N_26975,N_24501);
xor UO_421 (O_421,N_27869,N_25815);
or UO_422 (O_422,N_28045,N_28969);
and UO_423 (O_423,N_29287,N_26169);
and UO_424 (O_424,N_24654,N_28481);
nor UO_425 (O_425,N_26031,N_26930);
nand UO_426 (O_426,N_27882,N_25078);
nor UO_427 (O_427,N_29707,N_24556);
or UO_428 (O_428,N_24368,N_27294);
and UO_429 (O_429,N_29308,N_24561);
xor UO_430 (O_430,N_29088,N_24934);
and UO_431 (O_431,N_25276,N_26529);
nand UO_432 (O_432,N_26804,N_29012);
or UO_433 (O_433,N_27668,N_27163);
or UO_434 (O_434,N_26469,N_26233);
or UO_435 (O_435,N_25751,N_24815);
and UO_436 (O_436,N_27649,N_26886);
nand UO_437 (O_437,N_24384,N_24098);
or UO_438 (O_438,N_26480,N_29148);
nor UO_439 (O_439,N_24066,N_29166);
or UO_440 (O_440,N_25210,N_26043);
and UO_441 (O_441,N_29674,N_28841);
nor UO_442 (O_442,N_24321,N_25614);
xnor UO_443 (O_443,N_24203,N_26646);
and UO_444 (O_444,N_24875,N_26164);
nand UO_445 (O_445,N_26462,N_26748);
nand UO_446 (O_446,N_24861,N_24851);
xor UO_447 (O_447,N_26283,N_24308);
nor UO_448 (O_448,N_29694,N_25623);
nand UO_449 (O_449,N_26167,N_27843);
or UO_450 (O_450,N_27051,N_28054);
xor UO_451 (O_451,N_28300,N_29651);
nand UO_452 (O_452,N_27275,N_25607);
nor UO_453 (O_453,N_24822,N_28018);
nand UO_454 (O_454,N_29494,N_25133);
and UO_455 (O_455,N_27553,N_28069);
xor UO_456 (O_456,N_28370,N_27014);
nor UO_457 (O_457,N_27259,N_25893);
or UO_458 (O_458,N_25374,N_28493);
and UO_459 (O_459,N_26381,N_26416);
nand UO_460 (O_460,N_26158,N_27647);
nand UO_461 (O_461,N_28762,N_24332);
nand UO_462 (O_462,N_24980,N_25457);
and UO_463 (O_463,N_24911,N_29747);
and UO_464 (O_464,N_27634,N_29742);
nand UO_465 (O_465,N_28264,N_28862);
or UO_466 (O_466,N_26263,N_29103);
and UO_467 (O_467,N_29018,N_24884);
and UO_468 (O_468,N_25081,N_25910);
and UO_469 (O_469,N_24830,N_25314);
or UO_470 (O_470,N_24333,N_28776);
nand UO_471 (O_471,N_26753,N_25980);
nand UO_472 (O_472,N_28593,N_29650);
nor UO_473 (O_473,N_29975,N_25228);
nand UO_474 (O_474,N_28887,N_28764);
or UO_475 (O_475,N_28032,N_28452);
and UO_476 (O_476,N_25233,N_25249);
or UO_477 (O_477,N_25647,N_28736);
or UO_478 (O_478,N_27734,N_28206);
xor UO_479 (O_479,N_24202,N_24013);
and UO_480 (O_480,N_27220,N_27338);
xnor UO_481 (O_481,N_25411,N_24837);
and UO_482 (O_482,N_24216,N_28405);
and UO_483 (O_483,N_28965,N_28905);
or UO_484 (O_484,N_25885,N_29936);
or UO_485 (O_485,N_26578,N_29132);
xnor UO_486 (O_486,N_29865,N_25248);
nor UO_487 (O_487,N_27262,N_26163);
or UO_488 (O_488,N_26616,N_27525);
nor UO_489 (O_489,N_28036,N_28802);
and UO_490 (O_490,N_26527,N_24465);
nor UO_491 (O_491,N_27708,N_28063);
xor UO_492 (O_492,N_28001,N_24979);
nor UO_493 (O_493,N_28630,N_24816);
nor UO_494 (O_494,N_25919,N_25197);
xor UO_495 (O_495,N_25634,N_25481);
nor UO_496 (O_496,N_29258,N_24029);
or UO_497 (O_497,N_27038,N_28755);
xor UO_498 (O_498,N_25780,N_28504);
nor UO_499 (O_499,N_29373,N_24805);
nor UO_500 (O_500,N_28851,N_26841);
or UO_501 (O_501,N_25030,N_26401);
and UO_502 (O_502,N_26858,N_24161);
nand UO_503 (O_503,N_28664,N_29505);
or UO_504 (O_504,N_27638,N_28728);
xnor UO_505 (O_505,N_25051,N_29988);
or UO_506 (O_506,N_27476,N_29232);
nand UO_507 (O_507,N_26138,N_26092);
nand UO_508 (O_508,N_26242,N_27740);
and UO_509 (O_509,N_25788,N_25871);
nor UO_510 (O_510,N_26902,N_25728);
nand UO_511 (O_511,N_26551,N_27530);
and UO_512 (O_512,N_26605,N_28262);
nor UO_513 (O_513,N_24165,N_27080);
xnor UO_514 (O_514,N_28972,N_24494);
nand UO_515 (O_515,N_29691,N_28807);
nand UO_516 (O_516,N_27328,N_26074);
or UO_517 (O_517,N_27970,N_24554);
or UO_518 (O_518,N_28044,N_25500);
and UO_519 (O_519,N_29827,N_28506);
and UO_520 (O_520,N_24000,N_28308);
nor UO_521 (O_521,N_24694,N_29353);
nand UO_522 (O_522,N_26375,N_25432);
and UO_523 (O_523,N_27046,N_24747);
nand UO_524 (O_524,N_29660,N_25061);
nand UO_525 (O_525,N_25509,N_27602);
xor UO_526 (O_526,N_24180,N_25801);
nand UO_527 (O_527,N_27358,N_25409);
and UO_528 (O_528,N_27890,N_28337);
nand UO_529 (O_529,N_26635,N_25765);
nand UO_530 (O_530,N_28154,N_29325);
xnor UO_531 (O_531,N_29837,N_29562);
or UO_532 (O_532,N_26297,N_27133);
and UO_533 (O_533,N_27441,N_25483);
or UO_534 (O_534,N_24004,N_28275);
nor UO_535 (O_535,N_29962,N_28011);
nor UO_536 (O_536,N_27407,N_25042);
xor UO_537 (O_537,N_26035,N_29905);
nand UO_538 (O_538,N_29247,N_28971);
nand UO_539 (O_539,N_25166,N_24138);
nand UO_540 (O_540,N_29695,N_27627);
nand UO_541 (O_541,N_24942,N_27060);
or UO_542 (O_542,N_27600,N_28528);
and UO_543 (O_543,N_25399,N_28908);
nand UO_544 (O_544,N_28077,N_24039);
and UO_545 (O_545,N_28199,N_28748);
and UO_546 (O_546,N_24310,N_26270);
or UO_547 (O_547,N_29126,N_29058);
nand UO_548 (O_548,N_24318,N_28274);
and UO_549 (O_549,N_29039,N_28271);
nor UO_550 (O_550,N_26861,N_28519);
xor UO_551 (O_551,N_26293,N_25203);
nor UO_552 (O_552,N_25085,N_25951);
xor UO_553 (O_553,N_26750,N_27199);
or UO_554 (O_554,N_26517,N_28228);
and UO_555 (O_555,N_28474,N_28641);
and UO_556 (O_556,N_26014,N_29303);
nand UO_557 (O_557,N_25969,N_29803);
nand UO_558 (O_558,N_29646,N_27664);
nor UO_559 (O_559,N_25290,N_29642);
or UO_560 (O_560,N_27402,N_28864);
nand UO_561 (O_561,N_26542,N_25013);
xor UO_562 (O_562,N_24342,N_27534);
nor UO_563 (O_563,N_29359,N_24529);
nor UO_564 (O_564,N_28700,N_27596);
nor UO_565 (O_565,N_26740,N_26395);
nor UO_566 (O_566,N_25721,N_27209);
and UO_567 (O_567,N_29522,N_27528);
nand UO_568 (O_568,N_29969,N_27360);
nor UO_569 (O_569,N_29307,N_28981);
and UO_570 (O_570,N_28143,N_24157);
xnor UO_571 (O_571,N_26689,N_29224);
and UO_572 (O_572,N_26372,N_26928);
and UO_573 (O_573,N_28793,N_28800);
xnor UO_574 (O_574,N_24294,N_26402);
nor UO_575 (O_575,N_29109,N_26083);
xnor UO_576 (O_576,N_28838,N_28056);
nor UO_577 (O_577,N_27570,N_26883);
and UO_578 (O_578,N_27376,N_24821);
and UO_579 (O_579,N_29006,N_29388);
nor UO_580 (O_580,N_25413,N_27499);
or UO_581 (O_581,N_24734,N_26791);
and UO_582 (O_582,N_28672,N_26363);
and UO_583 (O_583,N_25244,N_28235);
or UO_584 (O_584,N_24023,N_28684);
or UO_585 (O_585,N_24580,N_26744);
and UO_586 (O_586,N_29178,N_24943);
and UO_587 (O_587,N_25918,N_25510);
and UO_588 (O_588,N_25736,N_29903);
nor UO_589 (O_589,N_29636,N_28034);
xnor UO_590 (O_590,N_26407,N_27430);
nor UO_591 (O_591,N_27830,N_24794);
and UO_592 (O_592,N_26772,N_25766);
or UO_593 (O_593,N_26271,N_29770);
xor UO_594 (O_594,N_24077,N_28723);
or UO_595 (O_595,N_24220,N_25339);
nor UO_596 (O_596,N_24448,N_29942);
and UO_597 (O_597,N_27802,N_27764);
or UO_598 (O_598,N_27564,N_26775);
and UO_599 (O_599,N_25445,N_27177);
nor UO_600 (O_600,N_27492,N_25063);
or UO_601 (O_601,N_25526,N_26576);
nand UO_602 (O_602,N_27989,N_29657);
xnor UO_603 (O_603,N_28284,N_28334);
and UO_604 (O_604,N_26595,N_29260);
nor UO_605 (O_605,N_27946,N_26580);
xnor UO_606 (O_606,N_27873,N_24237);
and UO_607 (O_607,N_27234,N_27420);
and UO_608 (O_608,N_26235,N_25804);
xnor UO_609 (O_609,N_24534,N_25629);
nand UO_610 (O_610,N_25841,N_28502);
or UO_611 (O_611,N_25492,N_25334);
nand UO_612 (O_612,N_25529,N_29343);
xnor UO_613 (O_613,N_29177,N_24423);
xnor UO_614 (O_614,N_25934,N_24367);
xnor UO_615 (O_615,N_29420,N_28645);
or UO_616 (O_616,N_28283,N_24083);
nor UO_617 (O_617,N_27257,N_29960);
or UO_618 (O_618,N_27140,N_25440);
xnor UO_619 (O_619,N_28551,N_29682);
nor UO_620 (O_620,N_24928,N_25964);
nor UO_621 (O_621,N_25164,N_27850);
xnor UO_622 (O_622,N_28174,N_24873);
nor UO_623 (O_623,N_24110,N_26682);
nor UO_624 (O_624,N_25195,N_27273);
nand UO_625 (O_625,N_26007,N_29098);
nand UO_626 (O_626,N_29422,N_28341);
xnor UO_627 (O_627,N_25764,N_27113);
or UO_628 (O_628,N_25840,N_29777);
nand UO_629 (O_629,N_27074,N_25496);
or UO_630 (O_630,N_26579,N_24876);
nor UO_631 (O_631,N_29016,N_24018);
and UO_632 (O_632,N_27502,N_29767);
or UO_633 (O_633,N_29471,N_25763);
nor UO_634 (O_634,N_24322,N_26913);
xnor UO_635 (O_635,N_27016,N_29576);
or UO_636 (O_636,N_25700,N_26658);
or UO_637 (O_637,N_25502,N_28002);
or UO_638 (O_638,N_28846,N_29568);
and UO_639 (O_639,N_26811,N_24596);
nor UO_640 (O_640,N_26102,N_25183);
nand UO_641 (O_641,N_24832,N_25477);
and UO_642 (O_642,N_27282,N_24718);
nor UO_643 (O_643,N_24329,N_25760);
nor UO_644 (O_644,N_25856,N_26986);
nor UO_645 (O_645,N_29835,N_27321);
or UO_646 (O_646,N_29331,N_28163);
nand UO_647 (O_647,N_24743,N_26572);
nand UO_648 (O_648,N_24758,N_25223);
and UO_649 (O_649,N_24439,N_25519);
xnor UO_650 (O_650,N_28156,N_25352);
and UO_651 (O_651,N_28378,N_26991);
and UO_652 (O_652,N_27305,N_29938);
nand UO_653 (O_653,N_27284,N_26086);
or UO_654 (O_654,N_25145,N_29344);
or UO_655 (O_655,N_25491,N_24735);
and UO_656 (O_656,N_25392,N_28900);
nor UO_657 (O_657,N_24027,N_24444);
and UO_658 (O_658,N_29670,N_24340);
xor UO_659 (O_659,N_24459,N_28797);
or UO_660 (O_660,N_27581,N_26571);
nor UO_661 (O_661,N_24228,N_29483);
or UO_662 (O_662,N_29643,N_25101);
or UO_663 (O_663,N_25859,N_26726);
nor UO_664 (O_664,N_28584,N_26743);
and UO_665 (O_665,N_29506,N_26042);
xor UO_666 (O_666,N_28535,N_26013);
and UO_667 (O_667,N_25317,N_26134);
and UO_668 (O_668,N_27383,N_26382);
nand UO_669 (O_669,N_25818,N_26188);
or UO_670 (O_670,N_24860,N_28881);
nand UO_671 (O_671,N_27945,N_26849);
and UO_672 (O_672,N_26850,N_24413);
or UO_673 (O_673,N_26617,N_29432);
and UO_674 (O_674,N_29035,N_24050);
xnor UO_675 (O_675,N_25676,N_29804);
or UO_676 (O_676,N_29187,N_27848);
nor UO_677 (O_677,N_28193,N_24242);
nand UO_678 (O_678,N_27977,N_25012);
xor UO_679 (O_679,N_28390,N_25070);
nor UO_680 (O_680,N_27719,N_29231);
xor UO_681 (O_681,N_27111,N_26767);
nand UO_682 (O_682,N_24594,N_25486);
nand UO_683 (O_683,N_25476,N_26620);
or UO_684 (O_684,N_26473,N_28290);
nor UO_685 (O_685,N_27340,N_25515);
nor UO_686 (O_686,N_26420,N_28331);
or UO_687 (O_687,N_24499,N_25066);
and UO_688 (O_688,N_28984,N_24303);
or UO_689 (O_689,N_26640,N_28467);
xnor UO_690 (O_690,N_29191,N_25875);
nand UO_691 (O_691,N_25888,N_26651);
nand UO_692 (O_692,N_24711,N_24052);
or UO_693 (O_693,N_25914,N_29479);
nor UO_694 (O_694,N_27243,N_28549);
xor UO_695 (O_695,N_29356,N_27232);
nor UO_696 (O_696,N_27671,N_24609);
or UO_697 (O_697,N_25048,N_28358);
xnor UO_698 (O_698,N_29404,N_24450);
nor UO_699 (O_699,N_28031,N_29796);
or UO_700 (O_700,N_25371,N_29705);
xnor UO_701 (O_701,N_25570,N_29405);
nand UO_702 (O_702,N_29424,N_27973);
nand UO_703 (O_703,N_29156,N_24143);
or UO_704 (O_704,N_28661,N_24998);
xor UO_705 (O_705,N_24054,N_24635);
xnor UO_706 (O_706,N_27333,N_27916);
nand UO_707 (O_707,N_29638,N_25908);
nand UO_708 (O_708,N_26144,N_24177);
nor UO_709 (O_709,N_24946,N_24486);
nand UO_710 (O_710,N_27810,N_29977);
or UO_711 (O_711,N_25180,N_28732);
nor UO_712 (O_712,N_28020,N_24786);
or UO_713 (O_713,N_26543,N_27968);
and UO_714 (O_714,N_25059,N_24941);
xor UO_715 (O_715,N_28316,N_29421);
or UO_716 (O_716,N_29160,N_27280);
and UO_717 (O_717,N_25937,N_24834);
and UO_718 (O_718,N_28395,N_29057);
and UO_719 (O_719,N_27246,N_24949);
nor UO_720 (O_720,N_29640,N_25786);
xnor UO_721 (O_721,N_24600,N_24009);
xnor UO_722 (O_722,N_26945,N_26786);
or UO_723 (O_723,N_25829,N_28412);
nor UO_724 (O_724,N_28169,N_29390);
xnor UO_725 (O_725,N_25582,N_25376);
xor UO_726 (O_726,N_25262,N_26510);
nand UO_727 (O_727,N_27903,N_29323);
nand UO_728 (O_728,N_29537,N_25664);
or UO_729 (O_729,N_25783,N_27795);
xnor UO_730 (O_730,N_24720,N_26349);
and UO_731 (O_731,N_28717,N_25665);
and UO_732 (O_732,N_26734,N_28788);
nand UO_733 (O_733,N_26457,N_25787);
xor UO_734 (O_734,N_26305,N_29759);
nor UO_735 (O_735,N_29139,N_29255);
nor UO_736 (O_736,N_25520,N_29310);
or UO_737 (O_737,N_24551,N_25299);
or UO_738 (O_738,N_28049,N_28244);
nand UO_739 (O_739,N_24201,N_29546);
xnor UO_740 (O_740,N_26071,N_27931);
and UO_741 (O_741,N_27184,N_24809);
nand UO_742 (O_742,N_26095,N_26114);
nand UO_743 (O_743,N_26237,N_26454);
or UO_744 (O_744,N_25658,N_27179);
nand UO_745 (O_745,N_25904,N_29737);
nor UO_746 (O_746,N_28161,N_26781);
nand UO_747 (O_747,N_29919,N_29632);
xnor UO_748 (O_748,N_28774,N_25558);
nor UO_749 (O_749,N_29267,N_27366);
and UO_750 (O_750,N_28624,N_28515);
or UO_751 (O_751,N_26497,N_27019);
and UO_752 (O_752,N_24434,N_28141);
nand UO_753 (O_753,N_26234,N_25584);
nor UO_754 (O_754,N_27365,N_28442);
nand UO_755 (O_755,N_29229,N_29800);
and UO_756 (O_756,N_27984,N_27283);
xnor UO_757 (O_757,N_28878,N_24730);
nand UO_758 (O_758,N_27497,N_29589);
nand UO_759 (O_759,N_24923,N_28996);
nor UO_760 (O_760,N_26768,N_26170);
nand UO_761 (O_761,N_26475,N_25324);
nor UO_762 (O_762,N_26568,N_29416);
or UO_763 (O_763,N_25564,N_29955);
nor UO_764 (O_764,N_25056,N_27875);
nand UO_765 (O_765,N_28867,N_29542);
or UO_766 (O_766,N_26481,N_29333);
and UO_767 (O_767,N_27937,N_24056);
xnor UO_768 (O_768,N_25107,N_26139);
nor UO_769 (O_769,N_27813,N_26780);
nor UO_770 (O_770,N_24032,N_27718);
or UO_771 (O_771,N_28604,N_24483);
nor UO_772 (O_772,N_29888,N_27972);
nand UO_773 (O_773,N_29524,N_27225);
xor UO_774 (O_774,N_26282,N_24563);
nand UO_775 (O_775,N_28781,N_27374);
and UO_776 (O_776,N_27722,N_28473);
nor UO_777 (O_777,N_27349,N_26403);
nor UO_778 (O_778,N_24835,N_25655);
xor UO_779 (O_779,N_29075,N_28131);
xor UO_780 (O_780,N_26716,N_25236);
nor UO_781 (O_781,N_24838,N_27847);
or UO_782 (O_782,N_25343,N_27622);
and UO_783 (O_783,N_27077,N_25426);
nand UO_784 (O_784,N_26717,N_27846);
and UO_785 (O_785,N_25744,N_24782);
and UO_786 (O_786,N_29815,N_27084);
and UO_787 (O_787,N_25444,N_26393);
nor UO_788 (O_788,N_28312,N_26671);
and UO_789 (O_789,N_25250,N_29115);
or UO_790 (O_790,N_26943,N_26967);
nand UO_791 (O_791,N_29013,N_27728);
nor UO_792 (O_792,N_29452,N_25258);
or UO_793 (O_793,N_27861,N_24533);
nor UO_794 (O_794,N_28310,N_24684);
and UO_795 (O_795,N_28768,N_28919);
xnor UO_796 (O_796,N_25813,N_25733);
nand UO_797 (O_797,N_25388,N_25695);
and UO_798 (O_798,N_27651,N_24965);
xnor UO_799 (O_799,N_28922,N_27770);
or UO_800 (O_800,N_29162,N_25593);
nor UO_801 (O_801,N_29981,N_24358);
xor UO_802 (O_802,N_26359,N_27212);
or UO_803 (O_803,N_25925,N_29611);
or UO_804 (O_804,N_26779,N_29180);
and UO_805 (O_805,N_28999,N_29560);
xor UO_806 (O_806,N_26688,N_28719);
xor UO_807 (O_807,N_28195,N_25775);
or UO_808 (O_808,N_29940,N_26039);
and UO_809 (O_809,N_27748,N_26919);
or UO_810 (O_810,N_27661,N_28157);
xnor UO_811 (O_811,N_25557,N_26837);
or UO_812 (O_812,N_29346,N_25866);
nor UO_813 (O_813,N_24991,N_28258);
nand UO_814 (O_814,N_27149,N_26437);
xnor UO_815 (O_815,N_26810,N_24001);
xor UO_816 (O_816,N_27829,N_25986);
or UO_817 (O_817,N_27552,N_25978);
and UO_818 (O_818,N_24108,N_29213);
nand UO_819 (O_819,N_26418,N_25028);
and UO_820 (O_820,N_29659,N_29547);
or UO_821 (O_821,N_29808,N_24854);
and UO_822 (O_822,N_25846,N_26323);
nor UO_823 (O_823,N_24859,N_24793);
xor UO_824 (O_824,N_28942,N_28414);
nand UO_825 (O_825,N_29204,N_26649);
nor UO_826 (O_826,N_25353,N_24336);
xor UO_827 (O_827,N_27147,N_27891);
nand UO_828 (O_828,N_25163,N_24723);
nor UO_829 (O_829,N_29899,N_29251);
nor UO_830 (O_830,N_26156,N_26970);
xor UO_831 (O_831,N_29429,N_25832);
and UO_832 (O_832,N_25361,N_26566);
nor UO_833 (O_833,N_28448,N_28983);
nor UO_834 (O_834,N_24538,N_26612);
and UO_835 (O_835,N_25691,N_27503);
xnor UO_836 (O_836,N_26160,N_24231);
and UO_837 (O_837,N_26383,N_26792);
and UO_838 (O_838,N_27994,N_26062);
nor UO_839 (O_839,N_26260,N_26018);
nand UO_840 (O_840,N_25313,N_26623);
xor UO_841 (O_841,N_27157,N_25087);
nor UO_842 (O_842,N_24028,N_28567);
and UO_843 (O_843,N_26392,N_27694);
xnor UO_844 (O_844,N_24286,N_28469);
xor UO_845 (O_845,N_27224,N_29915);
nand UO_846 (O_846,N_26895,N_25770);
xnor UO_847 (O_847,N_25199,N_25495);
and UO_848 (O_848,N_25058,N_26842);
nand UO_849 (O_849,N_28633,N_28426);
or UO_850 (O_850,N_27510,N_27299);
and UO_851 (O_851,N_25870,N_25458);
and UO_852 (O_852,N_28526,N_27227);
or UO_853 (O_853,N_28477,N_29025);
nor UO_854 (O_854,N_29335,N_27982);
nand UO_855 (O_855,N_27609,N_29579);
nor UO_856 (O_856,N_25828,N_24015);
and UO_857 (O_857,N_25709,N_27352);
or UO_858 (O_858,N_27192,N_28229);
nor UO_859 (O_859,N_28958,N_24064);
xor UO_860 (O_860,N_24645,N_25613);
nor UO_861 (O_861,N_27688,N_28421);
nand UO_862 (O_862,N_26472,N_27195);
nor UO_863 (O_863,N_25669,N_29084);
nand UO_864 (O_864,N_24802,N_26819);
xor UO_865 (O_865,N_25167,N_26933);
nand UO_866 (O_866,N_29832,N_28064);
nand UO_867 (O_867,N_25207,N_25659);
or UO_868 (O_868,N_25667,N_28030);
and UO_869 (O_869,N_26989,N_26695);
or UO_870 (O_870,N_26231,N_26766);
nor UO_871 (O_871,N_27469,N_29552);
nor UO_872 (O_872,N_25351,N_26366);
nand UO_873 (O_873,N_24158,N_29174);
and UO_874 (O_874,N_26956,N_29152);
nand UO_875 (O_875,N_28621,N_29882);
or UO_876 (O_876,N_29743,N_24750);
xnor UO_877 (O_877,N_24647,N_24206);
and UO_878 (O_878,N_28105,N_24767);
or UO_879 (O_879,N_28225,N_26505);
xnor UO_880 (O_880,N_26952,N_24883);
nand UO_881 (O_881,N_28766,N_26172);
xnor UO_882 (O_882,N_25820,N_24250);
nand UO_883 (O_883,N_24395,N_29850);
and UO_884 (O_884,N_29111,N_24789);
and UO_885 (O_885,N_26066,N_28514);
and UO_886 (O_886,N_29859,N_29246);
and UO_887 (O_887,N_26575,N_25346);
nand UO_888 (O_888,N_29288,N_27952);
and UO_889 (O_889,N_29355,N_28342);
nor UO_890 (O_890,N_25357,N_25971);
nand UO_891 (O_891,N_28738,N_24550);
xor UO_892 (O_892,N_26730,N_25996);
nand UO_893 (O_893,N_24994,N_24192);
nand UO_894 (O_894,N_29205,N_29970);
nand UO_895 (O_895,N_28658,N_25345);
or UO_896 (O_896,N_24620,N_29298);
xor UO_897 (O_897,N_26591,N_25219);
nor UO_898 (O_898,N_28086,N_25355);
nor UO_899 (O_899,N_25527,N_28688);
nor UO_900 (O_900,N_27944,N_29361);
or UO_901 (O_901,N_25741,N_29699);
nand UO_902 (O_902,N_24069,N_28560);
xnor UO_903 (O_903,N_26046,N_27561);
xor UO_904 (O_904,N_27832,N_24675);
nor UO_905 (O_905,N_24179,N_24140);
xor UO_906 (O_906,N_25480,N_29941);
and UO_907 (O_907,N_27698,N_24636);
nor UO_908 (O_908,N_29277,N_29393);
and UO_909 (O_909,N_24184,N_26805);
nor UO_910 (O_910,N_27712,N_27489);
nand UO_911 (O_911,N_25750,N_25661);
xor UO_912 (O_912,N_27645,N_28650);
nor UO_913 (O_913,N_24189,N_27166);
xnor UO_914 (O_914,N_24990,N_25191);
nand UO_915 (O_915,N_24191,N_24159);
nor UO_916 (O_916,N_24031,N_25790);
or UO_917 (O_917,N_25019,N_25148);
and UO_918 (O_918,N_29592,N_26476);
and UO_919 (O_919,N_26873,N_28591);
nor UO_920 (O_920,N_24921,N_25377);
nor UO_921 (O_921,N_28145,N_24285);
xnor UO_922 (O_922,N_29279,N_25464);
nor UO_923 (O_923,N_28581,N_25185);
and UO_924 (O_924,N_28557,N_26537);
nor UO_925 (O_925,N_29149,N_24260);
nand UO_926 (O_926,N_29839,N_26851);
xor UO_927 (O_927,N_24856,N_24892);
nor UO_928 (O_928,N_25631,N_24427);
and UO_929 (O_929,N_29578,N_25177);
or UO_930 (O_930,N_27607,N_24305);
xor UO_931 (O_931,N_25055,N_29851);
nand UO_932 (O_932,N_26036,N_25443);
and UO_933 (O_933,N_24870,N_29647);
xnor UO_934 (O_934,N_25895,N_29252);
nor UO_935 (O_935,N_26165,N_27716);
nand UO_936 (O_936,N_26002,N_29570);
xor UO_937 (O_937,N_25029,N_24210);
xor UO_938 (O_938,N_27081,N_26999);
or UO_939 (O_939,N_28106,N_26546);
and UO_940 (O_940,N_24474,N_26346);
and UO_941 (O_941,N_25112,N_25243);
and UO_942 (O_942,N_26932,N_26746);
xor UO_943 (O_943,N_29372,N_27432);
or UO_944 (O_944,N_24141,N_26757);
or UO_945 (O_945,N_26936,N_29413);
and UO_946 (O_946,N_29527,N_27006);
nor UO_947 (O_947,N_27771,N_24215);
or UO_948 (O_948,N_26448,N_24666);
nor UO_949 (O_949,N_26847,N_29516);
nand UO_950 (O_950,N_29273,N_26563);
xnor UO_951 (O_951,N_27219,N_24218);
and UO_952 (O_952,N_24710,N_29809);
or UO_953 (O_953,N_29226,N_24217);
or UO_954 (O_954,N_26141,N_28068);
xor UO_955 (O_955,N_25194,N_25900);
and UO_956 (O_956,N_27690,N_25381);
xor UO_957 (O_957,N_27290,N_29985);
nor UO_958 (O_958,N_24582,N_28946);
or UO_959 (O_959,N_29357,N_24703);
and UO_960 (O_960,N_27555,N_24724);
nor UO_961 (O_961,N_27344,N_24290);
xnor UO_962 (O_962,N_29854,N_25945);
nand UO_963 (O_963,N_29896,N_25847);
nand UO_964 (O_964,N_29771,N_27508);
nor UO_965 (O_965,N_27141,N_26754);
nor UO_966 (O_966,N_24008,N_28754);
or UO_967 (O_967,N_26972,N_25057);
and UO_968 (O_968,N_24924,N_25026);
xnor UO_969 (O_969,N_25316,N_27491);
and UO_970 (O_970,N_28246,N_28349);
nand UO_971 (O_971,N_29544,N_28932);
nor UO_972 (O_972,N_25241,N_27456);
and UO_973 (O_973,N_28697,N_26216);
nor UO_974 (O_974,N_28564,N_29312);
or UO_975 (O_975,N_24493,N_24044);
or UO_976 (O_976,N_27277,N_24798);
nor UO_977 (O_977,N_25420,N_28516);
and UO_978 (O_978,N_26098,N_24686);
or UO_979 (O_979,N_27911,N_24905);
nand UO_980 (O_980,N_28855,N_29751);
nor UO_981 (O_981,N_27175,N_27395);
xor UO_982 (O_982,N_25768,N_25049);
nor UO_983 (O_983,N_25889,N_26199);
and UO_984 (O_984,N_28991,N_29176);
nand UO_985 (O_985,N_28216,N_27901);
nand UO_986 (O_986,N_27821,N_27071);
nor UO_987 (O_987,N_27887,N_29883);
and UO_988 (O_988,N_29367,N_29470);
nor UO_989 (O_989,N_26220,N_26755);
or UO_990 (O_990,N_28110,N_25720);
xnor UO_991 (O_991,N_29814,N_25306);
and UO_992 (O_992,N_26254,N_29614);
xnor UO_993 (O_993,N_29681,N_25122);
and UO_994 (O_994,N_24472,N_24344);
and UO_995 (O_995,N_25911,N_26641);
nand UO_996 (O_996,N_27056,N_28575);
and UO_997 (O_997,N_24247,N_25090);
or UO_998 (O_998,N_24394,N_27386);
nor UO_999 (O_999,N_27130,N_24719);
and UO_1000 (O_1000,N_24567,N_25129);
nand UO_1001 (O_1001,N_29209,N_29856);
or UO_1002 (O_1002,N_25465,N_27702);
xnor UO_1003 (O_1003,N_26645,N_29118);
or UO_1004 (O_1004,N_28973,N_26915);
and UO_1005 (O_1005,N_27057,N_28410);
or UO_1006 (O_1006,N_25974,N_24513);
nand UO_1007 (O_1007,N_27151,N_25162);
nand UO_1008 (O_1008,N_28224,N_25020);
and UO_1009 (O_1009,N_28711,N_26684);
or UO_1010 (O_1010,N_29724,N_28201);
or UO_1011 (O_1011,N_25259,N_28941);
nor UO_1012 (O_1012,N_26876,N_26548);
and UO_1013 (O_1013,N_28212,N_26258);
xnor UO_1014 (O_1014,N_29490,N_27495);
or UO_1015 (O_1015,N_24913,N_26545);
and UO_1016 (O_1016,N_24678,N_26344);
nand UO_1017 (O_1017,N_28731,N_25938);
nand UO_1018 (O_1018,N_25493,N_29649);
nor UO_1019 (O_1019,N_29974,N_27853);
nand UO_1020 (O_1020,N_26508,N_28598);
and UO_1021 (O_1021,N_27957,N_26729);
xnor UO_1022 (O_1022,N_25547,N_28937);
nor UO_1023 (O_1023,N_28879,N_27818);
xor UO_1024 (O_1024,N_29487,N_24886);
xor UO_1025 (O_1025,N_25151,N_29015);
or UO_1026 (O_1026,N_26340,N_26751);
or UO_1027 (O_1027,N_24320,N_26072);
xnor UO_1028 (O_1028,N_26177,N_28569);
xor UO_1029 (O_1029,N_25684,N_26914);
or UO_1030 (O_1030,N_24757,N_26463);
nand UO_1031 (O_1031,N_29738,N_28587);
nand UO_1032 (O_1032,N_25511,N_29708);
or UO_1033 (O_1033,N_25930,N_24788);
and UO_1034 (O_1034,N_29094,N_26777);
nand UO_1035 (O_1035,N_29358,N_25307);
or UO_1036 (O_1036,N_26824,N_24407);
nand UO_1037 (O_1037,N_26843,N_29047);
xnor UO_1038 (O_1038,N_26644,N_24019);
or UO_1039 (O_1039,N_24602,N_28444);
and UO_1040 (O_1040,N_25111,N_28543);
or UO_1041 (O_1041,N_28429,N_24650);
nand UO_1042 (O_1042,N_25592,N_28057);
or UO_1043 (O_1043,N_25616,N_25416);
nand UO_1044 (O_1044,N_26501,N_27159);
xnor UO_1045 (O_1045,N_25902,N_27180);
nor UO_1046 (O_1046,N_24825,N_29197);
and UO_1047 (O_1047,N_26884,N_26982);
nand UO_1048 (O_1048,N_26676,N_26322);
xnor UO_1049 (O_1049,N_27144,N_24778);
xor UO_1050 (O_1050,N_25713,N_25300);
nand UO_1051 (O_1051,N_27924,N_29360);
or UO_1052 (O_1052,N_27595,N_29097);
and UO_1053 (O_1053,N_26672,N_28413);
nor UO_1054 (O_1054,N_27438,N_29005);
or UO_1055 (O_1055,N_25441,N_26877);
nor UO_1056 (O_1056,N_27210,N_24667);
nor UO_1057 (O_1057,N_24006,N_26983);
or UO_1058 (O_1058,N_28190,N_26709);
nand UO_1059 (O_1059,N_24833,N_28623);
nor UO_1060 (O_1060,N_29871,N_27474);
or UO_1061 (O_1061,N_26410,N_26533);
nor UO_1062 (O_1062,N_25641,N_28183);
xnor UO_1063 (O_1063,N_29384,N_27884);
xnor UO_1064 (O_1064,N_26756,N_24950);
or UO_1065 (O_1065,N_27457,N_26446);
xnor UO_1066 (O_1066,N_27537,N_26585);
or UO_1067 (O_1067,N_29216,N_26465);
or UO_1068 (O_1068,N_28799,N_27327);
nor UO_1069 (O_1069,N_28303,N_29818);
and UO_1070 (O_1070,N_26687,N_26715);
xor UO_1071 (O_1071,N_24451,N_28241);
or UO_1072 (O_1072,N_25127,N_24973);
nor UO_1073 (O_1073,N_29030,N_24282);
and UO_1074 (O_1074,N_24784,N_26866);
nor UO_1075 (O_1075,N_25672,N_26691);
or UO_1076 (O_1076,N_28089,N_28419);
xor UO_1077 (O_1077,N_27675,N_25835);
and UO_1078 (O_1078,N_26925,N_29824);
nor UO_1079 (O_1079,N_25278,N_26445);
and UO_1080 (O_1080,N_25404,N_28456);
or UO_1081 (O_1081,N_29082,N_27834);
and UO_1082 (O_1082,N_29199,N_24606);
and UO_1083 (O_1083,N_25235,N_26131);
nand UO_1084 (O_1084,N_28165,N_29010);
and UO_1085 (O_1085,N_27625,N_26301);
xnor UO_1086 (O_1086,N_26711,N_27908);
xor UO_1087 (O_1087,N_27640,N_24297);
xnor UO_1088 (O_1088,N_27486,N_28356);
xnor UO_1089 (O_1089,N_25192,N_24618);
or UO_1090 (O_1090,N_28281,N_29234);
or UO_1091 (O_1091,N_29048,N_24097);
nand UO_1092 (O_1092,N_25161,N_27465);
nand UO_1093 (O_1093,N_24096,N_27575);
xor UO_1094 (O_1094,N_27435,N_26435);
and UO_1095 (O_1095,N_26500,N_27413);
nand UO_1096 (O_1096,N_27172,N_24422);
xnor UO_1097 (O_1097,N_29833,N_24729);
xor UO_1098 (O_1098,N_26962,N_29569);
xnor UO_1099 (O_1099,N_28327,N_27298);
or UO_1100 (O_1100,N_25753,N_25093);
or UO_1101 (O_1101,N_28858,N_27868);
or UO_1102 (O_1102,N_28309,N_25099);
nand UO_1103 (O_1103,N_29230,N_29698);
and UO_1104 (O_1104,N_29290,N_25052);
nor UO_1105 (O_1105,N_25106,N_29543);
or UO_1106 (O_1106,N_29849,N_24167);
nand UO_1107 (O_1107,N_29475,N_29561);
or UO_1108 (O_1108,N_28234,N_25482);
or UO_1109 (O_1109,N_24887,N_27029);
nand UO_1110 (O_1110,N_24895,N_29710);
xor UO_1111 (O_1111,N_28827,N_25727);
nand UO_1112 (O_1112,N_27666,N_28849);
or UO_1113 (O_1113,N_24504,N_24591);
and UO_1114 (O_1114,N_28739,N_24553);
nor UO_1115 (O_1115,N_26316,N_27897);
nor UO_1116 (O_1116,N_29718,N_29518);
nand UO_1117 (O_1117,N_25833,N_25748);
nand UO_1118 (O_1118,N_24781,N_26397);
and UO_1119 (O_1119,N_25759,N_24721);
and UO_1120 (O_1120,N_28903,N_29023);
or UO_1121 (O_1121,N_28424,N_25861);
xnor UO_1122 (O_1122,N_29061,N_26484);
nor UO_1123 (O_1123,N_27660,N_28995);
nand UO_1124 (O_1124,N_24775,N_29669);
xor UO_1125 (O_1125,N_29510,N_24323);
and UO_1126 (O_1126,N_24590,N_29386);
nand UO_1127 (O_1127,N_24364,N_26076);
nor UO_1128 (O_1128,N_26314,N_26922);
nand UO_1129 (O_1129,N_26589,N_24983);
nand UO_1130 (O_1130,N_26386,N_28761);
nand UO_1131 (O_1131,N_28406,N_28730);
and UO_1132 (O_1132,N_28285,N_27419);
xor UO_1133 (O_1133,N_24902,N_28986);
and UO_1134 (O_1134,N_29122,N_24831);
xnor UO_1135 (O_1135,N_27752,N_28869);
nand UO_1136 (O_1136,N_28834,N_29711);
nand UO_1137 (O_1137,N_25238,N_29593);
and UO_1138 (O_1138,N_28127,N_28968);
nor UO_1139 (O_1139,N_25660,N_28423);
and UO_1140 (O_1140,N_29926,N_27035);
and UO_1141 (O_1141,N_27687,N_29313);
xnor UO_1142 (O_1142,N_25200,N_27058);
or UO_1143 (O_1143,N_28250,N_24071);
or UO_1144 (O_1144,N_24473,N_27440);
or UO_1145 (O_1145,N_25092,N_24457);
nor UO_1146 (O_1146,N_29945,N_28376);
xor UO_1147 (O_1147,N_24956,N_24485);
and UO_1148 (O_1148,N_29622,N_29293);
and UO_1149 (O_1149,N_27816,N_25405);
nand UO_1150 (O_1150,N_25625,N_27526);
and UO_1151 (O_1151,N_25033,N_28248);
or UO_1152 (O_1152,N_28789,N_24524);
xnor UO_1153 (O_1153,N_26513,N_29300);
nand UO_1154 (O_1154,N_27036,N_26582);
nand UO_1155 (O_1155,N_25677,N_27082);
and UO_1156 (O_1156,N_25598,N_28103);
nor UO_1157 (O_1157,N_24099,N_27473);
xnor UO_1158 (O_1158,N_26374,N_29129);
xnor UO_1159 (O_1159,N_26159,N_27477);
nor UO_1160 (O_1160,N_28631,N_27635);
and UO_1161 (O_1161,N_26162,N_27304);
and UO_1162 (O_1162,N_29715,N_24419);
or UO_1163 (O_1163,N_26878,N_24460);
nand UO_1164 (O_1164,N_25415,N_26453);
or UO_1165 (O_1165,N_28745,N_27482);
or UO_1166 (O_1166,N_26133,N_29530);
nand UO_1167 (O_1167,N_28313,N_26180);
nand UO_1168 (O_1168,N_25010,N_25378);
nor UO_1169 (O_1169,N_29842,N_29639);
and UO_1170 (O_1170,N_27254,N_29203);
xnor UO_1171 (O_1171,N_27146,N_29574);
nand UO_1172 (O_1172,N_29482,N_29055);
or UO_1173 (O_1173,N_29041,N_24101);
or UO_1174 (O_1174,N_25795,N_29998);
and UO_1175 (O_1175,N_29983,N_24689);
xnor UO_1176 (O_1176,N_28219,N_24489);
and UO_1177 (O_1177,N_29281,N_24571);
and UO_1178 (O_1178,N_24488,N_28562);
and UO_1179 (O_1179,N_28832,N_29445);
nor UO_1180 (O_1180,N_29020,N_27809);
or UO_1181 (O_1181,N_29996,N_24382);
nand UO_1182 (O_1182,N_28116,N_28523);
or UO_1183 (O_1183,N_26892,N_28636);
xor UO_1184 (O_1184,N_29170,N_25540);
or UO_1185 (O_1185,N_29829,N_24145);
nand UO_1186 (O_1186,N_27579,N_27950);
nor UO_1187 (O_1187,N_29485,N_28861);
nor UO_1188 (O_1188,N_28009,N_26974);
xnor UO_1189 (O_1189,N_24772,N_24370);
xnor UO_1190 (O_1190,N_27011,N_28252);
and UO_1191 (O_1191,N_26988,N_24593);
and UO_1192 (O_1192,N_28468,N_24699);
xnor UO_1193 (O_1193,N_26171,N_29297);
nor UO_1194 (O_1194,N_24519,N_27676);
and UO_1195 (O_1195,N_24214,N_28854);
and UO_1196 (O_1196,N_24693,N_28203);
nor UO_1197 (O_1197,N_28400,N_29438);
and UO_1198 (O_1198,N_25873,N_24560);
nor UO_1199 (O_1199,N_28885,N_28850);
nand UO_1200 (O_1200,N_26075,N_29140);
nand UO_1201 (O_1201,N_28307,N_24059);
nand UO_1202 (O_1202,N_26978,N_24055);
xor UO_1203 (O_1203,N_28437,N_25757);
and UO_1204 (O_1204,N_27824,N_24670);
or UO_1205 (O_1205,N_25329,N_26969);
nor UO_1206 (O_1206,N_28674,N_25453);
xnor UO_1207 (O_1207,N_29280,N_29541);
and UO_1208 (O_1208,N_27143,N_27249);
xnor UO_1209 (O_1209,N_29704,N_26882);
and UO_1210 (O_1210,N_25043,N_27726);
and UO_1211 (O_1211,N_28997,N_27379);
nand UO_1212 (O_1212,N_26570,N_26048);
or UO_1213 (O_1213,N_25807,N_28175);
xor UO_1214 (O_1214,N_24890,N_25802);
or UO_1215 (O_1215,N_24452,N_29120);
nand UO_1216 (O_1216,N_28696,N_27870);
nor UO_1217 (O_1217,N_26509,N_27064);
nand UO_1218 (O_1218,N_24507,N_27573);
nor UO_1219 (O_1219,N_29342,N_25468);
nor UO_1220 (O_1220,N_24545,N_29276);
xnor UO_1221 (O_1221,N_29810,N_26459);
or UO_1222 (O_1222,N_25688,N_25242);
or UO_1223 (O_1223,N_29836,N_26468);
xor UO_1224 (O_1224,N_27378,N_24289);
and UO_1225 (O_1225,N_25064,N_28028);
and UO_1226 (O_1226,N_28907,N_28257);
and UO_1227 (O_1227,N_25384,N_24378);
nor UO_1228 (O_1228,N_24541,N_24252);
nand UO_1229 (O_1229,N_24412,N_27987);
nand UO_1230 (O_1230,N_28484,N_26244);
xor UO_1231 (O_1231,N_25168,N_24592);
nand UO_1232 (O_1232,N_26425,N_28974);
or UO_1233 (O_1233,N_28648,N_27695);
xor UO_1234 (O_1234,N_24229,N_27251);
nand UO_1235 (O_1235,N_26600,N_25041);
nor UO_1236 (O_1236,N_24078,N_28635);
xor UO_1237 (O_1237,N_24665,N_26656);
nand UO_1238 (O_1238,N_28084,N_24154);
and UO_1239 (O_1239,N_29283,N_28100);
nor UO_1240 (O_1240,N_28295,N_27775);
nor UO_1241 (O_1241,N_26019,N_25456);
or UO_1242 (O_1242,N_26690,N_24897);
or UO_1243 (O_1243,N_25386,N_29101);
nand UO_1244 (O_1244,N_27194,N_24374);
nand UO_1245 (O_1245,N_28694,N_29419);
or UO_1246 (O_1246,N_27337,N_27576);
and UO_1247 (O_1247,N_25461,N_29067);
xor UO_1248 (O_1248,N_29274,N_26993);
nand UO_1249 (O_1249,N_24709,N_24685);
xor UO_1250 (O_1250,N_26526,N_24148);
or UO_1251 (O_1251,N_28019,N_29179);
nand UO_1252 (O_1252,N_29957,N_27451);
nand UO_1253 (O_1253,N_29588,N_29831);
nand UO_1254 (O_1254,N_29459,N_25252);
nand UO_1255 (O_1255,N_24627,N_26261);
and UO_1256 (O_1256,N_28058,N_28600);
xor UO_1257 (O_1257,N_26111,N_27738);
nor UO_1258 (O_1258,N_27446,N_26927);
nor UO_1259 (O_1259,N_29239,N_25940);
and UO_1260 (O_1260,N_28416,N_24559);
xnor UO_1261 (O_1261,N_24539,N_26512);
nand UO_1262 (O_1262,N_28439,N_26466);
or UO_1263 (O_1263,N_26219,N_24547);
xnor UO_1264 (O_1264,N_26835,N_29761);
nand UO_1265 (O_1265,N_28146,N_27724);
or UO_1266 (O_1266,N_25288,N_24525);
and UO_1267 (O_1267,N_28656,N_24092);
xnor UO_1268 (O_1268,N_28478,N_25851);
and UO_1269 (O_1269,N_26960,N_25060);
nor UO_1270 (O_1270,N_28906,N_27582);
and UO_1271 (O_1271,N_27654,N_28408);
xor UO_1272 (O_1272,N_25517,N_29533);
and UO_1273 (O_1273,N_27355,N_29992);
nand UO_1274 (O_1274,N_25521,N_24331);
nor UO_1275 (O_1275,N_26411,N_27757);
nand UO_1276 (O_1276,N_27992,N_29304);
and UO_1277 (O_1277,N_29150,N_29582);
or UO_1278 (O_1278,N_28652,N_25972);
nor UO_1279 (O_1279,N_24535,N_28749);
nor UO_1280 (O_1280,N_25045,N_29336);
or UO_1281 (O_1281,N_24366,N_28155);
nor UO_1282 (O_1282,N_26916,N_28286);
nand UO_1283 (O_1283,N_28476,N_25301);
nor UO_1284 (O_1284,N_27381,N_25845);
nand UO_1285 (O_1285,N_24981,N_27387);
nor UO_1286 (O_1286,N_26130,N_24753);
xor UO_1287 (O_1287,N_29049,N_24204);
nor UO_1288 (O_1288,N_27434,N_25499);
nor UO_1289 (O_1289,N_29107,N_26994);
nor UO_1290 (O_1290,N_24544,N_29773);
nor UO_1291 (O_1291,N_28826,N_29909);
or UO_1292 (O_1292,N_27490,N_24621);
nand UO_1293 (O_1293,N_25942,N_26890);
and UO_1294 (O_1294,N_25758,N_28726);
xor UO_1295 (O_1295,N_29022,N_24799);
or UO_1296 (O_1296,N_29052,N_24725);
nand UO_1297 (O_1297,N_28618,N_29212);
nor UO_1298 (O_1298,N_26471,N_26304);
nor UO_1299 (O_1299,N_27501,N_28808);
xnor UO_1300 (O_1300,N_29311,N_26507);
and UO_1301 (O_1301,N_25006,N_24293);
and UO_1302 (O_1302,N_24843,N_29566);
xor UO_1303 (O_1303,N_26795,N_26321);
or UO_1304 (O_1304,N_26846,N_28912);
nor UO_1305 (O_1305,N_29594,N_24392);
xnor UO_1306 (O_1306,N_29417,N_29687);
xor UO_1307 (O_1307,N_25610,N_27242);
xnor UO_1308 (O_1308,N_27426,N_24974);
and UO_1309 (O_1309,N_27986,N_29201);
nor UO_1310 (O_1310,N_25068,N_28489);
or UO_1311 (O_1311,N_27436,N_29598);
nand UO_1312 (O_1312,N_29468,N_29219);
xor UO_1313 (O_1313,N_26432,N_25184);
nand UO_1314 (O_1314,N_27735,N_24623);
nor UO_1315 (O_1315,N_27745,N_24150);
nor UO_1316 (O_1316,N_29678,N_25179);
or UO_1317 (O_1317,N_27574,N_24738);
nor UO_1318 (O_1318,N_24213,N_28757);
or UO_1319 (O_1319,N_25023,N_25717);
and UO_1320 (O_1320,N_26521,N_24836);
and UO_1321 (O_1321,N_27747,N_24993);
and UO_1322 (O_1322,N_29125,N_27500);
and UO_1323 (O_1323,N_25113,N_25640);
xnor UO_1324 (O_1324,N_28680,N_29846);
nor UO_1325 (O_1325,N_25878,N_27028);
and UO_1326 (O_1326,N_28718,N_24629);
nand UO_1327 (O_1327,N_24651,N_26985);
or UO_1328 (O_1328,N_27161,N_28060);
nor UO_1329 (O_1329,N_28078,N_24164);
xnor UO_1330 (O_1330,N_28122,N_25344);
nand UO_1331 (O_1331,N_28957,N_24061);
xor UO_1332 (O_1332,N_25812,N_26783);
nor UO_1333 (O_1333,N_26119,N_24076);
and UO_1334 (O_1334,N_29620,N_28333);
and UO_1335 (O_1335,N_25824,N_24568);
nand UO_1336 (O_1336,N_25430,N_26864);
or UO_1337 (O_1337,N_26361,N_24894);
xor UO_1338 (O_1338,N_25657,N_28417);
and UO_1339 (O_1339,N_29763,N_27443);
nand UO_1340 (O_1340,N_28052,N_24037);
or UO_1341 (O_1341,N_27558,N_25561);
and UO_1342 (O_1342,N_24603,N_29427);
nand UO_1343 (O_1343,N_28482,N_29736);
xor UO_1344 (O_1344,N_26400,N_24449);
nand UO_1345 (O_1345,N_25091,N_27895);
nor UO_1346 (O_1346,N_28462,N_28329);
and UO_1347 (O_1347,N_27800,N_27614);
xor UO_1348 (O_1348,N_24219,N_25229);
or UO_1349 (O_1349,N_28364,N_29194);
and UO_1350 (O_1350,N_28330,N_26215);
and UO_1351 (O_1351,N_26896,N_28050);
nor UO_1352 (O_1352,N_24611,N_29805);
nand UO_1353 (O_1353,N_25076,N_29324);
or UO_1354 (O_1354,N_27309,N_28345);
and UO_1355 (O_1355,N_24746,N_26554);
nand UO_1356 (O_1356,N_26451,N_28570);
nor UO_1357 (O_1357,N_24335,N_27681);
nor UO_1358 (O_1358,N_29884,N_26318);
nand UO_1359 (O_1359,N_29897,N_25675);
nand UO_1360 (O_1360,N_28121,N_28503);
nand UO_1361 (O_1361,N_25587,N_26590);
nand UO_1362 (O_1362,N_25761,N_26027);
nor UO_1363 (O_1363,N_28391,N_27343);
xor UO_1364 (O_1364,N_24774,N_25738);
xnor UO_1365 (O_1365,N_24024,N_25079);
and UO_1366 (O_1366,N_26308,N_26243);
nand UO_1367 (O_1367,N_28394,N_24572);
and UO_1368 (O_1368,N_28361,N_29151);
nor UO_1369 (O_1369,N_28572,N_27167);
and UO_1370 (O_1370,N_29625,N_25234);
nor UO_1371 (O_1371,N_26250,N_25124);
or UO_1372 (O_1372,N_25104,N_25158);
or UO_1373 (O_1373,N_29137,N_29168);
xor UO_1374 (O_1374,N_25039,N_26477);
and UO_1375 (O_1375,N_29679,N_28332);
nor UO_1376 (O_1376,N_29453,N_28269);
xor UO_1377 (O_1377,N_28403,N_26223);
nand UO_1378 (O_1378,N_28582,N_24139);
xnor UO_1379 (O_1379,N_25666,N_25067);
nand UO_1380 (O_1380,N_25146,N_25578);
and UO_1381 (O_1381,N_26732,N_24617);
nand UO_1382 (O_1382,N_25266,N_27137);
xor UO_1383 (O_1383,N_27504,N_28270);
nand UO_1384 (O_1384,N_25273,N_27898);
nor UO_1385 (O_1385,N_28464,N_24640);
nand UO_1386 (O_1386,N_27590,N_26946);
and UO_1387 (O_1387,N_28574,N_28892);
or UO_1388 (O_1388,N_28197,N_26541);
xor UO_1389 (O_1389,N_27287,N_25452);
xor UO_1390 (O_1390,N_28102,N_28117);
and UO_1391 (O_1391,N_27186,N_24940);
nor UO_1392 (O_1392,N_25985,N_24082);
nor UO_1393 (O_1393,N_29749,N_29512);
and UO_1394 (O_1394,N_27857,N_26078);
nor UO_1395 (O_1395,N_28198,N_28513);
xor UO_1396 (O_1396,N_27933,N_27700);
xor UO_1397 (O_1397,N_29781,N_25157);
or UO_1398 (O_1398,N_25272,N_29488);
or UO_1399 (O_1399,N_26256,N_26273);
nor UO_1400 (O_1400,N_25791,N_28453);
xor UO_1401 (O_1401,N_24880,N_25439);
and UO_1402 (O_1402,N_28542,N_27392);
or UO_1403 (O_1403,N_29302,N_24442);
xnor UO_1404 (O_1404,N_26797,N_29791);
or UO_1405 (O_1405,N_27538,N_26490);
and UO_1406 (O_1406,N_24326,N_24878);
or UO_1407 (O_1407,N_25035,N_28520);
and UO_1408 (O_1408,N_25016,N_27182);
xnor UO_1409 (O_1409,N_29464,N_29754);
nor UO_1410 (O_1410,N_29577,N_25618);
xor UO_1411 (O_1411,N_28676,N_28830);
or UO_1412 (O_1412,N_25488,N_26422);
nand UO_1413 (O_1413,N_27667,N_28014);
or UO_1414 (O_1414,N_26312,N_27996);
nand UO_1415 (O_1415,N_25327,N_27866);
nand UO_1416 (O_1416,N_28750,N_26683);
nor UO_1417 (O_1417,N_27418,N_24997);
and UO_1418 (O_1418,N_24871,N_27054);
xnor UO_1419 (O_1419,N_27471,N_25214);
nor UO_1420 (O_1420,N_25319,N_28741);
nand UO_1421 (O_1421,N_27131,N_28767);
or UO_1422 (O_1422,N_24443,N_26702);
xor UO_1423 (O_1423,N_29558,N_26012);
xnor UO_1424 (O_1424,N_25293,N_28377);
and UO_1425 (O_1425,N_24467,N_26390);
or UO_1426 (O_1426,N_29059,N_27765);
nor UO_1427 (O_1427,N_25811,N_27481);
xor UO_1428 (O_1428,N_29269,N_28871);
nor UO_1429 (O_1429,N_25286,N_26467);
or UO_1430 (O_1430,N_29920,N_25022);
nand UO_1431 (O_1431,N_28877,N_26630);
nand UO_1432 (O_1432,N_28763,N_25882);
and UO_1433 (O_1433,N_25342,N_25171);
and UO_1434 (O_1434,N_29021,N_27145);
and UO_1435 (O_1435,N_27042,N_25663);
and UO_1436 (O_1436,N_24352,N_29123);
nand UO_1437 (O_1437,N_29511,N_25328);
or UO_1438 (O_1438,N_29618,N_28960);
or UO_1439 (O_1439,N_28607,N_27760);
nor UO_1440 (O_1440,N_24728,N_27548);
nand UO_1441 (O_1441,N_26714,N_27715);
or UO_1442 (O_1442,N_25292,N_27189);
and UO_1443 (O_1443,N_27784,N_26249);
or UO_1444 (O_1444,N_27756,N_29292);
xnor UO_1445 (O_1445,N_26230,N_24464);
xor UO_1446 (O_1446,N_29240,N_24388);
or UO_1447 (O_1447,N_26391,N_25843);
nand UO_1448 (O_1448,N_26329,N_26610);
nor UO_1449 (O_1449,N_24111,N_25551);
xor UO_1450 (O_1450,N_24386,N_27013);
xnor UO_1451 (O_1451,N_25556,N_25588);
nor UO_1452 (O_1452,N_28743,N_25467);
or UO_1453 (O_1453,N_27644,N_27278);
nand UO_1454 (O_1454,N_28319,N_29181);
xor UO_1455 (O_1455,N_24707,N_24397);
xnor UO_1456 (O_1456,N_26430,N_24273);
or UO_1457 (O_1457,N_25395,N_25435);
or UO_1458 (O_1458,N_24197,N_25120);
and UO_1459 (O_1459,N_28856,N_26195);
nor UO_1460 (O_1460,N_27565,N_27302);
or UO_1461 (O_1461,N_24648,N_26583);
or UO_1462 (O_1462,N_29265,N_28355);
xnor UO_1463 (O_1463,N_28638,N_25612);
nand UO_1464 (O_1464,N_28992,N_29028);
or UO_1465 (O_1465,N_26692,N_29509);
nand UO_1466 (O_1466,N_25650,N_28833);
or UO_1467 (O_1467,N_29813,N_29171);
and UO_1468 (O_1468,N_28008,N_29702);
nor UO_1469 (O_1469,N_28352,N_24605);
nor UO_1470 (O_1470,N_26966,N_27026);
nand UO_1471 (O_1471,N_29655,N_26140);
nor UO_1472 (O_1472,N_24469,N_29192);
and UO_1473 (O_1473,N_29195,N_26987);
nor UO_1474 (O_1474,N_24124,N_29076);
or UO_1475 (O_1475,N_28434,N_24688);
nand UO_1476 (O_1476,N_28873,N_25110);
xor UO_1477 (O_1477,N_29858,N_28092);
xor UO_1478 (O_1478,N_25364,N_29881);
xor UO_1479 (O_1479,N_27518,N_27704);
nand UO_1480 (O_1480,N_27001,N_29056);
nand UO_1481 (O_1481,N_24114,N_24398);
xor UO_1482 (O_1482,N_27727,N_29317);
nand UO_1483 (O_1483,N_25285,N_24586);
or UO_1484 (O_1484,N_26654,N_26486);
nand UO_1485 (O_1485,N_24298,N_26051);
nor UO_1486 (O_1486,N_29159,N_27398);
xor UO_1487 (O_1487,N_28104,N_28095);
xnor UO_1488 (O_1488,N_28828,N_24796);
xor UO_1489 (O_1489,N_24299,N_24347);
nor UO_1490 (O_1490,N_24673,N_28843);
xor UO_1491 (O_1491,N_27458,N_26653);
or UO_1492 (O_1492,N_24420,N_25712);
and UO_1493 (O_1493,N_29282,N_28790);
xnor UO_1494 (O_1494,N_28642,N_24196);
and UO_1495 (O_1495,N_28510,N_26815);
or UO_1496 (O_1496,N_27311,N_26907);
xnor UO_1497 (O_1497,N_27803,N_24807);
and UO_1498 (O_1498,N_25652,N_24972);
nand UO_1499 (O_1499,N_24445,N_26150);
and UO_1500 (O_1500,N_25397,N_26705);
nor UO_1501 (O_1501,N_28893,N_29607);
nand UO_1502 (O_1502,N_24279,N_25644);
and UO_1503 (O_1503,N_29484,N_28933);
nand UO_1504 (O_1504,N_28287,N_25756);
and UO_1505 (O_1505,N_26065,N_24969);
nor UO_1506 (O_1506,N_24010,N_24337);
or UO_1507 (O_1507,N_26700,N_25771);
nand UO_1508 (O_1508,N_28565,N_29381);
xnor UO_1509 (O_1509,N_25498,N_24641);
xnor UO_1510 (O_1510,N_24947,N_26404);
nand UO_1511 (O_1511,N_29285,N_27656);
nor UO_1512 (O_1512,N_24697,N_26793);
nand UO_1513 (O_1513,N_27736,N_27047);
xnor UO_1514 (O_1514,N_29036,N_26003);
nor UO_1515 (O_1515,N_27751,N_25337);
or UO_1516 (O_1516,N_24233,N_27041);
and UO_1517 (O_1517,N_29652,N_28242);
nand UO_1518 (O_1518,N_28687,N_26253);
xnor UO_1519 (O_1519,N_27879,N_24812);
and UO_1520 (O_1520,N_24296,N_27154);
and UO_1521 (O_1521,N_28859,N_24608);
and UO_1522 (O_1522,N_25724,N_27859);
and UO_1523 (O_1523,N_29812,N_24936);
nor UO_1524 (O_1524,N_25747,N_26839);
and UO_1525 (O_1525,N_24853,N_29989);
and UO_1526 (O_1526,N_25926,N_26232);
and UO_1527 (O_1527,N_29802,N_29976);
and UO_1528 (O_1528,N_27329,N_29727);
and UO_1529 (O_1529,N_26926,N_29845);
nand UO_1530 (O_1530,N_26749,N_24599);
nor UO_1531 (O_1531,N_27345,N_28059);
nor UO_1532 (O_1532,N_28108,N_28742);
xor UO_1533 (O_1533,N_24090,N_28114);
and UO_1534 (O_1534,N_29726,N_24100);
nand UO_1535 (O_1535,N_25635,N_25359);
nor UO_1536 (O_1536,N_28880,N_25231);
nor UO_1537 (O_1537,N_27139,N_24127);
nor UO_1538 (O_1538,N_29002,N_27336);
xnor UO_1539 (O_1539,N_25698,N_27121);
and UO_1540 (O_1540,N_28787,N_28555);
xor UO_1541 (O_1541,N_27936,N_24839);
xor UO_1542 (O_1542,N_27148,N_24436);
nand UO_1543 (O_1543,N_26598,N_24847);
nand UO_1544 (O_1544,N_24811,N_25294);
nor UO_1545 (O_1545,N_24575,N_26115);
nor UO_1546 (O_1546,N_24803,N_27153);
or UO_1547 (O_1547,N_24072,N_25769);
nor UO_1548 (O_1548,N_28910,N_25221);
nand UO_1549 (O_1549,N_28943,N_25673);
or UO_1550 (O_1550,N_24301,N_28512);
and UO_1551 (O_1551,N_27828,N_25046);
xor UO_1552 (O_1552,N_26747,N_24330);
xnor UO_1553 (O_1553,N_24487,N_26026);
or UO_1554 (O_1554,N_27217,N_25174);
or UO_1555 (O_1555,N_28882,N_25857);
or UO_1556 (O_1556,N_28022,N_24146);
nand UO_1557 (O_1557,N_24683,N_26153);
nor UO_1558 (O_1558,N_24783,N_28682);
or UO_1559 (O_1559,N_27181,N_28948);
nand UO_1560 (O_1560,N_29766,N_26565);
xor UO_1561 (O_1561,N_27231,N_27761);
and UO_1562 (O_1562,N_29305,N_24269);
or UO_1563 (O_1563,N_25142,N_25116);
nand UO_1564 (O_1564,N_28328,N_27599);
xor UO_1565 (O_1565,N_28556,N_26319);
nor UO_1566 (O_1566,N_27822,N_27741);
or UO_1567 (O_1567,N_28994,N_28438);
xnor UO_1568 (O_1568,N_25941,N_26660);
nor UO_1569 (O_1569,N_27766,N_26450);
nor UO_1570 (O_1570,N_29994,N_28040);
xnor UO_1571 (O_1571,N_26006,N_26908);
xor UO_1572 (O_1572,N_29630,N_24864);
nor UO_1573 (O_1573,N_26614,N_25312);
xor UO_1574 (O_1574,N_29880,N_25865);
xnor UO_1575 (O_1575,N_27643,N_28187);
and UO_1576 (O_1576,N_29921,N_29486);
nand UO_1577 (O_1577,N_24869,N_27811);
nor UO_1578 (O_1578,N_28929,N_27174);
or UO_1579 (O_1579,N_27871,N_25367);
nand UO_1580 (O_1580,N_29217,N_24385);
xnor UO_1581 (O_1581,N_24103,N_25872);
nand UO_1582 (O_1582,N_27467,N_26948);
nand UO_1583 (O_1583,N_29662,N_24172);
xor UO_1584 (O_1584,N_28138,N_24126);
or UO_1585 (O_1585,N_28261,N_29834);
nor UO_1586 (O_1586,N_29895,N_25297);
nand UO_1587 (O_1587,N_29584,N_27849);
or UO_1588 (O_1588,N_27894,N_27844);
nand UO_1589 (O_1589,N_26557,N_29634);
nand UO_1590 (O_1590,N_27300,N_25115);
nor UO_1591 (O_1591,N_28055,N_26299);
xnor UO_1592 (O_1592,N_29712,N_25274);
xor UO_1593 (O_1593,N_28545,N_26368);
nand UO_1594 (O_1594,N_24200,N_28534);
xnor UO_1595 (O_1595,N_24806,N_28425);
xor UO_1596 (O_1596,N_29327,N_26082);
nand UO_1597 (O_1597,N_29188,N_28338);
nor UO_1598 (O_1598,N_27256,N_27271);
and UO_1599 (O_1599,N_25867,N_29227);
or UO_1600 (O_1600,N_27591,N_29370);
nand UO_1601 (O_1601,N_27799,N_28979);
or UO_1602 (O_1602,N_29428,N_28385);
nor UO_1603 (O_1603,N_29091,N_26038);
nand UO_1604 (O_1604,N_28888,N_24232);
nor UO_1605 (O_1605,N_26214,N_28485);
nor UO_1606 (O_1606,N_26355,N_28540);
xnor UO_1607 (O_1607,N_26424,N_28804);
and UO_1608 (O_1608,N_29605,N_29011);
and UO_1609 (O_1609,N_29722,N_29548);
or UO_1610 (O_1610,N_26515,N_27964);
and UO_1611 (O_1611,N_27587,N_29135);
nand UO_1612 (O_1612,N_28945,N_27588);
nor UO_1613 (O_1613,N_25671,N_27515);
xor UO_1614 (O_1614,N_26148,N_26255);
xor UO_1615 (O_1615,N_29658,N_27375);
xnor UO_1616 (O_1616,N_28214,N_26559);
nand UO_1617 (O_1617,N_24920,N_27959);
nor UO_1618 (O_1618,N_27935,N_24244);
or UO_1619 (O_1619,N_28220,N_28137);
or UO_1620 (O_1620,N_25946,N_29032);
or UO_1621 (O_1621,N_28525,N_26286);
or UO_1622 (O_1622,N_28347,N_27725);
and UO_1623 (O_1623,N_25354,N_25601);
or UO_1624 (O_1624,N_24402,N_29911);
nor UO_1625 (O_1625,N_26181,N_27389);
nor UO_1626 (O_1626,N_28374,N_24740);
or UO_1627 (O_1627,N_25553,N_29340);
nor UO_1628 (O_1628,N_27714,N_24978);
nor UO_1629 (O_1629,N_27002,N_29441);
nand UO_1630 (O_1630,N_28553,N_25884);
or UO_1631 (O_1631,N_26840,N_29134);
or UO_1632 (O_1632,N_27743,N_28675);
or UO_1633 (O_1633,N_24470,N_24679);
nand UO_1634 (O_1634,N_25734,N_28812);
xnor UO_1635 (O_1635,N_29575,N_29863);
or UO_1636 (O_1636,N_29563,N_25877);
xor UO_1637 (O_1637,N_29604,N_29291);
nand UO_1638 (O_1638,N_28940,N_27767);
nand UO_1639 (O_1639,N_28488,N_24628);
xor UO_1640 (O_1640,N_28119,N_24264);
xor UO_1641 (O_1641,N_24881,N_24917);
or UO_1642 (O_1642,N_26944,N_26599);
and UO_1643 (O_1643,N_24480,N_24183);
nand UO_1644 (O_1644,N_27075,N_28083);
nand UO_1645 (O_1645,N_26624,N_28685);
xor UO_1646 (O_1646,N_29697,N_26364);
xnor UO_1647 (O_1647,N_26953,N_24048);
or UO_1648 (O_1648,N_29806,N_25379);
nor UO_1649 (O_1649,N_24271,N_27633);
or UO_1650 (O_1650,N_28853,N_27488);
nand UO_1651 (O_1651,N_28164,N_24676);
or UO_1652 (O_1652,N_24634,N_27567);
nor UO_1653 (O_1653,N_26514,N_27646);
nor UO_1654 (O_1654,N_29031,N_29008);
xor UO_1655 (O_1655,N_24350,N_26950);
xor UO_1656 (O_1656,N_24849,N_24512);
nand UO_1657 (O_1657,N_27623,N_26317);
nand UO_1658 (O_1658,N_25518,N_26059);
or UO_1659 (O_1659,N_28251,N_29423);
and UO_1660 (O_1660,N_28460,N_25913);
nand UO_1661 (O_1661,N_24601,N_25094);
xor UO_1662 (O_1662,N_26204,N_29947);
nand UO_1663 (O_1663,N_26834,N_25189);
nor UO_1664 (O_1664,N_26487,N_28897);
xor UO_1665 (O_1665,N_27067,N_24415);
or UO_1666 (O_1666,N_29469,N_28647);
and UO_1667 (O_1667,N_29382,N_29780);
nand UO_1668 (O_1668,N_24800,N_27971);
nand UO_1669 (O_1669,N_25325,N_27778);
and UO_1670 (O_1670,N_28734,N_26669);
nor UO_1671 (O_1671,N_24992,N_27597);
xnor UO_1672 (O_1672,N_24595,N_25887);
nor UO_1673 (O_1673,N_29823,N_29667);
xnor UO_1674 (O_1674,N_27886,N_26384);
nor UO_1675 (O_1675,N_26118,N_25323);
and UO_1676 (O_1676,N_25333,N_28778);
nor UO_1677 (O_1677,N_28323,N_27425);
nor UO_1678 (O_1678,N_26120,N_25429);
xor UO_1679 (O_1679,N_25261,N_24117);
xor UO_1680 (O_1680,N_25886,N_26073);
and UO_1681 (O_1681,N_24453,N_27517);
nor UO_1682 (O_1682,N_27063,N_25594);
xnor UO_1683 (O_1683,N_27318,N_27463);
and UO_1684 (O_1684,N_27539,N_28614);
and UO_1685 (O_1685,N_26196,N_26530);
xnor UO_1686 (O_1686,N_29414,N_26593);
xnor UO_1687 (O_1687,N_27563,N_26191);
nor UO_1688 (O_1688,N_27368,N_29349);
or UO_1689 (O_1689,N_25602,N_25858);
xnor UO_1690 (O_1690,N_27611,N_24053);
and UO_1691 (O_1691,N_27437,N_26090);
xor UO_1692 (O_1692,N_29242,N_28359);
nor UO_1693 (O_1693,N_27350,N_28231);
xor UO_1694 (O_1694,N_28353,N_27975);
nor UO_1695 (O_1695,N_29768,N_27335);
nand UO_1696 (O_1696,N_25953,N_27511);
or UO_1697 (O_1697,N_29145,N_28204);
nand UO_1698 (O_1698,N_27744,N_24948);
and UO_1699 (O_1699,N_27923,N_24995);
or UO_1700 (O_1700,N_29108,N_29004);
and UO_1701 (O_1701,N_28870,N_27814);
or UO_1702 (O_1702,N_28038,N_29499);
nand UO_1703 (O_1703,N_24868,N_27165);
and UO_1704 (O_1704,N_28863,N_29463);
nand UO_1705 (O_1705,N_26964,N_27061);
xor UO_1706 (O_1706,N_24773,N_25137);
and UO_1707 (O_1707,N_26803,N_28362);
or UO_1708 (O_1708,N_27241,N_28491);
nand UO_1709 (O_1709,N_25819,N_29409);
and UO_1710 (O_1710,N_28956,N_26504);
or UO_1711 (O_1711,N_25973,N_25193);
or UO_1712 (O_1712,N_26185,N_28550);
xnor UO_1713 (O_1713,N_26483,N_29320);
or UO_1714 (O_1714,N_29893,N_28160);
and UO_1715 (O_1715,N_24033,N_25003);
xnor UO_1716 (O_1716,N_27185,N_27230);
or UO_1717 (O_1717,N_24046,N_27281);
or UO_1718 (O_1718,N_24429,N_24455);
xor UO_1719 (O_1719,N_25862,N_24025);
nor UO_1720 (O_1720,N_26764,N_29263);
and UO_1721 (O_1721,N_28949,N_26648);
nor UO_1722 (O_1722,N_27169,N_28944);
and UO_1723 (O_1723,N_28205,N_29673);
xor UO_1724 (O_1724,N_29493,N_25894);
or UO_1725 (O_1725,N_27585,N_29196);
nand UO_1726 (O_1726,N_28649,N_24908);
nand UO_1727 (O_1727,N_27820,N_29235);
and UO_1728 (O_1728,N_25532,N_26406);
or UO_1729 (O_1729,N_28669,N_26798);
or UO_1730 (O_1730,N_29245,N_26539);
or UO_1731 (O_1731,N_29497,N_24749);
or UO_1732 (O_1732,N_27112,N_25725);
nand UO_1733 (O_1733,N_24984,N_25943);
or UO_1734 (O_1734,N_26347,N_28752);
and UO_1735 (O_1735,N_28293,N_28568);
or UO_1736 (O_1736,N_25562,N_28839);
or UO_1737 (O_1737,N_27052,N_29840);
nor UO_1738 (O_1738,N_27099,N_24922);
nor UO_1739 (O_1739,N_28498,N_24171);
nor UO_1740 (O_1740,N_28866,N_24317);
nor UO_1741 (O_1741,N_25347,N_26942);
xor UO_1742 (O_1742,N_27865,N_26855);
xnor UO_1743 (O_1743,N_24270,N_27323);
nand UO_1744 (O_1744,N_24658,N_28959);
xor UO_1745 (O_1745,N_27808,N_29338);
or UO_1746 (O_1746,N_29973,N_26054);
and UO_1747 (O_1747,N_25789,N_25027);
xor UO_1748 (O_1748,N_27571,N_24523);
xnor UO_1749 (O_1749,N_29374,N_25263);
nor UO_1750 (O_1750,N_29425,N_25569);
or UO_1751 (O_1751,N_25208,N_25762);
or UO_1752 (O_1752,N_27976,N_26335);
nor UO_1753 (O_1753,N_25927,N_27296);
or UO_1754 (O_1754,N_26343,N_28619);
nand UO_1755 (O_1755,N_24741,N_28471);
xor UO_1756 (O_1756,N_25611,N_29867);
and UO_1757 (O_1757,N_29841,N_27851);
nand UO_1758 (O_1758,N_28988,N_24234);
nand UO_1759 (O_1759,N_26708,N_24377);
and UO_1760 (O_1760,N_24038,N_24867);
nand UO_1761 (O_1761,N_27837,N_29477);
and UO_1762 (O_1762,N_24327,N_25637);
nor UO_1763 (O_1763,N_26633,N_24341);
nand UO_1764 (O_1764,N_29073,N_24173);
xnor UO_1765 (O_1765,N_27639,N_28191);
or UO_1766 (O_1766,N_25240,N_27514);
nand UO_1767 (O_1767,N_24852,N_28371);
xor UO_1768 (O_1768,N_24909,N_24238);
or UO_1769 (O_1769,N_26502,N_24359);
xnor UO_1770 (O_1770,N_24633,N_27956);
nor UO_1771 (O_1771,N_27995,N_25178);
nor UO_1772 (O_1772,N_24589,N_28266);
nor UO_1773 (O_1773,N_28213,N_25489);
nor UO_1774 (O_1774,N_25574,N_25275);
nand UO_1775 (O_1775,N_29060,N_27498);
nand UO_1776 (O_1776,N_29600,N_26298);
nand UO_1777 (O_1777,N_28125,N_24360);
and UO_1778 (O_1778,N_26879,N_24254);
nand UO_1779 (O_1779,N_27068,N_24874);
and UO_1780 (O_1780,N_27650,N_24276);
and UO_1781 (O_1781,N_24962,N_27928);
nand UO_1782 (O_1782,N_26718,N_28921);
xor UO_1783 (O_1783,N_24314,N_25412);
or UO_1784 (O_1784,N_25767,N_27717);
nor UO_1785 (O_1785,N_26830,N_27774);
nor UO_1786 (O_1786,N_25230,N_29756);
and UO_1787 (O_1787,N_29641,N_29214);
nand UO_1788 (O_1788,N_28532,N_28842);
nor UO_1789 (O_1789,N_27999,N_29220);
and UO_1790 (O_1790,N_24888,N_28915);
and UO_1791 (O_1791,N_24999,N_27942);
or UO_1792 (O_1792,N_24840,N_25154);
or UO_1793 (O_1793,N_24672,N_26345);
nand UO_1794 (O_1794,N_29362,N_27173);
and UO_1795 (O_1795,N_25627,N_28428);
nand UO_1796 (O_1796,N_26396,N_27697);
nand UO_1797 (O_1797,N_27043,N_27461);
nand UO_1798 (O_1798,N_29946,N_29401);
nor UO_1799 (O_1799,N_27805,N_24116);
or UO_1800 (O_1800,N_26053,N_24708);
nor UO_1801 (O_1801,N_28848,N_26264);
nor UO_1802 (O_1802,N_26121,N_24926);
nor UO_1803 (O_1803,N_27780,N_29581);
nor UO_1804 (O_1804,N_24680,N_26652);
or UO_1805 (O_1805,N_26104,N_29066);
nor UO_1806 (O_1806,N_26288,N_27235);
nand UO_1807 (O_1807,N_25944,N_28245);
and UO_1808 (O_1808,N_29473,N_24841);
and UO_1809 (O_1809,N_25568,N_27044);
xnor UO_1810 (O_1810,N_24068,N_24240);
nor UO_1811 (O_1811,N_25988,N_24516);
nand UO_1812 (O_1812,N_24819,N_26592);
or UO_1813 (O_1813,N_25803,N_25131);
nor UO_1814 (O_1814,N_24278,N_28967);
or UO_1815 (O_1815,N_25998,N_29685);
and UO_1816 (O_1816,N_29316,N_26161);
nor UO_1817 (O_1817,N_27364,N_29202);
nand UO_1818 (O_1818,N_24079,N_28013);
nand UO_1819 (O_1819,N_25739,N_28090);
and UO_1820 (O_1820,N_28236,N_27445);
xor UO_1821 (O_1821,N_27370,N_26332);
nor UO_1822 (O_1822,N_24255,N_26016);
or UO_1823 (O_1823,N_25040,N_25550);
nor UO_1824 (O_1824,N_26325,N_25806);
nand UO_1825 (O_1825,N_28925,N_29329);
nor UO_1826 (O_1826,N_26491,N_29268);
and UO_1827 (O_1827,N_27543,N_24517);
xor UO_1828 (O_1828,N_25173,N_26348);
or UO_1829 (O_1829,N_29322,N_26901);
and UO_1830 (O_1830,N_26802,N_26940);
or UO_1831 (O_1831,N_26498,N_25009);
xor UO_1832 (O_1832,N_25425,N_24865);
nor UO_1833 (O_1833,N_28644,N_29218);
and UO_1834 (O_1834,N_24316,N_27000);
or UO_1835 (O_1835,N_25891,N_27777);
or UO_1836 (O_1836,N_24199,N_24225);
nand UO_1837 (O_1837,N_29392,N_27285);
and UO_1838 (O_1838,N_26137,N_29700);
nand UO_1839 (O_1839,N_29939,N_25649);
nand UO_1840 (O_1840,N_26796,N_27577);
nand UO_1841 (O_1841,N_24885,N_26784);
nand UO_1842 (O_1842,N_25202,N_24328);
nor UO_1843 (O_1843,N_25304,N_27798);
xnor UO_1844 (O_1844,N_25220,N_29000);
nor UO_1845 (O_1845,N_26350,N_26770);
or UO_1846 (O_1846,N_27520,N_24182);
nor UO_1847 (O_1847,N_27022,N_28904);
and UO_1848 (O_1848,N_27670,N_24638);
or UO_1849 (O_1849,N_29430,N_26093);
or UO_1850 (O_1850,N_29583,N_27289);
or UO_1851 (O_1851,N_29106,N_26812);
and UO_1852 (O_1852,N_26941,N_25982);
xor UO_1853 (O_1853,N_27568,N_29244);
xor UO_1854 (O_1854,N_29517,N_24404);
nand UO_1855 (O_1855,N_25837,N_25581);
xnor UO_1856 (O_1856,N_25752,N_27206);
or UO_1857 (O_1857,N_29157,N_27238);
and UO_1858 (O_1858,N_28126,N_29112);
and UO_1859 (O_1859,N_28896,N_28686);
nor UO_1860 (O_1860,N_26628,N_28292);
or UO_1861 (O_1861,N_27779,N_26070);
xor UO_1862 (O_1862,N_28365,N_29348);
xnor UO_1863 (O_1863,N_25295,N_28495);
and UO_1864 (O_1864,N_24855,N_29009);
or UO_1865 (O_1865,N_28012,N_29545);
nor UO_1866 (O_1866,N_26574,N_29621);
nand UO_1867 (O_1867,N_25375,N_25933);
nor UO_1868 (O_1868,N_28819,N_26414);
or UO_1869 (O_1869,N_27065,N_28920);
and UO_1870 (O_1870,N_28185,N_24300);
nor UO_1871 (O_1871,N_29557,N_26955);
or UO_1872 (O_1872,N_25169,N_29875);
nor UO_1873 (O_1873,N_24986,N_28608);
and UO_1874 (O_1874,N_29515,N_26801);
xor UO_1875 (O_1875,N_24632,N_26923);
nand UO_1876 (O_1876,N_28952,N_25450);
or UO_1877 (O_1877,N_28115,N_24002);
or UO_1878 (O_1878,N_27267,N_26190);
and UO_1879 (O_1879,N_24011,N_27692);
and UO_1880 (O_1880,N_28692,N_26561);
nand UO_1881 (O_1881,N_25970,N_26257);
xor UO_1882 (O_1882,N_24074,N_28101);
nand UO_1883 (O_1883,N_29719,N_26739);
nor UO_1884 (O_1884,N_26712,N_25793);
xor UO_1885 (O_1885,N_26664,N_27506);
or UO_1886 (O_1886,N_24346,N_25687);
xor UO_1887 (O_1887,N_28111,N_27706);
nand UO_1888 (O_1888,N_24466,N_25959);
and UO_1889 (O_1889,N_29130,N_25419);
nand UO_1890 (O_1890,N_28109,N_27034);
xor UO_1891 (O_1891,N_27076,N_24188);
xnor UO_1892 (O_1892,N_28415,N_28602);
nand UO_1893 (O_1893,N_24035,N_24151);
nand UO_1894 (O_1894,N_27954,N_27025);
and UO_1895 (O_1895,N_26022,N_26351);
xnor UO_1896 (O_1896,N_26248,N_29721);
nand UO_1897 (O_1897,N_28249,N_25975);
or UO_1898 (O_1898,N_25962,N_24771);
or UO_1899 (O_1899,N_24258,N_28074);
or UO_1900 (O_1900,N_27270,N_27991);
xor UO_1901 (O_1901,N_25994,N_29225);
nand UO_1902 (O_1902,N_24122,N_25298);
and UO_1903 (O_1903,N_24988,N_25360);
and UO_1904 (O_1904,N_26968,N_26269);
nand UO_1905 (O_1905,N_29315,N_27754);
nand UO_1906 (O_1906,N_24221,N_24573);
nor UO_1907 (O_1907,N_25096,N_24891);
xor UO_1908 (O_1908,N_28401,N_25949);
nor UO_1909 (O_1909,N_29816,N_29460);
and UO_1910 (O_1910,N_27686,N_29644);
xnor UO_1911 (O_1911,N_25400,N_26787);
nor UO_1912 (O_1912,N_24698,N_25798);
or UO_1913 (O_1913,N_28699,N_26921);
nor UO_1914 (O_1914,N_26588,N_24163);
and UO_1915 (O_1915,N_27363,N_24399);
xor UO_1916 (O_1916,N_27531,N_26667);
and UO_1917 (O_1917,N_29081,N_28701);
and UO_1918 (O_1918,N_27682,N_24577);
xnor UO_1919 (O_1919,N_27833,N_28585);
nor UO_1920 (O_1920,N_27852,N_24403);
and UO_1921 (O_1921,N_24162,N_24045);
xor UO_1922 (O_1922,N_27033,N_24546);
nor UO_1923 (O_1923,N_28128,N_24132);
or UO_1924 (O_1924,N_27632,N_29318);
xnor UO_1925 (O_1925,N_29243,N_28123);
nand UO_1926 (O_1926,N_28000,N_28643);
and UO_1927 (O_1927,N_24649,N_28712);
nor UO_1928 (O_1928,N_24503,N_24532);
or UO_1929 (O_1929,N_29443,N_28180);
nand UO_1930 (O_1930,N_29395,N_29825);
xor UO_1931 (O_1931,N_25222,N_28659);
or UO_1932 (O_1932,N_26971,N_29472);
nor UO_1933 (O_1933,N_29801,N_26520);
and UO_1934 (O_1934,N_26763,N_28296);
nand UO_1935 (O_1935,N_28226,N_25963);
and UO_1936 (O_1936,N_26303,N_25694);
and UO_1937 (O_1937,N_24454,N_27087);
nor UO_1938 (O_1938,N_25718,N_27101);
nor UO_1939 (O_1939,N_29755,N_25114);
xor UO_1940 (O_1940,N_28857,N_25254);
or UO_1941 (O_1941,N_26997,N_28490);
xor UO_1942 (O_1942,N_24371,N_27763);
and UO_1943 (O_1943,N_26021,N_27965);
nand UO_1944 (O_1944,N_26387,N_27412);
and UO_1945 (O_1945,N_24070,N_27796);
xnor UO_1946 (O_1946,N_28693,N_26033);
xor UO_1947 (O_1947,N_29590,N_24704);
xor UO_1948 (O_1948,N_25991,N_27594);
nor UO_1949 (O_1949,N_25826,N_26376);
and UO_1950 (O_1950,N_25617,N_25797);
or UO_1951 (O_1951,N_25662,N_24579);
nand UO_1952 (O_1952,N_25257,N_29795);
or UO_1953 (O_1953,N_25626,N_27603);
and UO_1954 (O_1954,N_25181,N_25004);
and UO_1955 (O_1955,N_29733,N_27155);
nand UO_1956 (O_1956,N_25159,N_25366);
nand UO_1957 (O_1957,N_27551,N_25535);
or UO_1958 (O_1958,N_29502,N_27496);
and UO_1959 (O_1959,N_27453,N_27509);
nor UO_1960 (O_1960,N_27244,N_25754);
or UO_1961 (O_1961,N_27479,N_27939);
and UO_1962 (O_1962,N_28402,N_29250);
or UO_1963 (O_1963,N_27790,N_28254);
xnor UO_1964 (O_1964,N_29271,N_26205);
and UO_1965 (O_1965,N_24484,N_28596);
nor UO_1966 (O_1966,N_25997,N_26247);
and UO_1967 (O_1967,N_28255,N_26534);
nor UO_1968 (O_1968,N_27158,N_27877);
nor UO_1969 (O_1969,N_29661,N_27310);
and UO_1970 (O_1970,N_28144,N_29498);
and UO_1971 (O_1971,N_26029,N_24187);
xnor UO_1972 (O_1972,N_24040,N_26831);
xnor UO_1973 (O_1973,N_26828,N_24284);
nor UO_1974 (O_1974,N_25653,N_28093);
nor UO_1975 (O_1975,N_29933,N_25960);
and UO_1976 (O_1976,N_29102,N_28326);
xnor UO_1977 (O_1977,N_24372,N_28716);
xor UO_1978 (O_1978,N_24955,N_25380);
xor UO_1979 (O_1979,N_27793,N_26276);
nand UO_1980 (O_1980,N_29272,N_25311);
or UO_1981 (O_1981,N_24817,N_28461);
nor UO_1982 (O_1982,N_25463,N_27322);
xor UO_1983 (O_1983,N_29937,N_27485);
nand UO_1984 (O_1984,N_29653,N_29507);
nor UO_1985 (O_1985,N_27693,N_24756);
and UO_1986 (O_1986,N_24862,N_24931);
nand UO_1987 (O_1987,N_29866,N_29228);
or UO_1988 (O_1988,N_25778,N_29714);
and UO_1989 (O_1989,N_29959,N_29793);
nand UO_1990 (O_1990,N_24879,N_25149);
or UO_1991 (O_1991,N_26306,N_28315);
or UO_1992 (O_1992,N_24823,N_29411);
xor UO_1993 (O_1993,N_29904,N_28457);
nor UO_1994 (O_1994,N_26736,N_24409);
and UO_1995 (O_1995,N_29965,N_24681);
nor UO_1996 (O_1996,N_29913,N_26562);
or UO_1997 (O_1997,N_24827,N_26675);
nor UO_1998 (O_1998,N_24642,N_25302);
nand UO_1999 (O_1999,N_24181,N_26821);
xnor UO_2000 (O_2000,N_27713,N_29929);
nand UO_2001 (O_2001,N_28132,N_28629);
and UO_2002 (O_2002,N_24585,N_28667);
or UO_2003 (O_2003,N_24235,N_24656);
and UO_2004 (O_2004,N_25808,N_28097);
nand UO_2005 (O_2005,N_24433,N_27550);
and UO_2006 (O_2006,N_25730,N_25505);
or UO_2007 (O_2007,N_26833,N_28411);
and UO_2008 (O_2008,N_25098,N_24792);
and UO_2009 (O_2009,N_27092,N_28993);
xor UO_2010 (O_2010,N_26826,N_24964);
xor UO_2011 (O_2011,N_29684,N_28232);
or UO_2012 (O_2012,N_25548,N_26596);
xor UO_2013 (O_2013,N_27024,N_27523);
xor UO_2014 (O_2014,N_26290,N_26677);
nor UO_2015 (O_2015,N_28196,N_26333);
and UO_2016 (O_2016,N_29559,N_27507);
nand UO_2017 (O_2017,N_28816,N_24361);
nand UO_2018 (O_2018,N_26327,N_28393);
and UO_2019 (O_2019,N_29447,N_28339);
or UO_2020 (O_2020,N_28397,N_27755);
nand UO_2021 (O_2021,N_26108,N_25567);
or UO_2022 (O_2022,N_28509,N_29113);
xnor UO_2023 (O_2023,N_29725,N_28299);
or UO_2024 (O_2024,N_26281,N_26262);
xor UO_2025 (O_2025,N_24007,N_29146);
and UO_2026 (O_2026,N_29233,N_24722);
nor UO_2027 (O_2027,N_27930,N_24727);
nor UO_2028 (O_2028,N_25279,N_24463);
or UO_2029 (O_2029,N_28048,N_27929);
nor UO_2030 (O_2030,N_25414,N_28824);
nand UO_2031 (O_2031,N_25523,N_29799);
nor UO_2032 (O_2032,N_26891,N_25992);
nand UO_2033 (O_2033,N_25305,N_26201);
nand UO_2034 (O_2034,N_25921,N_27396);
or UO_2035 (O_2035,N_27417,N_25172);
or UO_2036 (O_2036,N_25433,N_25072);
xor UO_2037 (O_2037,N_25455,N_28938);
nor UO_2038 (O_2038,N_29154,N_24581);
xor UO_2039 (O_2039,N_24637,N_28806);
nor UO_2040 (O_2040,N_29901,N_26217);
xor UO_2041 (O_2041,N_27685,N_26558);
xor UO_2042 (O_2042,N_24882,N_28153);
nor UO_2043 (O_2043,N_24205,N_25005);
and UO_2044 (O_2044,N_28179,N_27295);
and UO_2045 (O_2045,N_26443,N_25989);
xor UO_2046 (O_2046,N_28627,N_27228);
and UO_2047 (O_2047,N_27998,N_26741);
xnor UO_2048 (O_2048,N_24362,N_29033);
or UO_2049 (O_2049,N_24930,N_24348);
xor UO_2050 (O_2050,N_28758,N_26198);
nand UO_2051 (O_2051,N_28029,N_25001);
or UO_2052 (O_2052,N_28975,N_27885);
xor UO_2053 (O_2053,N_24147,N_24744);
nor UO_2054 (O_2054,N_28714,N_27753);
and UO_2055 (O_2055,N_26586,N_26485);
nand UO_2056 (O_2056,N_28070,N_28702);
and UO_2057 (O_2057,N_26132,N_28435);
xnor UO_2058 (O_2058,N_24047,N_25136);
and UO_2059 (O_2059,N_25449,N_26352);
or UO_2060 (O_2060,N_29034,N_28899);
or UO_2061 (O_2061,N_27721,N_29249);
nor UO_2062 (O_2062,N_26856,N_29426);
xnor UO_2063 (O_2063,N_26449,N_26506);
and UO_2064 (O_2064,N_26356,N_24543);
nor UO_2065 (O_2065,N_26049,N_25125);
xnor UO_2066 (O_2066,N_28665,N_25909);
xor UO_2067 (O_2067,N_27934,N_26034);
and UO_2068 (O_2068,N_26900,N_28450);
xor UO_2069 (O_2069,N_25825,N_28142);
or UO_2070 (O_2070,N_29730,N_27559);
or UO_2071 (O_2071,N_25251,N_28558);
and UO_2072 (O_2072,N_26428,N_27127);
nor UO_2073 (O_2073,N_26207,N_28539);
or UO_2074 (O_2074,N_27962,N_25961);
or UO_2075 (O_2075,N_24057,N_27512);
and UO_2076 (O_2076,N_26041,N_29319);
nor UO_2077 (O_2077,N_24702,N_29238);
or UO_2078 (O_2078,N_29377,N_27096);
nand UO_2079 (O_2079,N_27615,N_29556);
nor UO_2080 (O_2080,N_28653,N_29723);
xor UO_2081 (O_2081,N_25810,N_29394);
or UO_2082 (O_2082,N_24207,N_27069);
and UO_2083 (O_2083,N_25609,N_26552);
or UO_2084 (O_2084,N_26608,N_27094);
xnor UO_2085 (O_2085,N_28479,N_29337);
nor UO_2086 (O_2086,N_24953,N_27967);
nand UO_2087 (O_2087,N_25226,N_24319);
xor UO_2088 (O_2088,N_26127,N_27176);
or UO_2089 (O_2089,N_24797,N_27536);
nand UO_2090 (O_2090,N_27605,N_24613);
and UO_2091 (O_2091,N_26337,N_24615);
or UO_2092 (O_2092,N_26818,N_28170);
nand UO_2093 (O_2093,N_26055,N_29352);
or UO_2094 (O_2094,N_27566,N_26307);
nand UO_2095 (O_2095,N_29885,N_28278);
nand UO_2096 (O_2096,N_28239,N_28708);
xor UO_2097 (O_2097,N_27070,N_27556);
nand UO_2098 (O_2098,N_24152,N_27613);
nand UO_2099 (O_2099,N_24916,N_29591);
nand UO_2100 (O_2100,N_26182,N_26409);
nand UO_2101 (O_2101,N_28215,N_24652);
xnor UO_2102 (O_2102,N_26330,N_28617);
or UO_2103 (O_2103,N_27505,N_25999);
and UO_2104 (O_2104,N_27205,N_25315);
xor UO_2105 (O_2105,N_24075,N_24668);
nand UO_2106 (O_2106,N_29555,N_26569);
and UO_2107 (O_2107,N_25447,N_25566);
xnor UO_2108 (O_2108,N_25170,N_24858);
or UO_2109 (O_2109,N_28207,N_25513);
and UO_2110 (O_2110,N_27348,N_26674);
nand UO_2111 (O_2111,N_28616,N_26760);
nor UO_2112 (O_2112,N_29364,N_26920);
nand UO_2113 (O_2113,N_25083,N_25403);
nor UO_2114 (O_2114,N_28805,N_25868);
nand UO_2115 (O_2115,N_27699,N_26823);
nor UO_2116 (O_2116,N_28398,N_25155);
nand UO_2117 (O_2117,N_26179,N_28042);
or UO_2118 (O_2118,N_29910,N_29879);
and UO_2119 (O_2119,N_28923,N_28256);
xor UO_2120 (O_2120,N_28753,N_28891);
or UO_2121 (O_2121,N_29586,N_25842);
nor UO_2122 (O_2122,N_27272,N_29449);
nor UO_2123 (O_2123,N_29608,N_25308);
nand UO_2124 (O_2124,N_29365,N_25855);
or UO_2125 (O_2125,N_27888,N_24156);
nor UO_2126 (O_2126,N_28691,N_25773);
nand UO_2127 (O_2127,N_28496,N_27904);
or UO_2128 (O_2128,N_26313,N_27781);
and UO_2129 (O_2129,N_25369,N_29065);
and UO_2130 (O_2130,N_29521,N_28780);
or UO_2131 (O_2131,N_26045,N_24194);
xnor UO_2132 (O_2132,N_26929,N_27102);
and UO_2133 (O_2133,N_27253,N_29504);
or UO_2134 (O_2134,N_27889,N_27593);
nand UO_2135 (O_2135,N_29326,N_25864);
nor UO_2136 (O_2136,N_25038,N_27109);
or UO_2137 (O_2137,N_26581,N_24954);
or UO_2138 (O_2138,N_26278,N_29852);
or UO_2139 (O_2139,N_25571,N_24625);
nor UO_2140 (O_2140,N_26893,N_24814);
xor UO_2141 (O_2141,N_29637,N_27592);
nand UO_2142 (O_2142,N_29610,N_27658);
nor UO_2143 (O_2143,N_28379,N_24166);
nor UO_2144 (O_2144,N_24508,N_26745);
nor UO_2145 (O_2145,N_24907,N_24643);
or UO_2146 (O_2146,N_27470,N_26713);
or UO_2147 (O_2147,N_24578,N_26184);
nor UO_2148 (O_2148,N_26192,N_26069);
or UO_2149 (O_2149,N_26685,N_29765);
nor UO_2150 (O_2150,N_24509,N_26105);
nand UO_2151 (O_2151,N_25696,N_28801);
nor UO_2152 (O_2152,N_27341,N_24716);
or UO_2153 (O_2153,N_26176,N_28288);
nor UO_2154 (O_2154,N_25287,N_25674);
or UO_2155 (O_2155,N_24952,N_25303);
and UO_2156 (O_2156,N_25606,N_26109);
and UO_2157 (O_2157,N_29828,N_25310);
xor UO_2158 (O_2158,N_27083,N_24957);
nor UO_2159 (O_2159,N_28282,N_28947);
nor UO_2160 (O_2160,N_28033,N_26611);
nand UO_2161 (O_2161,N_26663,N_24119);
or UO_2162 (O_2162,N_29104,N_24375);
or UO_2163 (O_2163,N_29717,N_26662);
and UO_2164 (O_2164,N_27662,N_27197);
nand UO_2165 (O_2165,N_24338,N_25446);
nor UO_2166 (O_2166,N_25196,N_25212);
nand UO_2167 (O_2167,N_29857,N_26175);
and UO_2168 (O_2168,N_25745,N_27943);
nor UO_2169 (O_2169,N_24477,N_27710);
nand UO_2170 (O_2170,N_27652,N_29306);
nor UO_2171 (O_2171,N_27032,N_25427);
nor UO_2172 (O_2172,N_28821,N_25729);
or UO_2173 (O_2173,N_25431,N_25283);
and UO_2174 (O_2174,N_26992,N_28066);
or UO_2175 (O_2175,N_26295,N_25827);
nor UO_2176 (O_2176,N_29626,N_25134);
or UO_2177 (O_2177,N_25365,N_26194);
nor UO_2178 (O_2178,N_27027,N_26727);
nand UO_2179 (O_2179,N_24826,N_28384);
xnor UO_2180 (O_2180,N_29580,N_28521);
nor UO_2181 (O_2181,N_28930,N_25559);
and UO_2182 (O_2182,N_29029,N_24373);
nor UO_2183 (O_2183,N_24315,N_24966);
nor UO_2184 (O_2184,N_24185,N_25830);
xnor UO_2185 (O_2185,N_29666,N_27619);
nor UO_2186 (O_2186,N_25776,N_24748);
or UO_2187 (O_2187,N_29402,N_24307);
nand UO_2188 (O_2188,N_26447,N_29601);
and UO_2189 (O_2189,N_28041,N_27306);
nand UO_2190 (O_2190,N_26203,N_25714);
nor UO_2191 (O_2191,N_24475,N_26291);
and UO_2192 (O_2192,N_26091,N_29050);
and UO_2193 (O_2193,N_27097,N_27773);
or UO_2194 (O_2194,N_28601,N_25119);
or UO_2195 (O_2195,N_25370,N_25487);
or UO_2196 (O_2196,N_24135,N_27135);
nand UO_2197 (O_2197,N_27840,N_26371);
nor UO_2198 (O_2198,N_26889,N_27900);
nor UO_2199 (O_2199,N_24490,N_25047);
xor UO_2200 (O_2200,N_25512,N_29964);
nor UO_2201 (O_2201,N_25948,N_28099);
nand UO_2202 (O_2202,N_27171,N_28088);
nor UO_2203 (O_2203,N_27918,N_25393);
nor UO_2204 (O_2204,N_27769,N_29612);
or UO_2205 (O_2205,N_29686,N_24655);
nand UO_2206 (O_2206,N_24115,N_26464);
xor UO_2207 (O_2207,N_28760,N_27906);
and UO_2208 (O_2208,N_25742,N_26806);
xor UO_2209 (O_2209,N_26310,N_27003);
and UO_2210 (O_2210,N_28080,N_28713);
and UO_2211 (O_2211,N_28368,N_25007);
and UO_2212 (O_2212,N_26935,N_25408);
or UO_2213 (O_2213,N_26063,N_29169);
xnor UO_2214 (O_2214,N_24745,N_25954);
and UO_2215 (O_2215,N_25239,N_29925);
and UO_2216 (O_2216,N_26100,N_24659);
nand UO_2217 (O_2217,N_28822,N_25187);
nor UO_2218 (O_2218,N_24481,N_28811);
nor UO_2219 (O_2219,N_24769,N_26225);
xor UO_2220 (O_2220,N_24502,N_27198);
nor UO_2221 (O_2221,N_26735,N_26694);
xor UO_2222 (O_2222,N_29501,N_28681);
and UO_2223 (O_2223,N_29442,N_27048);
nor UO_2224 (O_2224,N_25608,N_28678);
or UO_2225 (O_2225,N_27007,N_28081);
nor UO_2226 (O_2226,N_24759,N_24736);
xor UO_2227 (O_2227,N_27762,N_25735);
nand UO_2228 (O_2228,N_26917,N_27838);
nand UO_2229 (O_2229,N_28238,N_27953);
nor UO_2230 (O_2230,N_27455,N_25848);
nand UO_2231 (O_2231,N_26544,N_29095);
nand UO_2232 (O_2232,N_24387,N_28230);
nor UO_2233 (O_2233,N_28620,N_28872);
xor UO_2234 (O_2234,N_26540,N_25062);
nor UO_2235 (O_2235,N_26495,N_28538);
nand UO_2236 (O_2236,N_24022,N_27679);
or UO_2237 (O_2237,N_27860,N_27100);
nand UO_2238 (O_2238,N_29861,N_25053);
or UO_2239 (O_2239,N_29257,N_25144);
xor UO_2240 (O_2240,N_28914,N_24976);
nand UO_2241 (O_2241,N_24400,N_26266);
nor UO_2242 (O_2242,N_24669,N_28026);
and UO_2243 (O_2243,N_27388,N_27819);
nor UO_2244 (O_2244,N_25271,N_25428);
nand UO_2245 (O_2245,N_24170,N_29330);
and UO_2246 (O_2246,N_26776,N_26898);
and UO_2247 (O_2247,N_28430,N_28536);
and UO_2248 (O_2248,N_27009,N_28706);
nand UO_2249 (O_2249,N_25336,N_29520);
or UO_2250 (O_2250,N_27239,N_26296);
or UO_2251 (O_2251,N_24349,N_25054);
or UO_2252 (O_2252,N_25368,N_29585);
nor UO_2253 (O_2253,N_28120,N_24893);
nor UO_2254 (O_2254,N_29284,N_27739);
and UO_2255 (O_2255,N_26037,N_26625);
or UO_2256 (O_2256,N_29182,N_28815);
nor UO_2257 (O_2257,N_28139,N_24687);
and UO_2258 (O_2258,N_28367,N_26771);
nor UO_2259 (O_2259,N_26679,N_24521);
or UO_2260 (O_2260,N_25237,N_26052);
nor UO_2261 (O_2261,N_24663,N_24846);
or UO_2262 (O_2262,N_24565,N_27037);
xor UO_2263 (O_2263,N_28898,N_24357);
nor UO_2264 (O_2264,N_27468,N_29071);
nand UO_2265 (O_2265,N_27017,N_25782);
nand UO_2266 (O_2266,N_27569,N_29045);
and UO_2267 (O_2267,N_26240,N_29444);
or UO_2268 (O_2268,N_29760,N_28527);
or UO_2269 (O_2269,N_28035,N_28015);
and UO_2270 (O_2270,N_29456,N_24288);
or UO_2271 (O_2271,N_24065,N_26638);
nor UO_2272 (O_2272,N_25225,N_24671);
and UO_2273 (O_2273,N_29462,N_25531);
nor UO_2274 (O_2274,N_28227,N_25965);
or UO_2275 (O_2275,N_29807,N_28773);
or UO_2276 (O_2276,N_26587,N_26577);
nand UO_2277 (O_2277,N_28118,N_24087);
nor UO_2278 (O_2278,N_27941,N_27156);
nor UO_2279 (O_2279,N_28259,N_29026);
nor UO_2280 (O_2280,N_28606,N_29183);
and UO_2281 (O_2281,N_29164,N_24631);
nand UO_2282 (O_2282,N_25924,N_27817);
nor UO_2283 (O_2283,N_24857,N_26149);
nand UO_2284 (O_2284,N_29328,N_27863);
or UO_2285 (O_2285,N_28786,N_24779);
xnor UO_2286 (O_2286,N_26328,N_29779);
xnor UO_2287 (O_2287,N_26681,N_27104);
or UO_2288 (O_2288,N_24569,N_28005);
and UO_2289 (O_2289,N_26888,N_28860);
xor UO_2290 (O_2290,N_29083,N_27095);
nand UO_2291 (O_2291,N_28451,N_29131);
nand UO_2292 (O_2292,N_27204,N_25071);
xor UO_2293 (O_2293,N_29478,N_26661);
nor UO_2294 (O_2294,N_26154,N_29467);
nor UO_2295 (O_2295,N_26251,N_24356);
nand UO_2296 (O_2296,N_27313,N_25508);
nand UO_2297 (O_2297,N_28135,N_28820);
and UO_2298 (O_2298,N_26287,N_29758);
nand UO_2299 (O_2299,N_24212,N_26535);
xor UO_2300 (O_2300,N_29175,N_26887);
or UO_2301 (O_2301,N_25201,N_28668);
or UO_2302 (O_2302,N_24195,N_28087);
nand UO_2303 (O_2303,N_26817,N_27749);
and UO_2304 (O_2304,N_28436,N_27385);
nor UO_2305 (O_2305,N_27960,N_25031);
nor UO_2306 (O_2306,N_25152,N_28809);
nand UO_2307 (O_2307,N_25390,N_26998);
xor UO_2308 (O_2308,N_24842,N_28964);
xnor UO_2309 (O_2309,N_27062,N_27527);
or UO_2310 (O_2310,N_26868,N_29826);
xor UO_2311 (O_2311,N_29332,N_29619);
nor UO_2312 (O_2312,N_27449,N_29675);
or UO_2313 (O_2313,N_24222,N_26331);
nand UO_2314 (O_2314,N_25880,N_25522);
and UO_2315 (O_2315,N_24428,N_24211);
xor UO_2316 (O_2316,N_27978,N_26899);
or UO_2317 (O_2317,N_28517,N_26996);
nor UO_2318 (O_2318,N_28375,N_24766);
nor UO_2319 (O_2319,N_25572,N_27030);
nor UO_2320 (O_2320,N_28475,N_28918);
xnor UO_2321 (O_2321,N_29354,N_26560);
or UO_2322 (O_2322,N_28221,N_27678);
nand UO_2323 (O_2323,N_29932,N_27696);
and UO_2324 (O_2324,N_28194,N_27415);
and UO_2325 (O_2325,N_26241,N_24576);
nor UO_2326 (O_2326,N_26790,N_26673);
or UO_2327 (O_2327,N_28626,N_26227);
nand UO_2328 (O_2328,N_29080,N_28657);
and UO_2329 (O_2329,N_28500,N_24570);
xnor UO_2330 (O_2330,N_27382,N_28939);
nand UO_2331 (O_2331,N_25176,N_29971);
nand UO_2332 (O_2332,N_29967,N_28124);
and UO_2333 (O_2333,N_26924,N_24754);
and UO_2334 (O_2334,N_26976,N_29301);
xor UO_2335 (O_2335,N_28583,N_26226);
xor UO_2336 (O_2336,N_29741,N_24505);
xnor UO_2337 (O_2337,N_29391,N_26113);
nand UO_2338 (O_2338,N_24737,N_29966);
nor UO_2339 (O_2339,N_27917,N_28381);
or UO_2340 (O_2340,N_26918,N_28837);
nor UO_2341 (O_2341,N_26412,N_24093);
nor UO_2342 (O_2342,N_25075,N_27367);
nor UO_2343 (O_2343,N_26168,N_24607);
xnor UO_2344 (O_2344,N_25135,N_24715);
nor UO_2345 (O_2345,N_26522,N_28980);
nand UO_2346 (O_2346,N_26385,N_24193);
or UO_2347 (O_2347,N_25990,N_24426);
or UO_2348 (O_2348,N_25264,N_29923);
and UO_2349 (O_2349,N_24391,N_27191);
or UO_2350 (O_2350,N_28724,N_29565);
and UO_2351 (O_2351,N_27226,N_26107);
xnor UO_2352 (O_2352,N_27580,N_24899);
xor UO_2353 (O_2353,N_29952,N_29489);
nand UO_2354 (O_2354,N_27346,N_28831);
nor UO_2355 (O_2355,N_25896,N_27759);
and UO_2356 (O_2356,N_28404,N_26084);
xor UO_2357 (O_2357,N_29278,N_27086);
and UO_2358 (O_2358,N_24425,N_24118);
xor UO_2359 (O_2359,N_24086,N_29211);
nand UO_2360 (O_2360,N_28152,N_28695);
or UO_2361 (O_2361,N_26186,N_25014);
and UO_2362 (O_2362,N_25628,N_26239);
xnor UO_2363 (O_2363,N_25542,N_28576);
nand UO_2364 (O_2364,N_26124,N_27730);
nor UO_2365 (O_2365,N_28449,N_26622);
xor UO_2366 (O_2366,N_29550,N_24795);
nor UO_2367 (O_2367,N_25182,N_28612);
nor UO_2368 (O_2368,N_26202,N_28172);
xnor UO_2369 (O_2369,N_24405,N_27258);
nor UO_2370 (O_2370,N_25680,N_29481);
nand UO_2371 (O_2371,N_24626,N_29167);
nor UO_2372 (O_2372,N_26394,N_24479);
or UO_2373 (O_2373,N_25289,N_29783);
or UO_2374 (O_2374,N_26564,N_28321);
and UO_2375 (O_2375,N_29496,N_28634);
xor UO_2376 (O_2376,N_25643,N_25779);
or UO_2377 (O_2377,N_28497,N_26135);
xnor UO_2378 (O_2378,N_29350,N_29794);
xnor UO_2379 (O_2379,N_28603,N_26011);
or UO_2380 (O_2380,N_27450,N_25638);
nand UO_2381 (O_2381,N_27250,N_29534);
nor UO_2382 (O_2382,N_26147,N_28590);
nand UO_2383 (O_2383,N_29876,N_29683);
or UO_2384 (O_2384,N_28561,N_27261);
nand UO_2385 (O_2385,N_25892,N_29133);
or UO_2386 (O_2386,N_28202,N_26369);
xnor UO_2387 (O_2387,N_29185,N_28673);
nand UO_2388 (O_2388,N_29665,N_27414);
nand UO_2389 (O_2389,N_27845,N_25394);
xor UO_2390 (O_2390,N_26338,N_26238);
xor UO_2391 (O_2391,N_24376,N_25642);
or UO_2392 (O_2392,N_25668,N_29720);
nor UO_2393 (O_2393,N_24850,N_26696);
nand UO_2394 (O_2394,N_29480,N_28886);
nor UO_2395 (O_2395,N_28998,N_25372);
and UO_2396 (O_2396,N_25928,N_27641);
nand UO_2397 (O_2397,N_26087,N_24209);
xor UO_2398 (O_2398,N_26373,N_25000);
xnor UO_2399 (O_2399,N_27393,N_25021);
nor UO_2400 (O_2400,N_25597,N_28168);
or UO_2401 (O_2401,N_27610,N_26494);
nand UO_2402 (O_2402,N_29991,N_28067);
nand UO_2403 (O_2403,N_25874,N_29948);
or UO_2404 (O_2404,N_29745,N_28690);
nor UO_2405 (O_2405,N_29455,N_27351);
xnor UO_2406 (O_2406,N_28813,N_29908);
or UO_2407 (O_2407,N_25792,N_28987);
and UO_2408 (O_2408,N_28431,N_24169);
xor UO_2409 (O_2409,N_24968,N_26959);
or UO_2410 (O_2410,N_26267,N_25204);
nand UO_2411 (O_2411,N_28963,N_25108);
nor UO_2412 (O_2412,N_27624,N_26211);
nor UO_2413 (O_2413,N_29688,N_27655);
nor UO_2414 (O_2414,N_24555,N_28876);
nand UO_2415 (O_2415,N_25472,N_24500);
nor UO_2416 (O_2416,N_24003,N_26862);
xnor UO_2417 (O_2417,N_24062,N_28670);
xnor UO_2418 (O_2418,N_24089,N_28277);
and UO_2419 (O_2419,N_26894,N_29868);
nor UO_2420 (O_2420,N_26458,N_29523);
or UO_2421 (O_2421,N_25555,N_28184);
or UO_2422 (O_2422,N_26370,N_25689);
or UO_2423 (O_2423,N_26245,N_25883);
xnor UO_2424 (O_2424,N_27478,N_25831);
and UO_2425 (O_2425,N_29017,N_26573);
or UO_2426 (O_2426,N_27106,N_25008);
xor UO_2427 (O_2427,N_24243,N_24552);
xnor UO_2428 (O_2428,N_26096,N_29142);
xnor UO_2429 (O_2429,N_27475,N_27988);
and UO_2430 (O_2430,N_29450,N_29902);
nand UO_2431 (O_2431,N_29525,N_28578);
or UO_2432 (O_2432,N_28409,N_28360);
or UO_2433 (O_2433,N_25034,N_26173);
nand UO_2434 (O_2434,N_26832,N_27410);
xor UO_2435 (O_2435,N_25679,N_28577);
nand UO_2436 (O_2436,N_28079,N_29603);
nor UO_2437 (O_2437,N_29914,N_25619);
nor UO_2438 (O_2438,N_24497,N_25544);
and UO_2439 (O_2439,N_27913,N_29890);
or UO_2440 (O_2440,N_29254,N_24910);
xor UO_2441 (O_2441,N_28325,N_27827);
nand UO_2442 (O_2442,N_28024,N_29351);
xnor UO_2443 (O_2443,N_26939,N_27787);
or UO_2444 (O_2444,N_25086,N_27292);
xnor UO_2445 (O_2445,N_26377,N_24263);
xnor UO_2446 (O_2446,N_26292,N_26415);
or UO_2447 (O_2447,N_28494,N_25165);
and UO_2448 (O_2448,N_25589,N_25560);
xor UO_2449 (O_2449,N_25206,N_24178);
xnor UO_2450 (O_2450,N_24714,N_26822);
nand UO_2451 (O_2451,N_26272,N_29072);
nand UO_2452 (O_2452,N_29886,N_26737);
nand UO_2453 (O_2453,N_29461,N_25716);
nor UO_2454 (O_2454,N_27669,N_27373);
xor UO_2455 (O_2455,N_28746,N_25050);
or UO_2456 (O_2456,N_25186,N_27703);
xor UO_2457 (O_2457,N_25406,N_25211);
and UO_2458 (O_2458,N_29752,N_27447);
nand UO_2459 (O_2459,N_29843,N_27535);
or UO_2460 (O_2460,N_24246,N_24026);
xor UO_2461 (O_2461,N_26603,N_24900);
xor UO_2462 (O_2462,N_28955,N_24828);
xor UO_2463 (O_2463,N_26274,N_26759);
nor UO_2464 (O_2464,N_29963,N_24958);
nor UO_2465 (O_2465,N_29147,N_25032);
or UO_2466 (O_2466,N_27021,N_26358);
xor UO_2467 (O_2467,N_27812,N_29064);
or UO_2468 (O_2468,N_25746,N_29786);
xnor UO_2469 (O_2469,N_29922,N_24408);
or UO_2470 (O_2470,N_29924,N_25402);
nand UO_2471 (O_2471,N_29270,N_26493);
nand UO_2472 (O_2472,N_24520,N_24506);
xor UO_2473 (O_2473,N_24067,N_25424);
xor UO_2474 (O_2474,N_25966,N_26538);
and UO_2475 (O_2475,N_29668,N_26621);
nand UO_2476 (O_2476,N_25349,N_28794);
nor UO_2477 (O_2477,N_27785,N_24967);
or UO_2478 (O_2478,N_27899,N_27826);
nand UO_2479 (O_2479,N_24584,N_27428);
or UO_2480 (O_2480,N_26905,N_28548);
or UO_2481 (O_2481,N_29431,N_28798);
and UO_2482 (O_2482,N_25646,N_24324);
or UO_2483 (O_2483,N_28961,N_27240);
xor UO_2484 (O_2484,N_29735,N_26183);
or UO_2485 (O_2485,N_24562,N_29830);
nor UO_2486 (O_2486,N_29163,N_28320);
nor UO_2487 (O_2487,N_27990,N_29986);
or UO_2488 (O_2488,N_28441,N_26326);
xor UO_2489 (O_2489,N_24982,N_27729);
nor UO_2490 (O_2490,N_28072,N_28989);
nand UO_2491 (O_2491,N_24583,N_27229);
nand UO_2492 (O_2492,N_25130,N_29713);
and UO_2493 (O_2493,N_26399,N_27521);
nor UO_2494 (O_2494,N_28836,N_29433);
nor UO_2495 (O_2495,N_27308,N_29535);
and UO_2496 (O_2496,N_27855,N_25270);
or UO_2497 (O_2497,N_24248,N_28747);
nor UO_2498 (O_2498,N_28744,N_25809);
or UO_2499 (O_2499,N_29602,N_27797);
nor UO_2500 (O_2500,N_24820,N_26693);
nand UO_2501 (O_2501,N_24751,N_27626);
and UO_2502 (O_2502,N_28392,N_26360);
nor UO_2503 (O_2503,N_29792,N_24355);
or UO_2504 (O_2504,N_28178,N_25407);
and UO_2505 (O_2505,N_27589,N_26419);
or UO_2506 (O_2506,N_26594,N_24536);
xor UO_2507 (O_2507,N_27423,N_24662);
or UO_2508 (O_2508,N_26367,N_26389);
xnor UO_2509 (O_2509,N_29053,N_26785);
xor UO_2510 (O_2510,N_25690,N_28594);
xnor UO_2511 (O_2511,N_24531,N_25984);
nand UO_2512 (O_2512,N_25719,N_28369);
nor UO_2513 (O_2513,N_28107,N_27325);
xnor UO_2514 (O_2514,N_26236,N_29573);
or UO_2515 (O_2515,N_24401,N_28075);
nand UO_2516 (O_2516,N_26193,N_28317);
and UO_2517 (O_2517,N_28466,N_26602);
nor UO_2518 (O_2518,N_29676,N_29119);
nor UO_2519 (O_2519,N_29339,N_28073);
nand UO_2520 (O_2520,N_24739,N_26110);
xnor UO_2521 (O_2521,N_26556,N_25077);
xnor UO_2522 (O_2522,N_27208,N_24049);
nand UO_2523 (O_2523,N_28505,N_28062);
or UO_2524 (O_2524,N_26854,N_28140);
nand UO_2525 (O_2525,N_26549,N_27160);
and UO_2526 (O_2526,N_29153,N_26088);
nand UO_2527 (O_2527,N_29887,N_27683);
nand UO_2528 (O_2528,N_27390,N_27794);
nand UO_2529 (O_2529,N_27583,N_29366);
or UO_2530 (O_2530,N_26099,N_25923);
and UO_2531 (O_2531,N_25539,N_26863);
or UO_2532 (O_2532,N_29817,N_27783);
nand UO_2533 (O_2533,N_29253,N_26979);
or UO_2534 (O_2534,N_27444,N_24765);
and UO_2535 (O_2535,N_28725,N_25838);
xnor UO_2536 (O_2536,N_27617,N_24106);
nor UO_2537 (O_2537,N_27601,N_24677);
nor UO_2538 (O_2538,N_25950,N_29787);
or UO_2539 (O_2539,N_28133,N_24253);
or UO_2540 (O_2540,N_28772,N_29927);
nand UO_2541 (O_2541,N_28791,N_28777);
and UO_2542 (O_2542,N_27196,N_29144);
nand UO_2543 (O_2543,N_28388,N_28829);
xnor UO_2544 (O_2544,N_25605,N_24396);
nor UO_2545 (O_2545,N_26606,N_25799);
and UO_2546 (O_2546,N_27120,N_26315);
nand UO_2547 (O_2547,N_26938,N_26844);
nand UO_2548 (O_2548,N_27152,N_29465);
or UO_2549 (O_2549,N_24458,N_25126);
nand UO_2550 (O_2550,N_27055,N_29874);
xor UO_2551 (O_2551,N_27720,N_27405);
or UO_2552 (O_2552,N_25153,N_24644);
or UO_2553 (O_2553,N_29931,N_29564);
xor UO_2554 (O_2554,N_25338,N_25860);
xor UO_2555 (O_2555,N_26977,N_25073);
xnor UO_2556 (O_2556,N_28609,N_28311);
xor UO_2557 (O_2557,N_28978,N_28818);
nor UO_2558 (O_2558,N_27431,N_26637);
nand UO_2559 (O_2559,N_25591,N_26532);
nor UO_2560 (O_2560,N_28289,N_29051);
and UO_2561 (O_2561,N_25685,N_25474);
xor UO_2562 (O_2562,N_29454,N_25348);
xnor UO_2563 (O_2563,N_24630,N_25473);
and UO_2564 (O_2564,N_29127,N_28703);
nor UO_2565 (O_2565,N_24813,N_24411);
or UO_2566 (O_2566,N_24274,N_24761);
nor UO_2567 (O_2567,N_28796,N_24564);
nand UO_2568 (O_2568,N_25501,N_27902);
or UO_2569 (O_2569,N_27665,N_24622);
xor UO_2570 (O_2570,N_25654,N_24363);
nor UO_2571 (O_2571,N_25816,N_28373);
and UO_2572 (O_2572,N_27245,N_29198);
nand UO_2573 (O_2573,N_24790,N_28346);
and UO_2574 (O_2574,N_26492,N_27586);
and UO_2575 (O_2575,N_28875,N_27427);
nor UO_2576 (O_2576,N_27947,N_27789);
nor UO_2577 (O_2577,N_27356,N_24963);
xor UO_2578 (O_2578,N_26050,N_27397);
or UO_2579 (O_2579,N_29407,N_29958);
and UO_2580 (O_2580,N_29797,N_25707);
xnor UO_2581 (O_2581,N_26431,N_27746);
and UO_2582 (O_2582,N_24801,N_27091);
xnor UO_2583 (O_2583,N_25554,N_25755);
and UO_2584 (O_2584,N_25082,N_24175);
nor UO_2585 (O_2585,N_26311,N_27400);
xor UO_2586 (O_2586,N_27409,N_29811);
xor UO_2587 (O_2587,N_25422,N_29956);
nand UO_2588 (O_2588,N_24283,N_26166);
and UO_2589 (O_2589,N_27132,N_28218);
nand UO_2590 (O_2590,N_26067,N_29529);
nor UO_2591 (O_2591,N_25800,N_26320);
nor UO_2592 (O_2592,N_29906,N_27353);
nor UO_2593 (O_2593,N_28913,N_28580);
or UO_2594 (O_2594,N_28655,N_29776);
or UO_2595 (O_2595,N_29629,N_26853);
or UO_2596 (O_2596,N_28046,N_27110);
and UO_2597 (O_2597,N_29086,N_25097);
or UO_2598 (O_2598,N_25284,N_24476);
nand UO_2599 (O_2599,N_26980,N_27788);
nor UO_2600 (O_2600,N_27008,N_29648);
nand UO_2601 (O_2601,N_26482,N_27424);
or UO_2602 (O_2602,N_27031,N_27260);
nand UO_2603 (O_2603,N_24527,N_24701);
and UO_2604 (O_2604,N_24417,N_29446);
nor UO_2605 (O_2605,N_25595,N_26686);
nor UO_2606 (O_2606,N_28025,N_28159);
xnor UO_2607 (O_2607,N_29528,N_26004);
xnor UO_2608 (O_2608,N_27854,N_28518);
and UO_2609 (O_2609,N_28935,N_25494);
nand UO_2610 (O_2610,N_25080,N_28463);
nor UO_2611 (O_2611,N_28911,N_25565);
nand UO_2612 (O_2612,N_29950,N_24726);
or UO_2613 (O_2613,N_26731,N_24945);
nor UO_2614 (O_2614,N_26909,N_28537);
or UO_2615 (O_2615,N_29412,N_24280);
nor UO_2616 (O_2616,N_27864,N_29855);
nor UO_2617 (O_2617,N_29068,N_26009);
and UO_2618 (O_2618,N_25469,N_28260);
nor UO_2619 (O_2619,N_27223,N_26028);
or UO_2620 (O_2620,N_27203,N_28301);
xnor UO_2621 (O_2621,N_24287,N_26809);
nor UO_2622 (O_2622,N_27404,N_27919);
nor UO_2623 (O_2623,N_29987,N_26040);
and UO_2624 (O_2624,N_27380,N_24682);
nor UO_2625 (O_2625,N_29596,N_27221);
nand UO_2626 (O_2626,N_26995,N_28874);
nor UO_2627 (O_2627,N_26958,N_24113);
or UO_2628 (O_2628,N_25318,N_25484);
nand UO_2629 (O_2629,N_27332,N_29396);
xnor UO_2630 (O_2630,N_25470,N_25903);
xor UO_2631 (O_2631,N_28544,N_29070);
and UO_2632 (O_2632,N_26354,N_24780);
nand UO_2633 (O_2633,N_29778,N_29690);
nor UO_2634 (O_2634,N_28047,N_28027);
or UO_2635 (O_2635,N_29769,N_28209);
or UO_2636 (O_2636,N_26309,N_29746);
xnor UO_2637 (O_2637,N_26005,N_28335);
or UO_2638 (O_2638,N_28756,N_29207);
or UO_2639 (O_2639,N_25391,N_29848);
nand UO_2640 (O_2640,N_24872,N_24418);
nor UO_2641 (O_2641,N_28348,N_25777);
and UO_2642 (O_2642,N_24256,N_27168);
nor UO_2643 (O_2643,N_28407,N_29680);
or UO_2644 (O_2644,N_25017,N_24381);
xor UO_2645 (O_2645,N_27215,N_24471);
xnor UO_2646 (O_2646,N_28589,N_26025);
nor UO_2647 (O_2647,N_28267,N_24020);
nand UO_2648 (O_2648,N_27616,N_24616);
nor UO_2649 (O_2649,N_25576,N_27545);
nor UO_2650 (O_2650,N_29953,N_24304);
or UO_2651 (O_2651,N_29526,N_28455);
or UO_2652 (O_2652,N_26128,N_29615);
nand UO_2653 (O_2653,N_27484,N_29513);
and UO_2654 (O_2654,N_29264,N_29753);
nand UO_2655 (O_2655,N_27362,N_27200);
xor UO_2656 (O_2656,N_24343,N_26224);
nor UO_2657 (O_2657,N_25190,N_28096);
and UO_2658 (O_2658,N_26659,N_24700);
nand UO_2659 (O_2659,N_27330,N_27317);
nand UO_2660 (O_2660,N_28113,N_27914);
and UO_2661 (O_2661,N_25579,N_26762);
xor UO_2662 (O_2662,N_27107,N_24302);
nand UO_2663 (O_2663,N_25706,N_29731);
nand UO_2664 (O_2664,N_29654,N_26719);
or UO_2665 (O_2665,N_29775,N_25490);
nor UO_2666 (O_2666,N_25599,N_27078);
and UO_2667 (O_2667,N_25686,N_28151);
nor UO_2668 (O_2668,N_29415,N_24030);
nor UO_2669 (O_2669,N_24430,N_25227);
or UO_2670 (O_2670,N_28632,N_25822);
and UO_2671 (O_2671,N_29259,N_29782);
nand UO_2672 (O_2672,N_25363,N_25915);
xor UO_2673 (O_2673,N_25128,N_29838);
and UO_2674 (O_2674,N_29943,N_29623);
or UO_2675 (O_2675,N_29951,N_24646);
or UO_2676 (O_2676,N_24091,N_24540);
and UO_2677 (O_2677,N_27276,N_26405);
nor UO_2678 (O_2678,N_27562,N_24223);
or UO_2679 (O_2679,N_26963,N_28322);
xnor UO_2680 (O_2680,N_28148,N_29476);
nand UO_2681 (O_2681,N_24128,N_28076);
and UO_2682 (O_2682,N_26129,N_26912);
nor UO_2683 (O_2683,N_27357,N_28446);
or UO_2684 (O_2684,N_28571,N_26499);
nor UO_2685 (O_2685,N_27951,N_24369);
and UO_2686 (O_2686,N_25246,N_29784);
and UO_2687 (O_2687,N_26937,N_27836);
nor UO_2688 (O_2688,N_28785,N_27233);
xor UO_2689 (O_2689,N_25454,N_24266);
nand UO_2690 (O_2690,N_28902,N_25175);
xnor UO_2691 (O_2691,N_26838,N_28279);
and UO_2692 (O_2692,N_26518,N_26421);
nor UO_2693 (O_2693,N_26470,N_29439);
nor UO_2694 (O_2694,N_29822,N_26178);
nand UO_2695 (O_2695,N_24021,N_25935);
nand UO_2696 (O_2696,N_28305,N_29764);
and UO_2697 (O_2697,N_26001,N_24334);
xor UO_2698 (O_2698,N_27955,N_28021);
and UO_2699 (O_2699,N_25681,N_26867);
and UO_2700 (O_2700,N_25417,N_24421);
xnor UO_2701 (O_2701,N_27247,N_29617);
or UO_2702 (O_2702,N_24597,N_28217);
nor UO_2703 (O_2703,N_27529,N_25678);
xnor UO_2704 (O_2704,N_27737,N_25995);
nor UO_2705 (O_2705,N_27637,N_25437);
or UO_2706 (O_2706,N_29117,N_24416);
and UO_2707 (O_2707,N_29208,N_25852);
nand UO_2708 (O_2708,N_24121,N_27892);
nand UO_2709 (O_2709,N_25466,N_27835);
nand UO_2710 (O_2710,N_24131,N_25385);
nor UO_2711 (O_2711,N_27546,N_27792);
or UO_2712 (O_2712,N_26765,N_28094);
nor UO_2713 (O_2713,N_27807,N_29406);
and UO_2714 (O_2714,N_25118,N_25503);
nand UO_2715 (O_2715,N_24393,N_28751);
xnor UO_2716 (O_2716,N_27316,N_27598);
nor UO_2717 (O_2717,N_27980,N_26280);
nand UO_2718 (O_2718,N_29672,N_28715);
and UO_2719 (O_2719,N_25105,N_26634);
nor UO_2720 (O_2720,N_26947,N_25711);
nand UO_2721 (O_2721,N_26097,N_29089);
and UO_2722 (O_2722,N_29334,N_25541);
and UO_2723 (O_2723,N_29378,N_26294);
nor UO_2724 (O_2724,N_29294,N_25332);
and UO_2725 (O_2725,N_29844,N_27872);
xnor UO_2726 (O_2726,N_25533,N_25772);
nor UO_2727 (O_2727,N_29155,N_27218);
nor UO_2728 (O_2728,N_26197,N_27905);
nand UO_2729 (O_2729,N_24731,N_25156);
nor UO_2730 (O_2730,N_28954,N_27314);
or UO_2731 (O_2731,N_28966,N_25563);
xnor UO_2732 (O_2732,N_27066,N_29790);
and UO_2733 (O_2733,N_24084,N_27216);
or UO_2734 (O_2734,N_28592,N_27907);
or UO_2735 (O_2735,N_25648,N_25326);
nor UO_2736 (O_2736,N_27134,N_27018);
nand UO_2737 (O_2737,N_27264,N_26064);
nand UO_2738 (O_2738,N_25936,N_27494);
or UO_2739 (O_2739,N_29907,N_29549);
or UO_2740 (O_2740,N_27938,N_28722);
and UO_2741 (O_2741,N_25702,N_27072);
nor UO_2742 (O_2742,N_29299,N_27731);
and UO_2743 (O_2743,N_25705,N_28306);
xnor UO_2744 (O_2744,N_24515,N_27547);
nor UO_2745 (O_2745,N_26813,N_29703);
xor UO_2746 (O_2746,N_26146,N_28294);
and UO_2747 (O_2747,N_25585,N_27584);
nand UO_2748 (O_2748,N_29440,N_28936);
nand UO_2749 (O_2749,N_26911,N_29934);
or UO_2750 (O_2750,N_27213,N_26699);
nand UO_2751 (O_2751,N_27572,N_25065);
and UO_2752 (O_2752,N_24389,N_27544);
nor UO_2753 (O_2753,N_24272,N_24261);
and UO_2754 (O_2754,N_28705,N_26300);
or UO_2755 (O_2755,N_28985,N_28182);
nor UO_2756 (O_2756,N_26820,N_29912);
nand UO_2757 (O_2757,N_28039,N_24944);
xor UO_2758 (O_2758,N_27331,N_26417);
nand UO_2759 (O_2759,N_27138,N_29044);
xnor UO_2760 (O_2760,N_24295,N_29862);
xnor UO_2761 (O_2761,N_26636,N_28324);
and UO_2762 (O_2762,N_25897,N_28318);
nand UO_2763 (O_2763,N_29739,N_25198);
nand UO_2764 (O_2764,N_28053,N_24236);
nand UO_2765 (O_2765,N_26657,N_28865);
nand UO_2766 (O_2766,N_26723,N_28599);
or UO_2767 (O_2767,N_24085,N_24190);
nand UO_2768 (O_2768,N_29631,N_24406);
or UO_2769 (O_2769,N_26516,N_29954);
or UO_2770 (O_2770,N_24929,N_25545);
nor UO_2771 (O_2771,N_28363,N_28387);
xor UO_2772 (O_2772,N_25839,N_27557);
or UO_2773 (O_2773,N_27010,N_25917);
xnor UO_2774 (O_2774,N_28522,N_25109);
nand UO_2775 (O_2775,N_24345,N_26906);
nand UO_2776 (O_2776,N_26910,N_26789);
nand UO_2777 (O_2777,N_24149,N_29457);
and UO_2778 (O_2778,N_29345,N_24379);
nand UO_2779 (O_2779,N_28840,N_25205);
nand UO_2780 (O_2780,N_27680,N_24311);
and UO_2781 (O_2781,N_29889,N_26145);
nand UO_2782 (O_2782,N_28459,N_25932);
or UO_2783 (O_2783,N_24390,N_25699);
and UO_2784 (O_2784,N_26904,N_25260);
nand UO_2785 (O_2785,N_27059,N_29900);
or UO_2786 (O_2786,N_26984,N_24898);
xor UO_2787 (O_2787,N_27711,N_24818);
and UO_2788 (O_2788,N_29400,N_24042);
and UO_2789 (O_2789,N_28759,N_24987);
nor UO_2790 (O_2790,N_24133,N_27921);
or UO_2791 (O_2791,N_25224,N_29261);
xor UO_2792 (O_2792,N_24462,N_27255);
nor UO_2793 (O_2793,N_28071,N_27187);
xor UO_2794 (O_2794,N_29385,N_27128);
and UO_2795 (O_2795,N_24034,N_28181);
and UO_2796 (O_2796,N_25321,N_26089);
or UO_2797 (O_2797,N_26816,N_26210);
and UO_2798 (O_2798,N_29696,N_24060);
nand UO_2799 (O_2799,N_29748,N_29380);
nor UO_2800 (O_2800,N_26733,N_25147);
and UO_2801 (O_2801,N_29165,N_28654);
and UO_2802 (O_2802,N_26339,N_25497);
or UO_2803 (O_2803,N_27005,N_27993);
nand UO_2804 (O_2804,N_29656,N_28112);
or UO_2805 (O_2805,N_26567,N_29740);
nor UO_2806 (O_2806,N_24257,N_28924);
and UO_2807 (O_2807,N_28433,N_29503);
nor UO_2808 (O_2808,N_25869,N_28237);
xor UO_2809 (O_2809,N_24478,N_25471);
nand UO_2810 (O_2810,N_27659,N_26085);
or UO_2811 (O_2811,N_26024,N_28508);
nand UO_2812 (O_2812,N_24692,N_25620);
and UO_2813 (O_2813,N_25583,N_27856);
xnor UO_2814 (O_2814,N_25957,N_24664);
nand UO_2815 (O_2815,N_29870,N_27315);
and UO_2816 (O_2816,N_27758,N_28901);
or UO_2817 (O_2817,N_26228,N_27291);
nand UO_2818 (O_2818,N_27252,N_27689);
xnor UO_2819 (O_2819,N_26808,N_24696);
nor UO_2820 (O_2820,N_24125,N_26000);
nand UO_2821 (O_2821,N_28149,N_29982);
or UO_2822 (O_2822,N_25710,N_29186);
and UO_2823 (O_2823,N_25216,N_27342);
nor UO_2824 (O_2824,N_28354,N_26474);
or UO_2825 (O_2825,N_27549,N_28934);
xor UO_2826 (O_2826,N_29371,N_26423);
nor UO_2827 (O_2827,N_27839,N_29663);
nand UO_2828 (O_2828,N_28628,N_27324);
nand UO_2829 (O_2829,N_25002,N_28977);
nor UO_2830 (O_2830,N_25069,N_24051);
or UO_2831 (O_2831,N_27831,N_29869);
xnor UO_2832 (O_2832,N_29403,N_26441);
xor UO_2833 (O_2833,N_27039,N_27791);
and UO_2834 (O_2834,N_28597,N_29266);
nor UO_2835 (O_2835,N_26647,N_26200);
or UO_2836 (O_2836,N_27429,N_27578);
nand UO_2837 (O_2837,N_26057,N_27825);
or UO_2838 (O_2838,N_25796,N_24277);
or UO_2839 (O_2839,N_27136,N_28595);
xnor UO_2840 (O_2840,N_29275,N_27401);
or UO_2841 (O_2841,N_26724,N_27958);
or UO_2842 (O_2842,N_29495,N_25615);
xor UO_2843 (O_2843,N_28302,N_26212);
nand UO_2844 (O_2844,N_26642,N_27606);
and UO_2845 (O_2845,N_25247,N_27448);
xnor UO_2846 (O_2846,N_26460,N_25396);
nor UO_2847 (O_2847,N_29693,N_25723);
nor UO_2848 (O_2848,N_29096,N_29063);
xnor UO_2849 (O_2849,N_28177,N_26774);
nor UO_2850 (O_2850,N_24136,N_27265);
nand UO_2851 (O_2851,N_29551,N_25138);
and UO_2852 (O_2852,N_26859,N_29387);
xnor UO_2853 (O_2853,N_29540,N_27815);
nor UO_2854 (O_2854,N_26213,N_29762);
xor UO_2855 (O_2855,N_28061,N_29878);
nand UO_2856 (O_2856,N_27049,N_29418);
nor UO_2857 (O_2857,N_28775,N_26728);
or UO_2858 (O_2858,N_25265,N_24041);
or UO_2859 (O_2859,N_29074,N_27519);
and UO_2860 (O_2860,N_24104,N_26523);
or UO_2861 (O_2861,N_26496,N_29437);
nor UO_2862 (O_2862,N_27487,N_28704);
xor UO_2863 (O_2863,N_25899,N_28733);
nor UO_2864 (O_2864,N_29587,N_29369);
or UO_2865 (O_2865,N_29873,N_26079);
nand UO_2866 (O_2866,N_29193,N_26773);
xor UO_2867 (O_2867,N_27732,N_27207);
and UO_2868 (O_2868,N_28171,N_28004);
nor UO_2869 (O_2869,N_27940,N_29864);
nor UO_2870 (O_2870,N_28710,N_24514);
or UO_2871 (O_2871,N_25291,N_29248);
nand UO_2872 (O_2872,N_25781,N_26869);
nor UO_2873 (O_2873,N_27454,N_26721);
and UO_2874 (O_2874,N_29105,N_25123);
nand UO_2875 (O_2875,N_29128,N_25737);
nand UO_2876 (O_2876,N_24424,N_29215);
nor UO_2877 (O_2877,N_26365,N_26289);
or UO_2878 (O_2878,N_28399,N_26528);
and UO_2879 (O_2879,N_24530,N_27079);
and UO_2880 (O_2880,N_26871,N_28162);
and UO_2881 (O_2881,N_24863,N_29492);
xnor UO_2882 (O_2882,N_26525,N_28465);
or UO_2883 (O_2883,N_26555,N_27707);
and UO_2884 (O_2884,N_27093,N_25967);
nor UO_2885 (O_2885,N_25844,N_25025);
or UO_2886 (O_2886,N_28472,N_26524);
nor UO_2887 (O_2887,N_26488,N_29928);
xnor UO_2888 (O_2888,N_24414,N_25898);
nand UO_2889 (O_2889,N_29200,N_25524);
and UO_2890 (O_2890,N_29435,N_25817);
and UO_2891 (O_2891,N_28792,N_25506);
or UO_2892 (O_2892,N_27709,N_26961);
xnor UO_2893 (O_2893,N_24088,N_24927);
nor UO_2894 (O_2894,N_26341,N_25356);
nand UO_2895 (O_2895,N_28709,N_28357);
nand UO_2896 (O_2896,N_26116,N_26020);
or UO_2897 (O_2897,N_26157,N_25448);
or UO_2898 (O_2898,N_24281,N_29606);
xnor UO_2899 (O_2899,N_26379,N_24437);
xnor UO_2900 (O_2900,N_28082,N_29571);
and UO_2901 (O_2901,N_29116,N_28492);
or UO_2902 (O_2902,N_24785,N_25462);
or UO_2903 (O_2903,N_24939,N_25309);
nand UO_2904 (O_2904,N_25656,N_28615);
or UO_2905 (O_2905,N_26015,N_25478);
or UO_2906 (O_2906,N_25267,N_29853);
nor UO_2907 (O_2907,N_28480,N_25955);
xor UO_2908 (O_2908,N_26426,N_26489);
nand UO_2909 (O_2909,N_28211,N_25876);
nand UO_2910 (O_2910,N_26957,N_24208);
xnor UO_2911 (O_2911,N_28130,N_27862);
xnor UO_2912 (O_2912,N_24619,N_24904);
nand UO_2913 (O_2913,N_27201,N_27263);
nor UO_2914 (O_2914,N_26742,N_27372);
or UO_2915 (O_2915,N_29701,N_29916);
or UO_2916 (O_2916,N_24312,N_27193);
nand UO_2917 (O_2917,N_27612,N_27691);
xor UO_2918 (O_2918,N_25504,N_25132);
nand UO_2919 (O_2919,N_25901,N_29314);
xor UO_2920 (O_2920,N_26857,N_28343);
xor UO_2921 (O_2921,N_24447,N_27126);
nand UO_2922 (O_2922,N_29821,N_29399);
nand UO_2923 (O_2923,N_25536,N_29295);
nor UO_2924 (O_2924,N_27997,N_24492);
xor UO_2925 (O_2925,N_29892,N_29894);
and UO_2926 (O_2926,N_25475,N_26479);
nand UO_2927 (O_2927,N_27116,N_27772);
or UO_2928 (O_2928,N_29458,N_27966);
xor UO_2929 (O_2929,N_29774,N_27705);
or UO_2930 (O_2930,N_27636,N_28422);
nand UO_2931 (O_2931,N_28916,N_24906);
nand UO_2932 (O_2932,N_25507,N_27522);
xnor UO_2933 (O_2933,N_26706,N_26698);
xnor UO_2934 (O_2934,N_29410,N_27452);
nand UO_2935 (O_2935,N_26604,N_28825);
nor UO_2936 (O_2936,N_29728,N_26439);
nand UO_2937 (O_2937,N_25881,N_25335);
nand UO_2938 (O_2938,N_27123,N_26697);
and UO_2939 (O_2939,N_28247,N_28926);
and UO_2940 (O_2940,N_29554,N_24777);
nand UO_2941 (O_2941,N_27012,N_24153);
xnor UO_2942 (O_2942,N_27391,N_27542);
nand UO_2943 (O_2943,N_28803,N_25600);
or UO_2944 (O_2944,N_25018,N_29448);
nand UO_2945 (O_2945,N_28176,N_26155);
nor UO_2946 (O_2946,N_28003,N_25645);
or UO_2947 (O_2947,N_28810,N_24624);
or UO_2948 (O_2948,N_24095,N_26455);
and UO_2949 (O_2949,N_28770,N_28192);
xor UO_2950 (O_2950,N_29019,N_26152);
and UO_2951 (O_2951,N_24306,N_27629);
and UO_2952 (O_2952,N_25534,N_28779);
and UO_2953 (O_2953,N_29664,N_28524);
or UO_2954 (O_2954,N_25682,N_28530);
and UO_2955 (O_2955,N_25692,N_29001);
xnor UO_2956 (O_2956,N_25296,N_25141);
nand UO_2957 (O_2957,N_28200,N_27876);
xor UO_2958 (O_2958,N_24094,N_25044);
and UO_2959 (O_2959,N_24528,N_25726);
nand UO_2960 (O_2960,N_28010,N_26872);
nand UO_2961 (O_2961,N_28679,N_29572);
nand UO_2962 (O_2962,N_25102,N_26433);
nand UO_2963 (O_2963,N_24137,N_28677);
nor UO_2964 (O_2964,N_27307,N_25836);
nand UO_2965 (O_2965,N_26752,N_24073);
nor UO_2966 (O_2966,N_26324,N_27170);
or UO_2967 (O_2967,N_26769,N_25633);
and UO_2968 (O_2968,N_29379,N_24824);
xnor UO_2969 (O_2969,N_29363,N_24292);
nor UO_2970 (O_2970,N_29616,N_25905);
nand UO_2971 (O_2971,N_24043,N_29918);
or UO_2972 (O_2972,N_29917,N_27776);
nor UO_2973 (O_2973,N_27023,N_25213);
and UO_2974 (O_2974,N_26827,N_28962);
nor UO_2975 (O_2975,N_24339,N_29223);
nor UO_2976 (O_2976,N_24598,N_27673);
nor UO_2977 (O_2977,N_28651,N_27040);
nand UO_2978 (O_2978,N_26208,N_28990);
xnor UO_2979 (O_2979,N_25890,N_27422);
nand UO_2980 (O_2980,N_26865,N_24014);
xor UO_2981 (O_2981,N_28894,N_25639);
or UO_2982 (O_2982,N_29434,N_25958);
nand UO_2983 (O_2983,N_24495,N_28737);
xnor UO_2984 (O_2984,N_24996,N_29519);
and UO_2985 (O_2985,N_28304,N_24717);
nand UO_2986 (O_2986,N_25362,N_24123);
nand UO_2987 (O_2987,N_29040,N_25011);
and UO_2988 (O_2988,N_26275,N_28298);
and UO_2989 (O_2989,N_25436,N_28646);
and UO_2990 (O_2990,N_29090,N_24120);
nor UO_2991 (O_2991,N_28835,N_26704);
xnor UO_2992 (O_2992,N_26852,N_26413);
or UO_2993 (O_2993,N_28389,N_27108);
or UO_2994 (O_2994,N_28541,N_25912);
nand UO_2995 (O_2995,N_27618,N_28098);
nor UO_2996 (O_2996,N_29567,N_25920);
and UO_2997 (O_2997,N_24518,N_24365);
xnor UO_2998 (O_2998,N_28547,N_24742);
nor UO_2999 (O_2999,N_29436,N_25269);
xor UO_3000 (O_3000,N_28408,N_26990);
and UO_3001 (O_3001,N_24065,N_26657);
nand UO_3002 (O_3002,N_28345,N_27936);
or UO_3003 (O_3003,N_25061,N_29701);
nor UO_3004 (O_3004,N_28351,N_28329);
and UO_3005 (O_3005,N_27678,N_29252);
and UO_3006 (O_3006,N_26835,N_25498);
or UO_3007 (O_3007,N_25451,N_29244);
nand UO_3008 (O_3008,N_27589,N_27835);
xnor UO_3009 (O_3009,N_25736,N_28939);
nor UO_3010 (O_3010,N_27329,N_25861);
nor UO_3011 (O_3011,N_28699,N_25798);
or UO_3012 (O_3012,N_25699,N_29347);
or UO_3013 (O_3013,N_25491,N_27517);
or UO_3014 (O_3014,N_25298,N_27161);
and UO_3015 (O_3015,N_25443,N_29659);
or UO_3016 (O_3016,N_29237,N_29768);
nand UO_3017 (O_3017,N_29167,N_28064);
and UO_3018 (O_3018,N_26872,N_29428);
nand UO_3019 (O_3019,N_27110,N_26146);
or UO_3020 (O_3020,N_26443,N_27140);
and UO_3021 (O_3021,N_24833,N_26899);
and UO_3022 (O_3022,N_28336,N_25810);
and UO_3023 (O_3023,N_28190,N_26321);
nand UO_3024 (O_3024,N_27276,N_28541);
nor UO_3025 (O_3025,N_25134,N_25527);
xnor UO_3026 (O_3026,N_26529,N_25322);
nor UO_3027 (O_3027,N_25308,N_25656);
and UO_3028 (O_3028,N_24749,N_29560);
or UO_3029 (O_3029,N_26699,N_27912);
xor UO_3030 (O_3030,N_29843,N_24427);
nor UO_3031 (O_3031,N_27493,N_26878);
xnor UO_3032 (O_3032,N_25359,N_27564);
nand UO_3033 (O_3033,N_25293,N_27845);
xor UO_3034 (O_3034,N_27284,N_27295);
and UO_3035 (O_3035,N_24297,N_26890);
or UO_3036 (O_3036,N_29743,N_29842);
xnor UO_3037 (O_3037,N_24817,N_29340);
xor UO_3038 (O_3038,N_25995,N_28212);
xnor UO_3039 (O_3039,N_28438,N_29168);
nand UO_3040 (O_3040,N_29200,N_25002);
and UO_3041 (O_3041,N_29305,N_25195);
or UO_3042 (O_3042,N_26866,N_24031);
nor UO_3043 (O_3043,N_25047,N_27314);
and UO_3044 (O_3044,N_24647,N_28391);
xnor UO_3045 (O_3045,N_24927,N_28731);
nand UO_3046 (O_3046,N_28851,N_28605);
or UO_3047 (O_3047,N_28943,N_24673);
nor UO_3048 (O_3048,N_26518,N_24858);
nor UO_3049 (O_3049,N_25811,N_24895);
and UO_3050 (O_3050,N_24615,N_26681);
xor UO_3051 (O_3051,N_26968,N_28279);
nand UO_3052 (O_3052,N_28148,N_28119);
nor UO_3053 (O_3053,N_26815,N_24005);
xor UO_3054 (O_3054,N_24255,N_24289);
or UO_3055 (O_3055,N_29461,N_28968);
nand UO_3056 (O_3056,N_27121,N_27871);
xnor UO_3057 (O_3057,N_24700,N_28284);
nand UO_3058 (O_3058,N_24307,N_24473);
nand UO_3059 (O_3059,N_27559,N_28230);
and UO_3060 (O_3060,N_27062,N_25721);
nor UO_3061 (O_3061,N_29099,N_25928);
and UO_3062 (O_3062,N_24754,N_27956);
xor UO_3063 (O_3063,N_24772,N_28706);
or UO_3064 (O_3064,N_28424,N_27766);
nor UO_3065 (O_3065,N_26249,N_29399);
and UO_3066 (O_3066,N_27062,N_24533);
or UO_3067 (O_3067,N_24206,N_26405);
nand UO_3068 (O_3068,N_25031,N_26042);
nor UO_3069 (O_3069,N_24667,N_24304);
and UO_3070 (O_3070,N_27001,N_26296);
and UO_3071 (O_3071,N_26019,N_28049);
nand UO_3072 (O_3072,N_26336,N_26191);
xnor UO_3073 (O_3073,N_24329,N_26002);
nand UO_3074 (O_3074,N_27463,N_27633);
nand UO_3075 (O_3075,N_25161,N_29372);
nand UO_3076 (O_3076,N_26952,N_29394);
nor UO_3077 (O_3077,N_24772,N_24259);
xnor UO_3078 (O_3078,N_24842,N_28015);
xnor UO_3079 (O_3079,N_29651,N_26451);
xnor UO_3080 (O_3080,N_29087,N_28449);
or UO_3081 (O_3081,N_28323,N_24621);
or UO_3082 (O_3082,N_25663,N_29892);
and UO_3083 (O_3083,N_27728,N_24418);
xnor UO_3084 (O_3084,N_28542,N_24991);
nor UO_3085 (O_3085,N_26647,N_25954);
nand UO_3086 (O_3086,N_28068,N_29728);
xor UO_3087 (O_3087,N_25648,N_29307);
or UO_3088 (O_3088,N_29218,N_28530);
xor UO_3089 (O_3089,N_27643,N_29204);
nand UO_3090 (O_3090,N_24382,N_26924);
nor UO_3091 (O_3091,N_27841,N_26779);
or UO_3092 (O_3092,N_28365,N_24487);
nand UO_3093 (O_3093,N_25340,N_24519);
xor UO_3094 (O_3094,N_24904,N_26740);
or UO_3095 (O_3095,N_26925,N_24059);
xor UO_3096 (O_3096,N_28104,N_29652);
and UO_3097 (O_3097,N_24871,N_25799);
or UO_3098 (O_3098,N_29682,N_28446);
xor UO_3099 (O_3099,N_26867,N_26882);
xnor UO_3100 (O_3100,N_27291,N_27855);
xor UO_3101 (O_3101,N_24633,N_28542);
or UO_3102 (O_3102,N_25572,N_24961);
nor UO_3103 (O_3103,N_24700,N_27269);
nor UO_3104 (O_3104,N_24058,N_26462);
nor UO_3105 (O_3105,N_27954,N_28397);
nor UO_3106 (O_3106,N_24473,N_27718);
xnor UO_3107 (O_3107,N_24036,N_24321);
xor UO_3108 (O_3108,N_27395,N_29947);
nor UO_3109 (O_3109,N_25256,N_25570);
or UO_3110 (O_3110,N_29237,N_25682);
nor UO_3111 (O_3111,N_24433,N_28497);
nor UO_3112 (O_3112,N_25735,N_28810);
xnor UO_3113 (O_3113,N_25890,N_29344);
nand UO_3114 (O_3114,N_29866,N_27039);
nor UO_3115 (O_3115,N_28244,N_26808);
nor UO_3116 (O_3116,N_24729,N_26566);
nor UO_3117 (O_3117,N_27121,N_26042);
or UO_3118 (O_3118,N_24692,N_26315);
and UO_3119 (O_3119,N_25021,N_29367);
and UO_3120 (O_3120,N_27143,N_24690);
nand UO_3121 (O_3121,N_27972,N_26027);
or UO_3122 (O_3122,N_25463,N_25925);
nand UO_3123 (O_3123,N_28191,N_28124);
and UO_3124 (O_3124,N_26485,N_24341);
and UO_3125 (O_3125,N_27514,N_28115);
xor UO_3126 (O_3126,N_26391,N_25746);
and UO_3127 (O_3127,N_24179,N_28176);
nor UO_3128 (O_3128,N_26901,N_25076);
nor UO_3129 (O_3129,N_24930,N_28556);
xnor UO_3130 (O_3130,N_25025,N_28419);
and UO_3131 (O_3131,N_24085,N_24232);
or UO_3132 (O_3132,N_24048,N_24999);
nor UO_3133 (O_3133,N_28144,N_24361);
and UO_3134 (O_3134,N_27308,N_27693);
or UO_3135 (O_3135,N_29487,N_28328);
and UO_3136 (O_3136,N_25580,N_29759);
nand UO_3137 (O_3137,N_29854,N_25743);
or UO_3138 (O_3138,N_28181,N_28831);
nor UO_3139 (O_3139,N_26857,N_28780);
or UO_3140 (O_3140,N_28839,N_29656);
xor UO_3141 (O_3141,N_27807,N_25631);
or UO_3142 (O_3142,N_25441,N_24939);
nand UO_3143 (O_3143,N_27160,N_28602);
or UO_3144 (O_3144,N_25588,N_26030);
and UO_3145 (O_3145,N_28069,N_28452);
nand UO_3146 (O_3146,N_24649,N_25425);
and UO_3147 (O_3147,N_24451,N_29462);
or UO_3148 (O_3148,N_24087,N_28142);
nor UO_3149 (O_3149,N_26115,N_27089);
or UO_3150 (O_3150,N_29246,N_26737);
and UO_3151 (O_3151,N_28786,N_27716);
nand UO_3152 (O_3152,N_24307,N_27738);
xnor UO_3153 (O_3153,N_26024,N_26463);
nand UO_3154 (O_3154,N_26054,N_29540);
and UO_3155 (O_3155,N_29367,N_29714);
xor UO_3156 (O_3156,N_27198,N_25155);
xor UO_3157 (O_3157,N_26313,N_24298);
xnor UO_3158 (O_3158,N_29194,N_26962);
nor UO_3159 (O_3159,N_25432,N_29225);
nand UO_3160 (O_3160,N_27005,N_29866);
xnor UO_3161 (O_3161,N_26171,N_25791);
xnor UO_3162 (O_3162,N_28138,N_25145);
and UO_3163 (O_3163,N_28476,N_24249);
nor UO_3164 (O_3164,N_26679,N_26972);
or UO_3165 (O_3165,N_27066,N_29158);
nor UO_3166 (O_3166,N_26629,N_26694);
and UO_3167 (O_3167,N_24437,N_27663);
nor UO_3168 (O_3168,N_29519,N_27941);
nand UO_3169 (O_3169,N_27313,N_26020);
xor UO_3170 (O_3170,N_26742,N_24759);
nor UO_3171 (O_3171,N_25649,N_29248);
nor UO_3172 (O_3172,N_28166,N_29380);
and UO_3173 (O_3173,N_24370,N_27212);
or UO_3174 (O_3174,N_24942,N_29015);
xnor UO_3175 (O_3175,N_26173,N_28389);
or UO_3176 (O_3176,N_29668,N_26626);
nand UO_3177 (O_3177,N_26306,N_27605);
and UO_3178 (O_3178,N_28654,N_27817);
and UO_3179 (O_3179,N_27657,N_27048);
and UO_3180 (O_3180,N_27261,N_29971);
nand UO_3181 (O_3181,N_28393,N_25854);
xor UO_3182 (O_3182,N_27094,N_27238);
and UO_3183 (O_3183,N_25719,N_29262);
nor UO_3184 (O_3184,N_29644,N_26500);
nand UO_3185 (O_3185,N_28411,N_29146);
or UO_3186 (O_3186,N_24940,N_28557);
nor UO_3187 (O_3187,N_26715,N_29578);
xor UO_3188 (O_3188,N_24731,N_25238);
xor UO_3189 (O_3189,N_27541,N_25081);
and UO_3190 (O_3190,N_27545,N_26538);
nor UO_3191 (O_3191,N_26443,N_27373);
and UO_3192 (O_3192,N_28002,N_25465);
nand UO_3193 (O_3193,N_24626,N_26997);
and UO_3194 (O_3194,N_24180,N_28786);
or UO_3195 (O_3195,N_28403,N_29048);
xnor UO_3196 (O_3196,N_24575,N_29310);
nand UO_3197 (O_3197,N_27926,N_28237);
and UO_3198 (O_3198,N_24144,N_29485);
nand UO_3199 (O_3199,N_26950,N_26624);
and UO_3200 (O_3200,N_29494,N_25851);
nand UO_3201 (O_3201,N_29132,N_24543);
xor UO_3202 (O_3202,N_28853,N_26117);
and UO_3203 (O_3203,N_27376,N_27805);
nand UO_3204 (O_3204,N_27288,N_24230);
nor UO_3205 (O_3205,N_27214,N_27793);
xor UO_3206 (O_3206,N_29854,N_26290);
or UO_3207 (O_3207,N_24707,N_25636);
nor UO_3208 (O_3208,N_25601,N_25048);
and UO_3209 (O_3209,N_25409,N_24170);
nor UO_3210 (O_3210,N_25898,N_26547);
and UO_3211 (O_3211,N_29545,N_25998);
nor UO_3212 (O_3212,N_29221,N_27654);
xnor UO_3213 (O_3213,N_28828,N_29729);
nand UO_3214 (O_3214,N_28761,N_29828);
nor UO_3215 (O_3215,N_26310,N_27453);
and UO_3216 (O_3216,N_24100,N_24002);
nand UO_3217 (O_3217,N_29068,N_29347);
nand UO_3218 (O_3218,N_26621,N_27139);
or UO_3219 (O_3219,N_27387,N_27352);
or UO_3220 (O_3220,N_26217,N_29465);
nor UO_3221 (O_3221,N_26003,N_24379);
or UO_3222 (O_3222,N_27097,N_29747);
nand UO_3223 (O_3223,N_29403,N_28644);
xor UO_3224 (O_3224,N_29763,N_24526);
nor UO_3225 (O_3225,N_25322,N_28940);
xor UO_3226 (O_3226,N_24710,N_26584);
nor UO_3227 (O_3227,N_28490,N_27753);
and UO_3228 (O_3228,N_25198,N_29726);
and UO_3229 (O_3229,N_28317,N_27379);
nor UO_3230 (O_3230,N_25016,N_29208);
and UO_3231 (O_3231,N_26973,N_28140);
or UO_3232 (O_3232,N_26879,N_25005);
and UO_3233 (O_3233,N_28256,N_26202);
or UO_3234 (O_3234,N_27527,N_24998);
nor UO_3235 (O_3235,N_28836,N_27607);
nor UO_3236 (O_3236,N_29224,N_28882);
or UO_3237 (O_3237,N_27589,N_28542);
nand UO_3238 (O_3238,N_26073,N_26647);
or UO_3239 (O_3239,N_29264,N_25960);
nand UO_3240 (O_3240,N_25200,N_25141);
xor UO_3241 (O_3241,N_28436,N_29795);
or UO_3242 (O_3242,N_28122,N_26830);
xor UO_3243 (O_3243,N_25125,N_29235);
nand UO_3244 (O_3244,N_25335,N_27698);
nand UO_3245 (O_3245,N_27536,N_26422);
or UO_3246 (O_3246,N_27478,N_24887);
nor UO_3247 (O_3247,N_29494,N_24731);
and UO_3248 (O_3248,N_28030,N_25359);
and UO_3249 (O_3249,N_28161,N_29483);
nor UO_3250 (O_3250,N_29973,N_26374);
xor UO_3251 (O_3251,N_26640,N_25133);
nor UO_3252 (O_3252,N_29924,N_29658);
nor UO_3253 (O_3253,N_28562,N_26109);
or UO_3254 (O_3254,N_24462,N_26432);
nor UO_3255 (O_3255,N_27911,N_27302);
xnor UO_3256 (O_3256,N_26358,N_27336);
nand UO_3257 (O_3257,N_27577,N_25415);
or UO_3258 (O_3258,N_25354,N_25528);
xor UO_3259 (O_3259,N_24372,N_26109);
xor UO_3260 (O_3260,N_27984,N_28976);
or UO_3261 (O_3261,N_26887,N_25148);
nor UO_3262 (O_3262,N_28133,N_29369);
nor UO_3263 (O_3263,N_29345,N_24621);
nor UO_3264 (O_3264,N_27297,N_29336);
or UO_3265 (O_3265,N_27028,N_28336);
xor UO_3266 (O_3266,N_24281,N_26954);
nor UO_3267 (O_3267,N_29531,N_27521);
and UO_3268 (O_3268,N_29083,N_29425);
or UO_3269 (O_3269,N_24279,N_25012);
nand UO_3270 (O_3270,N_25416,N_26584);
and UO_3271 (O_3271,N_26962,N_28945);
and UO_3272 (O_3272,N_29779,N_29216);
nor UO_3273 (O_3273,N_29867,N_29105);
xor UO_3274 (O_3274,N_26904,N_28492);
and UO_3275 (O_3275,N_24042,N_24748);
and UO_3276 (O_3276,N_28831,N_27355);
and UO_3277 (O_3277,N_29263,N_24658);
nand UO_3278 (O_3278,N_24602,N_28628);
nand UO_3279 (O_3279,N_26377,N_24094);
xnor UO_3280 (O_3280,N_24479,N_26971);
or UO_3281 (O_3281,N_26396,N_24480);
nand UO_3282 (O_3282,N_28758,N_29810);
xor UO_3283 (O_3283,N_29392,N_28584);
or UO_3284 (O_3284,N_28099,N_29215);
and UO_3285 (O_3285,N_28120,N_29661);
nor UO_3286 (O_3286,N_29266,N_28918);
nand UO_3287 (O_3287,N_26203,N_25963);
or UO_3288 (O_3288,N_25242,N_29794);
nor UO_3289 (O_3289,N_27119,N_28395);
xnor UO_3290 (O_3290,N_26221,N_29058);
and UO_3291 (O_3291,N_28462,N_26294);
and UO_3292 (O_3292,N_26063,N_26726);
nand UO_3293 (O_3293,N_26296,N_28720);
nor UO_3294 (O_3294,N_28985,N_24442);
or UO_3295 (O_3295,N_28381,N_28621);
nor UO_3296 (O_3296,N_24196,N_28041);
and UO_3297 (O_3297,N_27116,N_27167);
nand UO_3298 (O_3298,N_27204,N_24494);
nor UO_3299 (O_3299,N_24035,N_24459);
nor UO_3300 (O_3300,N_24692,N_24482);
and UO_3301 (O_3301,N_25096,N_26521);
nand UO_3302 (O_3302,N_28293,N_25507);
xor UO_3303 (O_3303,N_28314,N_25194);
or UO_3304 (O_3304,N_26056,N_28316);
xor UO_3305 (O_3305,N_26554,N_24468);
nor UO_3306 (O_3306,N_29900,N_25319);
nand UO_3307 (O_3307,N_27124,N_29058);
or UO_3308 (O_3308,N_25558,N_28279);
or UO_3309 (O_3309,N_24528,N_27100);
nand UO_3310 (O_3310,N_25312,N_25265);
xor UO_3311 (O_3311,N_26740,N_25912);
or UO_3312 (O_3312,N_25967,N_25322);
and UO_3313 (O_3313,N_27418,N_27228);
xnor UO_3314 (O_3314,N_25151,N_27016);
nor UO_3315 (O_3315,N_28754,N_25224);
or UO_3316 (O_3316,N_24748,N_26493);
nor UO_3317 (O_3317,N_29514,N_29188);
and UO_3318 (O_3318,N_27495,N_29571);
nand UO_3319 (O_3319,N_26484,N_25531);
xnor UO_3320 (O_3320,N_24140,N_24213);
xnor UO_3321 (O_3321,N_25428,N_29590);
and UO_3322 (O_3322,N_25590,N_29309);
or UO_3323 (O_3323,N_25983,N_24231);
nand UO_3324 (O_3324,N_24508,N_25691);
or UO_3325 (O_3325,N_29902,N_29571);
and UO_3326 (O_3326,N_25610,N_24292);
and UO_3327 (O_3327,N_24755,N_24967);
and UO_3328 (O_3328,N_27832,N_29694);
and UO_3329 (O_3329,N_29775,N_29236);
or UO_3330 (O_3330,N_25432,N_27349);
and UO_3331 (O_3331,N_27765,N_25456);
nor UO_3332 (O_3332,N_29239,N_28011);
nor UO_3333 (O_3333,N_25676,N_28988);
or UO_3334 (O_3334,N_26350,N_29250);
nor UO_3335 (O_3335,N_27540,N_24942);
and UO_3336 (O_3336,N_25064,N_26438);
and UO_3337 (O_3337,N_29550,N_28688);
xnor UO_3338 (O_3338,N_25865,N_27127);
nor UO_3339 (O_3339,N_24321,N_24976);
xnor UO_3340 (O_3340,N_29984,N_29986);
xnor UO_3341 (O_3341,N_25702,N_26540);
xnor UO_3342 (O_3342,N_26790,N_27607);
and UO_3343 (O_3343,N_28807,N_29009);
and UO_3344 (O_3344,N_25591,N_25695);
xnor UO_3345 (O_3345,N_24395,N_29035);
or UO_3346 (O_3346,N_28649,N_25528);
nor UO_3347 (O_3347,N_28435,N_27424);
nand UO_3348 (O_3348,N_29950,N_25879);
xor UO_3349 (O_3349,N_26663,N_28847);
xor UO_3350 (O_3350,N_24791,N_26388);
and UO_3351 (O_3351,N_25285,N_25301);
xnor UO_3352 (O_3352,N_29312,N_26213);
or UO_3353 (O_3353,N_25566,N_25283);
or UO_3354 (O_3354,N_27346,N_25544);
and UO_3355 (O_3355,N_29273,N_25671);
xor UO_3356 (O_3356,N_26612,N_24919);
xnor UO_3357 (O_3357,N_24659,N_27283);
and UO_3358 (O_3358,N_25223,N_24445);
nand UO_3359 (O_3359,N_24688,N_28866);
xor UO_3360 (O_3360,N_27670,N_29448);
xnor UO_3361 (O_3361,N_27125,N_26159);
nor UO_3362 (O_3362,N_29634,N_24145);
and UO_3363 (O_3363,N_29822,N_27102);
xnor UO_3364 (O_3364,N_28752,N_26029);
nor UO_3365 (O_3365,N_24269,N_29900);
nor UO_3366 (O_3366,N_25728,N_25099);
xnor UO_3367 (O_3367,N_26810,N_26344);
xor UO_3368 (O_3368,N_29718,N_27111);
and UO_3369 (O_3369,N_26619,N_26717);
xor UO_3370 (O_3370,N_26026,N_28776);
nand UO_3371 (O_3371,N_24750,N_29148);
or UO_3372 (O_3372,N_29839,N_25209);
nor UO_3373 (O_3373,N_28745,N_24954);
nand UO_3374 (O_3374,N_25830,N_25675);
and UO_3375 (O_3375,N_28542,N_25074);
and UO_3376 (O_3376,N_28193,N_27529);
and UO_3377 (O_3377,N_29350,N_25343);
and UO_3378 (O_3378,N_24091,N_25639);
or UO_3379 (O_3379,N_25299,N_29949);
or UO_3380 (O_3380,N_27048,N_25443);
xnor UO_3381 (O_3381,N_27209,N_28687);
nor UO_3382 (O_3382,N_28652,N_27549);
nor UO_3383 (O_3383,N_24460,N_28377);
and UO_3384 (O_3384,N_24624,N_26927);
xnor UO_3385 (O_3385,N_26288,N_26168);
xnor UO_3386 (O_3386,N_25970,N_24127);
xnor UO_3387 (O_3387,N_25725,N_25449);
and UO_3388 (O_3388,N_24630,N_26059);
or UO_3389 (O_3389,N_27485,N_26048);
or UO_3390 (O_3390,N_25464,N_28338);
nor UO_3391 (O_3391,N_25810,N_27543);
nor UO_3392 (O_3392,N_24011,N_24204);
xor UO_3393 (O_3393,N_25464,N_28642);
xnor UO_3394 (O_3394,N_26236,N_29242);
nand UO_3395 (O_3395,N_29116,N_28328);
or UO_3396 (O_3396,N_29868,N_24641);
xnor UO_3397 (O_3397,N_29287,N_29451);
nand UO_3398 (O_3398,N_24732,N_26225);
nor UO_3399 (O_3399,N_25698,N_25040);
nor UO_3400 (O_3400,N_24845,N_26919);
nand UO_3401 (O_3401,N_24103,N_29380);
xnor UO_3402 (O_3402,N_26207,N_26463);
nand UO_3403 (O_3403,N_25376,N_26492);
and UO_3404 (O_3404,N_24673,N_29211);
xor UO_3405 (O_3405,N_24176,N_26358);
and UO_3406 (O_3406,N_29828,N_27413);
xor UO_3407 (O_3407,N_27784,N_28881);
and UO_3408 (O_3408,N_24418,N_27921);
nor UO_3409 (O_3409,N_29469,N_27251);
nand UO_3410 (O_3410,N_26277,N_27932);
nand UO_3411 (O_3411,N_27650,N_29355);
or UO_3412 (O_3412,N_26623,N_25497);
nand UO_3413 (O_3413,N_29172,N_27503);
nand UO_3414 (O_3414,N_24478,N_28666);
or UO_3415 (O_3415,N_25848,N_25781);
and UO_3416 (O_3416,N_24906,N_28516);
and UO_3417 (O_3417,N_24516,N_25558);
nand UO_3418 (O_3418,N_25758,N_26114);
or UO_3419 (O_3419,N_26641,N_29144);
xnor UO_3420 (O_3420,N_28630,N_29922);
nor UO_3421 (O_3421,N_24382,N_26947);
and UO_3422 (O_3422,N_28652,N_26649);
nand UO_3423 (O_3423,N_26813,N_24209);
xnor UO_3424 (O_3424,N_27678,N_25237);
and UO_3425 (O_3425,N_28266,N_29086);
xnor UO_3426 (O_3426,N_27594,N_29631);
nand UO_3427 (O_3427,N_24257,N_29165);
xnor UO_3428 (O_3428,N_28097,N_26211);
nor UO_3429 (O_3429,N_26738,N_26063);
and UO_3430 (O_3430,N_28567,N_26887);
or UO_3431 (O_3431,N_28205,N_27250);
nor UO_3432 (O_3432,N_24004,N_29190);
and UO_3433 (O_3433,N_28188,N_26065);
xor UO_3434 (O_3434,N_27528,N_29073);
or UO_3435 (O_3435,N_25832,N_29302);
nor UO_3436 (O_3436,N_26751,N_29267);
nor UO_3437 (O_3437,N_26150,N_24769);
xnor UO_3438 (O_3438,N_28950,N_28041);
and UO_3439 (O_3439,N_26107,N_29846);
and UO_3440 (O_3440,N_27834,N_26357);
nor UO_3441 (O_3441,N_28348,N_25592);
nand UO_3442 (O_3442,N_25478,N_26863);
nor UO_3443 (O_3443,N_27450,N_27351);
nand UO_3444 (O_3444,N_26311,N_29998);
xnor UO_3445 (O_3445,N_28413,N_28174);
xor UO_3446 (O_3446,N_29812,N_29920);
nor UO_3447 (O_3447,N_27760,N_27126);
and UO_3448 (O_3448,N_26227,N_26270);
nor UO_3449 (O_3449,N_24023,N_27626);
nor UO_3450 (O_3450,N_28590,N_27633);
nor UO_3451 (O_3451,N_25805,N_25085);
or UO_3452 (O_3452,N_28677,N_25421);
and UO_3453 (O_3453,N_27338,N_27639);
and UO_3454 (O_3454,N_28483,N_26656);
and UO_3455 (O_3455,N_28111,N_28142);
nand UO_3456 (O_3456,N_29827,N_27741);
nor UO_3457 (O_3457,N_25390,N_29420);
or UO_3458 (O_3458,N_29718,N_26629);
and UO_3459 (O_3459,N_29975,N_28341);
nor UO_3460 (O_3460,N_28236,N_25288);
nand UO_3461 (O_3461,N_26326,N_28200);
nor UO_3462 (O_3462,N_25792,N_27209);
or UO_3463 (O_3463,N_28714,N_27466);
xnor UO_3464 (O_3464,N_27934,N_25347);
and UO_3465 (O_3465,N_29293,N_25922);
or UO_3466 (O_3466,N_29898,N_25411);
nand UO_3467 (O_3467,N_27376,N_24487);
nor UO_3468 (O_3468,N_24927,N_24153);
and UO_3469 (O_3469,N_27064,N_29495);
xnor UO_3470 (O_3470,N_29978,N_25331);
or UO_3471 (O_3471,N_24501,N_25468);
xor UO_3472 (O_3472,N_24148,N_25979);
or UO_3473 (O_3473,N_24037,N_25485);
xnor UO_3474 (O_3474,N_24715,N_28904);
nand UO_3475 (O_3475,N_27812,N_26410);
nand UO_3476 (O_3476,N_29172,N_28217);
xor UO_3477 (O_3477,N_29593,N_24983);
nor UO_3478 (O_3478,N_26175,N_25748);
and UO_3479 (O_3479,N_26248,N_25902);
nand UO_3480 (O_3480,N_25207,N_24542);
nor UO_3481 (O_3481,N_27920,N_27210);
nor UO_3482 (O_3482,N_26756,N_29012);
or UO_3483 (O_3483,N_26394,N_28591);
nand UO_3484 (O_3484,N_25942,N_24206);
nand UO_3485 (O_3485,N_26340,N_25864);
nor UO_3486 (O_3486,N_26653,N_27974);
xnor UO_3487 (O_3487,N_28297,N_28382);
nand UO_3488 (O_3488,N_26996,N_24988);
and UO_3489 (O_3489,N_26838,N_25633);
nor UO_3490 (O_3490,N_25143,N_28884);
and UO_3491 (O_3491,N_28052,N_24335);
xor UO_3492 (O_3492,N_24448,N_26768);
xnor UO_3493 (O_3493,N_26657,N_24071);
nand UO_3494 (O_3494,N_27890,N_27528);
nand UO_3495 (O_3495,N_27965,N_25404);
xnor UO_3496 (O_3496,N_27348,N_27701);
nor UO_3497 (O_3497,N_24389,N_29365);
nor UO_3498 (O_3498,N_29718,N_24284);
nor UO_3499 (O_3499,N_26211,N_25173);
endmodule