module basic_500_3000_500_5_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_20,In_80);
xnor U1 (N_1,In_42,In_464);
nand U2 (N_2,In_237,In_267);
nand U3 (N_3,In_454,In_384);
and U4 (N_4,In_248,In_32);
nor U5 (N_5,In_87,In_219);
nor U6 (N_6,In_220,In_240);
nor U7 (N_7,In_193,In_430);
nand U8 (N_8,In_132,In_272);
nand U9 (N_9,In_98,In_168);
nor U10 (N_10,In_497,In_301);
nor U11 (N_11,In_271,In_68);
and U12 (N_12,In_2,In_392);
and U13 (N_13,In_133,In_113);
nand U14 (N_14,In_289,In_177);
or U15 (N_15,In_474,In_286);
and U16 (N_16,In_189,In_35);
nor U17 (N_17,In_212,In_84);
nand U18 (N_18,In_163,In_231);
or U19 (N_19,In_122,In_103);
nand U20 (N_20,In_479,In_225);
and U21 (N_21,In_313,In_282);
and U22 (N_22,In_215,In_9);
or U23 (N_23,In_134,In_394);
or U24 (N_24,In_273,In_475);
or U25 (N_25,In_403,In_216);
or U26 (N_26,In_281,In_296);
and U27 (N_27,In_252,In_433);
or U28 (N_28,In_331,In_332);
nand U29 (N_29,In_81,In_438);
and U30 (N_30,In_310,In_445);
nand U31 (N_31,In_16,In_376);
and U32 (N_32,In_91,In_429);
or U33 (N_33,In_285,In_21);
or U34 (N_34,In_86,In_434);
nor U35 (N_35,In_211,In_339);
nor U36 (N_36,In_450,In_389);
or U37 (N_37,In_383,In_304);
or U38 (N_38,In_484,In_276);
xnor U39 (N_39,In_347,In_198);
nor U40 (N_40,In_493,In_19);
nand U41 (N_41,In_23,In_353);
nand U42 (N_42,In_184,In_302);
nor U43 (N_43,In_10,In_121);
and U44 (N_44,In_158,In_366);
nor U45 (N_45,In_314,In_204);
or U46 (N_46,In_473,In_238);
or U47 (N_47,In_130,In_49);
nor U48 (N_48,In_195,In_379);
nand U49 (N_49,In_264,In_357);
nor U50 (N_50,In_333,In_325);
nand U51 (N_51,In_48,In_170);
nand U52 (N_52,In_95,In_0);
nand U53 (N_53,In_171,In_254);
nand U54 (N_54,In_378,In_148);
and U55 (N_55,In_241,In_37);
or U56 (N_56,In_463,In_334);
nor U57 (N_57,In_190,In_259);
and U58 (N_58,In_387,In_415);
nor U59 (N_59,In_233,In_355);
nand U60 (N_60,In_70,In_230);
nand U61 (N_61,In_126,In_424);
and U62 (N_62,In_405,In_59);
nand U63 (N_63,In_185,In_476);
nor U64 (N_64,In_160,In_217);
and U65 (N_65,In_365,In_71);
and U66 (N_66,In_123,In_139);
nand U67 (N_67,In_27,In_459);
nor U68 (N_68,In_90,In_391);
and U69 (N_69,In_335,In_294);
or U70 (N_70,In_222,In_77);
nand U71 (N_71,In_316,In_323);
or U72 (N_72,In_181,In_38);
nand U73 (N_73,In_76,In_495);
and U74 (N_74,In_317,In_143);
or U75 (N_75,In_63,In_485);
nor U76 (N_76,In_480,In_109);
or U77 (N_77,In_441,In_440);
or U78 (N_78,In_402,In_174);
and U79 (N_79,In_477,In_371);
or U80 (N_80,In_196,In_102);
nor U81 (N_81,In_50,In_386);
nand U82 (N_82,In_208,In_421);
and U83 (N_83,In_53,In_266);
or U84 (N_84,In_187,In_299);
nor U85 (N_85,In_127,In_85);
and U86 (N_86,In_308,In_228);
nand U87 (N_87,In_437,In_253);
and U88 (N_88,In_446,In_283);
and U89 (N_89,In_428,In_342);
nor U90 (N_90,In_263,In_363);
nand U91 (N_91,In_93,In_239);
or U92 (N_92,In_360,In_256);
and U93 (N_93,In_72,In_277);
nand U94 (N_94,In_489,In_303);
and U95 (N_95,In_351,In_41);
nor U96 (N_96,In_447,In_456);
and U97 (N_97,In_169,In_206);
and U98 (N_98,In_369,In_186);
nand U99 (N_99,In_352,In_247);
and U100 (N_100,In_43,In_145);
or U101 (N_101,In_36,In_255);
nor U102 (N_102,In_461,In_468);
nor U103 (N_103,In_245,In_297);
nand U104 (N_104,In_11,In_292);
nand U105 (N_105,In_374,In_449);
or U106 (N_106,In_393,In_13);
nand U107 (N_107,In_124,In_406);
nor U108 (N_108,In_178,In_167);
nor U109 (N_109,In_452,In_107);
nand U110 (N_110,In_280,In_388);
nor U111 (N_111,In_492,In_201);
xnor U112 (N_112,In_229,In_131);
nand U113 (N_113,In_97,In_390);
or U114 (N_114,In_354,In_442);
and U115 (N_115,In_227,In_141);
and U116 (N_116,In_118,In_218);
or U117 (N_117,In_242,In_115);
and U118 (N_118,In_31,In_269);
and U119 (N_119,In_83,In_165);
or U120 (N_120,In_290,In_411);
or U121 (N_121,In_144,In_111);
and U122 (N_122,In_439,In_309);
nor U123 (N_123,In_375,In_419);
nor U124 (N_124,In_8,In_344);
nor U125 (N_125,In_60,In_47);
or U126 (N_126,In_108,In_359);
or U127 (N_127,In_65,In_75);
and U128 (N_128,In_129,In_96);
or U129 (N_129,In_346,In_451);
nor U130 (N_130,In_12,In_467);
and U131 (N_131,In_175,In_166);
and U132 (N_132,In_116,In_6);
nand U133 (N_133,In_343,In_491);
or U134 (N_134,In_172,In_135);
and U135 (N_135,In_457,In_82);
nand U136 (N_136,In_341,In_322);
and U137 (N_137,In_460,In_425);
nand U138 (N_138,In_396,In_268);
and U139 (N_139,In_194,In_100);
or U140 (N_140,In_223,In_173);
nor U141 (N_141,In_46,In_67);
or U142 (N_142,In_79,In_444);
nor U143 (N_143,In_104,In_338);
nor U144 (N_144,In_18,In_380);
nor U145 (N_145,In_156,In_221);
and U146 (N_146,In_210,In_400);
nand U147 (N_147,In_140,In_328);
nand U148 (N_148,In_407,In_370);
or U149 (N_149,In_398,In_182);
nand U150 (N_150,In_234,In_191);
or U151 (N_151,In_487,In_319);
nand U152 (N_152,In_136,In_284);
nand U153 (N_153,In_337,In_110);
nand U154 (N_154,In_404,In_436);
or U155 (N_155,In_348,In_496);
or U156 (N_156,In_51,In_279);
nor U157 (N_157,In_151,In_397);
or U158 (N_158,In_164,In_33);
or U159 (N_159,In_69,In_265);
nand U160 (N_160,In_57,In_327);
nand U161 (N_161,In_203,In_311);
nand U162 (N_162,In_312,In_270);
nand U163 (N_163,In_205,In_88);
and U164 (N_164,In_197,In_157);
or U165 (N_165,In_329,In_14);
nor U166 (N_166,In_5,In_249);
nand U167 (N_167,In_300,In_200);
or U168 (N_168,In_362,In_443);
and U169 (N_169,In_207,In_262);
nor U170 (N_170,In_154,In_209);
nand U171 (N_171,In_418,In_426);
and U172 (N_172,In_408,In_213);
nand U173 (N_173,In_305,In_431);
and U174 (N_174,In_306,In_120);
nor U175 (N_175,In_3,In_94);
nor U176 (N_176,In_260,In_64);
or U177 (N_177,In_89,In_448);
nand U178 (N_178,In_114,In_488);
or U179 (N_179,In_40,In_330);
nand U180 (N_180,In_192,In_326);
and U181 (N_181,In_432,In_138);
and U182 (N_182,In_202,In_368);
or U183 (N_183,In_364,In_412);
and U184 (N_184,In_482,In_416);
nor U185 (N_185,In_258,In_250);
nor U186 (N_186,In_56,In_410);
nand U187 (N_187,In_153,In_320);
nand U188 (N_188,In_24,In_382);
and U189 (N_189,In_414,In_128);
and U190 (N_190,In_350,In_4);
nand U191 (N_191,In_293,In_373);
nor U192 (N_192,In_427,In_490);
nand U193 (N_193,In_99,In_183);
or U194 (N_194,In_395,In_385);
nor U195 (N_195,In_261,In_498);
nand U196 (N_196,In_92,In_152);
or U197 (N_197,In_66,In_55);
and U198 (N_198,In_232,In_159);
or U199 (N_199,In_377,In_356);
and U200 (N_200,In_499,In_295);
nor U201 (N_201,In_214,In_17);
or U202 (N_202,In_176,In_150);
nor U203 (N_203,In_29,In_472);
or U204 (N_204,In_251,In_125);
nor U205 (N_205,In_453,In_161);
nand U206 (N_206,In_30,In_73);
or U207 (N_207,In_25,In_315);
and U208 (N_208,In_470,In_486);
nor U209 (N_209,In_149,In_288);
nor U210 (N_210,In_399,In_52);
nand U211 (N_211,In_147,In_44);
nand U212 (N_212,In_45,In_236);
nand U213 (N_213,In_455,In_469);
and U214 (N_214,In_22,In_318);
or U215 (N_215,In_275,In_119);
and U216 (N_216,In_381,In_137);
nor U217 (N_217,In_1,In_471);
nor U218 (N_218,In_349,In_243);
nand U219 (N_219,In_74,In_54);
or U220 (N_220,In_226,In_340);
or U221 (N_221,In_155,In_62);
nand U222 (N_222,In_324,In_291);
and U223 (N_223,In_34,In_117);
nor U224 (N_224,In_142,In_106);
nor U225 (N_225,In_78,In_101);
nor U226 (N_226,In_39,In_345);
nor U227 (N_227,In_105,In_199);
or U228 (N_228,In_26,In_257);
and U229 (N_229,In_478,In_28);
nand U230 (N_230,In_358,In_423);
nor U231 (N_231,In_361,In_298);
and U232 (N_232,In_235,In_417);
nor U233 (N_233,In_180,In_112);
and U234 (N_234,In_401,In_465);
and U235 (N_235,In_146,In_246);
and U236 (N_236,In_466,In_58);
and U237 (N_237,In_336,In_307);
and U238 (N_238,In_274,In_224);
nor U239 (N_239,In_179,In_458);
or U240 (N_240,In_7,In_244);
nor U241 (N_241,In_287,In_420);
nor U242 (N_242,In_422,In_367);
and U243 (N_243,In_481,In_483);
nand U244 (N_244,In_162,In_61);
nor U245 (N_245,In_409,In_494);
nand U246 (N_246,In_321,In_372);
nor U247 (N_247,In_278,In_435);
nor U248 (N_248,In_15,In_413);
and U249 (N_249,In_188,In_462);
or U250 (N_250,In_450,In_121);
and U251 (N_251,In_368,In_388);
and U252 (N_252,In_292,In_120);
and U253 (N_253,In_239,In_248);
or U254 (N_254,In_99,In_219);
or U255 (N_255,In_58,In_148);
nand U256 (N_256,In_240,In_299);
and U257 (N_257,In_373,In_130);
or U258 (N_258,In_490,In_261);
or U259 (N_259,In_326,In_203);
nand U260 (N_260,In_481,In_381);
nor U261 (N_261,In_15,In_287);
or U262 (N_262,In_391,In_127);
and U263 (N_263,In_418,In_249);
or U264 (N_264,In_426,In_347);
nand U265 (N_265,In_41,In_201);
nand U266 (N_266,In_279,In_225);
or U267 (N_267,In_315,In_217);
nor U268 (N_268,In_292,In_454);
nor U269 (N_269,In_424,In_119);
or U270 (N_270,In_251,In_236);
nor U271 (N_271,In_30,In_176);
or U272 (N_272,In_54,In_98);
nand U273 (N_273,In_239,In_131);
nor U274 (N_274,In_220,In_30);
nand U275 (N_275,In_312,In_376);
and U276 (N_276,In_379,In_312);
and U277 (N_277,In_390,In_304);
nor U278 (N_278,In_214,In_390);
or U279 (N_279,In_383,In_434);
nand U280 (N_280,In_236,In_343);
nor U281 (N_281,In_418,In_464);
and U282 (N_282,In_144,In_223);
nand U283 (N_283,In_241,In_220);
and U284 (N_284,In_207,In_431);
nand U285 (N_285,In_327,In_485);
nand U286 (N_286,In_54,In_13);
and U287 (N_287,In_155,In_348);
nor U288 (N_288,In_72,In_51);
and U289 (N_289,In_393,In_119);
nand U290 (N_290,In_32,In_367);
nand U291 (N_291,In_238,In_54);
or U292 (N_292,In_261,In_407);
nor U293 (N_293,In_148,In_282);
or U294 (N_294,In_327,In_232);
and U295 (N_295,In_25,In_403);
and U296 (N_296,In_289,In_323);
or U297 (N_297,In_398,In_278);
xnor U298 (N_298,In_457,In_400);
nand U299 (N_299,In_180,In_282);
or U300 (N_300,In_421,In_400);
nor U301 (N_301,In_302,In_487);
nor U302 (N_302,In_286,In_278);
and U303 (N_303,In_362,In_454);
nor U304 (N_304,In_445,In_48);
and U305 (N_305,In_200,In_417);
nand U306 (N_306,In_435,In_22);
or U307 (N_307,In_204,In_107);
nand U308 (N_308,In_125,In_375);
nor U309 (N_309,In_395,In_303);
nor U310 (N_310,In_387,In_329);
nor U311 (N_311,In_472,In_41);
and U312 (N_312,In_208,In_87);
and U313 (N_313,In_200,In_386);
and U314 (N_314,In_36,In_78);
nand U315 (N_315,In_18,In_61);
or U316 (N_316,In_261,In_265);
nand U317 (N_317,In_183,In_486);
nand U318 (N_318,In_466,In_387);
or U319 (N_319,In_208,In_79);
and U320 (N_320,In_255,In_258);
and U321 (N_321,In_126,In_495);
or U322 (N_322,In_351,In_278);
and U323 (N_323,In_492,In_129);
or U324 (N_324,In_194,In_328);
or U325 (N_325,In_191,In_300);
and U326 (N_326,In_32,In_3);
nor U327 (N_327,In_256,In_438);
nand U328 (N_328,In_29,In_367);
nand U329 (N_329,In_418,In_406);
and U330 (N_330,In_384,In_91);
nand U331 (N_331,In_119,In_182);
nand U332 (N_332,In_174,In_146);
or U333 (N_333,In_58,In_160);
nand U334 (N_334,In_478,In_244);
or U335 (N_335,In_327,In_437);
nand U336 (N_336,In_285,In_61);
nor U337 (N_337,In_196,In_142);
nor U338 (N_338,In_235,In_155);
nor U339 (N_339,In_274,In_479);
nand U340 (N_340,In_331,In_293);
and U341 (N_341,In_395,In_147);
or U342 (N_342,In_243,In_444);
nor U343 (N_343,In_486,In_10);
or U344 (N_344,In_247,In_35);
and U345 (N_345,In_437,In_105);
or U346 (N_346,In_188,In_432);
nand U347 (N_347,In_380,In_36);
nand U348 (N_348,In_103,In_377);
nor U349 (N_349,In_331,In_168);
nand U350 (N_350,In_343,In_98);
nand U351 (N_351,In_450,In_128);
nor U352 (N_352,In_308,In_487);
or U353 (N_353,In_153,In_26);
and U354 (N_354,In_335,In_422);
or U355 (N_355,In_337,In_42);
or U356 (N_356,In_321,In_45);
nor U357 (N_357,In_446,In_152);
xor U358 (N_358,In_242,In_405);
nand U359 (N_359,In_101,In_458);
and U360 (N_360,In_362,In_229);
or U361 (N_361,In_165,In_302);
and U362 (N_362,In_207,In_44);
and U363 (N_363,In_110,In_441);
nand U364 (N_364,In_161,In_155);
and U365 (N_365,In_180,In_297);
nand U366 (N_366,In_81,In_146);
and U367 (N_367,In_58,In_74);
nor U368 (N_368,In_355,In_287);
nand U369 (N_369,In_458,In_459);
or U370 (N_370,In_166,In_240);
or U371 (N_371,In_491,In_244);
nand U372 (N_372,In_372,In_404);
and U373 (N_373,In_258,In_431);
and U374 (N_374,In_366,In_389);
nor U375 (N_375,In_478,In_385);
nand U376 (N_376,In_457,In_418);
nand U377 (N_377,In_304,In_229);
nor U378 (N_378,In_331,In_31);
and U379 (N_379,In_48,In_377);
or U380 (N_380,In_235,In_326);
nor U381 (N_381,In_20,In_477);
and U382 (N_382,In_291,In_80);
or U383 (N_383,In_106,In_268);
nor U384 (N_384,In_83,In_406);
nand U385 (N_385,In_285,In_101);
or U386 (N_386,In_313,In_367);
nand U387 (N_387,In_67,In_385);
nand U388 (N_388,In_164,In_280);
nor U389 (N_389,In_434,In_99);
nand U390 (N_390,In_427,In_449);
nor U391 (N_391,In_369,In_43);
nand U392 (N_392,In_170,In_424);
and U393 (N_393,In_463,In_4);
or U394 (N_394,In_365,In_482);
or U395 (N_395,In_77,In_9);
nor U396 (N_396,In_260,In_43);
nor U397 (N_397,In_297,In_97);
nand U398 (N_398,In_8,In_379);
and U399 (N_399,In_96,In_300);
nor U400 (N_400,In_403,In_251);
nor U401 (N_401,In_405,In_245);
nand U402 (N_402,In_426,In_5);
and U403 (N_403,In_245,In_228);
nand U404 (N_404,In_363,In_350);
xnor U405 (N_405,In_348,In_182);
and U406 (N_406,In_18,In_344);
nor U407 (N_407,In_410,In_188);
and U408 (N_408,In_129,In_186);
nor U409 (N_409,In_308,In_474);
or U410 (N_410,In_444,In_450);
and U411 (N_411,In_485,In_232);
nand U412 (N_412,In_180,In_323);
nand U413 (N_413,In_483,In_223);
nor U414 (N_414,In_189,In_431);
nor U415 (N_415,In_264,In_165);
nand U416 (N_416,In_258,In_428);
nand U417 (N_417,In_288,In_485);
nor U418 (N_418,In_369,In_488);
or U419 (N_419,In_384,In_96);
and U420 (N_420,In_330,In_205);
and U421 (N_421,In_414,In_120);
nand U422 (N_422,In_300,In_62);
and U423 (N_423,In_225,In_342);
nand U424 (N_424,In_13,In_132);
or U425 (N_425,In_471,In_282);
and U426 (N_426,In_45,In_114);
or U427 (N_427,In_430,In_256);
nand U428 (N_428,In_289,In_132);
nand U429 (N_429,In_476,In_118);
or U430 (N_430,In_156,In_201);
and U431 (N_431,In_189,In_137);
and U432 (N_432,In_78,In_49);
nor U433 (N_433,In_212,In_145);
nand U434 (N_434,In_214,In_392);
nand U435 (N_435,In_175,In_177);
or U436 (N_436,In_119,In_338);
and U437 (N_437,In_1,In_108);
and U438 (N_438,In_144,In_8);
nor U439 (N_439,In_372,In_398);
nand U440 (N_440,In_274,In_219);
or U441 (N_441,In_48,In_499);
or U442 (N_442,In_470,In_217);
nor U443 (N_443,In_131,In_331);
or U444 (N_444,In_337,In_446);
and U445 (N_445,In_140,In_175);
and U446 (N_446,In_280,In_352);
or U447 (N_447,In_279,In_451);
or U448 (N_448,In_485,In_252);
or U449 (N_449,In_251,In_214);
nor U450 (N_450,In_115,In_361);
and U451 (N_451,In_209,In_185);
nand U452 (N_452,In_75,In_327);
nand U453 (N_453,In_7,In_243);
nor U454 (N_454,In_360,In_114);
and U455 (N_455,In_155,In_325);
or U456 (N_456,In_258,In_459);
or U457 (N_457,In_336,In_106);
or U458 (N_458,In_51,In_242);
and U459 (N_459,In_76,In_452);
or U460 (N_460,In_41,In_464);
and U461 (N_461,In_321,In_407);
nor U462 (N_462,In_321,In_25);
xor U463 (N_463,In_5,In_62);
or U464 (N_464,In_360,In_295);
or U465 (N_465,In_139,In_407);
nor U466 (N_466,In_239,In_394);
or U467 (N_467,In_229,In_225);
and U468 (N_468,In_45,In_312);
nor U469 (N_469,In_65,In_114);
or U470 (N_470,In_39,In_497);
and U471 (N_471,In_411,In_225);
nand U472 (N_472,In_431,In_378);
nand U473 (N_473,In_320,In_151);
nor U474 (N_474,In_62,In_81);
and U475 (N_475,In_215,In_229);
and U476 (N_476,In_345,In_270);
or U477 (N_477,In_286,In_241);
nand U478 (N_478,In_486,In_270);
nand U479 (N_479,In_50,In_437);
and U480 (N_480,In_481,In_428);
nor U481 (N_481,In_135,In_190);
nand U482 (N_482,In_448,In_146);
and U483 (N_483,In_327,In_38);
or U484 (N_484,In_140,In_139);
nor U485 (N_485,In_227,In_253);
nor U486 (N_486,In_268,In_113);
nor U487 (N_487,In_434,In_182);
or U488 (N_488,In_156,In_1);
nand U489 (N_489,In_452,In_326);
nand U490 (N_490,In_292,In_154);
nor U491 (N_491,In_409,In_288);
nor U492 (N_492,In_21,In_53);
or U493 (N_493,In_155,In_97);
nor U494 (N_494,In_346,In_389);
nand U495 (N_495,In_269,In_208);
and U496 (N_496,In_26,In_299);
or U497 (N_497,In_191,In_175);
nand U498 (N_498,In_125,In_462);
or U499 (N_499,In_329,In_431);
nand U500 (N_500,In_98,In_384);
or U501 (N_501,In_151,In_428);
and U502 (N_502,In_201,In_12);
and U503 (N_503,In_161,In_257);
and U504 (N_504,In_248,In_159);
nor U505 (N_505,In_261,In_410);
or U506 (N_506,In_334,In_159);
or U507 (N_507,In_84,In_159);
and U508 (N_508,In_169,In_87);
and U509 (N_509,In_328,In_450);
nand U510 (N_510,In_293,In_283);
or U511 (N_511,In_262,In_405);
and U512 (N_512,In_491,In_199);
and U513 (N_513,In_102,In_446);
xnor U514 (N_514,In_325,In_336);
and U515 (N_515,In_426,In_208);
and U516 (N_516,In_182,In_289);
or U517 (N_517,In_386,In_105);
and U518 (N_518,In_378,In_91);
or U519 (N_519,In_472,In_20);
and U520 (N_520,In_149,In_86);
nand U521 (N_521,In_326,In_379);
and U522 (N_522,In_257,In_119);
and U523 (N_523,In_165,In_361);
or U524 (N_524,In_97,In_417);
or U525 (N_525,In_94,In_172);
nand U526 (N_526,In_465,In_261);
nor U527 (N_527,In_370,In_252);
nor U528 (N_528,In_209,In_159);
nor U529 (N_529,In_51,In_494);
nand U530 (N_530,In_132,In_305);
nor U531 (N_531,In_226,In_434);
nand U532 (N_532,In_444,In_389);
or U533 (N_533,In_255,In_495);
and U534 (N_534,In_291,In_92);
and U535 (N_535,In_149,In_142);
nand U536 (N_536,In_298,In_28);
and U537 (N_537,In_223,In_161);
nor U538 (N_538,In_333,In_277);
or U539 (N_539,In_494,In_169);
or U540 (N_540,In_92,In_439);
nor U541 (N_541,In_463,In_57);
nor U542 (N_542,In_163,In_365);
and U543 (N_543,In_227,In_394);
nor U544 (N_544,In_157,In_227);
or U545 (N_545,In_420,In_3);
nor U546 (N_546,In_250,In_42);
or U547 (N_547,In_397,In_438);
nor U548 (N_548,In_6,In_145);
nor U549 (N_549,In_55,In_154);
nand U550 (N_550,In_341,In_364);
nor U551 (N_551,In_474,In_272);
nor U552 (N_552,In_112,In_287);
nor U553 (N_553,In_70,In_294);
or U554 (N_554,In_286,In_357);
nor U555 (N_555,In_433,In_465);
or U556 (N_556,In_8,In_420);
and U557 (N_557,In_143,In_398);
or U558 (N_558,In_149,In_244);
nand U559 (N_559,In_86,In_172);
nand U560 (N_560,In_104,In_186);
nand U561 (N_561,In_26,In_462);
nor U562 (N_562,In_304,In_130);
xor U563 (N_563,In_426,In_307);
nor U564 (N_564,In_50,In_48);
and U565 (N_565,In_300,In_72);
xnor U566 (N_566,In_239,In_198);
and U567 (N_567,In_264,In_482);
or U568 (N_568,In_120,In_41);
nand U569 (N_569,In_343,In_426);
nand U570 (N_570,In_321,In_196);
and U571 (N_571,In_193,In_474);
nor U572 (N_572,In_262,In_177);
nand U573 (N_573,In_115,In_480);
or U574 (N_574,In_232,In_335);
nor U575 (N_575,In_449,In_288);
and U576 (N_576,In_354,In_422);
nor U577 (N_577,In_475,In_373);
or U578 (N_578,In_379,In_132);
nor U579 (N_579,In_213,In_439);
and U580 (N_580,In_260,In_454);
and U581 (N_581,In_256,In_317);
nor U582 (N_582,In_463,In_379);
or U583 (N_583,In_278,In_41);
and U584 (N_584,In_233,In_250);
nand U585 (N_585,In_402,In_442);
nand U586 (N_586,In_95,In_283);
or U587 (N_587,In_402,In_216);
nor U588 (N_588,In_103,In_22);
nand U589 (N_589,In_75,In_98);
nor U590 (N_590,In_228,In_458);
and U591 (N_591,In_390,In_433);
or U592 (N_592,In_390,In_12);
xor U593 (N_593,In_248,In_483);
or U594 (N_594,In_50,In_337);
or U595 (N_595,In_283,In_64);
or U596 (N_596,In_383,In_73);
nor U597 (N_597,In_340,In_123);
nand U598 (N_598,In_487,In_461);
nor U599 (N_599,In_220,In_327);
or U600 (N_600,N_542,N_269);
nand U601 (N_601,N_107,N_285);
nand U602 (N_602,N_420,N_185);
or U603 (N_603,N_435,N_8);
and U604 (N_604,N_230,N_447);
nor U605 (N_605,N_2,N_385);
nand U606 (N_606,N_471,N_207);
and U607 (N_607,N_540,N_362);
nand U608 (N_608,N_551,N_556);
or U609 (N_609,N_375,N_358);
or U610 (N_610,N_498,N_562);
and U611 (N_611,N_227,N_328);
nor U612 (N_612,N_154,N_316);
and U613 (N_613,N_418,N_265);
or U614 (N_614,N_346,N_325);
nor U615 (N_615,N_522,N_514);
and U616 (N_616,N_436,N_569);
nand U617 (N_617,N_308,N_17);
or U618 (N_618,N_174,N_330);
or U619 (N_619,N_193,N_409);
nand U620 (N_620,N_88,N_527);
nand U621 (N_621,N_511,N_587);
and U622 (N_622,N_20,N_155);
and U623 (N_623,N_481,N_53);
and U624 (N_624,N_243,N_323);
nand U625 (N_625,N_79,N_4);
or U626 (N_626,N_93,N_239);
or U627 (N_627,N_386,N_242);
and U628 (N_628,N_581,N_566);
and U629 (N_629,N_177,N_283);
or U630 (N_630,N_156,N_90);
nor U631 (N_631,N_278,N_163);
or U632 (N_632,N_528,N_279);
or U633 (N_633,N_110,N_77);
and U634 (N_634,N_589,N_191);
nor U635 (N_635,N_403,N_27);
nor U636 (N_636,N_521,N_383);
nand U637 (N_637,N_5,N_422);
nor U638 (N_638,N_455,N_276);
or U639 (N_639,N_164,N_82);
or U640 (N_640,N_106,N_509);
and U641 (N_641,N_580,N_564);
nor U642 (N_642,N_475,N_359);
or U643 (N_643,N_459,N_99);
or U644 (N_644,N_554,N_329);
xnor U645 (N_645,N_439,N_275);
nand U646 (N_646,N_272,N_136);
and U647 (N_647,N_16,N_451);
nor U648 (N_648,N_371,N_264);
nand U649 (N_649,N_273,N_510);
nor U650 (N_650,N_468,N_121);
and U651 (N_651,N_132,N_263);
nand U652 (N_652,N_85,N_51);
nor U653 (N_653,N_573,N_181);
nand U654 (N_654,N_415,N_32);
and U655 (N_655,N_281,N_550);
nand U656 (N_656,N_526,N_476);
or U657 (N_657,N_582,N_496);
and U658 (N_658,N_478,N_280);
nor U659 (N_659,N_513,N_482);
nand U660 (N_660,N_389,N_404);
nand U661 (N_661,N_23,N_421);
nor U662 (N_662,N_341,N_261);
and U663 (N_663,N_55,N_312);
nor U664 (N_664,N_598,N_18);
nor U665 (N_665,N_240,N_424);
nor U666 (N_666,N_547,N_397);
nor U667 (N_667,N_247,N_348);
nor U668 (N_668,N_454,N_552);
or U669 (N_669,N_347,N_224);
and U670 (N_670,N_520,N_259);
and U671 (N_671,N_432,N_390);
or U672 (N_672,N_246,N_299);
and U673 (N_673,N_575,N_370);
and U674 (N_674,N_499,N_277);
nand U675 (N_675,N_119,N_599);
and U676 (N_676,N_146,N_548);
nand U677 (N_677,N_473,N_394);
nor U678 (N_678,N_512,N_203);
and U679 (N_679,N_34,N_402);
nor U680 (N_680,N_14,N_443);
or U681 (N_681,N_382,N_585);
and U682 (N_682,N_104,N_47);
and U683 (N_683,N_166,N_60);
and U684 (N_684,N_298,N_544);
nor U685 (N_685,N_322,N_423);
or U686 (N_686,N_135,N_15);
or U687 (N_687,N_66,N_398);
and U688 (N_688,N_376,N_452);
and U689 (N_689,N_315,N_306);
nand U690 (N_690,N_147,N_480);
nor U691 (N_691,N_0,N_334);
nand U692 (N_692,N_199,N_565);
and U693 (N_693,N_11,N_525);
or U694 (N_694,N_392,N_588);
xor U695 (N_695,N_39,N_568);
and U696 (N_696,N_217,N_180);
or U697 (N_697,N_142,N_595);
or U698 (N_698,N_405,N_364);
nand U699 (N_699,N_251,N_592);
nor U700 (N_700,N_108,N_558);
nor U701 (N_701,N_19,N_50);
nand U702 (N_702,N_296,N_326);
nor U703 (N_703,N_411,N_393);
or U704 (N_704,N_313,N_232);
and U705 (N_705,N_531,N_462);
nand U706 (N_706,N_95,N_293);
nand U707 (N_707,N_342,N_314);
and U708 (N_708,N_360,N_317);
nor U709 (N_709,N_6,N_324);
nand U710 (N_710,N_96,N_294);
and U711 (N_711,N_87,N_363);
xor U712 (N_712,N_225,N_429);
and U713 (N_713,N_152,N_428);
nor U714 (N_714,N_97,N_448);
nor U715 (N_715,N_593,N_42);
and U716 (N_716,N_523,N_101);
nand U717 (N_717,N_33,N_332);
nand U718 (N_718,N_461,N_67);
and U719 (N_719,N_352,N_37);
and U720 (N_720,N_190,N_367);
nor U721 (N_721,N_486,N_361);
or U722 (N_722,N_483,N_41);
nand U723 (N_723,N_305,N_576);
nand U724 (N_724,N_161,N_379);
or U725 (N_725,N_9,N_538);
or U726 (N_726,N_139,N_29);
and U727 (N_727,N_384,N_122);
nand U728 (N_728,N_501,N_216);
nand U729 (N_729,N_274,N_36);
and U730 (N_730,N_258,N_117);
or U731 (N_731,N_145,N_236);
nor U732 (N_732,N_515,N_215);
nand U733 (N_733,N_183,N_128);
nor U734 (N_734,N_453,N_338);
or U735 (N_735,N_380,N_237);
nand U736 (N_736,N_182,N_331);
nand U737 (N_737,N_49,N_65);
nand U738 (N_738,N_124,N_195);
nand U739 (N_739,N_86,N_68);
or U740 (N_740,N_201,N_416);
or U741 (N_741,N_333,N_408);
nand U742 (N_742,N_91,N_123);
and U743 (N_743,N_304,N_282);
or U744 (N_744,N_560,N_268);
nand U745 (N_745,N_433,N_572);
and U746 (N_746,N_151,N_175);
nor U747 (N_747,N_129,N_545);
or U748 (N_748,N_58,N_365);
and U749 (N_749,N_113,N_171);
and U750 (N_750,N_266,N_245);
nand U751 (N_751,N_30,N_488);
nand U752 (N_752,N_255,N_472);
nor U753 (N_753,N_596,N_319);
nor U754 (N_754,N_24,N_426);
nor U755 (N_755,N_143,N_541);
or U756 (N_756,N_44,N_109);
nor U757 (N_757,N_46,N_43);
and U758 (N_758,N_307,N_490);
nor U759 (N_759,N_149,N_45);
or U760 (N_760,N_396,N_343);
nand U761 (N_761,N_536,N_229);
nor U762 (N_762,N_223,N_226);
or U763 (N_763,N_355,N_178);
or U764 (N_764,N_549,N_484);
nor U765 (N_765,N_287,N_489);
nand U766 (N_766,N_208,N_137);
and U767 (N_767,N_374,N_567);
or U768 (N_768,N_546,N_102);
nor U769 (N_769,N_450,N_354);
or U770 (N_770,N_530,N_26);
or U771 (N_771,N_59,N_320);
nor U772 (N_772,N_406,N_284);
nor U773 (N_773,N_431,N_388);
nor U774 (N_774,N_463,N_464);
nor U775 (N_775,N_169,N_395);
nor U776 (N_776,N_532,N_209);
and U777 (N_777,N_500,N_543);
nand U778 (N_778,N_295,N_344);
nor U779 (N_779,N_414,N_114);
nor U780 (N_780,N_465,N_339);
and U781 (N_781,N_413,N_485);
and U782 (N_782,N_434,N_118);
nor U783 (N_783,N_503,N_130);
nor U784 (N_784,N_38,N_184);
nor U785 (N_785,N_148,N_73);
or U786 (N_786,N_368,N_63);
and U787 (N_787,N_577,N_539);
nor U788 (N_788,N_188,N_35);
or U789 (N_789,N_194,N_351);
nor U790 (N_790,N_336,N_52);
and U791 (N_791,N_12,N_92);
or U792 (N_792,N_591,N_494);
nor U793 (N_793,N_250,N_74);
or U794 (N_794,N_477,N_449);
nor U795 (N_795,N_189,N_288);
nand U796 (N_796,N_94,N_83);
and U797 (N_797,N_400,N_196);
nor U798 (N_798,N_357,N_378);
nand U799 (N_799,N_48,N_80);
and U800 (N_800,N_179,N_300);
or U801 (N_801,N_353,N_506);
nand U802 (N_802,N_535,N_310);
nand U803 (N_803,N_583,N_446);
nor U804 (N_804,N_249,N_231);
nand U805 (N_805,N_508,N_559);
and U806 (N_806,N_290,N_492);
nor U807 (N_807,N_377,N_356);
nor U808 (N_808,N_427,N_157);
nand U809 (N_809,N_369,N_241);
or U810 (N_810,N_211,N_441);
and U811 (N_811,N_252,N_248);
or U812 (N_812,N_103,N_141);
nand U813 (N_813,N_238,N_257);
and U814 (N_814,N_518,N_3);
nor U815 (N_815,N_574,N_25);
nor U816 (N_816,N_165,N_235);
or U817 (N_817,N_200,N_98);
and U818 (N_818,N_221,N_302);
nand U819 (N_819,N_271,N_430);
nor U820 (N_820,N_570,N_401);
nand U821 (N_821,N_586,N_366);
or U822 (N_822,N_140,N_407);
nand U823 (N_823,N_505,N_222);
and U824 (N_824,N_254,N_205);
or U825 (N_825,N_210,N_100);
nor U826 (N_826,N_197,N_286);
nor U827 (N_827,N_76,N_474);
and U828 (N_828,N_159,N_438);
and U829 (N_829,N_519,N_127);
nor U830 (N_830,N_318,N_218);
or U831 (N_831,N_469,N_84);
nand U832 (N_832,N_399,N_584);
nor U833 (N_833,N_534,N_69);
nor U834 (N_834,N_138,N_170);
nor U835 (N_835,N_31,N_557);
or U836 (N_836,N_213,N_524);
and U837 (N_837,N_105,N_78);
and U838 (N_838,N_311,N_204);
or U839 (N_839,N_244,N_457);
nor U840 (N_840,N_112,N_131);
nand U841 (N_841,N_187,N_202);
or U842 (N_842,N_21,N_479);
nand U843 (N_843,N_529,N_172);
nand U844 (N_844,N_289,N_168);
or U845 (N_845,N_440,N_228);
nand U846 (N_846,N_444,N_233);
and U847 (N_847,N_57,N_262);
nor U848 (N_848,N_10,N_167);
and U849 (N_849,N_340,N_160);
or U850 (N_850,N_301,N_186);
nor U851 (N_851,N_206,N_7);
nand U852 (N_852,N_192,N_212);
nand U853 (N_853,N_419,N_387);
or U854 (N_854,N_391,N_335);
nor U855 (N_855,N_111,N_350);
or U856 (N_856,N_62,N_253);
and U857 (N_857,N_497,N_516);
nor U858 (N_858,N_412,N_555);
and U859 (N_859,N_327,N_115);
nor U860 (N_860,N_561,N_75);
or U861 (N_861,N_495,N_153);
nor U862 (N_862,N_158,N_144);
or U863 (N_863,N_493,N_309);
or U864 (N_864,N_134,N_219);
or U865 (N_865,N_1,N_502);
nor U866 (N_866,N_597,N_198);
and U867 (N_867,N_456,N_291);
and U868 (N_868,N_40,N_260);
and U869 (N_869,N_491,N_173);
or U870 (N_870,N_89,N_56);
and U871 (N_871,N_533,N_270);
or U872 (N_872,N_64,N_220);
and U873 (N_873,N_571,N_578);
nor U874 (N_874,N_72,N_594);
or U875 (N_875,N_417,N_214);
nand U876 (N_876,N_256,N_553);
and U877 (N_877,N_458,N_297);
and U878 (N_878,N_71,N_321);
or U879 (N_879,N_442,N_517);
nor U880 (N_880,N_460,N_373);
or U881 (N_881,N_116,N_507);
nor U882 (N_882,N_345,N_61);
or U883 (N_883,N_425,N_579);
nor U884 (N_884,N_125,N_70);
nand U885 (N_885,N_133,N_590);
xor U886 (N_886,N_126,N_303);
nand U887 (N_887,N_267,N_504);
nand U888 (N_888,N_13,N_176);
and U889 (N_889,N_337,N_81);
and U890 (N_890,N_234,N_150);
nor U891 (N_891,N_470,N_410);
and U892 (N_892,N_120,N_563);
nor U893 (N_893,N_381,N_349);
or U894 (N_894,N_28,N_54);
nand U895 (N_895,N_537,N_292);
nor U896 (N_896,N_487,N_162);
and U897 (N_897,N_22,N_467);
nand U898 (N_898,N_445,N_437);
and U899 (N_899,N_372,N_466);
and U900 (N_900,N_216,N_530);
nand U901 (N_901,N_188,N_143);
nand U902 (N_902,N_359,N_547);
nand U903 (N_903,N_137,N_390);
nor U904 (N_904,N_238,N_44);
nor U905 (N_905,N_244,N_411);
nand U906 (N_906,N_414,N_591);
or U907 (N_907,N_60,N_397);
nand U908 (N_908,N_121,N_417);
or U909 (N_909,N_594,N_311);
nand U910 (N_910,N_177,N_440);
or U911 (N_911,N_210,N_82);
nand U912 (N_912,N_221,N_0);
and U913 (N_913,N_292,N_429);
and U914 (N_914,N_77,N_347);
nand U915 (N_915,N_158,N_587);
nor U916 (N_916,N_151,N_461);
nor U917 (N_917,N_180,N_500);
and U918 (N_918,N_382,N_470);
or U919 (N_919,N_23,N_154);
nand U920 (N_920,N_399,N_276);
nand U921 (N_921,N_358,N_521);
or U922 (N_922,N_200,N_545);
and U923 (N_923,N_215,N_224);
and U924 (N_924,N_572,N_285);
or U925 (N_925,N_12,N_194);
or U926 (N_926,N_104,N_251);
and U927 (N_927,N_495,N_145);
nand U928 (N_928,N_69,N_50);
or U929 (N_929,N_520,N_323);
nand U930 (N_930,N_484,N_139);
nand U931 (N_931,N_104,N_36);
nor U932 (N_932,N_506,N_137);
nand U933 (N_933,N_100,N_330);
and U934 (N_934,N_596,N_381);
nand U935 (N_935,N_97,N_490);
nor U936 (N_936,N_303,N_553);
and U937 (N_937,N_126,N_259);
or U938 (N_938,N_381,N_26);
and U939 (N_939,N_408,N_596);
nand U940 (N_940,N_141,N_109);
and U941 (N_941,N_238,N_576);
and U942 (N_942,N_146,N_534);
and U943 (N_943,N_551,N_307);
nand U944 (N_944,N_93,N_89);
or U945 (N_945,N_138,N_77);
nor U946 (N_946,N_62,N_93);
or U947 (N_947,N_65,N_415);
nor U948 (N_948,N_502,N_420);
and U949 (N_949,N_536,N_126);
nor U950 (N_950,N_270,N_280);
xor U951 (N_951,N_445,N_138);
nand U952 (N_952,N_133,N_481);
nand U953 (N_953,N_166,N_76);
xor U954 (N_954,N_319,N_17);
nor U955 (N_955,N_501,N_580);
nand U956 (N_956,N_333,N_364);
and U957 (N_957,N_165,N_553);
or U958 (N_958,N_470,N_446);
nor U959 (N_959,N_46,N_193);
nor U960 (N_960,N_206,N_392);
nor U961 (N_961,N_87,N_426);
or U962 (N_962,N_150,N_584);
nor U963 (N_963,N_348,N_494);
nor U964 (N_964,N_433,N_214);
or U965 (N_965,N_205,N_355);
and U966 (N_966,N_582,N_559);
or U967 (N_967,N_31,N_185);
and U968 (N_968,N_40,N_416);
nand U969 (N_969,N_550,N_321);
nand U970 (N_970,N_452,N_108);
nand U971 (N_971,N_229,N_49);
nand U972 (N_972,N_264,N_289);
nor U973 (N_973,N_170,N_456);
or U974 (N_974,N_1,N_410);
and U975 (N_975,N_80,N_97);
or U976 (N_976,N_67,N_415);
and U977 (N_977,N_323,N_193);
nor U978 (N_978,N_548,N_334);
and U979 (N_979,N_15,N_70);
and U980 (N_980,N_537,N_195);
and U981 (N_981,N_339,N_92);
or U982 (N_982,N_175,N_355);
nand U983 (N_983,N_385,N_81);
or U984 (N_984,N_69,N_84);
or U985 (N_985,N_450,N_0);
nor U986 (N_986,N_415,N_347);
or U987 (N_987,N_95,N_485);
and U988 (N_988,N_103,N_460);
or U989 (N_989,N_406,N_119);
nor U990 (N_990,N_71,N_379);
nand U991 (N_991,N_259,N_304);
or U992 (N_992,N_276,N_409);
or U993 (N_993,N_288,N_521);
nor U994 (N_994,N_215,N_227);
nor U995 (N_995,N_555,N_152);
and U996 (N_996,N_104,N_495);
nor U997 (N_997,N_450,N_215);
and U998 (N_998,N_144,N_470);
nand U999 (N_999,N_493,N_383);
nand U1000 (N_1000,N_261,N_506);
or U1001 (N_1001,N_413,N_385);
nor U1002 (N_1002,N_413,N_351);
nand U1003 (N_1003,N_99,N_178);
and U1004 (N_1004,N_302,N_77);
nor U1005 (N_1005,N_495,N_19);
or U1006 (N_1006,N_545,N_18);
and U1007 (N_1007,N_347,N_15);
or U1008 (N_1008,N_325,N_414);
nand U1009 (N_1009,N_528,N_577);
nor U1010 (N_1010,N_203,N_228);
and U1011 (N_1011,N_185,N_451);
and U1012 (N_1012,N_381,N_104);
nand U1013 (N_1013,N_285,N_472);
nand U1014 (N_1014,N_290,N_155);
nor U1015 (N_1015,N_142,N_176);
nor U1016 (N_1016,N_442,N_349);
and U1017 (N_1017,N_50,N_239);
or U1018 (N_1018,N_507,N_295);
nor U1019 (N_1019,N_64,N_185);
or U1020 (N_1020,N_284,N_262);
or U1021 (N_1021,N_122,N_389);
nand U1022 (N_1022,N_384,N_114);
nor U1023 (N_1023,N_344,N_57);
or U1024 (N_1024,N_473,N_323);
nor U1025 (N_1025,N_219,N_296);
or U1026 (N_1026,N_199,N_499);
nor U1027 (N_1027,N_539,N_511);
nand U1028 (N_1028,N_30,N_502);
and U1029 (N_1029,N_206,N_76);
or U1030 (N_1030,N_508,N_216);
nor U1031 (N_1031,N_489,N_372);
nand U1032 (N_1032,N_308,N_206);
nor U1033 (N_1033,N_539,N_515);
and U1034 (N_1034,N_117,N_543);
nand U1035 (N_1035,N_494,N_514);
or U1036 (N_1036,N_351,N_449);
nor U1037 (N_1037,N_286,N_46);
or U1038 (N_1038,N_478,N_486);
nor U1039 (N_1039,N_523,N_128);
nor U1040 (N_1040,N_315,N_182);
nor U1041 (N_1041,N_35,N_128);
nand U1042 (N_1042,N_354,N_81);
or U1043 (N_1043,N_529,N_389);
nor U1044 (N_1044,N_1,N_282);
or U1045 (N_1045,N_546,N_476);
nor U1046 (N_1046,N_497,N_539);
or U1047 (N_1047,N_199,N_130);
nand U1048 (N_1048,N_198,N_191);
nor U1049 (N_1049,N_393,N_210);
nor U1050 (N_1050,N_290,N_470);
or U1051 (N_1051,N_70,N_268);
and U1052 (N_1052,N_563,N_329);
nor U1053 (N_1053,N_277,N_357);
nand U1054 (N_1054,N_402,N_282);
nand U1055 (N_1055,N_215,N_405);
or U1056 (N_1056,N_138,N_504);
nand U1057 (N_1057,N_30,N_291);
or U1058 (N_1058,N_471,N_183);
or U1059 (N_1059,N_493,N_335);
nor U1060 (N_1060,N_263,N_397);
nand U1061 (N_1061,N_161,N_571);
nand U1062 (N_1062,N_273,N_94);
or U1063 (N_1063,N_427,N_593);
nand U1064 (N_1064,N_445,N_469);
nor U1065 (N_1065,N_85,N_289);
nor U1066 (N_1066,N_274,N_31);
xnor U1067 (N_1067,N_479,N_563);
or U1068 (N_1068,N_153,N_382);
or U1069 (N_1069,N_419,N_335);
and U1070 (N_1070,N_407,N_210);
nor U1071 (N_1071,N_518,N_37);
nand U1072 (N_1072,N_359,N_102);
or U1073 (N_1073,N_575,N_442);
or U1074 (N_1074,N_137,N_483);
or U1075 (N_1075,N_77,N_457);
and U1076 (N_1076,N_79,N_433);
and U1077 (N_1077,N_198,N_246);
nand U1078 (N_1078,N_190,N_38);
nand U1079 (N_1079,N_330,N_451);
and U1080 (N_1080,N_385,N_71);
or U1081 (N_1081,N_515,N_397);
or U1082 (N_1082,N_511,N_554);
nand U1083 (N_1083,N_505,N_314);
nor U1084 (N_1084,N_149,N_289);
or U1085 (N_1085,N_481,N_268);
or U1086 (N_1086,N_317,N_126);
or U1087 (N_1087,N_148,N_569);
nor U1088 (N_1088,N_288,N_346);
nand U1089 (N_1089,N_113,N_19);
nand U1090 (N_1090,N_350,N_7);
nand U1091 (N_1091,N_209,N_249);
nand U1092 (N_1092,N_238,N_129);
or U1093 (N_1093,N_338,N_301);
or U1094 (N_1094,N_350,N_190);
and U1095 (N_1095,N_387,N_26);
nand U1096 (N_1096,N_40,N_78);
nand U1097 (N_1097,N_48,N_375);
nand U1098 (N_1098,N_364,N_101);
and U1099 (N_1099,N_143,N_208);
nor U1100 (N_1100,N_544,N_158);
nand U1101 (N_1101,N_113,N_406);
and U1102 (N_1102,N_1,N_536);
nor U1103 (N_1103,N_227,N_585);
nor U1104 (N_1104,N_168,N_212);
nor U1105 (N_1105,N_375,N_202);
nand U1106 (N_1106,N_364,N_491);
and U1107 (N_1107,N_34,N_416);
and U1108 (N_1108,N_238,N_163);
nor U1109 (N_1109,N_217,N_143);
and U1110 (N_1110,N_435,N_59);
nor U1111 (N_1111,N_148,N_561);
nand U1112 (N_1112,N_1,N_532);
or U1113 (N_1113,N_343,N_112);
nor U1114 (N_1114,N_266,N_60);
nor U1115 (N_1115,N_570,N_83);
nand U1116 (N_1116,N_206,N_344);
and U1117 (N_1117,N_591,N_20);
and U1118 (N_1118,N_530,N_205);
or U1119 (N_1119,N_157,N_473);
nand U1120 (N_1120,N_15,N_263);
nand U1121 (N_1121,N_567,N_149);
and U1122 (N_1122,N_158,N_293);
nand U1123 (N_1123,N_463,N_5);
and U1124 (N_1124,N_184,N_146);
nand U1125 (N_1125,N_167,N_324);
or U1126 (N_1126,N_506,N_156);
nor U1127 (N_1127,N_79,N_279);
nand U1128 (N_1128,N_361,N_225);
nand U1129 (N_1129,N_508,N_134);
or U1130 (N_1130,N_223,N_13);
nand U1131 (N_1131,N_188,N_39);
nor U1132 (N_1132,N_520,N_288);
or U1133 (N_1133,N_575,N_6);
or U1134 (N_1134,N_208,N_9);
and U1135 (N_1135,N_90,N_598);
and U1136 (N_1136,N_188,N_15);
nand U1137 (N_1137,N_374,N_287);
or U1138 (N_1138,N_12,N_352);
and U1139 (N_1139,N_521,N_479);
nand U1140 (N_1140,N_542,N_125);
nor U1141 (N_1141,N_189,N_290);
nand U1142 (N_1142,N_480,N_239);
or U1143 (N_1143,N_38,N_536);
or U1144 (N_1144,N_355,N_585);
or U1145 (N_1145,N_276,N_61);
nor U1146 (N_1146,N_272,N_546);
and U1147 (N_1147,N_201,N_548);
nand U1148 (N_1148,N_169,N_276);
nor U1149 (N_1149,N_567,N_477);
nor U1150 (N_1150,N_144,N_572);
nor U1151 (N_1151,N_370,N_56);
and U1152 (N_1152,N_69,N_25);
nand U1153 (N_1153,N_476,N_219);
nor U1154 (N_1154,N_357,N_237);
and U1155 (N_1155,N_488,N_376);
or U1156 (N_1156,N_290,N_585);
nand U1157 (N_1157,N_250,N_414);
xnor U1158 (N_1158,N_579,N_175);
nor U1159 (N_1159,N_454,N_279);
nor U1160 (N_1160,N_28,N_257);
and U1161 (N_1161,N_358,N_508);
nor U1162 (N_1162,N_316,N_73);
nand U1163 (N_1163,N_289,N_415);
nor U1164 (N_1164,N_216,N_302);
and U1165 (N_1165,N_328,N_131);
nor U1166 (N_1166,N_505,N_31);
nor U1167 (N_1167,N_247,N_589);
and U1168 (N_1168,N_122,N_133);
nand U1169 (N_1169,N_128,N_107);
nand U1170 (N_1170,N_71,N_151);
or U1171 (N_1171,N_339,N_560);
nor U1172 (N_1172,N_302,N_279);
and U1173 (N_1173,N_96,N_175);
and U1174 (N_1174,N_588,N_402);
or U1175 (N_1175,N_12,N_588);
nor U1176 (N_1176,N_192,N_260);
or U1177 (N_1177,N_41,N_98);
nand U1178 (N_1178,N_423,N_479);
nor U1179 (N_1179,N_594,N_565);
and U1180 (N_1180,N_267,N_337);
or U1181 (N_1181,N_368,N_503);
nand U1182 (N_1182,N_305,N_101);
and U1183 (N_1183,N_284,N_563);
nor U1184 (N_1184,N_127,N_301);
and U1185 (N_1185,N_551,N_579);
nor U1186 (N_1186,N_197,N_120);
nand U1187 (N_1187,N_60,N_164);
and U1188 (N_1188,N_553,N_76);
nor U1189 (N_1189,N_174,N_123);
xor U1190 (N_1190,N_548,N_544);
nor U1191 (N_1191,N_585,N_321);
nor U1192 (N_1192,N_208,N_523);
and U1193 (N_1193,N_535,N_118);
xor U1194 (N_1194,N_428,N_366);
or U1195 (N_1195,N_255,N_269);
nand U1196 (N_1196,N_65,N_175);
or U1197 (N_1197,N_233,N_557);
or U1198 (N_1198,N_500,N_406);
nand U1199 (N_1199,N_539,N_362);
nand U1200 (N_1200,N_904,N_1030);
and U1201 (N_1201,N_1045,N_1129);
and U1202 (N_1202,N_816,N_844);
and U1203 (N_1203,N_622,N_885);
or U1204 (N_1204,N_800,N_940);
nor U1205 (N_1205,N_912,N_1152);
and U1206 (N_1206,N_714,N_1188);
and U1207 (N_1207,N_719,N_1011);
or U1208 (N_1208,N_664,N_968);
or U1209 (N_1209,N_1070,N_1115);
or U1210 (N_1210,N_626,N_846);
xnor U1211 (N_1211,N_717,N_644);
or U1212 (N_1212,N_1042,N_675);
and U1213 (N_1213,N_750,N_725);
nand U1214 (N_1214,N_1165,N_870);
nand U1215 (N_1215,N_1101,N_1123);
or U1216 (N_1216,N_720,N_908);
and U1217 (N_1217,N_722,N_740);
nand U1218 (N_1218,N_1155,N_753);
xor U1219 (N_1219,N_1046,N_1057);
nand U1220 (N_1220,N_774,N_918);
nor U1221 (N_1221,N_746,N_728);
nor U1222 (N_1222,N_1064,N_647);
and U1223 (N_1223,N_1060,N_701);
or U1224 (N_1224,N_996,N_933);
and U1225 (N_1225,N_919,N_741);
nor U1226 (N_1226,N_1172,N_752);
nor U1227 (N_1227,N_874,N_864);
nand U1228 (N_1228,N_1148,N_1110);
nor U1229 (N_1229,N_624,N_1062);
and U1230 (N_1230,N_687,N_814);
or U1231 (N_1231,N_681,N_869);
nor U1232 (N_1232,N_921,N_602);
or U1233 (N_1233,N_954,N_1161);
nand U1234 (N_1234,N_1008,N_713);
nor U1235 (N_1235,N_1053,N_1178);
or U1236 (N_1236,N_797,N_889);
and U1237 (N_1237,N_603,N_823);
nor U1238 (N_1238,N_1071,N_950);
nand U1239 (N_1239,N_1080,N_997);
or U1240 (N_1240,N_1088,N_831);
nor U1241 (N_1241,N_817,N_1028);
and U1242 (N_1242,N_936,N_1092);
nand U1243 (N_1243,N_977,N_1037);
and U1244 (N_1244,N_916,N_676);
nor U1245 (N_1245,N_821,N_866);
and U1246 (N_1246,N_615,N_994);
nor U1247 (N_1247,N_809,N_1035);
nand U1248 (N_1248,N_613,N_802);
and U1249 (N_1249,N_1009,N_951);
or U1250 (N_1250,N_652,N_839);
nor U1251 (N_1251,N_601,N_1108);
nor U1252 (N_1252,N_875,N_709);
nor U1253 (N_1253,N_989,N_1131);
xor U1254 (N_1254,N_893,N_1091);
nor U1255 (N_1255,N_892,N_653);
nor U1256 (N_1256,N_819,N_944);
nor U1257 (N_1257,N_837,N_779);
or U1258 (N_1258,N_682,N_739);
and U1259 (N_1259,N_804,N_1100);
and U1260 (N_1260,N_641,N_820);
nand U1261 (N_1261,N_833,N_1105);
and U1262 (N_1262,N_1089,N_679);
nand U1263 (N_1263,N_677,N_769);
nand U1264 (N_1264,N_632,N_1170);
or U1265 (N_1265,N_1066,N_790);
nand U1266 (N_1266,N_680,N_957);
nor U1267 (N_1267,N_1177,N_1087);
and U1268 (N_1268,N_886,N_777);
or U1269 (N_1269,N_818,N_668);
nor U1270 (N_1270,N_1039,N_995);
or U1271 (N_1271,N_1114,N_699);
nand U1272 (N_1272,N_964,N_662);
nand U1273 (N_1273,N_948,N_657);
nand U1274 (N_1274,N_648,N_1025);
or U1275 (N_1275,N_993,N_1168);
or U1276 (N_1276,N_1090,N_1140);
nor U1277 (N_1277,N_700,N_862);
and U1278 (N_1278,N_1079,N_941);
nor U1279 (N_1279,N_751,N_857);
nor U1280 (N_1280,N_1196,N_1132);
or U1281 (N_1281,N_1182,N_962);
nand U1282 (N_1282,N_934,N_1199);
and U1283 (N_1283,N_734,N_628);
nand U1284 (N_1284,N_903,N_898);
nand U1285 (N_1285,N_776,N_645);
nor U1286 (N_1286,N_860,N_946);
nand U1287 (N_1287,N_1160,N_929);
or U1288 (N_1288,N_651,N_1052);
or U1289 (N_1289,N_683,N_842);
nor U1290 (N_1290,N_609,N_959);
and U1291 (N_1291,N_983,N_785);
nand U1292 (N_1292,N_704,N_1067);
and U1293 (N_1293,N_1158,N_623);
and U1294 (N_1294,N_1026,N_876);
and U1295 (N_1295,N_963,N_690);
nor U1296 (N_1296,N_883,N_822);
and U1297 (N_1297,N_863,N_735);
nor U1298 (N_1298,N_640,N_1106);
nor U1299 (N_1299,N_770,N_911);
and U1300 (N_1300,N_654,N_1151);
or U1301 (N_1301,N_660,N_806);
or U1302 (N_1302,N_971,N_1063);
and U1303 (N_1303,N_1078,N_1163);
nor U1304 (N_1304,N_881,N_920);
or U1305 (N_1305,N_851,N_1098);
or U1306 (N_1306,N_1197,N_930);
nor U1307 (N_1307,N_656,N_1085);
or U1308 (N_1308,N_708,N_1022);
or U1309 (N_1309,N_991,N_1010);
or U1310 (N_1310,N_824,N_1166);
xnor U1311 (N_1311,N_793,N_917);
nor U1312 (N_1312,N_742,N_784);
nor U1313 (N_1313,N_686,N_754);
or U1314 (N_1314,N_634,N_1176);
nor U1315 (N_1315,N_1013,N_981);
or U1316 (N_1316,N_1107,N_765);
nand U1317 (N_1317,N_1136,N_829);
nor U1318 (N_1318,N_932,N_724);
and U1319 (N_1319,N_1034,N_1184);
nor U1320 (N_1320,N_845,N_812);
nand U1321 (N_1321,N_633,N_1116);
or U1322 (N_1322,N_858,N_1003);
nand U1323 (N_1323,N_772,N_1124);
and U1324 (N_1324,N_703,N_618);
or U1325 (N_1325,N_606,N_1093);
or U1326 (N_1326,N_848,N_763);
and U1327 (N_1327,N_1023,N_1084);
nand U1328 (N_1328,N_1137,N_1156);
and U1329 (N_1329,N_1012,N_672);
nor U1330 (N_1330,N_985,N_879);
or U1331 (N_1331,N_1000,N_878);
and U1332 (N_1332,N_1036,N_861);
and U1333 (N_1333,N_1058,N_961);
nand U1334 (N_1334,N_617,N_955);
or U1335 (N_1335,N_1065,N_853);
or U1336 (N_1336,N_678,N_1109);
nor U1337 (N_1337,N_937,N_1181);
nor U1338 (N_1338,N_1113,N_1146);
and U1339 (N_1339,N_610,N_670);
nor U1340 (N_1340,N_1002,N_1139);
or U1341 (N_1341,N_646,N_958);
or U1342 (N_1342,N_1051,N_859);
nand U1343 (N_1343,N_1024,N_808);
or U1344 (N_1344,N_1006,N_667);
nor U1345 (N_1345,N_674,N_608);
or U1346 (N_1346,N_1167,N_1133);
nor U1347 (N_1347,N_913,N_1171);
nor U1348 (N_1348,N_992,N_636);
nor U1349 (N_1349,N_1150,N_600);
and U1350 (N_1350,N_887,N_786);
nand U1351 (N_1351,N_1019,N_1047);
nor U1352 (N_1352,N_627,N_737);
and U1353 (N_1353,N_1141,N_1118);
and U1354 (N_1354,N_1162,N_673);
or U1355 (N_1355,N_743,N_854);
and U1356 (N_1356,N_909,N_1175);
or U1357 (N_1357,N_738,N_1198);
nand U1358 (N_1358,N_1130,N_745);
nand U1359 (N_1359,N_895,N_1083);
and U1360 (N_1360,N_935,N_1128);
and U1361 (N_1361,N_666,N_1159);
and U1362 (N_1362,N_1169,N_980);
nand U1363 (N_1363,N_787,N_1154);
and U1364 (N_1364,N_1021,N_639);
xor U1365 (N_1365,N_1174,N_947);
nor U1366 (N_1366,N_773,N_1072);
nor U1367 (N_1367,N_693,N_847);
nand U1368 (N_1368,N_972,N_710);
or U1369 (N_1369,N_688,N_924);
and U1370 (N_1370,N_1127,N_791);
nor U1371 (N_1371,N_1195,N_956);
nand U1372 (N_1372,N_852,N_1180);
or U1373 (N_1373,N_1001,N_794);
or U1374 (N_1374,N_1048,N_733);
or U1375 (N_1375,N_642,N_1094);
and U1376 (N_1376,N_755,N_718);
and U1377 (N_1377,N_905,N_1086);
and U1378 (N_1378,N_907,N_1186);
nor U1379 (N_1379,N_1044,N_730);
nand U1380 (N_1380,N_888,N_928);
nand U1381 (N_1381,N_1032,N_1068);
or U1382 (N_1382,N_894,N_960);
or U1383 (N_1383,N_988,N_760);
nor U1384 (N_1384,N_974,N_982);
or U1385 (N_1385,N_984,N_637);
or U1386 (N_1386,N_939,N_605);
and U1387 (N_1387,N_884,N_1027);
or U1388 (N_1388,N_1112,N_1015);
or U1389 (N_1389,N_1157,N_1153);
nand U1390 (N_1390,N_621,N_1031);
or U1391 (N_1391,N_872,N_943);
or U1392 (N_1392,N_1075,N_1143);
or U1393 (N_1393,N_1173,N_849);
and U1394 (N_1394,N_871,N_1193);
xnor U1395 (N_1395,N_635,N_611);
nor U1396 (N_1396,N_914,N_702);
nand U1397 (N_1397,N_1185,N_771);
nand U1398 (N_1398,N_973,N_938);
nand U1399 (N_1399,N_1033,N_783);
and U1400 (N_1400,N_727,N_868);
nand U1401 (N_1401,N_799,N_1061);
nor U1402 (N_1402,N_987,N_807);
nand U1403 (N_1403,N_840,N_828);
nand U1404 (N_1404,N_902,N_759);
and U1405 (N_1405,N_1102,N_1029);
nor U1406 (N_1406,N_761,N_877);
nand U1407 (N_1407,N_625,N_843);
nor U1408 (N_1408,N_744,N_890);
nand U1409 (N_1409,N_665,N_694);
and U1410 (N_1410,N_1004,N_1014);
and U1411 (N_1411,N_975,N_830);
and U1412 (N_1412,N_836,N_855);
or U1413 (N_1413,N_942,N_865);
nor U1414 (N_1414,N_798,N_1103);
and U1415 (N_1415,N_986,N_767);
and U1416 (N_1416,N_827,N_778);
and U1417 (N_1417,N_1142,N_1189);
nor U1418 (N_1418,N_614,N_813);
or U1419 (N_1419,N_1121,N_990);
nor U1420 (N_1420,N_825,N_1111);
nor U1421 (N_1421,N_669,N_923);
and U1422 (N_1422,N_970,N_792);
nor U1423 (N_1423,N_748,N_796);
nand U1424 (N_1424,N_705,N_910);
nor U1425 (N_1425,N_706,N_1179);
or U1426 (N_1426,N_795,N_834);
nor U1427 (N_1427,N_999,N_1095);
and U1428 (N_1428,N_1135,N_1040);
nor U1429 (N_1429,N_1122,N_1077);
and U1430 (N_1430,N_604,N_696);
nor U1431 (N_1431,N_707,N_780);
and U1432 (N_1432,N_1017,N_758);
or U1433 (N_1433,N_922,N_655);
nand U1434 (N_1434,N_1016,N_873);
or U1435 (N_1435,N_906,N_692);
nand U1436 (N_1436,N_965,N_882);
xnor U1437 (N_1437,N_749,N_1099);
nand U1438 (N_1438,N_1069,N_969);
or U1439 (N_1439,N_915,N_768);
nand U1440 (N_1440,N_901,N_1134);
nor U1441 (N_1441,N_1096,N_1081);
nand U1442 (N_1442,N_736,N_966);
nor U1443 (N_1443,N_880,N_1183);
nor U1444 (N_1444,N_619,N_1018);
and U1445 (N_1445,N_711,N_1117);
nand U1446 (N_1446,N_1138,N_630);
nand U1447 (N_1447,N_1145,N_867);
nand U1448 (N_1448,N_762,N_1076);
or U1449 (N_1449,N_659,N_649);
nand U1450 (N_1450,N_1149,N_1050);
nand U1451 (N_1451,N_689,N_756);
and U1452 (N_1452,N_732,N_1194);
or U1453 (N_1453,N_1074,N_1104);
nand U1454 (N_1454,N_897,N_695);
or U1455 (N_1455,N_967,N_927);
or U1456 (N_1456,N_1073,N_712);
xnor U1457 (N_1457,N_1038,N_1056);
nand U1458 (N_1458,N_926,N_826);
or U1459 (N_1459,N_1059,N_729);
nor U1460 (N_1460,N_978,N_684);
and U1461 (N_1461,N_841,N_1055);
nor U1462 (N_1462,N_976,N_715);
or U1463 (N_1463,N_764,N_661);
or U1464 (N_1464,N_1126,N_803);
and U1465 (N_1465,N_1097,N_896);
or U1466 (N_1466,N_629,N_616);
nor U1467 (N_1467,N_832,N_952);
nor U1468 (N_1468,N_945,N_731);
and U1469 (N_1469,N_1119,N_1020);
or U1470 (N_1470,N_638,N_810);
nand U1471 (N_1471,N_723,N_698);
and U1472 (N_1472,N_850,N_721);
nand U1473 (N_1473,N_1164,N_620);
nand U1474 (N_1474,N_757,N_979);
nand U1475 (N_1475,N_1192,N_716);
nand U1476 (N_1476,N_726,N_607);
and U1477 (N_1477,N_1120,N_1144);
nor U1478 (N_1478,N_1082,N_811);
and U1479 (N_1479,N_1049,N_856);
nand U1480 (N_1480,N_998,N_815);
or U1481 (N_1481,N_1007,N_1191);
nand U1482 (N_1482,N_781,N_1054);
and U1483 (N_1483,N_691,N_835);
nand U1484 (N_1484,N_891,N_1005);
nor U1485 (N_1485,N_663,N_900);
nand U1486 (N_1486,N_671,N_925);
and U1487 (N_1487,N_1187,N_801);
nand U1488 (N_1488,N_899,N_788);
nor U1489 (N_1489,N_953,N_631);
or U1490 (N_1490,N_643,N_1041);
and U1491 (N_1491,N_1147,N_685);
nor U1492 (N_1492,N_612,N_1190);
nor U1493 (N_1493,N_658,N_697);
nand U1494 (N_1494,N_650,N_931);
nor U1495 (N_1495,N_1125,N_805);
nor U1496 (N_1496,N_1043,N_838);
and U1497 (N_1497,N_949,N_789);
nor U1498 (N_1498,N_747,N_782);
nand U1499 (N_1499,N_766,N_775);
nand U1500 (N_1500,N_1093,N_937);
or U1501 (N_1501,N_754,N_704);
or U1502 (N_1502,N_1196,N_1136);
or U1503 (N_1503,N_964,N_945);
nor U1504 (N_1504,N_1180,N_665);
and U1505 (N_1505,N_1160,N_877);
nor U1506 (N_1506,N_682,N_772);
nor U1507 (N_1507,N_1089,N_1083);
nor U1508 (N_1508,N_1186,N_846);
or U1509 (N_1509,N_1025,N_842);
and U1510 (N_1510,N_1165,N_784);
nand U1511 (N_1511,N_966,N_770);
and U1512 (N_1512,N_827,N_955);
nor U1513 (N_1513,N_1002,N_1158);
or U1514 (N_1514,N_609,N_729);
or U1515 (N_1515,N_1041,N_1145);
and U1516 (N_1516,N_1012,N_820);
and U1517 (N_1517,N_740,N_703);
or U1518 (N_1518,N_1176,N_601);
and U1519 (N_1519,N_1172,N_820);
nor U1520 (N_1520,N_1180,N_1138);
and U1521 (N_1521,N_1163,N_1027);
nand U1522 (N_1522,N_1106,N_956);
nor U1523 (N_1523,N_834,N_835);
nor U1524 (N_1524,N_806,N_1015);
nor U1525 (N_1525,N_1051,N_929);
nand U1526 (N_1526,N_685,N_772);
or U1527 (N_1527,N_1168,N_916);
or U1528 (N_1528,N_1022,N_852);
nand U1529 (N_1529,N_821,N_639);
nand U1530 (N_1530,N_982,N_819);
nor U1531 (N_1531,N_1076,N_621);
or U1532 (N_1532,N_1140,N_837);
and U1533 (N_1533,N_1014,N_1112);
xor U1534 (N_1534,N_1094,N_747);
nand U1535 (N_1535,N_1052,N_922);
nand U1536 (N_1536,N_696,N_752);
and U1537 (N_1537,N_932,N_692);
nand U1538 (N_1538,N_669,N_797);
or U1539 (N_1539,N_1082,N_671);
nand U1540 (N_1540,N_1175,N_1119);
nand U1541 (N_1541,N_1120,N_1100);
or U1542 (N_1542,N_1098,N_1064);
nand U1543 (N_1543,N_674,N_682);
and U1544 (N_1544,N_821,N_607);
nand U1545 (N_1545,N_1054,N_702);
nor U1546 (N_1546,N_1171,N_867);
or U1547 (N_1547,N_844,N_805);
nand U1548 (N_1548,N_1059,N_801);
and U1549 (N_1549,N_807,N_676);
nand U1550 (N_1550,N_726,N_711);
or U1551 (N_1551,N_606,N_1083);
nor U1552 (N_1552,N_773,N_1199);
or U1553 (N_1553,N_1181,N_911);
nand U1554 (N_1554,N_994,N_1036);
nand U1555 (N_1555,N_760,N_1037);
nand U1556 (N_1556,N_758,N_606);
nand U1557 (N_1557,N_667,N_891);
and U1558 (N_1558,N_1114,N_1009);
and U1559 (N_1559,N_972,N_780);
nor U1560 (N_1560,N_1008,N_1049);
and U1561 (N_1561,N_1044,N_688);
nand U1562 (N_1562,N_1159,N_864);
nand U1563 (N_1563,N_825,N_1007);
or U1564 (N_1564,N_705,N_688);
xnor U1565 (N_1565,N_1179,N_1170);
or U1566 (N_1566,N_1057,N_974);
nand U1567 (N_1567,N_1035,N_1117);
nor U1568 (N_1568,N_717,N_608);
nor U1569 (N_1569,N_1027,N_1045);
and U1570 (N_1570,N_1084,N_1098);
nand U1571 (N_1571,N_858,N_628);
nand U1572 (N_1572,N_1192,N_776);
nand U1573 (N_1573,N_1103,N_1183);
or U1574 (N_1574,N_1025,N_732);
nand U1575 (N_1575,N_614,N_940);
and U1576 (N_1576,N_938,N_767);
and U1577 (N_1577,N_929,N_1116);
xnor U1578 (N_1578,N_1018,N_867);
nor U1579 (N_1579,N_645,N_723);
nand U1580 (N_1580,N_1095,N_1057);
or U1581 (N_1581,N_1027,N_1010);
and U1582 (N_1582,N_1127,N_873);
and U1583 (N_1583,N_671,N_1182);
nor U1584 (N_1584,N_824,N_905);
and U1585 (N_1585,N_859,N_879);
nand U1586 (N_1586,N_923,N_632);
or U1587 (N_1587,N_893,N_986);
nor U1588 (N_1588,N_769,N_731);
or U1589 (N_1589,N_1129,N_1128);
nand U1590 (N_1590,N_824,N_1179);
nor U1591 (N_1591,N_780,N_720);
and U1592 (N_1592,N_1002,N_1093);
nor U1593 (N_1593,N_667,N_947);
and U1594 (N_1594,N_1062,N_1009);
and U1595 (N_1595,N_1061,N_974);
nand U1596 (N_1596,N_891,N_781);
nand U1597 (N_1597,N_812,N_877);
or U1598 (N_1598,N_1174,N_1119);
and U1599 (N_1599,N_884,N_1078);
nor U1600 (N_1600,N_922,N_1143);
or U1601 (N_1601,N_635,N_1070);
or U1602 (N_1602,N_808,N_944);
or U1603 (N_1603,N_611,N_710);
nor U1604 (N_1604,N_848,N_952);
and U1605 (N_1605,N_1072,N_754);
or U1606 (N_1606,N_969,N_606);
or U1607 (N_1607,N_973,N_1046);
nor U1608 (N_1608,N_783,N_790);
nor U1609 (N_1609,N_748,N_1042);
nand U1610 (N_1610,N_1040,N_694);
nand U1611 (N_1611,N_994,N_956);
and U1612 (N_1612,N_748,N_1164);
and U1613 (N_1613,N_731,N_874);
nor U1614 (N_1614,N_853,N_886);
and U1615 (N_1615,N_856,N_859);
nand U1616 (N_1616,N_1007,N_1176);
nand U1617 (N_1617,N_659,N_946);
nor U1618 (N_1618,N_844,N_1199);
nor U1619 (N_1619,N_699,N_724);
nand U1620 (N_1620,N_745,N_883);
and U1621 (N_1621,N_671,N_883);
nand U1622 (N_1622,N_895,N_1122);
nand U1623 (N_1623,N_1047,N_885);
or U1624 (N_1624,N_858,N_1142);
nor U1625 (N_1625,N_1058,N_1124);
nand U1626 (N_1626,N_1084,N_1053);
nor U1627 (N_1627,N_1173,N_897);
nand U1628 (N_1628,N_759,N_922);
nor U1629 (N_1629,N_714,N_775);
and U1630 (N_1630,N_789,N_1093);
or U1631 (N_1631,N_908,N_1063);
nor U1632 (N_1632,N_744,N_696);
nand U1633 (N_1633,N_818,N_1195);
nand U1634 (N_1634,N_720,N_1126);
nand U1635 (N_1635,N_1177,N_769);
and U1636 (N_1636,N_816,N_994);
nand U1637 (N_1637,N_706,N_883);
and U1638 (N_1638,N_1139,N_1008);
or U1639 (N_1639,N_909,N_652);
or U1640 (N_1640,N_624,N_1011);
nor U1641 (N_1641,N_1137,N_646);
nand U1642 (N_1642,N_841,N_980);
nand U1643 (N_1643,N_919,N_927);
or U1644 (N_1644,N_891,N_1080);
and U1645 (N_1645,N_640,N_987);
and U1646 (N_1646,N_1170,N_618);
nand U1647 (N_1647,N_988,N_1199);
nor U1648 (N_1648,N_1143,N_850);
nand U1649 (N_1649,N_1145,N_1093);
or U1650 (N_1650,N_944,N_678);
nand U1651 (N_1651,N_1051,N_1092);
nor U1652 (N_1652,N_725,N_884);
or U1653 (N_1653,N_1148,N_695);
nor U1654 (N_1654,N_926,N_644);
nand U1655 (N_1655,N_665,N_1135);
and U1656 (N_1656,N_735,N_1169);
xnor U1657 (N_1657,N_1050,N_1032);
nand U1658 (N_1658,N_732,N_721);
nor U1659 (N_1659,N_744,N_896);
or U1660 (N_1660,N_1184,N_653);
nand U1661 (N_1661,N_1037,N_697);
nand U1662 (N_1662,N_1054,N_970);
or U1663 (N_1663,N_629,N_1199);
xor U1664 (N_1664,N_917,N_823);
nand U1665 (N_1665,N_1046,N_1109);
nor U1666 (N_1666,N_759,N_829);
nand U1667 (N_1667,N_751,N_1035);
or U1668 (N_1668,N_771,N_869);
and U1669 (N_1669,N_718,N_601);
and U1670 (N_1670,N_769,N_763);
nand U1671 (N_1671,N_869,N_1155);
or U1672 (N_1672,N_765,N_1141);
and U1673 (N_1673,N_1114,N_855);
and U1674 (N_1674,N_610,N_775);
and U1675 (N_1675,N_756,N_696);
nor U1676 (N_1676,N_786,N_855);
and U1677 (N_1677,N_707,N_774);
nor U1678 (N_1678,N_1160,N_1093);
nor U1679 (N_1679,N_643,N_1140);
or U1680 (N_1680,N_1065,N_966);
or U1681 (N_1681,N_943,N_974);
and U1682 (N_1682,N_913,N_803);
nor U1683 (N_1683,N_990,N_949);
or U1684 (N_1684,N_685,N_1005);
or U1685 (N_1685,N_898,N_657);
nand U1686 (N_1686,N_755,N_993);
nor U1687 (N_1687,N_1049,N_660);
or U1688 (N_1688,N_822,N_1072);
nor U1689 (N_1689,N_747,N_887);
nor U1690 (N_1690,N_1178,N_785);
nand U1691 (N_1691,N_982,N_796);
nand U1692 (N_1692,N_872,N_833);
and U1693 (N_1693,N_1179,N_876);
and U1694 (N_1694,N_1015,N_747);
or U1695 (N_1695,N_959,N_868);
or U1696 (N_1696,N_786,N_997);
nand U1697 (N_1697,N_920,N_1137);
and U1698 (N_1698,N_1104,N_796);
nand U1699 (N_1699,N_1151,N_834);
or U1700 (N_1700,N_972,N_1021);
or U1701 (N_1701,N_1052,N_783);
nor U1702 (N_1702,N_1160,N_1075);
or U1703 (N_1703,N_1015,N_954);
and U1704 (N_1704,N_844,N_789);
nor U1705 (N_1705,N_831,N_821);
and U1706 (N_1706,N_752,N_1016);
nor U1707 (N_1707,N_1039,N_646);
or U1708 (N_1708,N_827,N_1048);
nor U1709 (N_1709,N_800,N_721);
nand U1710 (N_1710,N_1135,N_720);
nand U1711 (N_1711,N_801,N_757);
and U1712 (N_1712,N_860,N_921);
nor U1713 (N_1713,N_656,N_949);
nor U1714 (N_1714,N_885,N_1134);
nand U1715 (N_1715,N_873,N_970);
nand U1716 (N_1716,N_676,N_914);
or U1717 (N_1717,N_677,N_963);
or U1718 (N_1718,N_744,N_974);
and U1719 (N_1719,N_959,N_1003);
or U1720 (N_1720,N_839,N_1116);
or U1721 (N_1721,N_961,N_812);
nand U1722 (N_1722,N_623,N_1091);
nand U1723 (N_1723,N_683,N_717);
or U1724 (N_1724,N_806,N_847);
and U1725 (N_1725,N_755,N_680);
nor U1726 (N_1726,N_709,N_1008);
or U1727 (N_1727,N_969,N_619);
or U1728 (N_1728,N_1159,N_898);
nand U1729 (N_1729,N_986,N_740);
nand U1730 (N_1730,N_1020,N_912);
nor U1731 (N_1731,N_1198,N_626);
and U1732 (N_1732,N_666,N_847);
or U1733 (N_1733,N_796,N_916);
or U1734 (N_1734,N_1077,N_915);
or U1735 (N_1735,N_694,N_980);
or U1736 (N_1736,N_619,N_1146);
and U1737 (N_1737,N_682,N_614);
nand U1738 (N_1738,N_950,N_688);
nand U1739 (N_1739,N_1090,N_745);
or U1740 (N_1740,N_864,N_899);
nor U1741 (N_1741,N_920,N_840);
nand U1742 (N_1742,N_1019,N_692);
and U1743 (N_1743,N_788,N_1100);
or U1744 (N_1744,N_818,N_983);
nor U1745 (N_1745,N_883,N_1114);
nand U1746 (N_1746,N_1194,N_723);
and U1747 (N_1747,N_1164,N_766);
nand U1748 (N_1748,N_1034,N_609);
and U1749 (N_1749,N_1146,N_789);
or U1750 (N_1750,N_965,N_989);
nor U1751 (N_1751,N_665,N_990);
nor U1752 (N_1752,N_786,N_1045);
nor U1753 (N_1753,N_631,N_622);
nand U1754 (N_1754,N_647,N_676);
nor U1755 (N_1755,N_812,N_999);
nand U1756 (N_1756,N_1157,N_1056);
xnor U1757 (N_1757,N_795,N_918);
nor U1758 (N_1758,N_676,N_1089);
xnor U1759 (N_1759,N_781,N_805);
or U1760 (N_1760,N_848,N_907);
or U1761 (N_1761,N_739,N_606);
or U1762 (N_1762,N_962,N_1098);
nor U1763 (N_1763,N_1173,N_1092);
nand U1764 (N_1764,N_721,N_750);
and U1765 (N_1765,N_1139,N_1015);
or U1766 (N_1766,N_673,N_1047);
or U1767 (N_1767,N_936,N_878);
nand U1768 (N_1768,N_666,N_855);
xnor U1769 (N_1769,N_1082,N_751);
or U1770 (N_1770,N_816,N_843);
or U1771 (N_1771,N_1087,N_1181);
and U1772 (N_1772,N_926,N_699);
and U1773 (N_1773,N_675,N_782);
and U1774 (N_1774,N_849,N_926);
or U1775 (N_1775,N_1025,N_948);
or U1776 (N_1776,N_724,N_810);
nand U1777 (N_1777,N_1115,N_716);
nand U1778 (N_1778,N_830,N_874);
or U1779 (N_1779,N_1023,N_716);
or U1780 (N_1780,N_864,N_1000);
nor U1781 (N_1781,N_706,N_1061);
or U1782 (N_1782,N_955,N_927);
or U1783 (N_1783,N_615,N_892);
nor U1784 (N_1784,N_909,N_1086);
or U1785 (N_1785,N_690,N_670);
and U1786 (N_1786,N_994,N_1176);
and U1787 (N_1787,N_687,N_730);
and U1788 (N_1788,N_814,N_870);
and U1789 (N_1789,N_755,N_963);
nand U1790 (N_1790,N_1064,N_899);
nand U1791 (N_1791,N_1181,N_989);
and U1792 (N_1792,N_1109,N_740);
or U1793 (N_1793,N_1095,N_749);
or U1794 (N_1794,N_1155,N_1105);
and U1795 (N_1795,N_954,N_1156);
nor U1796 (N_1796,N_839,N_996);
nor U1797 (N_1797,N_965,N_639);
nor U1798 (N_1798,N_865,N_834);
or U1799 (N_1799,N_683,N_878);
or U1800 (N_1800,N_1721,N_1406);
or U1801 (N_1801,N_1777,N_1476);
xnor U1802 (N_1802,N_1696,N_1401);
or U1803 (N_1803,N_1652,N_1384);
nand U1804 (N_1804,N_1786,N_1684);
and U1805 (N_1805,N_1290,N_1248);
and U1806 (N_1806,N_1782,N_1278);
and U1807 (N_1807,N_1667,N_1277);
or U1808 (N_1808,N_1269,N_1628);
nand U1809 (N_1809,N_1623,N_1718);
nor U1810 (N_1810,N_1456,N_1250);
and U1811 (N_1811,N_1375,N_1439);
and U1812 (N_1812,N_1580,N_1351);
nand U1813 (N_1813,N_1311,N_1585);
nand U1814 (N_1814,N_1722,N_1391);
and U1815 (N_1815,N_1230,N_1366);
and U1816 (N_1816,N_1238,N_1745);
or U1817 (N_1817,N_1335,N_1581);
nand U1818 (N_1818,N_1743,N_1697);
or U1819 (N_1819,N_1686,N_1307);
nor U1820 (N_1820,N_1685,N_1502);
nor U1821 (N_1821,N_1409,N_1261);
and U1822 (N_1822,N_1603,N_1668);
nand U1823 (N_1823,N_1450,N_1654);
nand U1824 (N_1824,N_1299,N_1280);
nand U1825 (N_1825,N_1732,N_1472);
nor U1826 (N_1826,N_1424,N_1267);
or U1827 (N_1827,N_1566,N_1759);
and U1828 (N_1828,N_1344,N_1320);
or U1829 (N_1829,N_1594,N_1694);
or U1830 (N_1830,N_1655,N_1631);
nand U1831 (N_1831,N_1239,N_1332);
nand U1832 (N_1832,N_1701,N_1610);
nand U1833 (N_1833,N_1491,N_1553);
and U1834 (N_1834,N_1474,N_1372);
nand U1835 (N_1835,N_1323,N_1303);
and U1836 (N_1836,N_1301,N_1708);
nor U1837 (N_1837,N_1750,N_1640);
and U1838 (N_1838,N_1659,N_1534);
or U1839 (N_1839,N_1243,N_1634);
nand U1840 (N_1840,N_1602,N_1369);
xor U1841 (N_1841,N_1312,N_1798);
and U1842 (N_1842,N_1785,N_1526);
nor U1843 (N_1843,N_1495,N_1263);
and U1844 (N_1844,N_1285,N_1377);
nor U1845 (N_1845,N_1609,N_1579);
nor U1846 (N_1846,N_1512,N_1264);
nand U1847 (N_1847,N_1359,N_1682);
or U1848 (N_1848,N_1229,N_1796);
nor U1849 (N_1849,N_1711,N_1547);
and U1850 (N_1850,N_1511,N_1317);
and U1851 (N_1851,N_1717,N_1309);
nor U1852 (N_1852,N_1557,N_1560);
and U1853 (N_1853,N_1220,N_1614);
nand U1854 (N_1854,N_1251,N_1225);
and U1855 (N_1855,N_1582,N_1712);
nand U1856 (N_1856,N_1328,N_1588);
and U1857 (N_1857,N_1428,N_1381);
nor U1858 (N_1858,N_1608,N_1630);
nor U1859 (N_1859,N_1574,N_1411);
or U1860 (N_1860,N_1425,N_1367);
or U1861 (N_1861,N_1447,N_1720);
nor U1862 (N_1862,N_1613,N_1397);
nand U1863 (N_1863,N_1200,N_1510);
nand U1864 (N_1864,N_1396,N_1597);
or U1865 (N_1865,N_1596,N_1246);
or U1866 (N_1866,N_1648,N_1653);
and U1867 (N_1867,N_1629,N_1212);
or U1868 (N_1868,N_1748,N_1679);
nand U1869 (N_1869,N_1733,N_1542);
or U1870 (N_1870,N_1504,N_1787);
and U1871 (N_1871,N_1780,N_1458);
nand U1872 (N_1872,N_1343,N_1237);
and U1873 (N_1873,N_1747,N_1546);
nand U1874 (N_1874,N_1778,N_1578);
and U1875 (N_1875,N_1434,N_1755);
nand U1876 (N_1876,N_1600,N_1673);
nor U1877 (N_1877,N_1693,N_1329);
nor U1878 (N_1878,N_1339,N_1656);
and U1879 (N_1879,N_1651,N_1440);
nand U1880 (N_1880,N_1775,N_1689);
or U1881 (N_1881,N_1501,N_1255);
or U1882 (N_1882,N_1625,N_1645);
nor U1883 (N_1883,N_1492,N_1498);
nor U1884 (N_1884,N_1342,N_1444);
nor U1885 (N_1885,N_1429,N_1486);
nor U1886 (N_1886,N_1292,N_1541);
or U1887 (N_1887,N_1616,N_1227);
or U1888 (N_1888,N_1618,N_1621);
or U1889 (N_1889,N_1347,N_1714);
nand U1890 (N_1890,N_1789,N_1410);
nor U1891 (N_1891,N_1567,N_1589);
nand U1892 (N_1892,N_1454,N_1724);
nand U1893 (N_1893,N_1738,N_1418);
or U1894 (N_1894,N_1240,N_1723);
or U1895 (N_1895,N_1296,N_1540);
nor U1896 (N_1896,N_1350,N_1284);
nor U1897 (N_1897,N_1306,N_1494);
nor U1898 (N_1898,N_1468,N_1270);
or U1899 (N_1899,N_1487,N_1515);
and U1900 (N_1900,N_1644,N_1352);
nor U1901 (N_1901,N_1680,N_1478);
or U1902 (N_1902,N_1271,N_1330);
nand U1903 (N_1903,N_1368,N_1247);
and U1904 (N_1904,N_1617,N_1314);
and U1905 (N_1905,N_1422,N_1666);
nand U1906 (N_1906,N_1399,N_1436);
nor U1907 (N_1907,N_1234,N_1346);
or U1908 (N_1908,N_1703,N_1531);
or U1909 (N_1909,N_1716,N_1216);
nor U1910 (N_1910,N_1683,N_1470);
and U1911 (N_1911,N_1387,N_1641);
xor U1912 (N_1912,N_1695,N_1275);
and U1913 (N_1913,N_1516,N_1606);
and U1914 (N_1914,N_1681,N_1767);
and U1915 (N_1915,N_1272,N_1287);
or U1916 (N_1916,N_1266,N_1671);
nand U1917 (N_1917,N_1336,N_1773);
and U1918 (N_1918,N_1662,N_1479);
nor U1919 (N_1919,N_1658,N_1788);
and U1920 (N_1920,N_1448,N_1799);
or U1921 (N_1921,N_1437,N_1783);
nor U1922 (N_1922,N_1611,N_1493);
nand U1923 (N_1923,N_1754,N_1242);
nand U1924 (N_1924,N_1626,N_1416);
and U1925 (N_1925,N_1549,N_1647);
nor U1926 (N_1926,N_1633,N_1518);
nand U1927 (N_1927,N_1371,N_1488);
and U1928 (N_1928,N_1550,N_1217);
and U1929 (N_1929,N_1457,N_1338);
or U1930 (N_1930,N_1548,N_1244);
nor U1931 (N_1931,N_1219,N_1643);
or U1932 (N_1932,N_1500,N_1354);
or U1933 (N_1933,N_1739,N_1279);
nand U1934 (N_1934,N_1768,N_1514);
xnor U1935 (N_1935,N_1706,N_1254);
nor U1936 (N_1936,N_1453,N_1532);
nor U1937 (N_1937,N_1459,N_1304);
nand U1938 (N_1938,N_1583,N_1252);
xnor U1939 (N_1939,N_1365,N_1333);
and U1940 (N_1940,N_1794,N_1520);
nor U1941 (N_1941,N_1402,N_1398);
nor U1942 (N_1942,N_1489,N_1624);
and U1943 (N_1943,N_1524,N_1283);
or U1944 (N_1944,N_1598,N_1506);
nand U1945 (N_1945,N_1664,N_1587);
nand U1946 (N_1946,N_1642,N_1360);
nor U1947 (N_1947,N_1779,N_1421);
or U1948 (N_1948,N_1528,N_1483);
and U1949 (N_1949,N_1282,N_1407);
and U1950 (N_1950,N_1509,N_1313);
and U1951 (N_1951,N_1210,N_1438);
or U1952 (N_1952,N_1576,N_1207);
nand U1953 (N_1953,N_1417,N_1527);
nand U1954 (N_1954,N_1341,N_1223);
nor U1955 (N_1955,N_1505,N_1233);
or U1956 (N_1956,N_1445,N_1568);
and U1957 (N_1957,N_1657,N_1393);
nand U1958 (N_1958,N_1321,N_1355);
and U1959 (N_1959,N_1373,N_1379);
nand U1960 (N_1960,N_1736,N_1559);
and U1961 (N_1961,N_1562,N_1432);
nand U1962 (N_1962,N_1357,N_1419);
nor U1963 (N_1963,N_1358,N_1334);
or U1964 (N_1964,N_1394,N_1431);
or U1965 (N_1965,N_1646,N_1764);
nor U1966 (N_1966,N_1464,N_1774);
nor U1967 (N_1967,N_1310,N_1403);
nand U1968 (N_1968,N_1563,N_1678);
nand U1969 (N_1969,N_1740,N_1363);
nor U1970 (N_1970,N_1412,N_1276);
or U1971 (N_1971,N_1291,N_1529);
or U1972 (N_1972,N_1298,N_1413);
nand U1973 (N_1973,N_1691,N_1762);
and U1974 (N_1974,N_1319,N_1776);
nor U1975 (N_1975,N_1218,N_1771);
or U1976 (N_1976,N_1496,N_1215);
or U1977 (N_1977,N_1388,N_1386);
nor U1978 (N_1978,N_1632,N_1665);
nand U1979 (N_1979,N_1537,N_1649);
nand U1980 (N_1980,N_1591,N_1620);
nand U1981 (N_1981,N_1224,N_1535);
or U1982 (N_1982,N_1258,N_1326);
and U1983 (N_1983,N_1715,N_1460);
or U1984 (N_1984,N_1622,N_1615);
nor U1985 (N_1985,N_1465,N_1577);
nor U1986 (N_1986,N_1390,N_1499);
or U1987 (N_1987,N_1385,N_1426);
nand U1988 (N_1988,N_1353,N_1348);
nand U1989 (N_1989,N_1294,N_1769);
and U1990 (N_1990,N_1265,N_1327);
and U1991 (N_1991,N_1710,N_1222);
nand U1992 (N_1992,N_1228,N_1677);
nor U1993 (N_1993,N_1268,N_1433);
nand U1994 (N_1994,N_1637,N_1538);
and U1995 (N_1995,N_1473,N_1451);
and U1996 (N_1996,N_1443,N_1204);
and U1997 (N_1997,N_1300,N_1719);
nor U1998 (N_1998,N_1430,N_1205);
nor U1999 (N_1999,N_1797,N_1727);
or U2000 (N_2000,N_1569,N_1395);
nor U2001 (N_2001,N_1232,N_1690);
nand U2002 (N_2002,N_1522,N_1584);
or U2003 (N_2003,N_1337,N_1249);
nor U2004 (N_2004,N_1760,N_1281);
or U2005 (N_2005,N_1211,N_1544);
or U2006 (N_2006,N_1262,N_1735);
and U2007 (N_2007,N_1675,N_1571);
nand U2008 (N_2008,N_1202,N_1517);
or U2009 (N_2009,N_1349,N_1392);
nand U2010 (N_2010,N_1525,N_1601);
nand U2011 (N_2011,N_1533,N_1700);
nor U2012 (N_2012,N_1383,N_1670);
nand U2013 (N_2013,N_1551,N_1452);
and U2014 (N_2014,N_1593,N_1374);
or U2015 (N_2015,N_1208,N_1556);
nor U2016 (N_2016,N_1400,N_1305);
nand U2017 (N_2017,N_1324,N_1235);
or U2018 (N_2018,N_1539,N_1378);
or U2019 (N_2019,N_1552,N_1751);
nand U2020 (N_2020,N_1639,N_1766);
and U2021 (N_2021,N_1519,N_1791);
nand U2022 (N_2022,N_1364,N_1586);
or U2023 (N_2023,N_1704,N_1757);
nor U2024 (N_2024,N_1592,N_1203);
and U2025 (N_2025,N_1302,N_1672);
nand U2026 (N_2026,N_1340,N_1441);
and U2027 (N_2027,N_1213,N_1484);
nand U2028 (N_2028,N_1555,N_1469);
nand U2029 (N_2029,N_1485,N_1536);
nand U2030 (N_2030,N_1362,N_1699);
or U2031 (N_2031,N_1245,N_1404);
nor U2032 (N_2032,N_1466,N_1753);
or U2033 (N_2033,N_1221,N_1761);
nor U2034 (N_2034,N_1236,N_1463);
nand U2035 (N_2035,N_1570,N_1669);
or U2036 (N_2036,N_1259,N_1607);
nand U2037 (N_2037,N_1763,N_1260);
nor U2038 (N_2038,N_1674,N_1705);
xor U2039 (N_2039,N_1380,N_1274);
nand U2040 (N_2040,N_1575,N_1565);
nand U2041 (N_2041,N_1523,N_1201);
and U2042 (N_2042,N_1731,N_1702);
or U2043 (N_2043,N_1461,N_1435);
nor U2044 (N_2044,N_1726,N_1605);
nor U2045 (N_2045,N_1661,N_1545);
and U2046 (N_2046,N_1638,N_1442);
nand U2047 (N_2047,N_1345,N_1572);
nand U2048 (N_2048,N_1734,N_1663);
nand U2049 (N_2049,N_1382,N_1627);
or U2050 (N_2050,N_1481,N_1286);
nand U2051 (N_2051,N_1325,N_1521);
or U2052 (N_2052,N_1530,N_1573);
or U2053 (N_2053,N_1737,N_1376);
nor U2054 (N_2054,N_1477,N_1729);
and U2055 (N_2055,N_1446,N_1257);
and U2056 (N_2056,N_1253,N_1503);
nand U2057 (N_2057,N_1784,N_1315);
or U2058 (N_2058,N_1513,N_1687);
nor U2059 (N_2059,N_1420,N_1467);
and U2060 (N_2060,N_1790,N_1793);
nand U2061 (N_2061,N_1742,N_1599);
nor U2062 (N_2062,N_1331,N_1497);
nor U2063 (N_2063,N_1698,N_1650);
nand U2064 (N_2064,N_1619,N_1709);
nor U2065 (N_2065,N_1765,N_1558);
and U2066 (N_2066,N_1564,N_1744);
nor U2067 (N_2067,N_1455,N_1770);
and U2068 (N_2068,N_1297,N_1741);
nor U2069 (N_2069,N_1728,N_1462);
or U2070 (N_2070,N_1590,N_1241);
or U2071 (N_2071,N_1356,N_1561);
or U2072 (N_2072,N_1389,N_1206);
and U2073 (N_2073,N_1756,N_1316);
or U2074 (N_2074,N_1322,N_1288);
nand U2075 (N_2075,N_1730,N_1414);
nor U2076 (N_2076,N_1449,N_1543);
nand U2077 (N_2077,N_1660,N_1595);
nor U2078 (N_2078,N_1772,N_1427);
nand U2079 (N_2079,N_1612,N_1507);
nor U2080 (N_2080,N_1749,N_1725);
nand U2081 (N_2081,N_1273,N_1209);
or U2082 (N_2082,N_1554,N_1508);
and U2083 (N_2083,N_1415,N_1713);
or U2084 (N_2084,N_1318,N_1781);
nand U2085 (N_2085,N_1370,N_1792);
nand U2086 (N_2086,N_1604,N_1676);
or U2087 (N_2087,N_1231,N_1293);
or U2088 (N_2088,N_1289,N_1226);
and U2089 (N_2089,N_1692,N_1635);
and U2090 (N_2090,N_1471,N_1688);
nor U2091 (N_2091,N_1295,N_1423);
nand U2092 (N_2092,N_1490,N_1408);
and U2093 (N_2093,N_1361,N_1214);
or U2094 (N_2094,N_1636,N_1752);
nor U2095 (N_2095,N_1795,N_1256);
or U2096 (N_2096,N_1475,N_1405);
nor U2097 (N_2097,N_1746,N_1482);
or U2098 (N_2098,N_1707,N_1308);
nor U2099 (N_2099,N_1480,N_1758);
and U2100 (N_2100,N_1603,N_1753);
and U2101 (N_2101,N_1426,N_1741);
or U2102 (N_2102,N_1277,N_1491);
or U2103 (N_2103,N_1637,N_1224);
nor U2104 (N_2104,N_1507,N_1568);
nor U2105 (N_2105,N_1263,N_1622);
nand U2106 (N_2106,N_1206,N_1537);
xnor U2107 (N_2107,N_1749,N_1365);
and U2108 (N_2108,N_1746,N_1765);
or U2109 (N_2109,N_1235,N_1450);
and U2110 (N_2110,N_1367,N_1717);
nor U2111 (N_2111,N_1384,N_1422);
or U2112 (N_2112,N_1347,N_1555);
nor U2113 (N_2113,N_1278,N_1737);
or U2114 (N_2114,N_1621,N_1574);
or U2115 (N_2115,N_1568,N_1254);
nand U2116 (N_2116,N_1745,N_1418);
and U2117 (N_2117,N_1630,N_1230);
or U2118 (N_2118,N_1211,N_1291);
nand U2119 (N_2119,N_1352,N_1241);
nand U2120 (N_2120,N_1703,N_1738);
and U2121 (N_2121,N_1423,N_1264);
nor U2122 (N_2122,N_1573,N_1591);
nor U2123 (N_2123,N_1703,N_1722);
nand U2124 (N_2124,N_1238,N_1413);
nand U2125 (N_2125,N_1691,N_1229);
and U2126 (N_2126,N_1481,N_1627);
or U2127 (N_2127,N_1765,N_1729);
or U2128 (N_2128,N_1552,N_1683);
nor U2129 (N_2129,N_1609,N_1787);
and U2130 (N_2130,N_1488,N_1367);
nand U2131 (N_2131,N_1232,N_1539);
nand U2132 (N_2132,N_1480,N_1356);
nor U2133 (N_2133,N_1273,N_1547);
or U2134 (N_2134,N_1781,N_1562);
nor U2135 (N_2135,N_1541,N_1210);
nor U2136 (N_2136,N_1296,N_1743);
and U2137 (N_2137,N_1330,N_1772);
nor U2138 (N_2138,N_1506,N_1563);
or U2139 (N_2139,N_1334,N_1373);
nand U2140 (N_2140,N_1259,N_1349);
or U2141 (N_2141,N_1536,N_1731);
nand U2142 (N_2142,N_1669,N_1417);
nor U2143 (N_2143,N_1504,N_1686);
nand U2144 (N_2144,N_1572,N_1445);
or U2145 (N_2145,N_1729,N_1751);
and U2146 (N_2146,N_1743,N_1368);
nor U2147 (N_2147,N_1305,N_1607);
nand U2148 (N_2148,N_1437,N_1220);
nand U2149 (N_2149,N_1391,N_1690);
nor U2150 (N_2150,N_1597,N_1588);
and U2151 (N_2151,N_1453,N_1780);
or U2152 (N_2152,N_1713,N_1220);
nor U2153 (N_2153,N_1500,N_1706);
or U2154 (N_2154,N_1662,N_1276);
and U2155 (N_2155,N_1742,N_1289);
nor U2156 (N_2156,N_1413,N_1463);
or U2157 (N_2157,N_1450,N_1547);
and U2158 (N_2158,N_1729,N_1766);
nand U2159 (N_2159,N_1541,N_1416);
or U2160 (N_2160,N_1289,N_1210);
nand U2161 (N_2161,N_1226,N_1475);
or U2162 (N_2162,N_1309,N_1618);
or U2163 (N_2163,N_1598,N_1760);
nor U2164 (N_2164,N_1581,N_1348);
or U2165 (N_2165,N_1591,N_1623);
and U2166 (N_2166,N_1398,N_1569);
or U2167 (N_2167,N_1611,N_1550);
and U2168 (N_2168,N_1215,N_1719);
nor U2169 (N_2169,N_1329,N_1581);
and U2170 (N_2170,N_1544,N_1687);
nor U2171 (N_2171,N_1600,N_1329);
or U2172 (N_2172,N_1476,N_1217);
and U2173 (N_2173,N_1585,N_1219);
or U2174 (N_2174,N_1501,N_1495);
and U2175 (N_2175,N_1645,N_1406);
or U2176 (N_2176,N_1666,N_1342);
nand U2177 (N_2177,N_1328,N_1255);
nor U2178 (N_2178,N_1383,N_1468);
nand U2179 (N_2179,N_1236,N_1547);
or U2180 (N_2180,N_1456,N_1500);
or U2181 (N_2181,N_1533,N_1494);
and U2182 (N_2182,N_1354,N_1321);
nand U2183 (N_2183,N_1451,N_1248);
nor U2184 (N_2184,N_1621,N_1623);
nor U2185 (N_2185,N_1346,N_1557);
and U2186 (N_2186,N_1440,N_1246);
nor U2187 (N_2187,N_1325,N_1248);
nor U2188 (N_2188,N_1420,N_1412);
nand U2189 (N_2189,N_1316,N_1674);
and U2190 (N_2190,N_1691,N_1426);
and U2191 (N_2191,N_1262,N_1656);
and U2192 (N_2192,N_1693,N_1318);
and U2193 (N_2193,N_1460,N_1593);
nand U2194 (N_2194,N_1706,N_1224);
nor U2195 (N_2195,N_1349,N_1669);
nor U2196 (N_2196,N_1631,N_1782);
nor U2197 (N_2197,N_1273,N_1777);
or U2198 (N_2198,N_1647,N_1565);
or U2199 (N_2199,N_1506,N_1591);
nor U2200 (N_2200,N_1259,N_1751);
nor U2201 (N_2201,N_1523,N_1244);
or U2202 (N_2202,N_1304,N_1799);
nor U2203 (N_2203,N_1470,N_1539);
and U2204 (N_2204,N_1792,N_1537);
nand U2205 (N_2205,N_1667,N_1281);
nor U2206 (N_2206,N_1433,N_1435);
and U2207 (N_2207,N_1619,N_1780);
and U2208 (N_2208,N_1798,N_1309);
nand U2209 (N_2209,N_1465,N_1248);
nand U2210 (N_2210,N_1277,N_1421);
and U2211 (N_2211,N_1448,N_1477);
or U2212 (N_2212,N_1788,N_1777);
and U2213 (N_2213,N_1567,N_1362);
nand U2214 (N_2214,N_1462,N_1402);
and U2215 (N_2215,N_1283,N_1709);
and U2216 (N_2216,N_1411,N_1587);
nor U2217 (N_2217,N_1291,N_1602);
and U2218 (N_2218,N_1592,N_1781);
nor U2219 (N_2219,N_1207,N_1256);
nand U2220 (N_2220,N_1443,N_1488);
or U2221 (N_2221,N_1752,N_1232);
or U2222 (N_2222,N_1669,N_1580);
or U2223 (N_2223,N_1524,N_1513);
and U2224 (N_2224,N_1439,N_1690);
and U2225 (N_2225,N_1662,N_1504);
nand U2226 (N_2226,N_1713,N_1497);
nand U2227 (N_2227,N_1636,N_1289);
and U2228 (N_2228,N_1369,N_1361);
and U2229 (N_2229,N_1468,N_1746);
or U2230 (N_2230,N_1738,N_1725);
nor U2231 (N_2231,N_1512,N_1211);
nand U2232 (N_2232,N_1544,N_1605);
and U2233 (N_2233,N_1761,N_1728);
xor U2234 (N_2234,N_1770,N_1486);
or U2235 (N_2235,N_1598,N_1562);
and U2236 (N_2236,N_1494,N_1789);
nor U2237 (N_2237,N_1494,N_1423);
nor U2238 (N_2238,N_1409,N_1747);
nor U2239 (N_2239,N_1651,N_1548);
or U2240 (N_2240,N_1678,N_1406);
nand U2241 (N_2241,N_1732,N_1343);
nor U2242 (N_2242,N_1383,N_1364);
or U2243 (N_2243,N_1506,N_1721);
or U2244 (N_2244,N_1416,N_1631);
or U2245 (N_2245,N_1548,N_1554);
nor U2246 (N_2246,N_1473,N_1433);
and U2247 (N_2247,N_1225,N_1487);
and U2248 (N_2248,N_1531,N_1575);
and U2249 (N_2249,N_1456,N_1252);
or U2250 (N_2250,N_1544,N_1668);
nor U2251 (N_2251,N_1720,N_1331);
and U2252 (N_2252,N_1268,N_1215);
and U2253 (N_2253,N_1379,N_1232);
or U2254 (N_2254,N_1659,N_1716);
or U2255 (N_2255,N_1203,N_1350);
or U2256 (N_2256,N_1769,N_1616);
nor U2257 (N_2257,N_1584,N_1757);
and U2258 (N_2258,N_1315,N_1347);
nand U2259 (N_2259,N_1766,N_1736);
nand U2260 (N_2260,N_1667,N_1377);
nand U2261 (N_2261,N_1456,N_1415);
and U2262 (N_2262,N_1340,N_1766);
or U2263 (N_2263,N_1673,N_1380);
and U2264 (N_2264,N_1391,N_1252);
or U2265 (N_2265,N_1507,N_1541);
or U2266 (N_2266,N_1425,N_1488);
nand U2267 (N_2267,N_1243,N_1477);
and U2268 (N_2268,N_1535,N_1731);
and U2269 (N_2269,N_1413,N_1419);
and U2270 (N_2270,N_1575,N_1777);
or U2271 (N_2271,N_1793,N_1740);
nand U2272 (N_2272,N_1418,N_1610);
or U2273 (N_2273,N_1664,N_1623);
xnor U2274 (N_2274,N_1356,N_1421);
or U2275 (N_2275,N_1733,N_1743);
and U2276 (N_2276,N_1396,N_1483);
nor U2277 (N_2277,N_1722,N_1321);
or U2278 (N_2278,N_1296,N_1587);
and U2279 (N_2279,N_1613,N_1715);
or U2280 (N_2280,N_1577,N_1528);
or U2281 (N_2281,N_1687,N_1484);
and U2282 (N_2282,N_1562,N_1532);
and U2283 (N_2283,N_1728,N_1291);
xor U2284 (N_2284,N_1674,N_1439);
or U2285 (N_2285,N_1706,N_1519);
nand U2286 (N_2286,N_1792,N_1406);
and U2287 (N_2287,N_1475,N_1202);
or U2288 (N_2288,N_1581,N_1318);
nand U2289 (N_2289,N_1474,N_1238);
nor U2290 (N_2290,N_1435,N_1569);
nand U2291 (N_2291,N_1362,N_1445);
nand U2292 (N_2292,N_1751,N_1705);
or U2293 (N_2293,N_1733,N_1282);
nor U2294 (N_2294,N_1454,N_1541);
and U2295 (N_2295,N_1532,N_1569);
nand U2296 (N_2296,N_1391,N_1577);
nor U2297 (N_2297,N_1779,N_1284);
and U2298 (N_2298,N_1602,N_1262);
nand U2299 (N_2299,N_1605,N_1720);
nand U2300 (N_2300,N_1361,N_1539);
nor U2301 (N_2301,N_1641,N_1499);
and U2302 (N_2302,N_1279,N_1258);
and U2303 (N_2303,N_1553,N_1265);
and U2304 (N_2304,N_1599,N_1384);
or U2305 (N_2305,N_1521,N_1519);
nor U2306 (N_2306,N_1454,N_1278);
nor U2307 (N_2307,N_1429,N_1625);
nand U2308 (N_2308,N_1476,N_1531);
or U2309 (N_2309,N_1557,N_1231);
and U2310 (N_2310,N_1521,N_1212);
nand U2311 (N_2311,N_1212,N_1247);
nand U2312 (N_2312,N_1311,N_1777);
xnor U2313 (N_2313,N_1651,N_1581);
or U2314 (N_2314,N_1479,N_1495);
nor U2315 (N_2315,N_1633,N_1619);
nor U2316 (N_2316,N_1582,N_1563);
nor U2317 (N_2317,N_1678,N_1495);
and U2318 (N_2318,N_1330,N_1625);
or U2319 (N_2319,N_1754,N_1617);
and U2320 (N_2320,N_1675,N_1405);
or U2321 (N_2321,N_1354,N_1341);
nand U2322 (N_2322,N_1214,N_1669);
nor U2323 (N_2323,N_1499,N_1689);
nor U2324 (N_2324,N_1601,N_1744);
nand U2325 (N_2325,N_1628,N_1314);
and U2326 (N_2326,N_1726,N_1206);
and U2327 (N_2327,N_1248,N_1437);
and U2328 (N_2328,N_1795,N_1482);
nor U2329 (N_2329,N_1680,N_1712);
nor U2330 (N_2330,N_1529,N_1245);
and U2331 (N_2331,N_1790,N_1780);
and U2332 (N_2332,N_1665,N_1310);
nor U2333 (N_2333,N_1205,N_1381);
nor U2334 (N_2334,N_1504,N_1769);
and U2335 (N_2335,N_1219,N_1405);
nor U2336 (N_2336,N_1209,N_1640);
or U2337 (N_2337,N_1220,N_1779);
nor U2338 (N_2338,N_1341,N_1683);
nor U2339 (N_2339,N_1459,N_1236);
and U2340 (N_2340,N_1206,N_1522);
nand U2341 (N_2341,N_1447,N_1305);
or U2342 (N_2342,N_1378,N_1625);
and U2343 (N_2343,N_1470,N_1544);
or U2344 (N_2344,N_1344,N_1735);
and U2345 (N_2345,N_1591,N_1460);
nand U2346 (N_2346,N_1266,N_1706);
nor U2347 (N_2347,N_1447,N_1773);
xor U2348 (N_2348,N_1240,N_1432);
nand U2349 (N_2349,N_1307,N_1233);
and U2350 (N_2350,N_1706,N_1462);
nor U2351 (N_2351,N_1534,N_1636);
nor U2352 (N_2352,N_1419,N_1348);
nand U2353 (N_2353,N_1309,N_1786);
nand U2354 (N_2354,N_1549,N_1311);
or U2355 (N_2355,N_1390,N_1494);
or U2356 (N_2356,N_1595,N_1657);
nor U2357 (N_2357,N_1438,N_1551);
or U2358 (N_2358,N_1348,N_1474);
nor U2359 (N_2359,N_1435,N_1444);
and U2360 (N_2360,N_1410,N_1700);
nor U2361 (N_2361,N_1770,N_1369);
or U2362 (N_2362,N_1332,N_1407);
and U2363 (N_2363,N_1640,N_1650);
nand U2364 (N_2364,N_1684,N_1478);
or U2365 (N_2365,N_1390,N_1693);
and U2366 (N_2366,N_1285,N_1733);
nor U2367 (N_2367,N_1221,N_1431);
or U2368 (N_2368,N_1353,N_1574);
nor U2369 (N_2369,N_1568,N_1583);
nand U2370 (N_2370,N_1438,N_1700);
or U2371 (N_2371,N_1684,N_1327);
or U2372 (N_2372,N_1220,N_1290);
nand U2373 (N_2373,N_1606,N_1549);
nor U2374 (N_2374,N_1458,N_1777);
nor U2375 (N_2375,N_1295,N_1782);
and U2376 (N_2376,N_1632,N_1649);
and U2377 (N_2377,N_1501,N_1517);
or U2378 (N_2378,N_1607,N_1647);
nor U2379 (N_2379,N_1243,N_1236);
and U2380 (N_2380,N_1291,N_1290);
nand U2381 (N_2381,N_1692,N_1628);
nand U2382 (N_2382,N_1258,N_1518);
or U2383 (N_2383,N_1661,N_1315);
or U2384 (N_2384,N_1329,N_1220);
nand U2385 (N_2385,N_1585,N_1272);
or U2386 (N_2386,N_1658,N_1453);
and U2387 (N_2387,N_1770,N_1688);
nand U2388 (N_2388,N_1462,N_1470);
nand U2389 (N_2389,N_1310,N_1656);
nor U2390 (N_2390,N_1683,N_1407);
and U2391 (N_2391,N_1647,N_1756);
and U2392 (N_2392,N_1780,N_1379);
or U2393 (N_2393,N_1606,N_1318);
or U2394 (N_2394,N_1798,N_1282);
nor U2395 (N_2395,N_1367,N_1686);
nand U2396 (N_2396,N_1347,N_1416);
and U2397 (N_2397,N_1484,N_1455);
nor U2398 (N_2398,N_1300,N_1299);
nor U2399 (N_2399,N_1430,N_1384);
nand U2400 (N_2400,N_2135,N_2275);
nor U2401 (N_2401,N_2394,N_2036);
nand U2402 (N_2402,N_2026,N_1993);
or U2403 (N_2403,N_1803,N_2029);
nand U2404 (N_2404,N_2309,N_1912);
and U2405 (N_2405,N_2189,N_2022);
and U2406 (N_2406,N_2058,N_2259);
nand U2407 (N_2407,N_1825,N_1844);
nand U2408 (N_2408,N_2395,N_2027);
nand U2409 (N_2409,N_2228,N_2114);
and U2410 (N_2410,N_2349,N_2177);
nand U2411 (N_2411,N_1963,N_2001);
nand U2412 (N_2412,N_1823,N_2168);
nor U2413 (N_2413,N_2186,N_2359);
nand U2414 (N_2414,N_2054,N_1967);
or U2415 (N_2415,N_2231,N_1816);
nand U2416 (N_2416,N_2223,N_2193);
nor U2417 (N_2417,N_2175,N_1918);
and U2418 (N_2418,N_1890,N_2315);
nand U2419 (N_2419,N_2295,N_2121);
nand U2420 (N_2420,N_1926,N_2269);
nand U2421 (N_2421,N_1853,N_1879);
or U2422 (N_2422,N_2200,N_2323);
or U2423 (N_2423,N_1812,N_1832);
and U2424 (N_2424,N_1835,N_2018);
and U2425 (N_2425,N_2093,N_2146);
or U2426 (N_2426,N_2075,N_2227);
and U2427 (N_2427,N_2131,N_2117);
nor U2428 (N_2428,N_2298,N_1884);
and U2429 (N_2429,N_2123,N_2381);
nor U2430 (N_2430,N_1839,N_2055);
nand U2431 (N_2431,N_2250,N_1834);
or U2432 (N_2432,N_1997,N_1917);
nor U2433 (N_2433,N_2377,N_2178);
or U2434 (N_2434,N_1973,N_2369);
nor U2435 (N_2435,N_2245,N_2097);
nor U2436 (N_2436,N_2110,N_2329);
or U2437 (N_2437,N_1856,N_2358);
and U2438 (N_2438,N_2328,N_2201);
nand U2439 (N_2439,N_2339,N_1907);
or U2440 (N_2440,N_2062,N_2282);
nand U2441 (N_2441,N_2089,N_2188);
nor U2442 (N_2442,N_2158,N_2324);
nand U2443 (N_2443,N_2287,N_1938);
nor U2444 (N_2444,N_2021,N_2370);
nor U2445 (N_2445,N_2336,N_2308);
and U2446 (N_2446,N_1897,N_1908);
nor U2447 (N_2447,N_1928,N_2101);
nor U2448 (N_2448,N_2144,N_2086);
and U2449 (N_2449,N_2399,N_2345);
or U2450 (N_2450,N_1802,N_2235);
nand U2451 (N_2451,N_2330,N_2078);
nand U2452 (N_2452,N_2127,N_2252);
nor U2453 (N_2453,N_2011,N_2007);
and U2454 (N_2454,N_2218,N_2139);
nand U2455 (N_2455,N_2073,N_2005);
or U2456 (N_2456,N_1910,N_2262);
and U2457 (N_2457,N_1877,N_2129);
and U2458 (N_2458,N_1849,N_2009);
nand U2459 (N_2459,N_1945,N_1871);
nand U2460 (N_2460,N_2348,N_2109);
or U2461 (N_2461,N_2130,N_1956);
and U2462 (N_2462,N_2289,N_2136);
nor U2463 (N_2463,N_2023,N_1954);
or U2464 (N_2464,N_2105,N_2331);
nor U2465 (N_2465,N_1914,N_2346);
nand U2466 (N_2466,N_1880,N_1970);
or U2467 (N_2467,N_2300,N_2068);
and U2468 (N_2468,N_1833,N_2085);
and U2469 (N_2469,N_2032,N_2003);
or U2470 (N_2470,N_2065,N_2080);
nor U2471 (N_2471,N_1957,N_2187);
nand U2472 (N_2472,N_2215,N_1920);
and U2473 (N_2473,N_2145,N_2050);
or U2474 (N_2474,N_2046,N_1903);
or U2475 (N_2475,N_2192,N_2041);
nand U2476 (N_2476,N_2334,N_1965);
or U2477 (N_2477,N_1894,N_2272);
nand U2478 (N_2478,N_2357,N_1846);
nand U2479 (N_2479,N_2142,N_1971);
nor U2480 (N_2480,N_1900,N_2154);
or U2481 (N_2481,N_2241,N_2035);
or U2482 (N_2482,N_1854,N_2364);
nand U2483 (N_2483,N_2389,N_2113);
or U2484 (N_2484,N_2179,N_2217);
nand U2485 (N_2485,N_2387,N_1818);
nor U2486 (N_2486,N_2350,N_1944);
and U2487 (N_2487,N_2354,N_1959);
nand U2488 (N_2488,N_2363,N_2040);
or U2489 (N_2489,N_2077,N_2224);
nand U2490 (N_2490,N_2102,N_1817);
nor U2491 (N_2491,N_2163,N_2081);
or U2492 (N_2492,N_2290,N_1909);
or U2493 (N_2493,N_2321,N_2061);
nand U2494 (N_2494,N_2320,N_1850);
nand U2495 (N_2495,N_2264,N_2118);
nor U2496 (N_2496,N_2184,N_1985);
nor U2497 (N_2497,N_2157,N_2010);
nor U2498 (N_2498,N_1981,N_2302);
nor U2499 (N_2499,N_2247,N_1898);
nor U2500 (N_2500,N_1919,N_2303);
nor U2501 (N_2501,N_2281,N_2197);
nand U2502 (N_2502,N_2216,N_2006);
or U2503 (N_2503,N_1896,N_1806);
xor U2504 (N_2504,N_2220,N_2014);
and U2505 (N_2505,N_2326,N_2286);
nor U2506 (N_2506,N_2292,N_1905);
and U2507 (N_2507,N_1949,N_1906);
nor U2508 (N_2508,N_1875,N_1838);
nand U2509 (N_2509,N_1888,N_2152);
nor U2510 (N_2510,N_2076,N_2088);
or U2511 (N_2511,N_1975,N_2053);
nor U2512 (N_2512,N_2033,N_1866);
xor U2513 (N_2513,N_2096,N_1827);
nor U2514 (N_2514,N_2258,N_2071);
nor U2515 (N_2515,N_2319,N_2148);
nor U2516 (N_2516,N_2393,N_2194);
nand U2517 (N_2517,N_1974,N_1976);
nand U2518 (N_2518,N_2316,N_1988);
nand U2519 (N_2519,N_1979,N_2276);
nor U2520 (N_2520,N_2052,N_2265);
nand U2521 (N_2521,N_2196,N_2383);
nor U2522 (N_2522,N_2362,N_2229);
nand U2523 (N_2523,N_2128,N_1994);
and U2524 (N_2524,N_1882,N_1881);
nand U2525 (N_2525,N_1961,N_2371);
nor U2526 (N_2526,N_2083,N_2043);
or U2527 (N_2527,N_2322,N_1969);
or U2528 (N_2528,N_2273,N_2103);
nor U2529 (N_2529,N_2238,N_1915);
and U2530 (N_2530,N_2256,N_2239);
xor U2531 (N_2531,N_2199,N_1980);
and U2532 (N_2532,N_2122,N_1810);
xnor U2533 (N_2533,N_2064,N_1822);
and U2534 (N_2534,N_2070,N_1901);
and U2535 (N_2535,N_2198,N_2310);
or U2536 (N_2536,N_2207,N_2341);
nand U2537 (N_2537,N_1960,N_2291);
or U2538 (N_2538,N_2260,N_1916);
or U2539 (N_2539,N_2045,N_1962);
or U2540 (N_2540,N_2051,N_2047);
or U2541 (N_2541,N_2398,N_2133);
nor U2542 (N_2542,N_2222,N_2351);
or U2543 (N_2543,N_2016,N_2283);
and U2544 (N_2544,N_2376,N_2185);
nor U2545 (N_2545,N_1902,N_2211);
nand U2546 (N_2546,N_1865,N_2367);
nand U2547 (N_2547,N_2072,N_2174);
and U2548 (N_2548,N_2237,N_1984);
nor U2549 (N_2549,N_2195,N_1851);
nand U2550 (N_2550,N_1872,N_2297);
and U2551 (N_2551,N_1932,N_1996);
nand U2552 (N_2552,N_1936,N_1927);
and U2553 (N_2553,N_2056,N_2249);
nor U2554 (N_2554,N_2327,N_2049);
or U2555 (N_2555,N_1892,N_1977);
and U2556 (N_2556,N_1828,N_1899);
and U2557 (N_2557,N_2268,N_2396);
nor U2558 (N_2558,N_1930,N_1941);
and U2559 (N_2559,N_2380,N_1830);
nor U2560 (N_2560,N_2385,N_1840);
or U2561 (N_2561,N_2312,N_2244);
or U2562 (N_2562,N_1887,N_2079);
nand U2563 (N_2563,N_1943,N_1942);
and U2564 (N_2564,N_2203,N_2378);
nand U2565 (N_2565,N_2277,N_1804);
or U2566 (N_2566,N_2301,N_2388);
nor U2567 (N_2567,N_2391,N_2095);
and U2568 (N_2568,N_2280,N_2221);
nor U2569 (N_2569,N_2119,N_1931);
nor U2570 (N_2570,N_1955,N_2180);
or U2571 (N_2571,N_1847,N_1911);
and U2572 (N_2572,N_2156,N_2008);
nand U2573 (N_2573,N_2125,N_2274);
or U2574 (N_2574,N_1968,N_2164);
or U2575 (N_2575,N_2074,N_2147);
or U2576 (N_2576,N_1859,N_2210);
or U2577 (N_2577,N_1992,N_1893);
nand U2578 (N_2578,N_1815,N_1870);
nor U2579 (N_2579,N_1958,N_2155);
nor U2580 (N_2580,N_2138,N_2090);
nand U2581 (N_2581,N_2373,N_2299);
and U2582 (N_2582,N_2150,N_1950);
or U2583 (N_2583,N_2233,N_2000);
or U2584 (N_2584,N_2342,N_2332);
or U2585 (N_2585,N_2304,N_1998);
and U2586 (N_2586,N_2356,N_2360);
nor U2587 (N_2587,N_2368,N_1867);
or U2588 (N_2588,N_2335,N_2031);
or U2589 (N_2589,N_2165,N_1852);
nand U2590 (N_2590,N_2205,N_2104);
or U2591 (N_2591,N_1952,N_2116);
and U2592 (N_2592,N_2271,N_1857);
nand U2593 (N_2593,N_2325,N_2167);
and U2594 (N_2594,N_2037,N_1821);
xnor U2595 (N_2595,N_1824,N_2170);
nor U2596 (N_2596,N_1819,N_2253);
or U2597 (N_2597,N_2248,N_1841);
and U2598 (N_2598,N_2162,N_2028);
or U2599 (N_2599,N_2171,N_2025);
nor U2600 (N_2600,N_2375,N_2153);
nand U2601 (N_2601,N_2202,N_2151);
or U2602 (N_2602,N_1869,N_1904);
and U2603 (N_2603,N_1972,N_2161);
or U2604 (N_2604,N_1883,N_1935);
or U2605 (N_2605,N_1885,N_2063);
nand U2606 (N_2606,N_2020,N_2232);
and U2607 (N_2607,N_2115,N_1923);
nand U2608 (N_2608,N_2019,N_2038);
and U2609 (N_2609,N_2172,N_2206);
nand U2610 (N_2610,N_2160,N_1999);
nand U2611 (N_2611,N_2182,N_1836);
and U2612 (N_2612,N_1820,N_2100);
nand U2613 (N_2613,N_1826,N_1929);
or U2614 (N_2614,N_2243,N_2106);
and U2615 (N_2615,N_2317,N_2034);
and U2616 (N_2616,N_2374,N_2313);
or U2617 (N_2617,N_2091,N_2296);
or U2618 (N_2618,N_2213,N_1829);
or U2619 (N_2619,N_2107,N_1807);
nor U2620 (N_2620,N_1939,N_1966);
or U2621 (N_2621,N_2181,N_2285);
or U2622 (N_2622,N_1874,N_1922);
nand U2623 (N_2623,N_1845,N_2191);
and U2624 (N_2624,N_2352,N_2343);
or U2625 (N_2625,N_2112,N_2379);
and U2626 (N_2626,N_2386,N_1940);
or U2627 (N_2627,N_2306,N_2390);
or U2628 (N_2628,N_2099,N_1895);
or U2629 (N_2629,N_1933,N_2270);
and U2630 (N_2630,N_2209,N_1991);
nor U2631 (N_2631,N_2242,N_2084);
or U2632 (N_2632,N_2126,N_1862);
or U2633 (N_2633,N_2208,N_1814);
nand U2634 (N_2634,N_1937,N_2057);
nor U2635 (N_2635,N_2044,N_2149);
or U2636 (N_2636,N_2340,N_2366);
nor U2637 (N_2637,N_1953,N_2318);
nor U2638 (N_2638,N_2344,N_1990);
nor U2639 (N_2639,N_1855,N_2307);
nor U2640 (N_2640,N_1987,N_2353);
or U2641 (N_2641,N_2267,N_2013);
and U2642 (N_2642,N_2042,N_2048);
nand U2643 (N_2643,N_2240,N_2060);
or U2644 (N_2644,N_2212,N_2294);
nand U2645 (N_2645,N_1848,N_2255);
or U2646 (N_2646,N_2012,N_2002);
or U2647 (N_2647,N_2134,N_2278);
or U2648 (N_2648,N_2069,N_2214);
nand U2649 (N_2649,N_2173,N_2365);
or U2650 (N_2650,N_2392,N_2166);
nand U2651 (N_2651,N_1837,N_2355);
or U2652 (N_2652,N_1864,N_2284);
nand U2653 (N_2653,N_1964,N_2311);
nand U2654 (N_2654,N_1989,N_2293);
or U2655 (N_2655,N_1876,N_1891);
or U2656 (N_2656,N_2132,N_2257);
nor U2657 (N_2657,N_2141,N_2059);
or U2658 (N_2658,N_2082,N_1878);
and U2659 (N_2659,N_2382,N_2124);
and U2660 (N_2660,N_2024,N_2372);
nor U2661 (N_2661,N_1808,N_1858);
nor U2662 (N_2662,N_2030,N_2333);
and U2663 (N_2663,N_2169,N_1800);
and U2664 (N_2664,N_1925,N_2183);
nand U2665 (N_2665,N_2225,N_2279);
nand U2666 (N_2666,N_1913,N_1843);
and U2667 (N_2667,N_1809,N_1983);
and U2668 (N_2668,N_2263,N_1947);
nor U2669 (N_2669,N_1842,N_2015);
and U2670 (N_2670,N_2067,N_2087);
and U2671 (N_2671,N_1889,N_2337);
and U2672 (N_2672,N_2159,N_1995);
nor U2673 (N_2673,N_2288,N_2219);
nand U2674 (N_2674,N_1946,N_2098);
or U2675 (N_2675,N_1831,N_1982);
nand U2676 (N_2676,N_1978,N_1805);
or U2677 (N_2677,N_2246,N_1863);
nor U2678 (N_2678,N_2004,N_1886);
xor U2679 (N_2679,N_2120,N_1924);
and U2680 (N_2680,N_2230,N_2236);
nor U2681 (N_2681,N_2397,N_1811);
and U2682 (N_2682,N_1801,N_2039);
or U2683 (N_2683,N_1934,N_2266);
nor U2684 (N_2684,N_2384,N_2251);
nand U2685 (N_2685,N_2137,N_1873);
and U2686 (N_2686,N_1986,N_2226);
and U2687 (N_2687,N_1948,N_2176);
nand U2688 (N_2688,N_1951,N_2314);
and U2689 (N_2689,N_2143,N_2108);
and U2690 (N_2690,N_2094,N_2347);
and U2691 (N_2691,N_2361,N_1868);
or U2692 (N_2692,N_2066,N_2140);
or U2693 (N_2693,N_2234,N_1860);
nor U2694 (N_2694,N_2204,N_2338);
or U2695 (N_2695,N_2111,N_1921);
nor U2696 (N_2696,N_2254,N_2305);
or U2697 (N_2697,N_2092,N_2017);
or U2698 (N_2698,N_1861,N_2190);
and U2699 (N_2699,N_2261,N_1813);
or U2700 (N_2700,N_2308,N_2196);
or U2701 (N_2701,N_2298,N_2225);
and U2702 (N_2702,N_2185,N_1861);
or U2703 (N_2703,N_1894,N_2100);
and U2704 (N_2704,N_2057,N_2267);
nand U2705 (N_2705,N_1856,N_2024);
or U2706 (N_2706,N_1846,N_2282);
nor U2707 (N_2707,N_2315,N_1944);
and U2708 (N_2708,N_2211,N_2278);
nand U2709 (N_2709,N_2307,N_2071);
nand U2710 (N_2710,N_1920,N_1824);
or U2711 (N_2711,N_1980,N_2326);
or U2712 (N_2712,N_2353,N_2019);
or U2713 (N_2713,N_2326,N_1800);
or U2714 (N_2714,N_2269,N_2262);
nand U2715 (N_2715,N_2258,N_1820);
nor U2716 (N_2716,N_1991,N_1937);
or U2717 (N_2717,N_1907,N_2294);
nand U2718 (N_2718,N_2349,N_2366);
nand U2719 (N_2719,N_2177,N_2078);
nand U2720 (N_2720,N_2102,N_2012);
or U2721 (N_2721,N_2086,N_1876);
and U2722 (N_2722,N_1957,N_2383);
nor U2723 (N_2723,N_2136,N_2120);
or U2724 (N_2724,N_1984,N_2091);
nand U2725 (N_2725,N_2359,N_2221);
or U2726 (N_2726,N_2203,N_2186);
or U2727 (N_2727,N_2304,N_2291);
nor U2728 (N_2728,N_2087,N_1864);
or U2729 (N_2729,N_1848,N_2342);
or U2730 (N_2730,N_2381,N_2394);
nand U2731 (N_2731,N_2333,N_1937);
and U2732 (N_2732,N_2028,N_2325);
and U2733 (N_2733,N_1928,N_2151);
nor U2734 (N_2734,N_2396,N_2314);
nor U2735 (N_2735,N_1970,N_1876);
nand U2736 (N_2736,N_2283,N_2192);
nor U2737 (N_2737,N_2261,N_1955);
nand U2738 (N_2738,N_2306,N_1875);
nand U2739 (N_2739,N_2257,N_1853);
nand U2740 (N_2740,N_2155,N_2213);
or U2741 (N_2741,N_2038,N_1983);
or U2742 (N_2742,N_2337,N_1845);
nand U2743 (N_2743,N_1828,N_1966);
nand U2744 (N_2744,N_2011,N_1865);
nor U2745 (N_2745,N_2237,N_2294);
or U2746 (N_2746,N_1866,N_2202);
or U2747 (N_2747,N_2162,N_2380);
nand U2748 (N_2748,N_2162,N_2187);
and U2749 (N_2749,N_2101,N_2139);
xnor U2750 (N_2750,N_2200,N_2203);
nand U2751 (N_2751,N_2350,N_2319);
nor U2752 (N_2752,N_1803,N_1826);
nand U2753 (N_2753,N_2309,N_1900);
and U2754 (N_2754,N_2289,N_2385);
and U2755 (N_2755,N_1996,N_1801);
and U2756 (N_2756,N_1902,N_1841);
nand U2757 (N_2757,N_2303,N_2054);
and U2758 (N_2758,N_2000,N_2297);
nand U2759 (N_2759,N_1885,N_1851);
nor U2760 (N_2760,N_1813,N_2125);
and U2761 (N_2761,N_2391,N_2368);
nor U2762 (N_2762,N_1946,N_2359);
nor U2763 (N_2763,N_1942,N_2112);
nor U2764 (N_2764,N_2081,N_2143);
xor U2765 (N_2765,N_1950,N_1999);
nor U2766 (N_2766,N_1987,N_1915);
nor U2767 (N_2767,N_2292,N_2091);
xor U2768 (N_2768,N_1831,N_2132);
or U2769 (N_2769,N_2235,N_1858);
nor U2770 (N_2770,N_2106,N_2249);
nand U2771 (N_2771,N_2224,N_1805);
and U2772 (N_2772,N_1943,N_2090);
nor U2773 (N_2773,N_2360,N_1978);
or U2774 (N_2774,N_2160,N_1870);
nand U2775 (N_2775,N_2351,N_2140);
and U2776 (N_2776,N_2287,N_1828);
and U2777 (N_2777,N_2374,N_1934);
and U2778 (N_2778,N_2254,N_2160);
or U2779 (N_2779,N_1934,N_1887);
nand U2780 (N_2780,N_1854,N_2369);
nor U2781 (N_2781,N_2089,N_2208);
or U2782 (N_2782,N_2160,N_1829);
and U2783 (N_2783,N_2060,N_2235);
or U2784 (N_2784,N_1862,N_2033);
nor U2785 (N_2785,N_1831,N_2178);
nor U2786 (N_2786,N_2318,N_1885);
and U2787 (N_2787,N_1881,N_2363);
nand U2788 (N_2788,N_2376,N_2215);
or U2789 (N_2789,N_1854,N_2263);
nand U2790 (N_2790,N_2054,N_2024);
nor U2791 (N_2791,N_2066,N_1980);
and U2792 (N_2792,N_2157,N_1852);
or U2793 (N_2793,N_2241,N_1950);
nand U2794 (N_2794,N_1819,N_2001);
nor U2795 (N_2795,N_2321,N_1957);
nand U2796 (N_2796,N_2059,N_2138);
and U2797 (N_2797,N_2043,N_1938);
or U2798 (N_2798,N_2204,N_2340);
nor U2799 (N_2799,N_1832,N_2033);
and U2800 (N_2800,N_1863,N_2393);
nand U2801 (N_2801,N_2204,N_2295);
nand U2802 (N_2802,N_2081,N_2012);
and U2803 (N_2803,N_2149,N_2269);
and U2804 (N_2804,N_1979,N_1976);
and U2805 (N_2805,N_2056,N_2096);
or U2806 (N_2806,N_1876,N_2058);
nor U2807 (N_2807,N_2364,N_2360);
nor U2808 (N_2808,N_1898,N_2319);
or U2809 (N_2809,N_2232,N_2360);
and U2810 (N_2810,N_1947,N_1934);
or U2811 (N_2811,N_2364,N_1873);
or U2812 (N_2812,N_2218,N_2299);
nor U2813 (N_2813,N_1979,N_2166);
and U2814 (N_2814,N_1876,N_2330);
and U2815 (N_2815,N_2251,N_2135);
nor U2816 (N_2816,N_2110,N_2399);
nor U2817 (N_2817,N_2119,N_2208);
nor U2818 (N_2818,N_2212,N_2243);
or U2819 (N_2819,N_2397,N_2242);
nor U2820 (N_2820,N_2030,N_2147);
and U2821 (N_2821,N_2056,N_2105);
and U2822 (N_2822,N_2206,N_2232);
nor U2823 (N_2823,N_1894,N_1846);
and U2824 (N_2824,N_1923,N_2311);
and U2825 (N_2825,N_2037,N_2251);
nor U2826 (N_2826,N_2146,N_1933);
nand U2827 (N_2827,N_2061,N_2126);
and U2828 (N_2828,N_1958,N_2161);
and U2829 (N_2829,N_2280,N_2067);
or U2830 (N_2830,N_1951,N_1839);
nand U2831 (N_2831,N_1912,N_2294);
or U2832 (N_2832,N_2145,N_2026);
and U2833 (N_2833,N_2185,N_1919);
nand U2834 (N_2834,N_1977,N_2208);
nor U2835 (N_2835,N_2227,N_1941);
and U2836 (N_2836,N_2075,N_1821);
and U2837 (N_2837,N_1876,N_2231);
nand U2838 (N_2838,N_1927,N_1966);
and U2839 (N_2839,N_2096,N_1899);
nor U2840 (N_2840,N_2281,N_1990);
or U2841 (N_2841,N_1975,N_2396);
nor U2842 (N_2842,N_2302,N_2135);
nor U2843 (N_2843,N_2005,N_1992);
nand U2844 (N_2844,N_1803,N_2361);
and U2845 (N_2845,N_1978,N_2233);
nand U2846 (N_2846,N_2109,N_1941);
nand U2847 (N_2847,N_2365,N_2264);
nand U2848 (N_2848,N_2131,N_2191);
and U2849 (N_2849,N_1819,N_1812);
nor U2850 (N_2850,N_2305,N_2355);
nand U2851 (N_2851,N_2381,N_2322);
and U2852 (N_2852,N_2276,N_2208);
or U2853 (N_2853,N_2047,N_1846);
and U2854 (N_2854,N_1857,N_2066);
nand U2855 (N_2855,N_2152,N_1990);
or U2856 (N_2856,N_2091,N_2346);
nor U2857 (N_2857,N_2112,N_1937);
or U2858 (N_2858,N_1889,N_2159);
or U2859 (N_2859,N_2059,N_1910);
nand U2860 (N_2860,N_2010,N_2036);
nand U2861 (N_2861,N_2306,N_2318);
nor U2862 (N_2862,N_2174,N_2123);
nand U2863 (N_2863,N_2038,N_2167);
and U2864 (N_2864,N_2063,N_2282);
or U2865 (N_2865,N_2072,N_1984);
nor U2866 (N_2866,N_2045,N_2332);
nand U2867 (N_2867,N_2335,N_2175);
nand U2868 (N_2868,N_1852,N_1882);
nand U2869 (N_2869,N_1874,N_2017);
and U2870 (N_2870,N_2150,N_1868);
and U2871 (N_2871,N_2264,N_1984);
nand U2872 (N_2872,N_1860,N_2326);
nand U2873 (N_2873,N_1956,N_1902);
nand U2874 (N_2874,N_1931,N_2063);
and U2875 (N_2875,N_2334,N_1837);
nand U2876 (N_2876,N_2013,N_2381);
nor U2877 (N_2877,N_2165,N_2111);
or U2878 (N_2878,N_1803,N_2295);
nand U2879 (N_2879,N_2098,N_2191);
and U2880 (N_2880,N_1872,N_2280);
and U2881 (N_2881,N_2017,N_2187);
or U2882 (N_2882,N_1961,N_2366);
nand U2883 (N_2883,N_1923,N_2099);
nand U2884 (N_2884,N_2172,N_1980);
nand U2885 (N_2885,N_2346,N_1831);
and U2886 (N_2886,N_1863,N_2370);
or U2887 (N_2887,N_2121,N_1884);
nor U2888 (N_2888,N_1963,N_1952);
nand U2889 (N_2889,N_2279,N_1824);
and U2890 (N_2890,N_1807,N_1840);
or U2891 (N_2891,N_1994,N_2266);
nand U2892 (N_2892,N_2001,N_1960);
and U2893 (N_2893,N_1803,N_2144);
nand U2894 (N_2894,N_1804,N_1953);
nand U2895 (N_2895,N_1938,N_2177);
nand U2896 (N_2896,N_2250,N_1801);
nor U2897 (N_2897,N_1882,N_2144);
and U2898 (N_2898,N_2326,N_2384);
nand U2899 (N_2899,N_2135,N_2276);
or U2900 (N_2900,N_1959,N_2178);
nand U2901 (N_2901,N_2209,N_1837);
or U2902 (N_2902,N_2154,N_2030);
nor U2903 (N_2903,N_1939,N_2136);
nor U2904 (N_2904,N_1855,N_2178);
or U2905 (N_2905,N_1900,N_2292);
or U2906 (N_2906,N_1873,N_2396);
and U2907 (N_2907,N_1990,N_2010);
nand U2908 (N_2908,N_2131,N_2318);
or U2909 (N_2909,N_2372,N_2327);
and U2910 (N_2910,N_2016,N_1974);
and U2911 (N_2911,N_2298,N_2204);
nor U2912 (N_2912,N_2261,N_1990);
nand U2913 (N_2913,N_2225,N_2241);
nor U2914 (N_2914,N_1890,N_2259);
nor U2915 (N_2915,N_2184,N_1973);
nor U2916 (N_2916,N_2163,N_1995);
and U2917 (N_2917,N_2177,N_2306);
nor U2918 (N_2918,N_2135,N_2270);
and U2919 (N_2919,N_1944,N_2183);
nor U2920 (N_2920,N_1805,N_2087);
nor U2921 (N_2921,N_2094,N_1823);
nor U2922 (N_2922,N_2284,N_1863);
and U2923 (N_2923,N_2234,N_2212);
nor U2924 (N_2924,N_1868,N_2296);
nand U2925 (N_2925,N_2226,N_2285);
nand U2926 (N_2926,N_2106,N_2013);
xor U2927 (N_2927,N_2171,N_2173);
nor U2928 (N_2928,N_2283,N_2181);
nand U2929 (N_2929,N_2292,N_2298);
nor U2930 (N_2930,N_1881,N_2138);
or U2931 (N_2931,N_2150,N_2258);
nor U2932 (N_2932,N_2257,N_2217);
and U2933 (N_2933,N_2287,N_2051);
nor U2934 (N_2934,N_2333,N_1983);
nand U2935 (N_2935,N_1826,N_1853);
and U2936 (N_2936,N_2205,N_1845);
or U2937 (N_2937,N_1948,N_1943);
nor U2938 (N_2938,N_1945,N_2292);
nand U2939 (N_2939,N_1902,N_1800);
or U2940 (N_2940,N_2054,N_2324);
nand U2941 (N_2941,N_2138,N_2243);
nand U2942 (N_2942,N_2162,N_2278);
xor U2943 (N_2943,N_1882,N_1991);
nand U2944 (N_2944,N_1838,N_2105);
or U2945 (N_2945,N_1809,N_2284);
nand U2946 (N_2946,N_2104,N_1985);
and U2947 (N_2947,N_2000,N_2286);
nand U2948 (N_2948,N_2146,N_1806);
nand U2949 (N_2949,N_2305,N_2317);
and U2950 (N_2950,N_1831,N_2282);
nor U2951 (N_2951,N_2370,N_2301);
or U2952 (N_2952,N_1852,N_2369);
nor U2953 (N_2953,N_2238,N_1857);
nor U2954 (N_2954,N_2333,N_1869);
or U2955 (N_2955,N_2278,N_1843);
nor U2956 (N_2956,N_2173,N_2221);
and U2957 (N_2957,N_2206,N_1868);
and U2958 (N_2958,N_2044,N_1959);
or U2959 (N_2959,N_2317,N_2371);
or U2960 (N_2960,N_2158,N_1979);
nand U2961 (N_2961,N_1831,N_2101);
and U2962 (N_2962,N_1996,N_2072);
nor U2963 (N_2963,N_1951,N_2269);
nor U2964 (N_2964,N_2164,N_1998);
nor U2965 (N_2965,N_1904,N_2266);
or U2966 (N_2966,N_2070,N_2249);
and U2967 (N_2967,N_2220,N_2390);
or U2968 (N_2968,N_2168,N_2155);
and U2969 (N_2969,N_2156,N_2103);
and U2970 (N_2970,N_2107,N_2068);
and U2971 (N_2971,N_2378,N_1850);
or U2972 (N_2972,N_2350,N_2133);
and U2973 (N_2973,N_2188,N_2029);
or U2974 (N_2974,N_1815,N_1994);
nor U2975 (N_2975,N_2280,N_1812);
or U2976 (N_2976,N_1988,N_1830);
nor U2977 (N_2977,N_1830,N_1973);
nand U2978 (N_2978,N_2099,N_2077);
nor U2979 (N_2979,N_1975,N_1865);
or U2980 (N_2980,N_2068,N_1954);
nand U2981 (N_2981,N_1841,N_2159);
nand U2982 (N_2982,N_1917,N_2239);
and U2983 (N_2983,N_1941,N_2013);
or U2984 (N_2984,N_2170,N_2188);
nand U2985 (N_2985,N_1805,N_2315);
and U2986 (N_2986,N_1928,N_2118);
nand U2987 (N_2987,N_2161,N_2374);
and U2988 (N_2988,N_1893,N_2106);
or U2989 (N_2989,N_1978,N_2100);
or U2990 (N_2990,N_2234,N_2328);
nand U2991 (N_2991,N_2170,N_2374);
and U2992 (N_2992,N_1844,N_2068);
nand U2993 (N_2993,N_2323,N_2147);
nor U2994 (N_2994,N_1871,N_2265);
or U2995 (N_2995,N_2375,N_2135);
or U2996 (N_2996,N_2136,N_2314);
or U2997 (N_2997,N_2008,N_2395);
nor U2998 (N_2998,N_2331,N_1954);
and U2999 (N_2999,N_2211,N_2303);
nand UO_0 (O_0,N_2810,N_2579);
nand UO_1 (O_1,N_2791,N_2696);
nor UO_2 (O_2,N_2801,N_2650);
or UO_3 (O_3,N_2774,N_2482);
and UO_4 (O_4,N_2449,N_2707);
or UO_5 (O_5,N_2597,N_2499);
nor UO_6 (O_6,N_2450,N_2785);
and UO_7 (O_7,N_2563,N_2637);
nand UO_8 (O_8,N_2625,N_2840);
nand UO_9 (O_9,N_2535,N_2910);
and UO_10 (O_10,N_2870,N_2755);
and UO_11 (O_11,N_2610,N_2849);
and UO_12 (O_12,N_2583,N_2505);
nand UO_13 (O_13,N_2880,N_2997);
nand UO_14 (O_14,N_2585,N_2802);
and UO_15 (O_15,N_2770,N_2458);
nand UO_16 (O_16,N_2846,N_2768);
nand UO_17 (O_17,N_2565,N_2575);
nand UO_18 (O_18,N_2715,N_2541);
and UO_19 (O_19,N_2558,N_2963);
or UO_20 (O_20,N_2589,N_2699);
nand UO_21 (O_21,N_2488,N_2772);
and UO_22 (O_22,N_2649,N_2968);
nor UO_23 (O_23,N_2987,N_2468);
and UO_24 (O_24,N_2540,N_2994);
or UO_25 (O_25,N_2518,N_2821);
xnor UO_26 (O_26,N_2847,N_2553);
nand UO_27 (O_27,N_2977,N_2662);
nand UO_28 (O_28,N_2722,N_2783);
and UO_29 (O_29,N_2651,N_2947);
or UO_30 (O_30,N_2559,N_2412);
nor UO_31 (O_31,N_2995,N_2401);
or UO_32 (O_32,N_2764,N_2964);
nor UO_33 (O_33,N_2591,N_2477);
xnor UO_34 (O_34,N_2430,N_2684);
or UO_35 (O_35,N_2714,N_2506);
and UO_36 (O_36,N_2823,N_2492);
or UO_37 (O_37,N_2570,N_2984);
or UO_38 (O_38,N_2421,N_2965);
nor UO_39 (O_39,N_2648,N_2655);
or UO_40 (O_40,N_2415,N_2989);
or UO_41 (O_41,N_2920,N_2627);
or UO_42 (O_42,N_2786,N_2456);
and UO_43 (O_43,N_2544,N_2400);
or UO_44 (O_44,N_2685,N_2760);
and UO_45 (O_45,N_2673,N_2659);
nor UO_46 (O_46,N_2891,N_2854);
nor UO_47 (O_47,N_2527,N_2517);
nor UO_48 (O_48,N_2717,N_2639);
and UO_49 (O_49,N_2466,N_2879);
and UO_50 (O_50,N_2614,N_2773);
nor UO_51 (O_51,N_2915,N_2682);
nand UO_52 (O_52,N_2694,N_2473);
nor UO_53 (O_53,N_2554,N_2633);
nand UO_54 (O_54,N_2749,N_2405);
and UO_55 (O_55,N_2660,N_2720);
nor UO_56 (O_56,N_2729,N_2586);
or UO_57 (O_57,N_2798,N_2873);
or UO_58 (O_58,N_2726,N_2958);
nor UO_59 (O_59,N_2936,N_2413);
and UO_60 (O_60,N_2676,N_2919);
and UO_61 (O_61,N_2519,N_2538);
or UO_62 (O_62,N_2738,N_2868);
nor UO_63 (O_63,N_2446,N_2561);
and UO_64 (O_64,N_2512,N_2489);
nand UO_65 (O_65,N_2767,N_2551);
and UO_66 (O_66,N_2668,N_2797);
nor UO_67 (O_67,N_2467,N_2486);
and UO_68 (O_68,N_2463,N_2858);
and UO_69 (O_69,N_2776,N_2719);
nor UO_70 (O_70,N_2441,N_2562);
or UO_71 (O_71,N_2874,N_2971);
nand UO_72 (O_72,N_2885,N_2941);
or UO_73 (O_73,N_2713,N_2951);
nand UO_74 (O_74,N_2686,N_2698);
or UO_75 (O_75,N_2602,N_2679);
nand UO_76 (O_76,N_2761,N_2702);
nand UO_77 (O_77,N_2646,N_2611);
and UO_78 (O_78,N_2769,N_2864);
or UO_79 (O_79,N_2745,N_2624);
or UO_80 (O_80,N_2934,N_2661);
nor UO_81 (O_81,N_2582,N_2804);
nand UO_82 (O_82,N_2520,N_2740);
or UO_83 (O_83,N_2911,N_2432);
or UO_84 (O_84,N_2833,N_2800);
nand UO_85 (O_85,N_2688,N_2571);
and UO_86 (O_86,N_2931,N_2781);
and UO_87 (O_87,N_2572,N_2929);
nand UO_88 (O_88,N_2612,N_2855);
and UO_89 (O_89,N_2594,N_2683);
nor UO_90 (O_90,N_2875,N_2939);
or UO_91 (O_91,N_2792,N_2407);
nor UO_92 (O_92,N_2727,N_2427);
nor UO_93 (O_93,N_2710,N_2613);
and UO_94 (O_94,N_2657,N_2495);
and UO_95 (O_95,N_2852,N_2498);
and UO_96 (O_96,N_2771,N_2440);
or UO_97 (O_97,N_2724,N_2998);
and UO_98 (O_98,N_2895,N_2690);
and UO_99 (O_99,N_2990,N_2819);
or UO_100 (O_100,N_2905,N_2952);
nor UO_101 (O_101,N_2595,N_2453);
nor UO_102 (O_102,N_2568,N_2681);
or UO_103 (O_103,N_2652,N_2493);
nand UO_104 (O_104,N_2967,N_2513);
nor UO_105 (O_105,N_2887,N_2590);
or UO_106 (O_106,N_2872,N_2787);
and UO_107 (O_107,N_2675,N_2593);
and UO_108 (O_108,N_2983,N_2985);
or UO_109 (O_109,N_2451,N_2937);
and UO_110 (O_110,N_2414,N_2835);
nor UO_111 (O_111,N_2403,N_2548);
nand UO_112 (O_112,N_2539,N_2980);
and UO_113 (O_113,N_2481,N_2496);
nor UO_114 (O_114,N_2617,N_2596);
and UO_115 (O_115,N_2999,N_2973);
nand UO_116 (O_116,N_2647,N_2507);
nor UO_117 (O_117,N_2629,N_2842);
nand UO_118 (O_118,N_2577,N_2991);
or UO_119 (O_119,N_2645,N_2634);
or UO_120 (O_120,N_2922,N_2908);
nor UO_121 (O_121,N_2871,N_2938);
or UO_122 (O_122,N_2461,N_2763);
nand UO_123 (O_123,N_2457,N_2981);
nor UO_124 (O_124,N_2547,N_2709);
nor UO_125 (O_125,N_2643,N_2423);
and UO_126 (O_126,N_2788,N_2689);
nor UO_127 (O_127,N_2896,N_2912);
nor UO_128 (O_128,N_2509,N_2424);
and UO_129 (O_129,N_2946,N_2902);
or UO_130 (O_130,N_2530,N_2808);
and UO_131 (O_131,N_2824,N_2460);
and UO_132 (O_132,N_2913,N_2867);
or UO_133 (O_133,N_2670,N_2826);
nand UO_134 (O_134,N_2916,N_2529);
or UO_135 (O_135,N_2576,N_2433);
or UO_136 (O_136,N_2564,N_2925);
and UO_137 (O_137,N_2497,N_2806);
xor UO_138 (O_138,N_2567,N_2812);
or UO_139 (O_139,N_2669,N_2472);
and UO_140 (O_140,N_2628,N_2584);
and UO_141 (O_141,N_2494,N_2933);
nand UO_142 (O_142,N_2705,N_2532);
or UO_143 (O_143,N_2526,N_2704);
or UO_144 (O_144,N_2741,N_2831);
nor UO_145 (O_145,N_2502,N_2618);
nand UO_146 (O_146,N_2569,N_2932);
and UO_147 (O_147,N_2695,N_2664);
nor UO_148 (O_148,N_2779,N_2439);
and UO_149 (O_149,N_2654,N_2816);
nand UO_150 (O_150,N_2483,N_2436);
and UO_151 (O_151,N_2886,N_2703);
or UO_152 (O_152,N_2678,N_2969);
or UO_153 (O_153,N_2665,N_2795);
and UO_154 (O_154,N_2574,N_2743);
and UO_155 (O_155,N_2537,N_2863);
and UO_156 (O_156,N_2803,N_2817);
nand UO_157 (O_157,N_2438,N_2636);
and UO_158 (O_158,N_2600,N_2723);
or UO_159 (O_159,N_2543,N_2970);
or UO_160 (O_160,N_2511,N_2578);
and UO_161 (O_161,N_2815,N_2860);
nor UO_162 (O_162,N_2504,N_2974);
and UO_163 (O_163,N_2666,N_2924);
nand UO_164 (O_164,N_2807,N_2701);
and UO_165 (O_165,N_2419,N_2672);
nand UO_166 (O_166,N_2663,N_2805);
nand UO_167 (O_167,N_2844,N_2728);
nor UO_168 (O_168,N_2443,N_2884);
nand UO_169 (O_169,N_2428,N_2982);
or UO_170 (O_170,N_2640,N_2603);
nand UO_171 (O_171,N_2573,N_2918);
and UO_172 (O_172,N_2988,N_2956);
and UO_173 (O_173,N_2725,N_2623);
or UO_174 (O_174,N_2914,N_2992);
nand UO_175 (O_175,N_2406,N_2978);
or UO_176 (O_176,N_2853,N_2533);
and UO_177 (O_177,N_2876,N_2927);
and UO_178 (O_178,N_2903,N_2746);
nor UO_179 (O_179,N_2954,N_2587);
nand UO_180 (O_180,N_2471,N_2751);
or UO_181 (O_181,N_2750,N_2524);
and UO_182 (O_182,N_2889,N_2455);
nand UO_183 (O_183,N_2829,N_2976);
and UO_184 (O_184,N_2893,N_2881);
nand UO_185 (O_185,N_2656,N_2671);
nor UO_186 (O_186,N_2957,N_2930);
or UO_187 (O_187,N_2712,N_2437);
and UO_188 (O_188,N_2869,N_2510);
xor UO_189 (O_189,N_2818,N_2598);
and UO_190 (O_190,N_2516,N_2757);
nand UO_191 (O_191,N_2474,N_2491);
nand UO_192 (O_192,N_2476,N_2566);
nor UO_193 (O_193,N_2475,N_2759);
nor UO_194 (O_194,N_2462,N_2429);
or UO_195 (O_195,N_2777,N_2861);
or UO_196 (O_196,N_2850,N_2878);
nor UO_197 (O_197,N_2626,N_2638);
nand UO_198 (O_198,N_2422,N_2503);
nor UO_199 (O_199,N_2445,N_2906);
nor UO_200 (O_200,N_2425,N_2907);
nor UO_201 (O_201,N_2448,N_2811);
or UO_202 (O_202,N_2856,N_2465);
nor UO_203 (O_203,N_2827,N_2555);
nor UO_204 (O_204,N_2882,N_2635);
and UO_205 (O_205,N_2653,N_2747);
and UO_206 (O_206,N_2809,N_2545);
and UO_207 (O_207,N_2848,N_2528);
nor UO_208 (O_208,N_2888,N_2644);
or UO_209 (O_209,N_2828,N_2814);
xor UO_210 (O_210,N_2744,N_2851);
or UO_211 (O_211,N_2962,N_2490);
nand UO_212 (O_212,N_2834,N_2825);
nor UO_213 (O_213,N_2841,N_2836);
or UO_214 (O_214,N_2959,N_2732);
or UO_215 (O_215,N_2616,N_2478);
nand UO_216 (O_216,N_2753,N_2556);
nor UO_217 (O_217,N_2758,N_2630);
and UO_218 (O_218,N_2961,N_2549);
nand UO_219 (O_219,N_2716,N_2859);
and UO_220 (O_220,N_2742,N_2687);
or UO_221 (O_221,N_2677,N_2960);
or UO_222 (O_222,N_2601,N_2609);
or UO_223 (O_223,N_2560,N_2935);
nor UO_224 (O_224,N_2754,N_2793);
and UO_225 (O_225,N_2546,N_2706);
nand UO_226 (O_226,N_2459,N_2837);
and UO_227 (O_227,N_2508,N_2950);
and UO_228 (O_228,N_2838,N_2890);
xor UO_229 (O_229,N_2975,N_2944);
and UO_230 (O_230,N_2730,N_2447);
and UO_231 (O_231,N_2943,N_2845);
or UO_232 (O_232,N_2622,N_2408);
and UO_233 (O_233,N_2531,N_2940);
nand UO_234 (O_234,N_2464,N_2923);
nor UO_235 (O_235,N_2733,N_2514);
nor UO_236 (O_236,N_2796,N_2945);
nand UO_237 (O_237,N_2454,N_2409);
or UO_238 (O_238,N_2799,N_2621);
nand UO_239 (O_239,N_2892,N_2708);
nor UO_240 (O_240,N_2862,N_2718);
or UO_241 (O_241,N_2550,N_2865);
and UO_242 (O_242,N_2909,N_2731);
and UO_243 (O_243,N_2452,N_2500);
and UO_244 (O_244,N_2700,N_2789);
and UO_245 (O_245,N_2592,N_2697);
nand UO_246 (O_246,N_2748,N_2955);
nand UO_247 (O_247,N_2608,N_2928);
nor UO_248 (O_248,N_2739,N_2900);
nor UO_249 (O_249,N_2658,N_2479);
and UO_250 (O_250,N_2534,N_2417);
or UO_251 (O_251,N_2894,N_2917);
or UO_252 (O_252,N_2735,N_2469);
and UO_253 (O_253,N_2953,N_2790);
nand UO_254 (O_254,N_2766,N_2484);
nor UO_255 (O_255,N_2680,N_2599);
and UO_256 (O_256,N_2813,N_2993);
and UO_257 (O_257,N_2536,N_2921);
nand UO_258 (O_258,N_2604,N_2515);
and UO_259 (O_259,N_2442,N_2866);
nor UO_260 (O_260,N_2605,N_2480);
or UO_261 (O_261,N_2431,N_2552);
nand UO_262 (O_262,N_2557,N_2752);
or UO_263 (O_263,N_2619,N_2667);
nor UO_264 (O_264,N_2691,N_2784);
nand UO_265 (O_265,N_2418,N_2607);
nor UO_266 (O_266,N_2435,N_2734);
nand UO_267 (O_267,N_2822,N_2765);
or UO_268 (O_268,N_2883,N_2404);
or UO_269 (O_269,N_2780,N_2402);
nor UO_270 (O_270,N_2948,N_2966);
nor UO_271 (O_271,N_2487,N_2501);
and UO_272 (O_272,N_2641,N_2820);
nand UO_273 (O_273,N_2642,N_2711);
and UO_274 (O_274,N_2426,N_2420);
or UO_275 (O_275,N_2839,N_2778);
and UO_276 (O_276,N_2606,N_2721);
or UO_277 (O_277,N_2444,N_2411);
or UO_278 (O_278,N_2762,N_2899);
or UO_279 (O_279,N_2736,N_2525);
nand UO_280 (O_280,N_2904,N_2832);
nor UO_281 (O_281,N_2897,N_2470);
and UO_282 (O_282,N_2615,N_2692);
and UO_283 (O_283,N_2523,N_2581);
nand UO_284 (O_284,N_2737,N_2631);
nor UO_285 (O_285,N_2620,N_2986);
nor UO_286 (O_286,N_2674,N_2830);
or UO_287 (O_287,N_2521,N_2756);
and UO_288 (O_288,N_2901,N_2996);
nand UO_289 (O_289,N_2949,N_2972);
nand UO_290 (O_290,N_2588,N_2632);
or UO_291 (O_291,N_2693,N_2857);
nand UO_292 (O_292,N_2979,N_2782);
nand UO_293 (O_293,N_2843,N_2794);
nand UO_294 (O_294,N_2416,N_2434);
and UO_295 (O_295,N_2542,N_2898);
and UO_296 (O_296,N_2522,N_2580);
xnor UO_297 (O_297,N_2926,N_2942);
or UO_298 (O_298,N_2485,N_2877);
nor UO_299 (O_299,N_2410,N_2775);
or UO_300 (O_300,N_2664,N_2940);
nand UO_301 (O_301,N_2922,N_2439);
nor UO_302 (O_302,N_2789,N_2847);
and UO_303 (O_303,N_2470,N_2443);
or UO_304 (O_304,N_2653,N_2554);
nor UO_305 (O_305,N_2407,N_2480);
nor UO_306 (O_306,N_2459,N_2978);
and UO_307 (O_307,N_2427,N_2920);
and UO_308 (O_308,N_2918,N_2799);
or UO_309 (O_309,N_2733,N_2421);
nor UO_310 (O_310,N_2549,N_2684);
nor UO_311 (O_311,N_2743,N_2878);
nand UO_312 (O_312,N_2834,N_2933);
nand UO_313 (O_313,N_2808,N_2416);
nor UO_314 (O_314,N_2807,N_2620);
or UO_315 (O_315,N_2839,N_2540);
nor UO_316 (O_316,N_2729,N_2430);
or UO_317 (O_317,N_2679,N_2794);
nand UO_318 (O_318,N_2510,N_2698);
nand UO_319 (O_319,N_2714,N_2869);
nand UO_320 (O_320,N_2597,N_2682);
or UO_321 (O_321,N_2499,N_2945);
or UO_322 (O_322,N_2938,N_2695);
or UO_323 (O_323,N_2651,N_2635);
and UO_324 (O_324,N_2491,N_2760);
and UO_325 (O_325,N_2499,N_2899);
or UO_326 (O_326,N_2529,N_2670);
nand UO_327 (O_327,N_2820,N_2828);
and UO_328 (O_328,N_2618,N_2498);
and UO_329 (O_329,N_2540,N_2747);
nor UO_330 (O_330,N_2940,N_2598);
nand UO_331 (O_331,N_2851,N_2614);
nand UO_332 (O_332,N_2809,N_2683);
nor UO_333 (O_333,N_2464,N_2917);
and UO_334 (O_334,N_2933,N_2885);
nand UO_335 (O_335,N_2608,N_2589);
xor UO_336 (O_336,N_2552,N_2476);
or UO_337 (O_337,N_2439,N_2423);
or UO_338 (O_338,N_2970,N_2666);
or UO_339 (O_339,N_2945,N_2850);
and UO_340 (O_340,N_2859,N_2627);
nand UO_341 (O_341,N_2867,N_2691);
nor UO_342 (O_342,N_2712,N_2523);
and UO_343 (O_343,N_2554,N_2881);
and UO_344 (O_344,N_2823,N_2478);
nand UO_345 (O_345,N_2718,N_2498);
nand UO_346 (O_346,N_2939,N_2700);
or UO_347 (O_347,N_2481,N_2931);
nand UO_348 (O_348,N_2731,N_2911);
nor UO_349 (O_349,N_2555,N_2593);
or UO_350 (O_350,N_2906,N_2446);
nand UO_351 (O_351,N_2506,N_2851);
and UO_352 (O_352,N_2936,N_2500);
or UO_353 (O_353,N_2971,N_2612);
nor UO_354 (O_354,N_2939,N_2955);
nor UO_355 (O_355,N_2861,N_2543);
nor UO_356 (O_356,N_2781,N_2800);
nand UO_357 (O_357,N_2712,N_2807);
and UO_358 (O_358,N_2790,N_2664);
and UO_359 (O_359,N_2501,N_2867);
nand UO_360 (O_360,N_2536,N_2490);
nor UO_361 (O_361,N_2972,N_2920);
and UO_362 (O_362,N_2435,N_2489);
nand UO_363 (O_363,N_2974,N_2474);
nor UO_364 (O_364,N_2613,N_2960);
nor UO_365 (O_365,N_2477,N_2900);
and UO_366 (O_366,N_2444,N_2753);
nor UO_367 (O_367,N_2659,N_2633);
or UO_368 (O_368,N_2546,N_2480);
nor UO_369 (O_369,N_2610,N_2652);
nor UO_370 (O_370,N_2575,N_2673);
and UO_371 (O_371,N_2469,N_2850);
nor UO_372 (O_372,N_2723,N_2689);
or UO_373 (O_373,N_2766,N_2780);
nor UO_374 (O_374,N_2501,N_2445);
and UO_375 (O_375,N_2943,N_2477);
and UO_376 (O_376,N_2756,N_2608);
nand UO_377 (O_377,N_2424,N_2985);
nor UO_378 (O_378,N_2736,N_2915);
or UO_379 (O_379,N_2639,N_2755);
or UO_380 (O_380,N_2453,N_2735);
nand UO_381 (O_381,N_2485,N_2866);
and UO_382 (O_382,N_2777,N_2917);
or UO_383 (O_383,N_2426,N_2775);
nand UO_384 (O_384,N_2848,N_2516);
nor UO_385 (O_385,N_2911,N_2975);
and UO_386 (O_386,N_2581,N_2760);
xor UO_387 (O_387,N_2729,N_2762);
nor UO_388 (O_388,N_2602,N_2982);
or UO_389 (O_389,N_2856,N_2943);
nand UO_390 (O_390,N_2742,N_2525);
and UO_391 (O_391,N_2952,N_2887);
nand UO_392 (O_392,N_2577,N_2909);
nor UO_393 (O_393,N_2615,N_2551);
nor UO_394 (O_394,N_2628,N_2664);
nor UO_395 (O_395,N_2629,N_2789);
and UO_396 (O_396,N_2637,N_2615);
and UO_397 (O_397,N_2419,N_2457);
nand UO_398 (O_398,N_2757,N_2512);
nor UO_399 (O_399,N_2580,N_2941);
or UO_400 (O_400,N_2888,N_2856);
and UO_401 (O_401,N_2887,N_2815);
or UO_402 (O_402,N_2426,N_2731);
or UO_403 (O_403,N_2693,N_2482);
and UO_404 (O_404,N_2849,N_2559);
or UO_405 (O_405,N_2929,N_2529);
nor UO_406 (O_406,N_2538,N_2923);
nand UO_407 (O_407,N_2947,N_2432);
and UO_408 (O_408,N_2516,N_2939);
and UO_409 (O_409,N_2895,N_2457);
or UO_410 (O_410,N_2596,N_2567);
or UO_411 (O_411,N_2748,N_2781);
and UO_412 (O_412,N_2936,N_2614);
nor UO_413 (O_413,N_2709,N_2920);
nor UO_414 (O_414,N_2975,N_2558);
or UO_415 (O_415,N_2786,N_2933);
nand UO_416 (O_416,N_2972,N_2463);
nor UO_417 (O_417,N_2767,N_2944);
nand UO_418 (O_418,N_2817,N_2572);
nand UO_419 (O_419,N_2779,N_2701);
or UO_420 (O_420,N_2831,N_2716);
nor UO_421 (O_421,N_2811,N_2457);
or UO_422 (O_422,N_2668,N_2596);
nand UO_423 (O_423,N_2407,N_2496);
and UO_424 (O_424,N_2643,N_2429);
nand UO_425 (O_425,N_2883,N_2780);
xnor UO_426 (O_426,N_2929,N_2800);
nand UO_427 (O_427,N_2819,N_2693);
and UO_428 (O_428,N_2993,N_2567);
nand UO_429 (O_429,N_2971,N_2553);
or UO_430 (O_430,N_2507,N_2620);
and UO_431 (O_431,N_2622,N_2843);
nor UO_432 (O_432,N_2400,N_2538);
and UO_433 (O_433,N_2721,N_2886);
nor UO_434 (O_434,N_2673,N_2927);
nand UO_435 (O_435,N_2961,N_2408);
and UO_436 (O_436,N_2533,N_2560);
and UO_437 (O_437,N_2893,N_2453);
nand UO_438 (O_438,N_2444,N_2759);
nand UO_439 (O_439,N_2994,N_2806);
and UO_440 (O_440,N_2808,N_2876);
and UO_441 (O_441,N_2781,N_2866);
and UO_442 (O_442,N_2909,N_2748);
nor UO_443 (O_443,N_2838,N_2997);
nor UO_444 (O_444,N_2505,N_2848);
or UO_445 (O_445,N_2787,N_2559);
and UO_446 (O_446,N_2514,N_2728);
nand UO_447 (O_447,N_2594,N_2785);
or UO_448 (O_448,N_2598,N_2680);
and UO_449 (O_449,N_2493,N_2418);
nand UO_450 (O_450,N_2660,N_2566);
or UO_451 (O_451,N_2790,N_2523);
nand UO_452 (O_452,N_2509,N_2981);
and UO_453 (O_453,N_2894,N_2973);
or UO_454 (O_454,N_2772,N_2949);
and UO_455 (O_455,N_2976,N_2447);
or UO_456 (O_456,N_2818,N_2535);
nor UO_457 (O_457,N_2915,N_2920);
nand UO_458 (O_458,N_2409,N_2462);
and UO_459 (O_459,N_2888,N_2831);
nor UO_460 (O_460,N_2808,N_2834);
nand UO_461 (O_461,N_2454,N_2895);
nor UO_462 (O_462,N_2527,N_2492);
and UO_463 (O_463,N_2719,N_2815);
nand UO_464 (O_464,N_2465,N_2632);
and UO_465 (O_465,N_2487,N_2415);
nor UO_466 (O_466,N_2540,N_2864);
nor UO_467 (O_467,N_2712,N_2619);
and UO_468 (O_468,N_2904,N_2930);
and UO_469 (O_469,N_2843,N_2675);
nor UO_470 (O_470,N_2983,N_2924);
and UO_471 (O_471,N_2977,N_2507);
and UO_472 (O_472,N_2868,N_2947);
or UO_473 (O_473,N_2882,N_2480);
nand UO_474 (O_474,N_2538,N_2933);
nand UO_475 (O_475,N_2439,N_2738);
nor UO_476 (O_476,N_2751,N_2514);
nand UO_477 (O_477,N_2858,N_2648);
or UO_478 (O_478,N_2478,N_2786);
and UO_479 (O_479,N_2865,N_2615);
nor UO_480 (O_480,N_2994,N_2473);
nor UO_481 (O_481,N_2857,N_2459);
nor UO_482 (O_482,N_2744,N_2472);
nor UO_483 (O_483,N_2805,N_2614);
nand UO_484 (O_484,N_2775,N_2771);
and UO_485 (O_485,N_2529,N_2579);
nand UO_486 (O_486,N_2965,N_2683);
and UO_487 (O_487,N_2979,N_2680);
and UO_488 (O_488,N_2717,N_2518);
or UO_489 (O_489,N_2415,N_2717);
nand UO_490 (O_490,N_2476,N_2533);
nand UO_491 (O_491,N_2460,N_2849);
or UO_492 (O_492,N_2637,N_2568);
and UO_493 (O_493,N_2774,N_2958);
nor UO_494 (O_494,N_2707,N_2800);
or UO_495 (O_495,N_2798,N_2484);
nor UO_496 (O_496,N_2599,N_2677);
and UO_497 (O_497,N_2429,N_2519);
xnor UO_498 (O_498,N_2464,N_2646);
and UO_499 (O_499,N_2643,N_2693);
endmodule