module basic_500_3000_500_40_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_471,In_97);
xnor U1 (N_1,In_53,In_461);
nand U2 (N_2,In_380,In_98);
nand U3 (N_3,In_448,In_379);
nor U4 (N_4,In_355,In_356);
nor U5 (N_5,In_319,In_308);
nand U6 (N_6,In_101,In_124);
nand U7 (N_7,In_298,In_175);
and U8 (N_8,In_77,In_72);
or U9 (N_9,In_20,In_265);
nand U10 (N_10,In_40,In_107);
and U11 (N_11,In_6,In_256);
nor U12 (N_12,In_400,In_62);
nor U13 (N_13,In_132,In_499);
and U14 (N_14,In_34,In_223);
or U15 (N_15,In_146,In_255);
nor U16 (N_16,In_38,In_393);
nor U17 (N_17,In_164,In_83);
nand U18 (N_18,In_18,In_154);
nand U19 (N_19,In_392,In_15);
or U20 (N_20,In_197,In_160);
or U21 (N_21,In_496,In_424);
nand U22 (N_22,In_112,In_188);
and U23 (N_23,In_231,In_141);
xnor U24 (N_24,In_269,In_353);
nor U25 (N_25,In_486,In_429);
xnor U26 (N_26,In_252,In_297);
xnor U27 (N_27,In_19,In_365);
or U28 (N_28,In_236,In_158);
and U29 (N_29,In_17,In_412);
nand U30 (N_30,In_117,In_389);
xnor U31 (N_31,In_456,In_162);
and U32 (N_32,In_425,In_327);
and U33 (N_33,In_396,In_428);
nor U34 (N_34,In_320,In_270);
xnor U35 (N_35,In_364,In_470);
or U36 (N_36,In_481,In_90);
and U37 (N_37,In_346,In_55);
xnor U38 (N_38,In_415,In_94);
xnor U39 (N_39,In_445,In_488);
and U40 (N_40,In_113,In_23);
or U41 (N_41,In_86,In_193);
nor U42 (N_42,In_221,In_292);
xnor U43 (N_43,In_64,In_63);
nand U44 (N_44,In_110,In_242);
xor U45 (N_45,In_174,In_430);
and U46 (N_46,In_244,In_225);
nand U47 (N_47,In_479,In_247);
or U48 (N_48,In_281,In_120);
or U49 (N_49,In_105,In_200);
nand U50 (N_50,In_167,In_119);
and U51 (N_51,In_104,In_33);
nand U52 (N_52,In_227,In_378);
or U53 (N_53,In_84,In_208);
nand U54 (N_54,In_21,In_377);
or U55 (N_55,In_280,In_368);
nor U56 (N_56,In_182,In_3);
xnor U57 (N_57,In_142,In_16);
and U58 (N_58,In_246,In_135);
nand U59 (N_59,In_226,In_65);
nand U60 (N_60,In_399,In_183);
xnor U61 (N_61,In_59,In_358);
or U62 (N_62,In_68,In_12);
or U63 (N_63,In_152,In_279);
and U64 (N_64,In_264,In_395);
xor U65 (N_65,In_230,In_274);
nand U66 (N_66,In_473,In_345);
and U67 (N_67,In_204,In_179);
nand U68 (N_68,In_70,In_422);
nor U69 (N_69,In_307,In_245);
nand U70 (N_70,In_491,In_317);
or U71 (N_71,In_439,In_216);
xnor U72 (N_72,In_166,In_344);
nand U73 (N_73,In_10,In_219);
nor U74 (N_74,In_293,In_277);
and U75 (N_75,In_258,N_10);
nand U76 (N_76,In_35,In_8);
xnor U77 (N_77,In_420,N_43);
or U78 (N_78,In_433,In_138);
or U79 (N_79,In_478,In_447);
nor U80 (N_80,In_139,In_347);
nor U81 (N_81,In_343,In_272);
or U82 (N_82,In_467,N_52);
nand U83 (N_83,In_390,N_24);
or U84 (N_84,In_44,In_351);
and U85 (N_85,In_143,In_100);
xor U86 (N_86,In_176,N_47);
and U87 (N_87,In_335,In_475);
nand U88 (N_88,In_39,In_386);
or U89 (N_89,In_432,In_304);
xnor U90 (N_90,In_76,In_81);
or U91 (N_91,In_26,N_27);
xnor U92 (N_92,In_338,In_29);
or U93 (N_93,In_329,N_21);
or U94 (N_94,In_214,In_136);
xnor U95 (N_95,In_14,In_66);
or U96 (N_96,In_299,In_106);
xor U97 (N_97,In_383,In_462);
or U98 (N_98,In_318,In_239);
nand U99 (N_99,In_212,N_63);
xor U100 (N_100,In_257,In_263);
or U101 (N_101,In_178,In_248);
nand U102 (N_102,In_238,In_476);
nand U103 (N_103,In_91,N_48);
nor U104 (N_104,N_29,N_20);
and U105 (N_105,In_454,In_303);
nand U106 (N_106,In_401,In_170);
nor U107 (N_107,In_316,In_144);
xnor U108 (N_108,In_67,In_87);
nand U109 (N_109,In_131,In_349);
or U110 (N_110,In_122,In_165);
and U111 (N_111,In_275,In_213);
nor U112 (N_112,In_410,In_13);
or U113 (N_113,In_427,In_434);
nor U114 (N_114,In_169,In_443);
xor U115 (N_115,In_357,In_177);
nor U116 (N_116,In_235,In_171);
nor U117 (N_117,In_133,In_321);
xnor U118 (N_118,In_184,In_114);
nor U119 (N_119,N_58,N_2);
xor U120 (N_120,In_46,In_331);
or U121 (N_121,In_421,N_8);
nand U122 (N_122,In_49,N_60);
nor U123 (N_123,In_123,In_237);
nand U124 (N_124,In_134,In_414);
xnor U125 (N_125,In_56,In_294);
and U126 (N_126,In_283,In_449);
nor U127 (N_127,In_472,In_350);
and U128 (N_128,In_373,In_157);
xnor U129 (N_129,In_352,In_41);
xor U130 (N_130,In_376,In_147);
nand U131 (N_131,In_480,In_413);
or U132 (N_132,In_103,In_334);
nand U133 (N_133,In_145,In_498);
nor U134 (N_134,N_0,In_451);
xnor U135 (N_135,In_69,In_385);
nand U136 (N_136,In_116,In_27);
nor U137 (N_137,In_28,In_375);
xnor U138 (N_138,N_41,In_42);
and U139 (N_139,In_191,In_418);
or U140 (N_140,N_67,In_95);
or U141 (N_141,In_58,In_228);
xnor U142 (N_142,In_232,In_2);
and U143 (N_143,In_423,In_207);
xnor U144 (N_144,In_79,N_50);
xnor U145 (N_145,In_489,In_52);
and U146 (N_146,N_70,In_394);
or U147 (N_147,In_286,In_465);
nor U148 (N_148,In_487,In_111);
or U149 (N_149,In_115,In_366);
xnor U150 (N_150,In_306,In_71);
or U151 (N_151,In_497,In_267);
xnor U152 (N_152,In_495,In_431);
and U153 (N_153,N_46,In_9);
nor U154 (N_154,N_130,In_458);
xnor U155 (N_155,In_173,N_42);
nand U156 (N_156,N_113,In_483);
or U157 (N_157,In_240,In_253);
xor U158 (N_158,In_450,In_367);
or U159 (N_159,In_382,In_397);
and U160 (N_160,In_436,In_140);
xnor U161 (N_161,In_354,N_40);
or U162 (N_162,In_322,In_45);
nor U163 (N_163,N_106,In_150);
xnor U164 (N_164,In_201,N_116);
or U165 (N_165,N_6,N_31);
and U166 (N_166,In_159,N_51);
and U167 (N_167,In_61,In_477);
or U168 (N_168,N_16,In_282);
and U169 (N_169,In_254,N_139);
or U170 (N_170,In_296,N_69);
nor U171 (N_171,N_120,In_36);
xnor U172 (N_172,N_57,N_38);
or U173 (N_173,N_128,In_57);
nand U174 (N_174,In_129,In_340);
and U175 (N_175,N_1,In_339);
and U176 (N_176,In_305,In_371);
xor U177 (N_177,In_287,N_115);
xnor U178 (N_178,N_81,In_5);
nand U179 (N_179,In_215,In_222);
nand U180 (N_180,In_342,N_98);
nand U181 (N_181,N_99,In_192);
and U182 (N_182,In_493,In_217);
nor U183 (N_183,N_118,In_468);
xor U184 (N_184,N_92,N_97);
nand U185 (N_185,In_315,N_17);
and U186 (N_186,N_64,N_5);
and U187 (N_187,In_126,In_348);
or U188 (N_188,N_103,In_407);
or U189 (N_189,In_250,In_388);
nand U190 (N_190,N_143,N_33);
nor U191 (N_191,N_7,In_234);
and U192 (N_192,In_130,In_1);
xnor U193 (N_193,N_62,In_482);
or U194 (N_194,N_137,N_91);
or U195 (N_195,N_124,In_446);
or U196 (N_196,In_336,In_220);
or U197 (N_197,In_198,In_474);
and U198 (N_198,In_73,N_77);
and U199 (N_199,In_185,In_440);
nand U200 (N_200,N_14,N_121);
nor U201 (N_201,In_459,In_205);
or U202 (N_202,In_466,N_100);
nand U203 (N_203,N_66,In_121);
nand U204 (N_204,In_54,In_241);
or U205 (N_205,N_148,In_455);
nand U206 (N_206,In_300,In_47);
xnor U207 (N_207,In_156,In_374);
nor U208 (N_208,N_68,N_19);
or U209 (N_209,In_469,N_127);
nor U210 (N_210,In_289,N_26);
or U211 (N_211,N_30,In_404);
nor U212 (N_212,N_75,N_104);
and U213 (N_213,N_12,N_3);
or U214 (N_214,N_83,In_22);
xnor U215 (N_215,N_56,N_78);
and U216 (N_216,In_80,N_35);
and U217 (N_217,N_126,In_332);
and U218 (N_218,In_43,In_271);
or U219 (N_219,N_108,In_288);
xor U220 (N_220,N_133,N_119);
nand U221 (N_221,In_457,N_144);
xnor U222 (N_222,In_259,In_312);
xnor U223 (N_223,In_333,In_437);
nor U224 (N_224,In_261,In_187);
nor U225 (N_225,In_359,In_24);
and U226 (N_226,N_28,N_150);
nand U227 (N_227,In_416,N_192);
xnor U228 (N_228,N_175,In_381);
xnor U229 (N_229,In_196,In_361);
or U230 (N_230,In_209,In_181);
nand U231 (N_231,N_190,In_309);
nor U232 (N_232,In_484,In_278);
nor U233 (N_233,N_138,In_224);
xnor U234 (N_234,N_72,In_118);
or U235 (N_235,N_90,N_125);
nand U236 (N_236,N_188,In_453);
nor U237 (N_237,In_11,N_209);
nand U238 (N_238,N_171,N_217);
xor U239 (N_239,N_193,In_202);
nand U240 (N_240,In_60,In_92);
nor U241 (N_241,N_155,In_89);
xnor U242 (N_242,In_464,N_179);
xnor U243 (N_243,N_15,N_87);
nor U244 (N_244,In_243,N_189);
and U245 (N_245,N_154,In_441);
and U246 (N_246,In_444,In_324);
or U247 (N_247,In_108,N_22);
xor U248 (N_248,N_37,N_145);
and U249 (N_249,N_55,In_328);
xnor U250 (N_250,N_210,N_167);
xor U251 (N_251,N_13,In_51);
nand U252 (N_252,In_128,N_214);
and U253 (N_253,In_85,N_84);
xnor U254 (N_254,N_95,In_326);
or U255 (N_255,N_174,In_249);
nand U256 (N_256,N_219,In_161);
xor U257 (N_257,N_76,N_177);
and U258 (N_258,N_39,In_7);
nor U259 (N_259,In_408,In_229);
nor U260 (N_260,In_180,In_251);
or U261 (N_261,N_223,In_284);
nand U262 (N_262,N_152,N_156);
nand U263 (N_263,N_94,N_169);
and U264 (N_264,N_122,N_135);
xnor U265 (N_265,In_194,In_463);
or U266 (N_266,In_302,N_82);
and U267 (N_267,N_186,In_4);
xnor U268 (N_268,N_172,In_30);
nor U269 (N_269,In_426,In_206);
and U270 (N_270,N_23,N_45);
or U271 (N_271,N_102,In_403);
xor U272 (N_272,N_224,In_337);
or U273 (N_273,N_65,N_149);
and U274 (N_274,In_50,In_25);
or U275 (N_275,In_262,N_25);
or U276 (N_276,N_197,In_93);
and U277 (N_277,N_85,N_221);
and U278 (N_278,In_301,In_78);
and U279 (N_279,N_178,In_273);
and U280 (N_280,N_134,In_186);
or U281 (N_281,In_37,N_153);
and U282 (N_282,N_140,In_411);
and U283 (N_283,In_266,In_387);
nand U284 (N_284,N_18,In_363);
xor U285 (N_285,N_61,In_360);
or U286 (N_286,N_213,N_205);
nand U287 (N_287,N_117,N_142);
nor U288 (N_288,N_206,N_114);
and U289 (N_289,In_492,In_460);
or U290 (N_290,N_129,In_153);
or U291 (N_291,In_406,N_123);
and U292 (N_292,N_89,N_44);
and U293 (N_293,In_88,In_438);
or U294 (N_294,In_452,N_105);
and U295 (N_295,N_191,In_137);
or U296 (N_296,In_211,N_36);
xor U297 (N_297,N_200,N_161);
or U298 (N_298,N_173,N_162);
nand U299 (N_299,N_147,In_260);
nor U300 (N_300,N_146,N_255);
or U301 (N_301,N_215,N_227);
xnor U302 (N_302,N_298,N_234);
xnor U303 (N_303,N_112,N_246);
nor U304 (N_304,N_244,N_159);
nor U305 (N_305,In_370,In_310);
or U306 (N_306,In_311,N_53);
and U307 (N_307,N_208,N_262);
xnor U308 (N_308,In_74,N_252);
nor U309 (N_309,N_131,In_151);
or U310 (N_310,N_218,In_405);
or U311 (N_311,N_254,N_243);
nand U312 (N_312,In_190,In_314);
or U313 (N_313,N_277,In_485);
and U314 (N_314,In_494,In_127);
nor U315 (N_315,N_107,N_198);
nand U316 (N_316,N_250,N_185);
nor U317 (N_317,N_73,In_82);
or U318 (N_318,N_261,N_9);
or U319 (N_319,N_279,N_34);
nor U320 (N_320,In_168,N_111);
nand U321 (N_321,N_222,N_291);
xor U322 (N_322,N_168,N_212);
nor U323 (N_323,In_295,N_11);
xnor U324 (N_324,N_253,In_48);
xnor U325 (N_325,N_267,In_398);
or U326 (N_326,N_54,N_204);
or U327 (N_327,N_225,In_233);
and U328 (N_328,N_180,In_409);
nand U329 (N_329,N_59,N_258);
nor U330 (N_330,In_323,N_290);
xor U331 (N_331,N_226,In_313);
or U332 (N_332,N_271,In_442);
or U333 (N_333,N_293,N_266);
nand U334 (N_334,In_325,In_341);
and U335 (N_335,N_249,In_210);
nand U336 (N_336,N_264,N_201);
or U337 (N_337,In_435,N_287);
or U338 (N_338,N_182,N_229);
or U339 (N_339,N_141,In_163);
nand U340 (N_340,In_419,N_211);
or U341 (N_341,N_181,In_330);
nor U342 (N_342,N_288,N_248);
xnor U343 (N_343,N_158,N_284);
xor U344 (N_344,In_372,In_0);
and U345 (N_345,N_196,N_269);
or U346 (N_346,In_218,N_263);
nand U347 (N_347,In_32,N_282);
or U348 (N_348,N_136,N_260);
nand U349 (N_349,N_259,N_203);
or U350 (N_350,N_183,N_207);
xor U351 (N_351,In_96,N_166);
or U352 (N_352,N_285,N_170);
and U353 (N_353,N_110,N_245);
xor U354 (N_354,N_251,In_268);
xnor U355 (N_355,N_79,In_149);
nor U356 (N_356,N_299,N_231);
and U357 (N_357,N_93,In_291);
xor U358 (N_358,N_151,N_195);
and U359 (N_359,N_278,N_74);
or U360 (N_360,N_132,In_195);
xor U361 (N_361,N_4,In_490);
xor U362 (N_362,In_369,N_236);
nor U363 (N_363,In_362,N_165);
nor U364 (N_364,In_285,In_417);
and U365 (N_365,N_160,N_164);
and U366 (N_366,N_86,N_199);
nor U367 (N_367,N_296,N_272);
nand U368 (N_368,N_71,N_295);
nor U369 (N_369,In_276,N_157);
and U370 (N_370,In_155,N_256);
or U371 (N_371,N_235,N_265);
or U372 (N_372,N_292,In_31);
xnor U373 (N_373,In_203,N_233);
or U374 (N_374,N_281,N_280);
or U375 (N_375,N_366,N_335);
and U376 (N_376,N_317,N_333);
xor U377 (N_377,N_300,N_276);
or U378 (N_378,N_220,N_228);
xor U379 (N_379,N_237,N_216);
xnor U380 (N_380,N_247,N_321);
nor U381 (N_381,In_290,N_325);
and U382 (N_382,N_242,N_313);
xor U383 (N_383,N_320,N_338);
nand U384 (N_384,N_374,In_199);
or U385 (N_385,N_273,N_314);
and U386 (N_386,N_337,N_329);
xor U387 (N_387,N_289,N_328);
or U388 (N_388,N_326,N_257);
nor U389 (N_389,In_172,N_354);
or U390 (N_390,N_306,N_318);
nor U391 (N_391,N_348,N_294);
or U392 (N_392,N_372,N_330);
nor U393 (N_393,N_304,N_315);
nand U394 (N_394,N_96,N_240);
xor U395 (N_395,N_80,N_283);
nor U396 (N_396,N_344,N_305);
nand U397 (N_397,N_230,N_49);
xnor U398 (N_398,N_238,N_367);
nand U399 (N_399,N_343,N_345);
or U400 (N_400,N_322,N_327);
nor U401 (N_401,N_349,N_324);
or U402 (N_402,N_308,N_307);
or U403 (N_403,N_297,In_99);
and U404 (N_404,N_303,N_163);
nand U405 (N_405,N_301,In_75);
or U406 (N_406,N_339,N_350);
nor U407 (N_407,N_309,In_109);
or U408 (N_408,N_359,N_347);
and U409 (N_409,N_353,N_371);
or U410 (N_410,N_232,N_351);
nor U411 (N_411,N_176,N_336);
nand U412 (N_412,N_365,N_184);
nand U413 (N_413,N_239,In_125);
nand U414 (N_414,N_342,N_270);
nand U415 (N_415,N_241,In_102);
xor U416 (N_416,N_274,N_202);
xor U417 (N_417,N_355,N_361);
or U418 (N_418,N_332,N_358);
nand U419 (N_419,N_357,N_370);
nand U420 (N_420,N_316,N_352);
or U421 (N_421,N_268,N_362);
nand U422 (N_422,N_88,N_311);
xnor U423 (N_423,N_331,N_346);
and U424 (N_424,In_391,N_373);
and U425 (N_425,N_369,N_341);
xor U426 (N_426,N_319,In_148);
nor U427 (N_427,N_187,N_368);
or U428 (N_428,N_310,N_364);
xor U429 (N_429,In_189,In_402);
nand U430 (N_430,N_360,N_286);
xor U431 (N_431,N_275,N_356);
or U432 (N_432,N_101,N_194);
xnor U433 (N_433,N_312,N_363);
and U434 (N_434,N_109,N_323);
nand U435 (N_435,N_32,N_302);
and U436 (N_436,N_334,N_340);
and U437 (N_437,In_384,N_342);
and U438 (N_438,N_268,N_303);
nand U439 (N_439,N_311,N_347);
or U440 (N_440,N_202,N_342);
or U441 (N_441,N_316,N_348);
xor U442 (N_442,N_372,N_232);
xnor U443 (N_443,N_305,N_329);
or U444 (N_444,N_101,N_339);
or U445 (N_445,N_239,N_347);
nand U446 (N_446,In_75,N_351);
nor U447 (N_447,N_345,N_350);
nand U448 (N_448,N_187,N_372);
nand U449 (N_449,In_290,N_328);
xnor U450 (N_450,N_411,N_405);
nand U451 (N_451,N_439,N_418);
nor U452 (N_452,N_429,N_426);
xnor U453 (N_453,N_432,N_392);
nor U454 (N_454,N_416,N_384);
and U455 (N_455,N_417,N_383);
or U456 (N_456,N_391,N_400);
xnor U457 (N_457,N_395,N_427);
nand U458 (N_458,N_385,N_413);
nand U459 (N_459,N_423,N_397);
and U460 (N_460,N_446,N_390);
nor U461 (N_461,N_447,N_376);
and U462 (N_462,N_377,N_424);
nand U463 (N_463,N_394,N_403);
and U464 (N_464,N_441,N_382);
and U465 (N_465,N_420,N_409);
nor U466 (N_466,N_388,N_379);
xnor U467 (N_467,N_414,N_437);
or U468 (N_468,N_378,N_375);
or U469 (N_469,N_444,N_407);
xnor U470 (N_470,N_440,N_415);
nor U471 (N_471,N_422,N_419);
or U472 (N_472,N_386,N_436);
or U473 (N_473,N_402,N_421);
nor U474 (N_474,N_381,N_438);
and U475 (N_475,N_410,N_389);
or U476 (N_476,N_408,N_406);
nand U477 (N_477,N_399,N_443);
or U478 (N_478,N_412,N_431);
nor U479 (N_479,N_398,N_425);
xnor U480 (N_480,N_434,N_393);
and U481 (N_481,N_449,N_448);
xor U482 (N_482,N_442,N_445);
or U483 (N_483,N_387,N_401);
nand U484 (N_484,N_380,N_396);
nand U485 (N_485,N_433,N_435);
or U486 (N_486,N_430,N_404);
or U487 (N_487,N_428,N_397);
or U488 (N_488,N_416,N_434);
or U489 (N_489,N_395,N_398);
and U490 (N_490,N_415,N_392);
nor U491 (N_491,N_415,N_405);
or U492 (N_492,N_421,N_405);
or U493 (N_493,N_403,N_425);
xnor U494 (N_494,N_442,N_430);
or U495 (N_495,N_413,N_441);
nor U496 (N_496,N_398,N_443);
xor U497 (N_497,N_411,N_441);
xnor U498 (N_498,N_405,N_403);
nor U499 (N_499,N_387,N_410);
nor U500 (N_500,N_382,N_444);
or U501 (N_501,N_448,N_399);
nand U502 (N_502,N_440,N_402);
nor U503 (N_503,N_407,N_423);
or U504 (N_504,N_394,N_395);
nor U505 (N_505,N_446,N_382);
nor U506 (N_506,N_409,N_402);
xnor U507 (N_507,N_427,N_429);
or U508 (N_508,N_444,N_413);
or U509 (N_509,N_411,N_418);
nand U510 (N_510,N_449,N_394);
or U511 (N_511,N_424,N_392);
xnor U512 (N_512,N_385,N_440);
nand U513 (N_513,N_444,N_441);
nor U514 (N_514,N_427,N_396);
nor U515 (N_515,N_405,N_442);
or U516 (N_516,N_428,N_439);
or U517 (N_517,N_445,N_413);
and U518 (N_518,N_435,N_382);
nor U519 (N_519,N_447,N_378);
and U520 (N_520,N_398,N_396);
xor U521 (N_521,N_421,N_382);
and U522 (N_522,N_434,N_436);
and U523 (N_523,N_400,N_381);
nor U524 (N_524,N_444,N_376);
nand U525 (N_525,N_503,N_479);
nand U526 (N_526,N_450,N_502);
and U527 (N_527,N_456,N_495);
and U528 (N_528,N_510,N_470);
xnor U529 (N_529,N_457,N_455);
and U530 (N_530,N_474,N_480);
and U531 (N_531,N_461,N_499);
xor U532 (N_532,N_498,N_522);
and U533 (N_533,N_523,N_519);
nor U534 (N_534,N_467,N_452);
nand U535 (N_535,N_516,N_489);
and U536 (N_536,N_464,N_500);
and U537 (N_537,N_453,N_488);
nor U538 (N_538,N_496,N_486);
nand U539 (N_539,N_505,N_472);
nor U540 (N_540,N_492,N_459);
or U541 (N_541,N_484,N_478);
and U542 (N_542,N_515,N_477);
nor U543 (N_543,N_476,N_497);
or U544 (N_544,N_506,N_471);
and U545 (N_545,N_513,N_465);
xnor U546 (N_546,N_491,N_468);
or U547 (N_547,N_462,N_487);
xor U548 (N_548,N_518,N_520);
xnor U549 (N_549,N_509,N_469);
nand U550 (N_550,N_508,N_514);
and U551 (N_551,N_494,N_521);
nand U552 (N_552,N_463,N_501);
nor U553 (N_553,N_517,N_524);
and U554 (N_554,N_511,N_473);
and U555 (N_555,N_493,N_483);
and U556 (N_556,N_475,N_482);
and U557 (N_557,N_507,N_504);
or U558 (N_558,N_454,N_458);
or U559 (N_559,N_512,N_466);
nand U560 (N_560,N_451,N_485);
nand U561 (N_561,N_481,N_490);
or U562 (N_562,N_460,N_507);
nand U563 (N_563,N_474,N_485);
nand U564 (N_564,N_471,N_454);
nor U565 (N_565,N_511,N_484);
or U566 (N_566,N_456,N_494);
and U567 (N_567,N_452,N_482);
xor U568 (N_568,N_501,N_500);
nor U569 (N_569,N_490,N_480);
or U570 (N_570,N_502,N_488);
nand U571 (N_571,N_473,N_487);
and U572 (N_572,N_462,N_498);
or U573 (N_573,N_516,N_492);
nand U574 (N_574,N_502,N_492);
nand U575 (N_575,N_511,N_504);
nand U576 (N_576,N_493,N_475);
nor U577 (N_577,N_501,N_518);
nand U578 (N_578,N_514,N_505);
and U579 (N_579,N_497,N_452);
and U580 (N_580,N_524,N_486);
xnor U581 (N_581,N_493,N_472);
or U582 (N_582,N_458,N_502);
nand U583 (N_583,N_514,N_501);
or U584 (N_584,N_490,N_473);
xnor U585 (N_585,N_452,N_468);
and U586 (N_586,N_484,N_510);
xor U587 (N_587,N_501,N_511);
nor U588 (N_588,N_467,N_455);
and U589 (N_589,N_494,N_480);
or U590 (N_590,N_524,N_470);
or U591 (N_591,N_473,N_517);
nand U592 (N_592,N_515,N_473);
xor U593 (N_593,N_465,N_455);
or U594 (N_594,N_485,N_479);
xor U595 (N_595,N_465,N_524);
nand U596 (N_596,N_520,N_462);
or U597 (N_597,N_474,N_524);
nand U598 (N_598,N_484,N_523);
nand U599 (N_599,N_487,N_480);
and U600 (N_600,N_551,N_577);
xnor U601 (N_601,N_571,N_566);
and U602 (N_602,N_598,N_584);
nor U603 (N_603,N_587,N_583);
or U604 (N_604,N_592,N_550);
nor U605 (N_605,N_575,N_533);
or U606 (N_606,N_525,N_539);
or U607 (N_607,N_588,N_562);
xnor U608 (N_608,N_585,N_563);
nand U609 (N_609,N_579,N_530);
nand U610 (N_610,N_581,N_567);
or U611 (N_611,N_543,N_527);
nor U612 (N_612,N_560,N_559);
nor U613 (N_613,N_547,N_534);
nor U614 (N_614,N_558,N_596);
xor U615 (N_615,N_552,N_554);
and U616 (N_616,N_549,N_594);
nor U617 (N_617,N_576,N_580);
or U618 (N_618,N_564,N_572);
nand U619 (N_619,N_574,N_546);
and U620 (N_620,N_589,N_536);
and U621 (N_621,N_542,N_528);
or U622 (N_622,N_597,N_570);
nor U623 (N_623,N_529,N_553);
or U624 (N_624,N_593,N_537);
nand U625 (N_625,N_544,N_595);
nor U626 (N_626,N_541,N_591);
and U627 (N_627,N_535,N_582);
nor U628 (N_628,N_545,N_532);
nand U629 (N_629,N_540,N_561);
nor U630 (N_630,N_538,N_555);
nand U631 (N_631,N_526,N_578);
xnor U632 (N_632,N_586,N_531);
xor U633 (N_633,N_590,N_599);
xnor U634 (N_634,N_548,N_556);
and U635 (N_635,N_569,N_573);
nand U636 (N_636,N_568,N_557);
xor U637 (N_637,N_565,N_590);
or U638 (N_638,N_555,N_595);
xnor U639 (N_639,N_541,N_593);
or U640 (N_640,N_588,N_582);
or U641 (N_641,N_530,N_576);
and U642 (N_642,N_533,N_597);
xnor U643 (N_643,N_526,N_587);
nand U644 (N_644,N_559,N_588);
or U645 (N_645,N_567,N_527);
or U646 (N_646,N_595,N_572);
nor U647 (N_647,N_568,N_566);
and U648 (N_648,N_532,N_554);
nor U649 (N_649,N_534,N_538);
or U650 (N_650,N_596,N_535);
xor U651 (N_651,N_527,N_526);
nor U652 (N_652,N_547,N_535);
and U653 (N_653,N_527,N_596);
or U654 (N_654,N_566,N_547);
nand U655 (N_655,N_558,N_527);
nand U656 (N_656,N_536,N_533);
nand U657 (N_657,N_573,N_580);
nand U658 (N_658,N_587,N_537);
and U659 (N_659,N_535,N_549);
nor U660 (N_660,N_569,N_587);
and U661 (N_661,N_560,N_585);
nand U662 (N_662,N_536,N_586);
and U663 (N_663,N_553,N_573);
xnor U664 (N_664,N_525,N_557);
nand U665 (N_665,N_531,N_559);
and U666 (N_666,N_587,N_595);
or U667 (N_667,N_561,N_589);
nor U668 (N_668,N_592,N_534);
and U669 (N_669,N_573,N_570);
nor U670 (N_670,N_588,N_598);
or U671 (N_671,N_546,N_593);
and U672 (N_672,N_538,N_568);
and U673 (N_673,N_596,N_554);
nor U674 (N_674,N_588,N_541);
xor U675 (N_675,N_668,N_619);
xnor U676 (N_676,N_638,N_609);
nand U677 (N_677,N_602,N_644);
or U678 (N_678,N_648,N_606);
and U679 (N_679,N_600,N_640);
nor U680 (N_680,N_651,N_641);
xnor U681 (N_681,N_604,N_634);
or U682 (N_682,N_613,N_601);
nand U683 (N_683,N_616,N_653);
nand U684 (N_684,N_612,N_656);
or U685 (N_685,N_623,N_626);
and U686 (N_686,N_658,N_662);
nor U687 (N_687,N_660,N_642);
nand U688 (N_688,N_652,N_671);
or U689 (N_689,N_615,N_607);
nand U690 (N_690,N_643,N_614);
xnor U691 (N_691,N_639,N_620);
or U692 (N_692,N_674,N_666);
or U693 (N_693,N_608,N_637);
or U694 (N_694,N_654,N_631);
nor U695 (N_695,N_625,N_605);
nor U696 (N_696,N_627,N_617);
nand U697 (N_697,N_633,N_645);
nor U698 (N_698,N_670,N_610);
or U699 (N_699,N_611,N_657);
or U700 (N_700,N_635,N_650);
or U701 (N_701,N_630,N_647);
or U702 (N_702,N_624,N_636);
and U703 (N_703,N_663,N_646);
or U704 (N_704,N_664,N_661);
nor U705 (N_705,N_603,N_618);
or U706 (N_706,N_655,N_649);
nand U707 (N_707,N_667,N_629);
xor U708 (N_708,N_659,N_632);
nand U709 (N_709,N_672,N_673);
or U710 (N_710,N_622,N_665);
nand U711 (N_711,N_628,N_669);
nor U712 (N_712,N_621,N_613);
and U713 (N_713,N_632,N_615);
or U714 (N_714,N_630,N_640);
nand U715 (N_715,N_624,N_635);
nor U716 (N_716,N_613,N_657);
xnor U717 (N_717,N_663,N_618);
xor U718 (N_718,N_625,N_649);
nand U719 (N_719,N_613,N_630);
nand U720 (N_720,N_664,N_606);
or U721 (N_721,N_619,N_666);
and U722 (N_722,N_611,N_658);
and U723 (N_723,N_605,N_673);
or U724 (N_724,N_656,N_653);
and U725 (N_725,N_618,N_657);
and U726 (N_726,N_655,N_631);
nor U727 (N_727,N_653,N_632);
xor U728 (N_728,N_655,N_651);
or U729 (N_729,N_636,N_627);
nand U730 (N_730,N_606,N_666);
and U731 (N_731,N_673,N_630);
xor U732 (N_732,N_650,N_668);
xnor U733 (N_733,N_647,N_654);
nand U734 (N_734,N_635,N_653);
nand U735 (N_735,N_645,N_671);
xor U736 (N_736,N_625,N_611);
nor U737 (N_737,N_664,N_635);
xnor U738 (N_738,N_617,N_646);
xnor U739 (N_739,N_640,N_669);
nor U740 (N_740,N_602,N_632);
and U741 (N_741,N_662,N_646);
and U742 (N_742,N_605,N_633);
xnor U743 (N_743,N_648,N_612);
nand U744 (N_744,N_600,N_663);
xnor U745 (N_745,N_605,N_657);
or U746 (N_746,N_613,N_637);
xor U747 (N_747,N_633,N_642);
nand U748 (N_748,N_624,N_634);
and U749 (N_749,N_610,N_659);
xor U750 (N_750,N_702,N_716);
or U751 (N_751,N_734,N_740);
nor U752 (N_752,N_694,N_675);
xnor U753 (N_753,N_738,N_700);
xor U754 (N_754,N_709,N_717);
and U755 (N_755,N_723,N_744);
and U756 (N_756,N_699,N_685);
and U757 (N_757,N_728,N_726);
nor U758 (N_758,N_721,N_747);
nor U759 (N_759,N_695,N_707);
xor U760 (N_760,N_745,N_718);
nand U761 (N_761,N_746,N_682);
xnor U762 (N_762,N_749,N_686);
nor U763 (N_763,N_680,N_687);
nand U764 (N_764,N_698,N_711);
nand U765 (N_765,N_732,N_706);
xor U766 (N_766,N_715,N_724);
nand U767 (N_767,N_722,N_684);
nand U768 (N_768,N_708,N_679);
nand U769 (N_769,N_704,N_743);
and U770 (N_770,N_677,N_696);
and U771 (N_771,N_689,N_727);
or U772 (N_772,N_720,N_678);
xor U773 (N_773,N_737,N_733);
and U774 (N_774,N_705,N_741);
or U775 (N_775,N_693,N_714);
xnor U776 (N_776,N_701,N_710);
or U777 (N_777,N_692,N_739);
and U778 (N_778,N_681,N_736);
xnor U779 (N_779,N_731,N_735);
or U780 (N_780,N_703,N_729);
nor U781 (N_781,N_683,N_719);
and U782 (N_782,N_748,N_691);
nor U783 (N_783,N_697,N_742);
xnor U784 (N_784,N_690,N_725);
nor U785 (N_785,N_712,N_713);
nor U786 (N_786,N_676,N_730);
nor U787 (N_787,N_688,N_697);
or U788 (N_788,N_741,N_736);
xnor U789 (N_789,N_728,N_736);
nand U790 (N_790,N_742,N_720);
or U791 (N_791,N_688,N_734);
and U792 (N_792,N_743,N_696);
and U793 (N_793,N_735,N_700);
nor U794 (N_794,N_741,N_684);
and U795 (N_795,N_685,N_715);
xor U796 (N_796,N_732,N_748);
or U797 (N_797,N_722,N_699);
and U798 (N_798,N_676,N_746);
nor U799 (N_799,N_697,N_731);
or U800 (N_800,N_738,N_749);
xor U801 (N_801,N_741,N_698);
xnor U802 (N_802,N_681,N_698);
xor U803 (N_803,N_737,N_690);
and U804 (N_804,N_718,N_710);
nand U805 (N_805,N_717,N_707);
nor U806 (N_806,N_694,N_682);
nand U807 (N_807,N_709,N_682);
nand U808 (N_808,N_709,N_739);
nor U809 (N_809,N_675,N_679);
nor U810 (N_810,N_705,N_686);
xnor U811 (N_811,N_716,N_706);
nor U812 (N_812,N_719,N_736);
and U813 (N_813,N_701,N_747);
and U814 (N_814,N_706,N_720);
or U815 (N_815,N_723,N_748);
nand U816 (N_816,N_720,N_728);
nor U817 (N_817,N_706,N_708);
and U818 (N_818,N_727,N_741);
xor U819 (N_819,N_736,N_748);
xor U820 (N_820,N_743,N_711);
and U821 (N_821,N_718,N_740);
nand U822 (N_822,N_713,N_678);
and U823 (N_823,N_713,N_738);
or U824 (N_824,N_746,N_740);
xor U825 (N_825,N_777,N_754);
nand U826 (N_826,N_817,N_787);
nand U827 (N_827,N_803,N_776);
nor U828 (N_828,N_810,N_758);
nand U829 (N_829,N_797,N_761);
or U830 (N_830,N_792,N_790);
or U831 (N_831,N_768,N_812);
or U832 (N_832,N_808,N_769);
or U833 (N_833,N_814,N_757);
and U834 (N_834,N_794,N_766);
nor U835 (N_835,N_752,N_764);
nor U836 (N_836,N_785,N_760);
xor U837 (N_837,N_772,N_782);
or U838 (N_838,N_818,N_798);
xor U839 (N_839,N_813,N_774);
and U840 (N_840,N_802,N_793);
nor U841 (N_841,N_801,N_823);
nand U842 (N_842,N_784,N_789);
and U843 (N_843,N_775,N_816);
or U844 (N_844,N_750,N_778);
or U845 (N_845,N_796,N_751);
nand U846 (N_846,N_788,N_773);
and U847 (N_847,N_771,N_781);
nor U848 (N_848,N_804,N_806);
nor U849 (N_849,N_824,N_799);
or U850 (N_850,N_822,N_765);
xor U851 (N_851,N_809,N_759);
and U852 (N_852,N_795,N_786);
nand U853 (N_853,N_819,N_779);
xor U854 (N_854,N_756,N_800);
nor U855 (N_855,N_767,N_815);
nor U856 (N_856,N_821,N_807);
nor U857 (N_857,N_811,N_762);
nand U858 (N_858,N_780,N_791);
xnor U859 (N_859,N_805,N_755);
or U860 (N_860,N_770,N_753);
nand U861 (N_861,N_763,N_820);
or U862 (N_862,N_783,N_819);
or U863 (N_863,N_824,N_770);
and U864 (N_864,N_794,N_778);
or U865 (N_865,N_786,N_768);
or U866 (N_866,N_812,N_754);
nand U867 (N_867,N_824,N_821);
nand U868 (N_868,N_807,N_814);
nand U869 (N_869,N_824,N_778);
xnor U870 (N_870,N_781,N_769);
xor U871 (N_871,N_774,N_801);
xnor U872 (N_872,N_817,N_811);
or U873 (N_873,N_780,N_798);
nor U874 (N_874,N_809,N_818);
and U875 (N_875,N_816,N_758);
nand U876 (N_876,N_794,N_819);
nand U877 (N_877,N_782,N_757);
nor U878 (N_878,N_755,N_798);
and U879 (N_879,N_757,N_750);
and U880 (N_880,N_799,N_784);
nor U881 (N_881,N_809,N_821);
nand U882 (N_882,N_808,N_770);
and U883 (N_883,N_773,N_779);
nand U884 (N_884,N_810,N_753);
xor U885 (N_885,N_783,N_799);
and U886 (N_886,N_797,N_808);
or U887 (N_887,N_822,N_788);
nand U888 (N_888,N_812,N_777);
or U889 (N_889,N_760,N_824);
xor U890 (N_890,N_757,N_761);
nor U891 (N_891,N_764,N_767);
nand U892 (N_892,N_758,N_752);
or U893 (N_893,N_801,N_754);
nor U894 (N_894,N_786,N_773);
nor U895 (N_895,N_766,N_778);
and U896 (N_896,N_816,N_811);
nor U897 (N_897,N_801,N_798);
or U898 (N_898,N_810,N_802);
and U899 (N_899,N_813,N_807);
xor U900 (N_900,N_898,N_884);
and U901 (N_901,N_893,N_885);
and U902 (N_902,N_868,N_837);
or U903 (N_903,N_886,N_848);
nor U904 (N_904,N_858,N_840);
and U905 (N_905,N_883,N_859);
or U906 (N_906,N_846,N_829);
xnor U907 (N_907,N_861,N_851);
xor U908 (N_908,N_878,N_863);
nor U909 (N_909,N_891,N_879);
nor U910 (N_910,N_889,N_874);
nor U911 (N_911,N_890,N_852);
nand U912 (N_912,N_877,N_860);
or U913 (N_913,N_827,N_896);
xor U914 (N_914,N_841,N_867);
xor U915 (N_915,N_869,N_871);
nand U916 (N_916,N_880,N_873);
nand U917 (N_917,N_838,N_899);
and U918 (N_918,N_864,N_866);
and U919 (N_919,N_865,N_857);
nand U920 (N_920,N_881,N_854);
nand U921 (N_921,N_853,N_836);
and U922 (N_922,N_830,N_872);
and U923 (N_923,N_826,N_847);
nor U924 (N_924,N_850,N_882);
nor U925 (N_925,N_844,N_895);
nand U926 (N_926,N_870,N_876);
nor U927 (N_927,N_875,N_842);
nor U928 (N_928,N_828,N_845);
nor U929 (N_929,N_849,N_831);
xor U930 (N_930,N_856,N_888);
and U931 (N_931,N_855,N_825);
nor U932 (N_932,N_843,N_834);
or U933 (N_933,N_832,N_862);
xnor U934 (N_934,N_887,N_833);
nand U935 (N_935,N_897,N_892);
nand U936 (N_936,N_839,N_835);
and U937 (N_937,N_894,N_884);
nor U938 (N_938,N_878,N_899);
and U939 (N_939,N_869,N_876);
nor U940 (N_940,N_870,N_868);
and U941 (N_941,N_879,N_850);
or U942 (N_942,N_892,N_882);
xor U943 (N_943,N_841,N_865);
xor U944 (N_944,N_849,N_852);
and U945 (N_945,N_882,N_890);
and U946 (N_946,N_863,N_855);
or U947 (N_947,N_833,N_841);
nor U948 (N_948,N_890,N_870);
nand U949 (N_949,N_856,N_829);
and U950 (N_950,N_870,N_845);
nand U951 (N_951,N_873,N_869);
nand U952 (N_952,N_856,N_893);
nand U953 (N_953,N_846,N_868);
nor U954 (N_954,N_845,N_841);
and U955 (N_955,N_879,N_887);
xor U956 (N_956,N_827,N_898);
and U957 (N_957,N_833,N_865);
or U958 (N_958,N_879,N_871);
xnor U959 (N_959,N_862,N_873);
or U960 (N_960,N_868,N_836);
nand U961 (N_961,N_873,N_867);
xor U962 (N_962,N_899,N_857);
or U963 (N_963,N_881,N_884);
nor U964 (N_964,N_874,N_853);
nor U965 (N_965,N_873,N_858);
nand U966 (N_966,N_858,N_855);
and U967 (N_967,N_897,N_866);
or U968 (N_968,N_862,N_855);
nor U969 (N_969,N_835,N_856);
nor U970 (N_970,N_849,N_847);
or U971 (N_971,N_843,N_833);
xnor U972 (N_972,N_843,N_878);
xnor U973 (N_973,N_831,N_848);
nand U974 (N_974,N_893,N_859);
nor U975 (N_975,N_940,N_941);
or U976 (N_976,N_967,N_974);
nor U977 (N_977,N_954,N_957);
nand U978 (N_978,N_907,N_920);
nand U979 (N_979,N_928,N_903);
xor U980 (N_980,N_924,N_964);
nor U981 (N_981,N_962,N_926);
nor U982 (N_982,N_968,N_905);
xnor U983 (N_983,N_931,N_952);
nor U984 (N_984,N_919,N_972);
xnor U985 (N_985,N_916,N_901);
nor U986 (N_986,N_947,N_965);
or U987 (N_987,N_961,N_910);
nor U988 (N_988,N_922,N_960);
nand U989 (N_989,N_966,N_902);
and U990 (N_990,N_939,N_937);
nor U991 (N_991,N_904,N_900);
nand U992 (N_992,N_932,N_914);
nor U993 (N_993,N_963,N_930);
xnor U994 (N_994,N_945,N_948);
nor U995 (N_995,N_959,N_912);
or U996 (N_996,N_929,N_949);
nor U997 (N_997,N_918,N_927);
nand U998 (N_998,N_913,N_944);
xor U999 (N_999,N_970,N_933);
or U1000 (N_1000,N_955,N_971);
xnor U1001 (N_1001,N_943,N_951);
or U1002 (N_1002,N_946,N_909);
nand U1003 (N_1003,N_935,N_908);
or U1004 (N_1004,N_911,N_958);
or U1005 (N_1005,N_921,N_938);
nand U1006 (N_1006,N_973,N_934);
xnor U1007 (N_1007,N_950,N_942);
or U1008 (N_1008,N_956,N_969);
xor U1009 (N_1009,N_906,N_923);
xnor U1010 (N_1010,N_915,N_917);
or U1011 (N_1011,N_936,N_953);
or U1012 (N_1012,N_925,N_922);
and U1013 (N_1013,N_911,N_926);
xor U1014 (N_1014,N_940,N_929);
nor U1015 (N_1015,N_955,N_911);
nor U1016 (N_1016,N_962,N_947);
nor U1017 (N_1017,N_971,N_966);
nand U1018 (N_1018,N_934,N_972);
xnor U1019 (N_1019,N_917,N_900);
nand U1020 (N_1020,N_922,N_917);
xor U1021 (N_1021,N_905,N_913);
nor U1022 (N_1022,N_935,N_901);
and U1023 (N_1023,N_970,N_964);
and U1024 (N_1024,N_913,N_940);
or U1025 (N_1025,N_940,N_916);
nand U1026 (N_1026,N_912,N_972);
nand U1027 (N_1027,N_938,N_914);
nor U1028 (N_1028,N_951,N_939);
nand U1029 (N_1029,N_948,N_925);
or U1030 (N_1030,N_916,N_933);
and U1031 (N_1031,N_904,N_907);
nor U1032 (N_1032,N_937,N_907);
nand U1033 (N_1033,N_928,N_935);
nor U1034 (N_1034,N_937,N_962);
xnor U1035 (N_1035,N_906,N_900);
xor U1036 (N_1036,N_908,N_956);
nor U1037 (N_1037,N_956,N_973);
xnor U1038 (N_1038,N_971,N_938);
nand U1039 (N_1039,N_905,N_958);
or U1040 (N_1040,N_957,N_942);
nand U1041 (N_1041,N_954,N_970);
and U1042 (N_1042,N_925,N_903);
nand U1043 (N_1043,N_913,N_962);
nand U1044 (N_1044,N_930,N_940);
nand U1045 (N_1045,N_973,N_908);
or U1046 (N_1046,N_927,N_923);
nand U1047 (N_1047,N_914,N_931);
or U1048 (N_1048,N_920,N_923);
xor U1049 (N_1049,N_949,N_936);
or U1050 (N_1050,N_1001,N_1034);
and U1051 (N_1051,N_982,N_1006);
nor U1052 (N_1052,N_977,N_978);
nor U1053 (N_1053,N_1010,N_1008);
nor U1054 (N_1054,N_1035,N_981);
or U1055 (N_1055,N_1011,N_1007);
xnor U1056 (N_1056,N_983,N_1040);
or U1057 (N_1057,N_1030,N_1004);
nor U1058 (N_1058,N_1049,N_1017);
nand U1059 (N_1059,N_990,N_979);
or U1060 (N_1060,N_1039,N_1029);
nor U1061 (N_1061,N_1016,N_1043);
nor U1062 (N_1062,N_988,N_997);
or U1063 (N_1063,N_1037,N_1024);
nor U1064 (N_1064,N_985,N_995);
or U1065 (N_1065,N_1048,N_1031);
nand U1066 (N_1066,N_986,N_1041);
xnor U1067 (N_1067,N_1038,N_1005);
or U1068 (N_1068,N_1044,N_1012);
and U1069 (N_1069,N_1003,N_1014);
or U1070 (N_1070,N_1026,N_1021);
nand U1071 (N_1071,N_1032,N_1015);
nand U1072 (N_1072,N_1013,N_993);
xnor U1073 (N_1073,N_1027,N_1046);
nand U1074 (N_1074,N_994,N_1042);
or U1075 (N_1075,N_1033,N_987);
and U1076 (N_1076,N_1045,N_1020);
nor U1077 (N_1077,N_999,N_976);
xor U1078 (N_1078,N_996,N_1002);
nor U1079 (N_1079,N_991,N_1023);
and U1080 (N_1080,N_1018,N_980);
nor U1081 (N_1081,N_1022,N_984);
and U1082 (N_1082,N_989,N_1009);
xor U1083 (N_1083,N_998,N_1036);
nor U1084 (N_1084,N_1028,N_1019);
and U1085 (N_1085,N_1025,N_975);
and U1086 (N_1086,N_1047,N_992);
nor U1087 (N_1087,N_1000,N_1008);
nor U1088 (N_1088,N_995,N_993);
nand U1089 (N_1089,N_996,N_1031);
and U1090 (N_1090,N_1022,N_1034);
or U1091 (N_1091,N_1037,N_1043);
nor U1092 (N_1092,N_1017,N_1048);
and U1093 (N_1093,N_1024,N_1018);
or U1094 (N_1094,N_998,N_989);
and U1095 (N_1095,N_983,N_1009);
nand U1096 (N_1096,N_1027,N_1023);
xor U1097 (N_1097,N_1008,N_980);
nor U1098 (N_1098,N_1023,N_999);
and U1099 (N_1099,N_1013,N_1008);
nand U1100 (N_1100,N_989,N_988);
nand U1101 (N_1101,N_978,N_1035);
or U1102 (N_1102,N_1018,N_995);
nand U1103 (N_1103,N_999,N_1047);
and U1104 (N_1104,N_1023,N_1048);
xnor U1105 (N_1105,N_992,N_1036);
xnor U1106 (N_1106,N_978,N_984);
and U1107 (N_1107,N_1044,N_1029);
xor U1108 (N_1108,N_1010,N_1047);
nor U1109 (N_1109,N_987,N_1006);
and U1110 (N_1110,N_1006,N_1001);
and U1111 (N_1111,N_1047,N_1037);
and U1112 (N_1112,N_995,N_984);
xor U1113 (N_1113,N_1003,N_1039);
nand U1114 (N_1114,N_1015,N_1049);
or U1115 (N_1115,N_1018,N_1046);
or U1116 (N_1116,N_1003,N_986);
and U1117 (N_1117,N_1035,N_1034);
xnor U1118 (N_1118,N_1044,N_1019);
xor U1119 (N_1119,N_1032,N_1044);
xor U1120 (N_1120,N_994,N_982);
and U1121 (N_1121,N_1010,N_1029);
nor U1122 (N_1122,N_1003,N_979);
nand U1123 (N_1123,N_996,N_1037);
nand U1124 (N_1124,N_978,N_1029);
xnor U1125 (N_1125,N_1110,N_1109);
nand U1126 (N_1126,N_1077,N_1091);
or U1127 (N_1127,N_1074,N_1124);
nand U1128 (N_1128,N_1061,N_1100);
nor U1129 (N_1129,N_1057,N_1104);
nand U1130 (N_1130,N_1114,N_1055);
or U1131 (N_1131,N_1073,N_1087);
or U1132 (N_1132,N_1101,N_1076);
and U1133 (N_1133,N_1107,N_1081);
xor U1134 (N_1134,N_1070,N_1062);
xor U1135 (N_1135,N_1058,N_1112);
nor U1136 (N_1136,N_1095,N_1105);
nor U1137 (N_1137,N_1052,N_1096);
xor U1138 (N_1138,N_1050,N_1106);
and U1139 (N_1139,N_1118,N_1088);
xnor U1140 (N_1140,N_1066,N_1054);
and U1141 (N_1141,N_1060,N_1080);
or U1142 (N_1142,N_1085,N_1072);
nor U1143 (N_1143,N_1093,N_1084);
or U1144 (N_1144,N_1090,N_1068);
nor U1145 (N_1145,N_1078,N_1098);
nor U1146 (N_1146,N_1111,N_1115);
or U1147 (N_1147,N_1122,N_1071);
nor U1148 (N_1148,N_1092,N_1119);
nand U1149 (N_1149,N_1056,N_1075);
nand U1150 (N_1150,N_1099,N_1102);
nor U1151 (N_1151,N_1123,N_1086);
or U1152 (N_1152,N_1094,N_1121);
or U1153 (N_1153,N_1116,N_1083);
nor U1154 (N_1154,N_1097,N_1108);
nand U1155 (N_1155,N_1053,N_1120);
and U1156 (N_1156,N_1082,N_1063);
xor U1157 (N_1157,N_1051,N_1064);
and U1158 (N_1158,N_1067,N_1113);
xnor U1159 (N_1159,N_1065,N_1059);
nand U1160 (N_1160,N_1103,N_1079);
or U1161 (N_1161,N_1069,N_1089);
xor U1162 (N_1162,N_1117,N_1052);
or U1163 (N_1163,N_1121,N_1052);
nor U1164 (N_1164,N_1094,N_1058);
or U1165 (N_1165,N_1071,N_1072);
nor U1166 (N_1166,N_1093,N_1056);
or U1167 (N_1167,N_1056,N_1114);
nand U1168 (N_1168,N_1077,N_1095);
nor U1169 (N_1169,N_1109,N_1107);
nor U1170 (N_1170,N_1111,N_1093);
or U1171 (N_1171,N_1118,N_1111);
and U1172 (N_1172,N_1065,N_1069);
nand U1173 (N_1173,N_1116,N_1061);
xor U1174 (N_1174,N_1121,N_1071);
xnor U1175 (N_1175,N_1116,N_1115);
and U1176 (N_1176,N_1112,N_1077);
and U1177 (N_1177,N_1056,N_1078);
and U1178 (N_1178,N_1098,N_1050);
and U1179 (N_1179,N_1116,N_1058);
nand U1180 (N_1180,N_1120,N_1050);
xnor U1181 (N_1181,N_1096,N_1066);
and U1182 (N_1182,N_1059,N_1088);
or U1183 (N_1183,N_1103,N_1115);
and U1184 (N_1184,N_1117,N_1050);
nor U1185 (N_1185,N_1094,N_1085);
nor U1186 (N_1186,N_1072,N_1118);
or U1187 (N_1187,N_1111,N_1071);
and U1188 (N_1188,N_1079,N_1086);
and U1189 (N_1189,N_1113,N_1087);
xnor U1190 (N_1190,N_1075,N_1116);
or U1191 (N_1191,N_1090,N_1124);
nor U1192 (N_1192,N_1052,N_1068);
nor U1193 (N_1193,N_1084,N_1114);
nor U1194 (N_1194,N_1069,N_1119);
or U1195 (N_1195,N_1061,N_1081);
xnor U1196 (N_1196,N_1085,N_1084);
nand U1197 (N_1197,N_1094,N_1086);
or U1198 (N_1198,N_1079,N_1109);
or U1199 (N_1199,N_1111,N_1063);
xor U1200 (N_1200,N_1142,N_1147);
nand U1201 (N_1201,N_1156,N_1136);
nand U1202 (N_1202,N_1159,N_1199);
nor U1203 (N_1203,N_1198,N_1184);
nand U1204 (N_1204,N_1126,N_1133);
and U1205 (N_1205,N_1158,N_1146);
or U1206 (N_1206,N_1153,N_1144);
or U1207 (N_1207,N_1185,N_1154);
nor U1208 (N_1208,N_1188,N_1148);
nor U1209 (N_1209,N_1194,N_1173);
nor U1210 (N_1210,N_1130,N_1165);
nand U1211 (N_1211,N_1171,N_1138);
nand U1212 (N_1212,N_1191,N_1127);
or U1213 (N_1213,N_1190,N_1134);
nor U1214 (N_1214,N_1141,N_1167);
nor U1215 (N_1215,N_1183,N_1170);
and U1216 (N_1216,N_1187,N_1157);
xor U1217 (N_1217,N_1131,N_1161);
xnor U1218 (N_1218,N_1151,N_1140);
nand U1219 (N_1219,N_1145,N_1179);
or U1220 (N_1220,N_1177,N_1139);
nor U1221 (N_1221,N_1143,N_1128);
nor U1222 (N_1222,N_1168,N_1129);
or U1223 (N_1223,N_1192,N_1181);
xor U1224 (N_1224,N_1150,N_1166);
and U1225 (N_1225,N_1169,N_1160);
and U1226 (N_1226,N_1137,N_1125);
nand U1227 (N_1227,N_1149,N_1196);
xor U1228 (N_1228,N_1186,N_1164);
nor U1229 (N_1229,N_1178,N_1152);
or U1230 (N_1230,N_1195,N_1189);
nor U1231 (N_1231,N_1132,N_1175);
nor U1232 (N_1232,N_1162,N_1163);
or U1233 (N_1233,N_1174,N_1197);
or U1234 (N_1234,N_1180,N_1155);
nor U1235 (N_1235,N_1176,N_1193);
xor U1236 (N_1236,N_1135,N_1182);
xnor U1237 (N_1237,N_1172,N_1195);
or U1238 (N_1238,N_1163,N_1182);
nand U1239 (N_1239,N_1132,N_1176);
nor U1240 (N_1240,N_1128,N_1142);
xnor U1241 (N_1241,N_1171,N_1181);
or U1242 (N_1242,N_1142,N_1184);
nand U1243 (N_1243,N_1148,N_1157);
or U1244 (N_1244,N_1157,N_1189);
or U1245 (N_1245,N_1171,N_1140);
or U1246 (N_1246,N_1190,N_1197);
or U1247 (N_1247,N_1165,N_1151);
xor U1248 (N_1248,N_1167,N_1142);
and U1249 (N_1249,N_1143,N_1162);
nor U1250 (N_1250,N_1125,N_1196);
nand U1251 (N_1251,N_1186,N_1189);
and U1252 (N_1252,N_1153,N_1188);
and U1253 (N_1253,N_1181,N_1133);
nand U1254 (N_1254,N_1155,N_1177);
nor U1255 (N_1255,N_1159,N_1197);
and U1256 (N_1256,N_1166,N_1170);
nor U1257 (N_1257,N_1148,N_1140);
and U1258 (N_1258,N_1133,N_1194);
xnor U1259 (N_1259,N_1135,N_1148);
or U1260 (N_1260,N_1188,N_1194);
or U1261 (N_1261,N_1131,N_1154);
nand U1262 (N_1262,N_1177,N_1143);
xor U1263 (N_1263,N_1176,N_1169);
or U1264 (N_1264,N_1190,N_1128);
or U1265 (N_1265,N_1142,N_1139);
and U1266 (N_1266,N_1181,N_1126);
nor U1267 (N_1267,N_1187,N_1183);
nor U1268 (N_1268,N_1187,N_1160);
nor U1269 (N_1269,N_1152,N_1130);
and U1270 (N_1270,N_1193,N_1151);
or U1271 (N_1271,N_1145,N_1171);
nand U1272 (N_1272,N_1154,N_1187);
xnor U1273 (N_1273,N_1193,N_1125);
and U1274 (N_1274,N_1175,N_1142);
xnor U1275 (N_1275,N_1250,N_1265);
xor U1276 (N_1276,N_1262,N_1229);
xnor U1277 (N_1277,N_1243,N_1259);
and U1278 (N_1278,N_1249,N_1258);
nor U1279 (N_1279,N_1268,N_1242);
nor U1280 (N_1280,N_1226,N_1236);
or U1281 (N_1281,N_1273,N_1251);
or U1282 (N_1282,N_1256,N_1223);
or U1283 (N_1283,N_1238,N_1216);
nand U1284 (N_1284,N_1246,N_1206);
xor U1285 (N_1285,N_1213,N_1247);
or U1286 (N_1286,N_1266,N_1255);
or U1287 (N_1287,N_1221,N_1231);
xor U1288 (N_1288,N_1203,N_1244);
and U1289 (N_1289,N_1211,N_1234);
nand U1290 (N_1290,N_1267,N_1245);
nor U1291 (N_1291,N_1269,N_1207);
nand U1292 (N_1292,N_1228,N_1227);
or U1293 (N_1293,N_1230,N_1210);
nor U1294 (N_1294,N_1261,N_1260);
nand U1295 (N_1295,N_1209,N_1224);
and U1296 (N_1296,N_1270,N_1263);
and U1297 (N_1297,N_1212,N_1257);
nor U1298 (N_1298,N_1264,N_1205);
nand U1299 (N_1299,N_1200,N_1214);
nor U1300 (N_1300,N_1217,N_1252);
and U1301 (N_1301,N_1241,N_1237);
xnor U1302 (N_1302,N_1271,N_1232);
or U1303 (N_1303,N_1235,N_1201);
or U1304 (N_1304,N_1272,N_1208);
xor U1305 (N_1305,N_1220,N_1239);
or U1306 (N_1306,N_1204,N_1240);
or U1307 (N_1307,N_1222,N_1248);
and U1308 (N_1308,N_1254,N_1225);
or U1309 (N_1309,N_1202,N_1274);
nand U1310 (N_1310,N_1215,N_1218);
nor U1311 (N_1311,N_1253,N_1233);
and U1312 (N_1312,N_1219,N_1230);
nor U1313 (N_1313,N_1250,N_1258);
nor U1314 (N_1314,N_1264,N_1225);
nand U1315 (N_1315,N_1203,N_1242);
or U1316 (N_1316,N_1228,N_1256);
xnor U1317 (N_1317,N_1228,N_1234);
and U1318 (N_1318,N_1260,N_1223);
nor U1319 (N_1319,N_1266,N_1226);
nand U1320 (N_1320,N_1273,N_1220);
xnor U1321 (N_1321,N_1274,N_1241);
or U1322 (N_1322,N_1201,N_1216);
or U1323 (N_1323,N_1256,N_1242);
or U1324 (N_1324,N_1231,N_1268);
xnor U1325 (N_1325,N_1265,N_1262);
or U1326 (N_1326,N_1257,N_1258);
nor U1327 (N_1327,N_1236,N_1212);
and U1328 (N_1328,N_1263,N_1258);
xor U1329 (N_1329,N_1262,N_1215);
xor U1330 (N_1330,N_1251,N_1238);
or U1331 (N_1331,N_1211,N_1218);
xor U1332 (N_1332,N_1264,N_1249);
xnor U1333 (N_1333,N_1230,N_1238);
or U1334 (N_1334,N_1273,N_1264);
nand U1335 (N_1335,N_1238,N_1208);
xor U1336 (N_1336,N_1264,N_1274);
and U1337 (N_1337,N_1213,N_1212);
xor U1338 (N_1338,N_1268,N_1213);
and U1339 (N_1339,N_1238,N_1233);
nor U1340 (N_1340,N_1245,N_1228);
nor U1341 (N_1341,N_1266,N_1254);
nand U1342 (N_1342,N_1223,N_1257);
nand U1343 (N_1343,N_1225,N_1235);
and U1344 (N_1344,N_1250,N_1251);
nor U1345 (N_1345,N_1251,N_1243);
xnor U1346 (N_1346,N_1258,N_1240);
nand U1347 (N_1347,N_1203,N_1221);
xnor U1348 (N_1348,N_1236,N_1262);
or U1349 (N_1349,N_1214,N_1201);
or U1350 (N_1350,N_1285,N_1292);
xor U1351 (N_1351,N_1349,N_1344);
nand U1352 (N_1352,N_1331,N_1329);
xnor U1353 (N_1353,N_1347,N_1288);
or U1354 (N_1354,N_1281,N_1312);
and U1355 (N_1355,N_1295,N_1315);
nor U1356 (N_1356,N_1317,N_1325);
or U1357 (N_1357,N_1313,N_1326);
nand U1358 (N_1358,N_1301,N_1286);
nor U1359 (N_1359,N_1324,N_1342);
nand U1360 (N_1360,N_1335,N_1305);
xor U1361 (N_1361,N_1333,N_1336);
nor U1362 (N_1362,N_1328,N_1334);
nor U1363 (N_1363,N_1345,N_1340);
nand U1364 (N_1364,N_1307,N_1287);
nand U1365 (N_1365,N_1294,N_1296);
xor U1366 (N_1366,N_1346,N_1337);
nand U1367 (N_1367,N_1297,N_1290);
and U1368 (N_1368,N_1322,N_1323);
nand U1369 (N_1369,N_1291,N_1278);
or U1370 (N_1370,N_1303,N_1284);
or U1371 (N_1371,N_1338,N_1277);
nor U1372 (N_1372,N_1289,N_1275);
or U1373 (N_1373,N_1280,N_1343);
nand U1374 (N_1374,N_1320,N_1304);
or U1375 (N_1375,N_1299,N_1348);
xnor U1376 (N_1376,N_1283,N_1309);
or U1377 (N_1377,N_1330,N_1319);
and U1378 (N_1378,N_1306,N_1311);
nand U1379 (N_1379,N_1318,N_1279);
xnor U1380 (N_1380,N_1321,N_1276);
and U1381 (N_1381,N_1327,N_1341);
nor U1382 (N_1382,N_1339,N_1302);
nand U1383 (N_1383,N_1282,N_1293);
or U1384 (N_1384,N_1308,N_1310);
nand U1385 (N_1385,N_1298,N_1332);
and U1386 (N_1386,N_1314,N_1300);
or U1387 (N_1387,N_1316,N_1325);
or U1388 (N_1388,N_1331,N_1295);
or U1389 (N_1389,N_1305,N_1309);
and U1390 (N_1390,N_1327,N_1277);
nand U1391 (N_1391,N_1300,N_1324);
or U1392 (N_1392,N_1325,N_1338);
nor U1393 (N_1393,N_1313,N_1331);
and U1394 (N_1394,N_1289,N_1340);
and U1395 (N_1395,N_1340,N_1306);
xnor U1396 (N_1396,N_1302,N_1282);
or U1397 (N_1397,N_1341,N_1303);
nand U1398 (N_1398,N_1314,N_1315);
nor U1399 (N_1399,N_1281,N_1328);
and U1400 (N_1400,N_1316,N_1337);
nand U1401 (N_1401,N_1324,N_1345);
nor U1402 (N_1402,N_1298,N_1285);
nand U1403 (N_1403,N_1324,N_1349);
or U1404 (N_1404,N_1349,N_1335);
nand U1405 (N_1405,N_1315,N_1343);
nor U1406 (N_1406,N_1278,N_1289);
nor U1407 (N_1407,N_1316,N_1297);
and U1408 (N_1408,N_1298,N_1324);
nand U1409 (N_1409,N_1308,N_1283);
nand U1410 (N_1410,N_1317,N_1307);
and U1411 (N_1411,N_1341,N_1324);
nor U1412 (N_1412,N_1312,N_1332);
nor U1413 (N_1413,N_1280,N_1331);
and U1414 (N_1414,N_1307,N_1288);
nor U1415 (N_1415,N_1341,N_1334);
nor U1416 (N_1416,N_1295,N_1289);
and U1417 (N_1417,N_1336,N_1302);
nand U1418 (N_1418,N_1306,N_1281);
nor U1419 (N_1419,N_1295,N_1327);
nor U1420 (N_1420,N_1324,N_1276);
xor U1421 (N_1421,N_1339,N_1279);
or U1422 (N_1422,N_1327,N_1323);
nand U1423 (N_1423,N_1307,N_1344);
and U1424 (N_1424,N_1286,N_1288);
and U1425 (N_1425,N_1369,N_1411);
or U1426 (N_1426,N_1356,N_1372);
xor U1427 (N_1427,N_1379,N_1399);
nor U1428 (N_1428,N_1405,N_1381);
nand U1429 (N_1429,N_1362,N_1375);
xnor U1430 (N_1430,N_1397,N_1365);
nor U1431 (N_1431,N_1413,N_1368);
and U1432 (N_1432,N_1412,N_1387);
nand U1433 (N_1433,N_1376,N_1419);
nor U1434 (N_1434,N_1370,N_1407);
nor U1435 (N_1435,N_1390,N_1416);
nor U1436 (N_1436,N_1400,N_1359);
nand U1437 (N_1437,N_1406,N_1360);
and U1438 (N_1438,N_1377,N_1363);
and U1439 (N_1439,N_1367,N_1364);
or U1440 (N_1440,N_1366,N_1373);
and U1441 (N_1441,N_1361,N_1418);
nor U1442 (N_1442,N_1391,N_1380);
nand U1443 (N_1443,N_1395,N_1424);
or U1444 (N_1444,N_1351,N_1410);
or U1445 (N_1445,N_1396,N_1389);
or U1446 (N_1446,N_1353,N_1355);
or U1447 (N_1447,N_1393,N_1422);
nor U1448 (N_1448,N_1382,N_1352);
xor U1449 (N_1449,N_1378,N_1420);
and U1450 (N_1450,N_1408,N_1388);
nand U1451 (N_1451,N_1358,N_1386);
nor U1452 (N_1452,N_1357,N_1417);
nor U1453 (N_1453,N_1392,N_1402);
nand U1454 (N_1454,N_1374,N_1404);
xnor U1455 (N_1455,N_1409,N_1394);
nor U1456 (N_1456,N_1401,N_1398);
xnor U1457 (N_1457,N_1385,N_1414);
or U1458 (N_1458,N_1350,N_1354);
xor U1459 (N_1459,N_1403,N_1415);
or U1460 (N_1460,N_1383,N_1384);
xor U1461 (N_1461,N_1371,N_1423);
and U1462 (N_1462,N_1421,N_1399);
nand U1463 (N_1463,N_1399,N_1402);
or U1464 (N_1464,N_1389,N_1392);
nand U1465 (N_1465,N_1356,N_1362);
or U1466 (N_1466,N_1397,N_1414);
nor U1467 (N_1467,N_1371,N_1415);
or U1468 (N_1468,N_1381,N_1350);
nor U1469 (N_1469,N_1350,N_1382);
and U1470 (N_1470,N_1383,N_1393);
or U1471 (N_1471,N_1378,N_1373);
nand U1472 (N_1472,N_1364,N_1359);
nand U1473 (N_1473,N_1359,N_1355);
nor U1474 (N_1474,N_1374,N_1367);
xnor U1475 (N_1475,N_1415,N_1413);
or U1476 (N_1476,N_1358,N_1407);
nor U1477 (N_1477,N_1419,N_1374);
nor U1478 (N_1478,N_1401,N_1414);
xnor U1479 (N_1479,N_1367,N_1379);
nor U1480 (N_1480,N_1390,N_1375);
or U1481 (N_1481,N_1391,N_1359);
or U1482 (N_1482,N_1386,N_1355);
or U1483 (N_1483,N_1378,N_1357);
xnor U1484 (N_1484,N_1422,N_1370);
xnor U1485 (N_1485,N_1422,N_1411);
nand U1486 (N_1486,N_1384,N_1424);
or U1487 (N_1487,N_1358,N_1412);
and U1488 (N_1488,N_1398,N_1393);
xor U1489 (N_1489,N_1416,N_1364);
or U1490 (N_1490,N_1354,N_1423);
nand U1491 (N_1491,N_1388,N_1420);
xnor U1492 (N_1492,N_1403,N_1372);
and U1493 (N_1493,N_1399,N_1391);
nor U1494 (N_1494,N_1362,N_1388);
and U1495 (N_1495,N_1413,N_1350);
nor U1496 (N_1496,N_1378,N_1411);
nor U1497 (N_1497,N_1411,N_1396);
nand U1498 (N_1498,N_1389,N_1350);
and U1499 (N_1499,N_1373,N_1406);
nand U1500 (N_1500,N_1436,N_1481);
nand U1501 (N_1501,N_1455,N_1497);
and U1502 (N_1502,N_1470,N_1464);
nand U1503 (N_1503,N_1443,N_1458);
nor U1504 (N_1504,N_1426,N_1451);
nand U1505 (N_1505,N_1449,N_1468);
or U1506 (N_1506,N_1485,N_1486);
nor U1507 (N_1507,N_1431,N_1433);
and U1508 (N_1508,N_1496,N_1459);
xor U1509 (N_1509,N_1489,N_1452);
xnor U1510 (N_1510,N_1440,N_1479);
nand U1511 (N_1511,N_1435,N_1494);
and U1512 (N_1512,N_1471,N_1465);
or U1513 (N_1513,N_1487,N_1476);
and U1514 (N_1514,N_1457,N_1491);
nand U1515 (N_1515,N_1429,N_1444);
or U1516 (N_1516,N_1472,N_1447);
nor U1517 (N_1517,N_1441,N_1484);
or U1518 (N_1518,N_1450,N_1483);
xor U1519 (N_1519,N_1434,N_1493);
xnor U1520 (N_1520,N_1446,N_1478);
xnor U1521 (N_1521,N_1438,N_1492);
nor U1522 (N_1522,N_1454,N_1430);
nor U1523 (N_1523,N_1425,N_1428);
nand U1524 (N_1524,N_1453,N_1469);
or U1525 (N_1525,N_1467,N_1475);
nand U1526 (N_1526,N_1495,N_1461);
xnor U1527 (N_1527,N_1442,N_1448);
or U1528 (N_1528,N_1462,N_1480);
xnor U1529 (N_1529,N_1490,N_1460);
and U1530 (N_1530,N_1439,N_1499);
nand U1531 (N_1531,N_1466,N_1488);
and U1532 (N_1532,N_1474,N_1482);
or U1533 (N_1533,N_1445,N_1427);
nand U1534 (N_1534,N_1477,N_1456);
nor U1535 (N_1535,N_1432,N_1437);
xor U1536 (N_1536,N_1473,N_1498);
or U1537 (N_1537,N_1463,N_1445);
or U1538 (N_1538,N_1439,N_1444);
nand U1539 (N_1539,N_1465,N_1425);
nand U1540 (N_1540,N_1482,N_1426);
and U1541 (N_1541,N_1435,N_1471);
xnor U1542 (N_1542,N_1428,N_1469);
or U1543 (N_1543,N_1481,N_1455);
or U1544 (N_1544,N_1492,N_1496);
and U1545 (N_1545,N_1443,N_1453);
and U1546 (N_1546,N_1462,N_1450);
nor U1547 (N_1547,N_1463,N_1479);
nand U1548 (N_1548,N_1476,N_1453);
or U1549 (N_1549,N_1482,N_1446);
nand U1550 (N_1550,N_1488,N_1479);
nor U1551 (N_1551,N_1498,N_1496);
and U1552 (N_1552,N_1449,N_1475);
xnor U1553 (N_1553,N_1489,N_1480);
or U1554 (N_1554,N_1491,N_1452);
nand U1555 (N_1555,N_1498,N_1433);
or U1556 (N_1556,N_1492,N_1452);
nand U1557 (N_1557,N_1451,N_1494);
or U1558 (N_1558,N_1462,N_1441);
and U1559 (N_1559,N_1496,N_1464);
nand U1560 (N_1560,N_1469,N_1474);
and U1561 (N_1561,N_1494,N_1483);
xor U1562 (N_1562,N_1432,N_1499);
nand U1563 (N_1563,N_1482,N_1456);
nor U1564 (N_1564,N_1485,N_1491);
or U1565 (N_1565,N_1460,N_1449);
nor U1566 (N_1566,N_1470,N_1441);
nand U1567 (N_1567,N_1489,N_1498);
xnor U1568 (N_1568,N_1483,N_1439);
or U1569 (N_1569,N_1445,N_1497);
nand U1570 (N_1570,N_1427,N_1473);
nand U1571 (N_1571,N_1425,N_1483);
or U1572 (N_1572,N_1469,N_1459);
nor U1573 (N_1573,N_1447,N_1497);
or U1574 (N_1574,N_1470,N_1479);
xnor U1575 (N_1575,N_1533,N_1564);
nand U1576 (N_1576,N_1552,N_1511);
xnor U1577 (N_1577,N_1561,N_1542);
nand U1578 (N_1578,N_1507,N_1543);
xnor U1579 (N_1579,N_1562,N_1569);
xor U1580 (N_1580,N_1522,N_1534);
and U1581 (N_1581,N_1519,N_1501);
or U1582 (N_1582,N_1538,N_1549);
nor U1583 (N_1583,N_1546,N_1550);
and U1584 (N_1584,N_1528,N_1506);
or U1585 (N_1585,N_1539,N_1568);
or U1586 (N_1586,N_1535,N_1508);
nand U1587 (N_1587,N_1515,N_1572);
xor U1588 (N_1588,N_1523,N_1527);
nand U1589 (N_1589,N_1521,N_1525);
or U1590 (N_1590,N_1545,N_1532);
or U1591 (N_1591,N_1557,N_1555);
nand U1592 (N_1592,N_1553,N_1560);
nand U1593 (N_1593,N_1503,N_1529);
and U1594 (N_1594,N_1547,N_1505);
nand U1595 (N_1595,N_1556,N_1517);
and U1596 (N_1596,N_1500,N_1551);
xor U1597 (N_1597,N_1536,N_1558);
nand U1598 (N_1598,N_1537,N_1518);
or U1599 (N_1599,N_1520,N_1574);
or U1600 (N_1600,N_1541,N_1530);
and U1601 (N_1601,N_1571,N_1566);
nor U1602 (N_1602,N_1516,N_1544);
and U1603 (N_1603,N_1559,N_1524);
nor U1604 (N_1604,N_1509,N_1565);
xor U1605 (N_1605,N_1548,N_1531);
nand U1606 (N_1606,N_1502,N_1554);
nor U1607 (N_1607,N_1510,N_1513);
and U1608 (N_1608,N_1504,N_1526);
nor U1609 (N_1609,N_1563,N_1512);
or U1610 (N_1610,N_1570,N_1540);
xor U1611 (N_1611,N_1514,N_1567);
and U1612 (N_1612,N_1573,N_1537);
xor U1613 (N_1613,N_1514,N_1547);
or U1614 (N_1614,N_1573,N_1560);
nor U1615 (N_1615,N_1552,N_1564);
and U1616 (N_1616,N_1569,N_1555);
and U1617 (N_1617,N_1531,N_1558);
and U1618 (N_1618,N_1530,N_1512);
xor U1619 (N_1619,N_1521,N_1544);
nand U1620 (N_1620,N_1550,N_1525);
nor U1621 (N_1621,N_1532,N_1564);
xor U1622 (N_1622,N_1546,N_1524);
nand U1623 (N_1623,N_1522,N_1560);
xor U1624 (N_1624,N_1500,N_1509);
and U1625 (N_1625,N_1514,N_1510);
or U1626 (N_1626,N_1524,N_1529);
xor U1627 (N_1627,N_1546,N_1502);
xnor U1628 (N_1628,N_1513,N_1563);
xor U1629 (N_1629,N_1555,N_1546);
nor U1630 (N_1630,N_1570,N_1562);
or U1631 (N_1631,N_1502,N_1547);
nor U1632 (N_1632,N_1566,N_1512);
xor U1633 (N_1633,N_1554,N_1572);
xor U1634 (N_1634,N_1505,N_1529);
and U1635 (N_1635,N_1553,N_1566);
xnor U1636 (N_1636,N_1521,N_1545);
nand U1637 (N_1637,N_1538,N_1502);
nor U1638 (N_1638,N_1505,N_1568);
nor U1639 (N_1639,N_1562,N_1572);
and U1640 (N_1640,N_1516,N_1519);
xnor U1641 (N_1641,N_1506,N_1517);
or U1642 (N_1642,N_1537,N_1539);
nand U1643 (N_1643,N_1553,N_1527);
or U1644 (N_1644,N_1516,N_1548);
nand U1645 (N_1645,N_1509,N_1549);
nor U1646 (N_1646,N_1504,N_1572);
nand U1647 (N_1647,N_1562,N_1571);
xor U1648 (N_1648,N_1515,N_1516);
nor U1649 (N_1649,N_1519,N_1569);
or U1650 (N_1650,N_1613,N_1589);
and U1651 (N_1651,N_1624,N_1579);
and U1652 (N_1652,N_1646,N_1623);
nand U1653 (N_1653,N_1578,N_1593);
or U1654 (N_1654,N_1591,N_1620);
nor U1655 (N_1655,N_1631,N_1626);
xor U1656 (N_1656,N_1585,N_1607);
nor U1657 (N_1657,N_1598,N_1599);
and U1658 (N_1658,N_1602,N_1600);
xor U1659 (N_1659,N_1629,N_1605);
nand U1660 (N_1660,N_1606,N_1609);
and U1661 (N_1661,N_1581,N_1628);
and U1662 (N_1662,N_1587,N_1616);
nand U1663 (N_1663,N_1618,N_1643);
nor U1664 (N_1664,N_1635,N_1642);
nor U1665 (N_1665,N_1621,N_1638);
or U1666 (N_1666,N_1641,N_1644);
nor U1667 (N_1667,N_1576,N_1590);
and U1668 (N_1668,N_1625,N_1634);
xnor U1669 (N_1669,N_1604,N_1630);
nor U1670 (N_1670,N_1610,N_1594);
nand U1671 (N_1671,N_1582,N_1597);
nand U1672 (N_1672,N_1633,N_1612);
xor U1673 (N_1673,N_1603,N_1637);
and U1674 (N_1674,N_1577,N_1645);
or U1675 (N_1675,N_1575,N_1583);
nor U1676 (N_1676,N_1619,N_1586);
nor U1677 (N_1677,N_1580,N_1595);
nor U1678 (N_1678,N_1632,N_1611);
xnor U1679 (N_1679,N_1596,N_1588);
nand U1680 (N_1680,N_1592,N_1608);
or U1681 (N_1681,N_1615,N_1640);
and U1682 (N_1682,N_1622,N_1614);
and U1683 (N_1683,N_1649,N_1636);
and U1684 (N_1684,N_1648,N_1647);
or U1685 (N_1685,N_1584,N_1639);
xor U1686 (N_1686,N_1627,N_1601);
or U1687 (N_1687,N_1617,N_1599);
xnor U1688 (N_1688,N_1581,N_1608);
nand U1689 (N_1689,N_1636,N_1617);
nor U1690 (N_1690,N_1644,N_1623);
nor U1691 (N_1691,N_1577,N_1590);
nor U1692 (N_1692,N_1614,N_1645);
xor U1693 (N_1693,N_1611,N_1628);
and U1694 (N_1694,N_1612,N_1640);
or U1695 (N_1695,N_1602,N_1576);
nor U1696 (N_1696,N_1626,N_1596);
nor U1697 (N_1697,N_1631,N_1602);
nor U1698 (N_1698,N_1618,N_1587);
and U1699 (N_1699,N_1579,N_1634);
or U1700 (N_1700,N_1599,N_1605);
and U1701 (N_1701,N_1616,N_1632);
or U1702 (N_1702,N_1627,N_1602);
nor U1703 (N_1703,N_1626,N_1584);
nand U1704 (N_1704,N_1622,N_1591);
nor U1705 (N_1705,N_1591,N_1623);
nor U1706 (N_1706,N_1584,N_1622);
or U1707 (N_1707,N_1613,N_1602);
xnor U1708 (N_1708,N_1618,N_1617);
xnor U1709 (N_1709,N_1623,N_1602);
and U1710 (N_1710,N_1584,N_1576);
nand U1711 (N_1711,N_1625,N_1579);
and U1712 (N_1712,N_1621,N_1626);
or U1713 (N_1713,N_1590,N_1585);
nor U1714 (N_1714,N_1644,N_1592);
and U1715 (N_1715,N_1601,N_1618);
xnor U1716 (N_1716,N_1586,N_1629);
xnor U1717 (N_1717,N_1608,N_1600);
xnor U1718 (N_1718,N_1597,N_1589);
nor U1719 (N_1719,N_1605,N_1575);
nor U1720 (N_1720,N_1580,N_1623);
nand U1721 (N_1721,N_1618,N_1631);
and U1722 (N_1722,N_1622,N_1624);
nor U1723 (N_1723,N_1637,N_1619);
or U1724 (N_1724,N_1617,N_1584);
or U1725 (N_1725,N_1680,N_1676);
and U1726 (N_1726,N_1683,N_1691);
xor U1727 (N_1727,N_1708,N_1652);
xnor U1728 (N_1728,N_1677,N_1703);
nand U1729 (N_1729,N_1720,N_1696);
xor U1730 (N_1730,N_1684,N_1670);
and U1731 (N_1731,N_1660,N_1663);
nor U1732 (N_1732,N_1657,N_1679);
nor U1733 (N_1733,N_1713,N_1711);
and U1734 (N_1734,N_1685,N_1658);
nor U1735 (N_1735,N_1673,N_1689);
nand U1736 (N_1736,N_1669,N_1653);
xor U1737 (N_1737,N_1714,N_1695);
nand U1738 (N_1738,N_1724,N_1717);
or U1739 (N_1739,N_1665,N_1710);
xnor U1740 (N_1740,N_1706,N_1681);
xnor U1741 (N_1741,N_1697,N_1661);
or U1742 (N_1742,N_1721,N_1707);
nand U1743 (N_1743,N_1723,N_1664);
nor U1744 (N_1744,N_1716,N_1671);
nand U1745 (N_1745,N_1662,N_1659);
and U1746 (N_1746,N_1651,N_1678);
nand U1747 (N_1747,N_1672,N_1655);
nand U1748 (N_1748,N_1666,N_1694);
and U1749 (N_1749,N_1698,N_1699);
nor U1750 (N_1750,N_1668,N_1700);
or U1751 (N_1751,N_1718,N_1674);
nand U1752 (N_1752,N_1688,N_1715);
and U1753 (N_1753,N_1687,N_1650);
nand U1754 (N_1754,N_1693,N_1690);
and U1755 (N_1755,N_1686,N_1692);
or U1756 (N_1756,N_1705,N_1656);
and U1757 (N_1757,N_1709,N_1712);
nand U1758 (N_1758,N_1682,N_1704);
and U1759 (N_1759,N_1722,N_1675);
nand U1760 (N_1760,N_1667,N_1701);
nor U1761 (N_1761,N_1702,N_1654);
nor U1762 (N_1762,N_1719,N_1660);
nor U1763 (N_1763,N_1668,N_1678);
and U1764 (N_1764,N_1722,N_1665);
nor U1765 (N_1765,N_1657,N_1650);
nand U1766 (N_1766,N_1661,N_1713);
or U1767 (N_1767,N_1692,N_1652);
nor U1768 (N_1768,N_1684,N_1672);
and U1769 (N_1769,N_1711,N_1679);
nand U1770 (N_1770,N_1651,N_1666);
xor U1771 (N_1771,N_1685,N_1714);
or U1772 (N_1772,N_1662,N_1664);
xnor U1773 (N_1773,N_1720,N_1716);
nor U1774 (N_1774,N_1699,N_1654);
nand U1775 (N_1775,N_1723,N_1710);
nand U1776 (N_1776,N_1687,N_1671);
xnor U1777 (N_1777,N_1697,N_1683);
and U1778 (N_1778,N_1705,N_1694);
xor U1779 (N_1779,N_1700,N_1715);
nor U1780 (N_1780,N_1700,N_1697);
xnor U1781 (N_1781,N_1694,N_1652);
nand U1782 (N_1782,N_1721,N_1716);
xor U1783 (N_1783,N_1666,N_1665);
xor U1784 (N_1784,N_1654,N_1697);
and U1785 (N_1785,N_1714,N_1686);
nor U1786 (N_1786,N_1653,N_1654);
and U1787 (N_1787,N_1685,N_1686);
or U1788 (N_1788,N_1696,N_1676);
or U1789 (N_1789,N_1721,N_1652);
nand U1790 (N_1790,N_1683,N_1677);
and U1791 (N_1791,N_1656,N_1707);
nor U1792 (N_1792,N_1663,N_1693);
and U1793 (N_1793,N_1720,N_1686);
and U1794 (N_1794,N_1713,N_1691);
nor U1795 (N_1795,N_1721,N_1671);
or U1796 (N_1796,N_1704,N_1674);
or U1797 (N_1797,N_1706,N_1673);
nor U1798 (N_1798,N_1662,N_1666);
and U1799 (N_1799,N_1709,N_1693);
nand U1800 (N_1800,N_1776,N_1730);
xnor U1801 (N_1801,N_1792,N_1795);
nor U1802 (N_1802,N_1751,N_1745);
nor U1803 (N_1803,N_1747,N_1741);
nand U1804 (N_1804,N_1740,N_1727);
and U1805 (N_1805,N_1791,N_1739);
xor U1806 (N_1806,N_1726,N_1769);
and U1807 (N_1807,N_1733,N_1781);
nand U1808 (N_1808,N_1799,N_1771);
or U1809 (N_1809,N_1756,N_1763);
or U1810 (N_1810,N_1744,N_1794);
nand U1811 (N_1811,N_1759,N_1762);
and U1812 (N_1812,N_1789,N_1790);
nor U1813 (N_1813,N_1787,N_1784);
or U1814 (N_1814,N_1752,N_1788);
and U1815 (N_1815,N_1742,N_1778);
or U1816 (N_1816,N_1764,N_1725);
xor U1817 (N_1817,N_1780,N_1754);
or U1818 (N_1818,N_1774,N_1758);
and U1819 (N_1819,N_1743,N_1796);
nor U1820 (N_1820,N_1729,N_1782);
nor U1821 (N_1821,N_1765,N_1777);
nand U1822 (N_1822,N_1793,N_1779);
nand U1823 (N_1823,N_1732,N_1783);
nand U1824 (N_1824,N_1748,N_1753);
and U1825 (N_1825,N_1767,N_1761);
or U1826 (N_1826,N_1750,N_1728);
or U1827 (N_1827,N_1734,N_1735);
or U1828 (N_1828,N_1773,N_1797);
nor U1829 (N_1829,N_1770,N_1772);
nor U1830 (N_1830,N_1798,N_1786);
nor U1831 (N_1831,N_1736,N_1775);
or U1832 (N_1832,N_1746,N_1766);
nand U1833 (N_1833,N_1768,N_1785);
and U1834 (N_1834,N_1749,N_1755);
xor U1835 (N_1835,N_1731,N_1737);
or U1836 (N_1836,N_1757,N_1760);
and U1837 (N_1837,N_1738,N_1788);
or U1838 (N_1838,N_1767,N_1736);
and U1839 (N_1839,N_1771,N_1778);
and U1840 (N_1840,N_1790,N_1760);
nand U1841 (N_1841,N_1775,N_1786);
nand U1842 (N_1842,N_1790,N_1771);
and U1843 (N_1843,N_1773,N_1761);
or U1844 (N_1844,N_1733,N_1788);
and U1845 (N_1845,N_1793,N_1788);
and U1846 (N_1846,N_1749,N_1734);
and U1847 (N_1847,N_1764,N_1780);
nor U1848 (N_1848,N_1753,N_1772);
nor U1849 (N_1849,N_1772,N_1768);
and U1850 (N_1850,N_1787,N_1739);
or U1851 (N_1851,N_1746,N_1787);
xor U1852 (N_1852,N_1751,N_1775);
nand U1853 (N_1853,N_1775,N_1782);
xor U1854 (N_1854,N_1748,N_1727);
xor U1855 (N_1855,N_1783,N_1747);
or U1856 (N_1856,N_1799,N_1786);
or U1857 (N_1857,N_1741,N_1767);
or U1858 (N_1858,N_1759,N_1792);
or U1859 (N_1859,N_1739,N_1759);
nand U1860 (N_1860,N_1776,N_1748);
nor U1861 (N_1861,N_1759,N_1726);
xnor U1862 (N_1862,N_1752,N_1766);
and U1863 (N_1863,N_1743,N_1778);
xor U1864 (N_1864,N_1740,N_1787);
or U1865 (N_1865,N_1745,N_1769);
nor U1866 (N_1866,N_1745,N_1728);
xor U1867 (N_1867,N_1726,N_1755);
nand U1868 (N_1868,N_1729,N_1733);
nand U1869 (N_1869,N_1785,N_1737);
xnor U1870 (N_1870,N_1730,N_1787);
nand U1871 (N_1871,N_1765,N_1750);
nor U1872 (N_1872,N_1796,N_1779);
or U1873 (N_1873,N_1785,N_1777);
nor U1874 (N_1874,N_1732,N_1733);
or U1875 (N_1875,N_1861,N_1852);
nor U1876 (N_1876,N_1837,N_1812);
and U1877 (N_1877,N_1846,N_1826);
nand U1878 (N_1878,N_1820,N_1828);
nor U1879 (N_1879,N_1853,N_1854);
and U1880 (N_1880,N_1813,N_1844);
nand U1881 (N_1881,N_1838,N_1867);
and U1882 (N_1882,N_1830,N_1810);
nand U1883 (N_1883,N_1816,N_1834);
and U1884 (N_1884,N_1849,N_1872);
nor U1885 (N_1885,N_1802,N_1845);
nand U1886 (N_1886,N_1835,N_1855);
nand U1887 (N_1887,N_1868,N_1831);
xnor U1888 (N_1888,N_1848,N_1829);
and U1889 (N_1889,N_1808,N_1839);
and U1890 (N_1890,N_1807,N_1858);
nor U1891 (N_1891,N_1817,N_1825);
or U1892 (N_1892,N_1842,N_1869);
and U1893 (N_1893,N_1822,N_1864);
nand U1894 (N_1894,N_1823,N_1818);
and U1895 (N_1895,N_1851,N_1860);
and U1896 (N_1896,N_1832,N_1859);
nor U1897 (N_1897,N_1803,N_1806);
xor U1898 (N_1898,N_1870,N_1836);
nor U1899 (N_1899,N_1865,N_1833);
nand U1900 (N_1900,N_1850,N_1871);
nor U1901 (N_1901,N_1840,N_1847);
nand U1902 (N_1902,N_1811,N_1819);
nand U1903 (N_1903,N_1874,N_1821);
nand U1904 (N_1904,N_1809,N_1805);
nand U1905 (N_1905,N_1827,N_1801);
nand U1906 (N_1906,N_1863,N_1804);
or U1907 (N_1907,N_1824,N_1843);
nor U1908 (N_1908,N_1841,N_1800);
and U1909 (N_1909,N_1815,N_1873);
nand U1910 (N_1910,N_1856,N_1814);
or U1911 (N_1911,N_1866,N_1857);
xnor U1912 (N_1912,N_1862,N_1811);
and U1913 (N_1913,N_1851,N_1857);
nor U1914 (N_1914,N_1872,N_1838);
or U1915 (N_1915,N_1805,N_1817);
or U1916 (N_1916,N_1817,N_1843);
xnor U1917 (N_1917,N_1855,N_1828);
or U1918 (N_1918,N_1871,N_1809);
xnor U1919 (N_1919,N_1806,N_1864);
xnor U1920 (N_1920,N_1862,N_1866);
nand U1921 (N_1921,N_1861,N_1800);
xnor U1922 (N_1922,N_1820,N_1813);
nand U1923 (N_1923,N_1826,N_1809);
nor U1924 (N_1924,N_1844,N_1832);
or U1925 (N_1925,N_1814,N_1845);
xor U1926 (N_1926,N_1817,N_1854);
xor U1927 (N_1927,N_1812,N_1841);
xor U1928 (N_1928,N_1836,N_1847);
nor U1929 (N_1929,N_1843,N_1868);
xnor U1930 (N_1930,N_1825,N_1827);
and U1931 (N_1931,N_1827,N_1839);
or U1932 (N_1932,N_1813,N_1822);
or U1933 (N_1933,N_1826,N_1870);
nand U1934 (N_1934,N_1863,N_1843);
and U1935 (N_1935,N_1859,N_1866);
xor U1936 (N_1936,N_1830,N_1854);
xnor U1937 (N_1937,N_1872,N_1837);
xnor U1938 (N_1938,N_1831,N_1871);
nor U1939 (N_1939,N_1821,N_1863);
xor U1940 (N_1940,N_1820,N_1824);
nand U1941 (N_1941,N_1815,N_1866);
nand U1942 (N_1942,N_1873,N_1821);
and U1943 (N_1943,N_1871,N_1868);
and U1944 (N_1944,N_1802,N_1815);
nor U1945 (N_1945,N_1840,N_1819);
and U1946 (N_1946,N_1871,N_1865);
or U1947 (N_1947,N_1869,N_1866);
xnor U1948 (N_1948,N_1849,N_1812);
or U1949 (N_1949,N_1852,N_1847);
xor U1950 (N_1950,N_1913,N_1903);
and U1951 (N_1951,N_1882,N_1908);
nor U1952 (N_1952,N_1883,N_1923);
xnor U1953 (N_1953,N_1932,N_1930);
and U1954 (N_1954,N_1916,N_1898);
nand U1955 (N_1955,N_1921,N_1943);
and U1956 (N_1956,N_1905,N_1899);
nand U1957 (N_1957,N_1926,N_1875);
and U1958 (N_1958,N_1909,N_1942);
nor U1959 (N_1959,N_1933,N_1922);
xor U1960 (N_1960,N_1887,N_1890);
or U1961 (N_1961,N_1907,N_1888);
or U1962 (N_1962,N_1928,N_1936);
nor U1963 (N_1963,N_1878,N_1893);
nand U1964 (N_1964,N_1881,N_1876);
or U1965 (N_1965,N_1929,N_1897);
and U1966 (N_1966,N_1925,N_1891);
nor U1967 (N_1967,N_1938,N_1892);
or U1968 (N_1968,N_1895,N_1917);
or U1969 (N_1969,N_1920,N_1889);
or U1970 (N_1970,N_1877,N_1906);
nor U1971 (N_1971,N_1941,N_1915);
or U1972 (N_1972,N_1885,N_1948);
nor U1973 (N_1973,N_1896,N_1886);
and U1974 (N_1974,N_1894,N_1919);
nor U1975 (N_1975,N_1901,N_1912);
xnor U1976 (N_1976,N_1946,N_1934);
nand U1977 (N_1977,N_1914,N_1935);
xnor U1978 (N_1978,N_1939,N_1902);
xor U1979 (N_1979,N_1911,N_1949);
nor U1980 (N_1980,N_1918,N_1910);
xnor U1981 (N_1981,N_1884,N_1944);
nand U1982 (N_1982,N_1931,N_1940);
xor U1983 (N_1983,N_1947,N_1879);
or U1984 (N_1984,N_1900,N_1937);
nand U1985 (N_1985,N_1904,N_1927);
xor U1986 (N_1986,N_1880,N_1945);
and U1987 (N_1987,N_1924,N_1929);
or U1988 (N_1988,N_1922,N_1876);
and U1989 (N_1989,N_1904,N_1930);
xor U1990 (N_1990,N_1879,N_1883);
xnor U1991 (N_1991,N_1928,N_1878);
and U1992 (N_1992,N_1927,N_1895);
and U1993 (N_1993,N_1906,N_1928);
xnor U1994 (N_1994,N_1938,N_1914);
and U1995 (N_1995,N_1913,N_1926);
nor U1996 (N_1996,N_1910,N_1879);
nand U1997 (N_1997,N_1922,N_1881);
nand U1998 (N_1998,N_1936,N_1929);
and U1999 (N_1999,N_1880,N_1883);
xor U2000 (N_2000,N_1884,N_1901);
nand U2001 (N_2001,N_1898,N_1946);
or U2002 (N_2002,N_1926,N_1902);
and U2003 (N_2003,N_1910,N_1901);
nand U2004 (N_2004,N_1904,N_1910);
or U2005 (N_2005,N_1878,N_1916);
or U2006 (N_2006,N_1883,N_1906);
nand U2007 (N_2007,N_1895,N_1905);
or U2008 (N_2008,N_1889,N_1948);
or U2009 (N_2009,N_1933,N_1903);
and U2010 (N_2010,N_1945,N_1930);
nor U2011 (N_2011,N_1919,N_1913);
nand U2012 (N_2012,N_1888,N_1894);
or U2013 (N_2013,N_1934,N_1878);
and U2014 (N_2014,N_1912,N_1942);
nor U2015 (N_2015,N_1897,N_1917);
nor U2016 (N_2016,N_1875,N_1919);
nor U2017 (N_2017,N_1890,N_1885);
nor U2018 (N_2018,N_1918,N_1892);
or U2019 (N_2019,N_1940,N_1887);
xor U2020 (N_2020,N_1906,N_1909);
or U2021 (N_2021,N_1925,N_1928);
nand U2022 (N_2022,N_1897,N_1945);
nand U2023 (N_2023,N_1885,N_1888);
nor U2024 (N_2024,N_1921,N_1887);
or U2025 (N_2025,N_1994,N_2017);
nand U2026 (N_2026,N_1978,N_1992);
nor U2027 (N_2027,N_2002,N_1993);
or U2028 (N_2028,N_1966,N_2007);
and U2029 (N_2029,N_1961,N_1985);
or U2030 (N_2030,N_1998,N_1964);
nor U2031 (N_2031,N_1958,N_2019);
xnor U2032 (N_2032,N_1975,N_2003);
nand U2033 (N_2033,N_1988,N_1957);
and U2034 (N_2034,N_2018,N_1974);
nand U2035 (N_2035,N_1963,N_2010);
nor U2036 (N_2036,N_2015,N_1971);
and U2037 (N_2037,N_2014,N_1987);
and U2038 (N_2038,N_1997,N_1996);
nor U2039 (N_2039,N_1983,N_1977);
and U2040 (N_2040,N_2020,N_2009);
or U2041 (N_2041,N_2005,N_2013);
nand U2042 (N_2042,N_1999,N_1965);
xnor U2043 (N_2043,N_2000,N_2016);
xnor U2044 (N_2044,N_1959,N_1953);
or U2045 (N_2045,N_1991,N_1956);
or U2046 (N_2046,N_1982,N_1976);
and U2047 (N_2047,N_2008,N_1955);
nor U2048 (N_2048,N_1984,N_2022);
or U2049 (N_2049,N_2012,N_2001);
or U2050 (N_2050,N_1962,N_1981);
or U2051 (N_2051,N_2023,N_1972);
and U2052 (N_2052,N_1951,N_1995);
and U2053 (N_2053,N_2011,N_1980);
nor U2054 (N_2054,N_2004,N_1950);
and U2055 (N_2055,N_1986,N_1989);
nand U2056 (N_2056,N_1969,N_2024);
or U2057 (N_2057,N_1952,N_2006);
nor U2058 (N_2058,N_1970,N_1954);
or U2059 (N_2059,N_1990,N_2021);
nor U2060 (N_2060,N_1973,N_1960);
xor U2061 (N_2061,N_1967,N_1979);
nand U2062 (N_2062,N_1968,N_2001);
and U2063 (N_2063,N_2016,N_1987);
or U2064 (N_2064,N_1980,N_2022);
nand U2065 (N_2065,N_2005,N_1977);
nor U2066 (N_2066,N_2004,N_1964);
nor U2067 (N_2067,N_2015,N_1978);
or U2068 (N_2068,N_1965,N_2000);
nor U2069 (N_2069,N_1993,N_2014);
and U2070 (N_2070,N_1981,N_1989);
nand U2071 (N_2071,N_1956,N_1966);
and U2072 (N_2072,N_1968,N_1975);
and U2073 (N_2073,N_1986,N_2013);
xnor U2074 (N_2074,N_1960,N_1963);
nor U2075 (N_2075,N_1994,N_1989);
xnor U2076 (N_2076,N_1990,N_2011);
and U2077 (N_2077,N_1973,N_2016);
and U2078 (N_2078,N_1972,N_1991);
or U2079 (N_2079,N_2022,N_1954);
nand U2080 (N_2080,N_2006,N_1986);
or U2081 (N_2081,N_1976,N_2007);
nor U2082 (N_2082,N_1958,N_1992);
xor U2083 (N_2083,N_1985,N_1980);
nand U2084 (N_2084,N_2022,N_1951);
xnor U2085 (N_2085,N_1990,N_1962);
and U2086 (N_2086,N_1991,N_1979);
or U2087 (N_2087,N_1957,N_1953);
nor U2088 (N_2088,N_2017,N_1978);
and U2089 (N_2089,N_1955,N_1990);
and U2090 (N_2090,N_2010,N_1967);
nor U2091 (N_2091,N_1983,N_1976);
xor U2092 (N_2092,N_1975,N_1974);
and U2093 (N_2093,N_2011,N_1995);
nor U2094 (N_2094,N_1986,N_2010);
xnor U2095 (N_2095,N_1964,N_1971);
nor U2096 (N_2096,N_1973,N_1953);
or U2097 (N_2097,N_2016,N_1957);
nand U2098 (N_2098,N_1976,N_2010);
or U2099 (N_2099,N_1974,N_1969);
nor U2100 (N_2100,N_2055,N_2095);
nand U2101 (N_2101,N_2059,N_2044);
or U2102 (N_2102,N_2079,N_2060);
or U2103 (N_2103,N_2091,N_2031);
xnor U2104 (N_2104,N_2083,N_2038);
nor U2105 (N_2105,N_2094,N_2043);
nand U2106 (N_2106,N_2075,N_2026);
and U2107 (N_2107,N_2051,N_2065);
nand U2108 (N_2108,N_2097,N_2081);
xnor U2109 (N_2109,N_2086,N_2082);
xor U2110 (N_2110,N_2099,N_2061);
nand U2111 (N_2111,N_2037,N_2069);
and U2112 (N_2112,N_2071,N_2089);
or U2113 (N_2113,N_2025,N_2087);
xor U2114 (N_2114,N_2035,N_2053);
xor U2115 (N_2115,N_2050,N_2080);
and U2116 (N_2116,N_2056,N_2058);
nand U2117 (N_2117,N_2027,N_2064);
nand U2118 (N_2118,N_2032,N_2029);
or U2119 (N_2119,N_2047,N_2049);
xor U2120 (N_2120,N_2054,N_2090);
nor U2121 (N_2121,N_2093,N_2052);
nand U2122 (N_2122,N_2077,N_2040);
nand U2123 (N_2123,N_2042,N_2068);
xnor U2124 (N_2124,N_2062,N_2098);
nor U2125 (N_2125,N_2092,N_2030);
xnor U2126 (N_2126,N_2084,N_2045);
xor U2127 (N_2127,N_2096,N_2085);
or U2128 (N_2128,N_2046,N_2041);
and U2129 (N_2129,N_2073,N_2070);
nor U2130 (N_2130,N_2028,N_2033);
nand U2131 (N_2131,N_2034,N_2063);
nor U2132 (N_2132,N_2072,N_2066);
xor U2133 (N_2133,N_2088,N_2057);
xnor U2134 (N_2134,N_2067,N_2078);
nor U2135 (N_2135,N_2074,N_2076);
nand U2136 (N_2136,N_2036,N_2039);
nand U2137 (N_2137,N_2048,N_2096);
and U2138 (N_2138,N_2039,N_2044);
or U2139 (N_2139,N_2035,N_2070);
or U2140 (N_2140,N_2070,N_2049);
nor U2141 (N_2141,N_2063,N_2071);
nand U2142 (N_2142,N_2078,N_2056);
or U2143 (N_2143,N_2093,N_2067);
and U2144 (N_2144,N_2035,N_2066);
nor U2145 (N_2145,N_2025,N_2094);
xnor U2146 (N_2146,N_2038,N_2078);
nand U2147 (N_2147,N_2092,N_2063);
xor U2148 (N_2148,N_2076,N_2073);
nand U2149 (N_2149,N_2041,N_2028);
and U2150 (N_2150,N_2087,N_2046);
nand U2151 (N_2151,N_2055,N_2039);
xor U2152 (N_2152,N_2088,N_2046);
or U2153 (N_2153,N_2096,N_2029);
nor U2154 (N_2154,N_2027,N_2033);
or U2155 (N_2155,N_2030,N_2097);
nand U2156 (N_2156,N_2046,N_2032);
xnor U2157 (N_2157,N_2087,N_2080);
nor U2158 (N_2158,N_2069,N_2059);
nand U2159 (N_2159,N_2072,N_2058);
nor U2160 (N_2160,N_2044,N_2050);
and U2161 (N_2161,N_2037,N_2081);
nor U2162 (N_2162,N_2057,N_2045);
or U2163 (N_2163,N_2035,N_2098);
nor U2164 (N_2164,N_2060,N_2096);
nand U2165 (N_2165,N_2069,N_2094);
xnor U2166 (N_2166,N_2072,N_2095);
nor U2167 (N_2167,N_2097,N_2059);
nor U2168 (N_2168,N_2080,N_2037);
nand U2169 (N_2169,N_2089,N_2076);
nand U2170 (N_2170,N_2091,N_2082);
nand U2171 (N_2171,N_2039,N_2066);
nor U2172 (N_2172,N_2098,N_2041);
or U2173 (N_2173,N_2045,N_2074);
nand U2174 (N_2174,N_2035,N_2031);
nor U2175 (N_2175,N_2133,N_2115);
nand U2176 (N_2176,N_2111,N_2174);
nand U2177 (N_2177,N_2150,N_2131);
nand U2178 (N_2178,N_2124,N_2167);
or U2179 (N_2179,N_2162,N_2142);
xor U2180 (N_2180,N_2101,N_2117);
nor U2181 (N_2181,N_2168,N_2104);
nand U2182 (N_2182,N_2173,N_2156);
and U2183 (N_2183,N_2108,N_2149);
xor U2184 (N_2184,N_2135,N_2103);
xor U2185 (N_2185,N_2118,N_2107);
nand U2186 (N_2186,N_2132,N_2136);
nand U2187 (N_2187,N_2161,N_2163);
nand U2188 (N_2188,N_2139,N_2155);
or U2189 (N_2189,N_2147,N_2110);
or U2190 (N_2190,N_2127,N_2170);
or U2191 (N_2191,N_2144,N_2113);
or U2192 (N_2192,N_2128,N_2130);
and U2193 (N_2193,N_2112,N_2125);
xor U2194 (N_2194,N_2169,N_2116);
xnor U2195 (N_2195,N_2114,N_2151);
xnor U2196 (N_2196,N_2123,N_2122);
and U2197 (N_2197,N_2157,N_2126);
or U2198 (N_2198,N_2129,N_2120);
and U2199 (N_2199,N_2153,N_2164);
or U2200 (N_2200,N_2145,N_2137);
and U2201 (N_2201,N_2105,N_2143);
xor U2202 (N_2202,N_2106,N_2102);
or U2203 (N_2203,N_2152,N_2141);
xor U2204 (N_2204,N_2158,N_2159);
nand U2205 (N_2205,N_2121,N_2154);
and U2206 (N_2206,N_2172,N_2109);
nand U2207 (N_2207,N_2100,N_2138);
xor U2208 (N_2208,N_2140,N_2119);
nand U2209 (N_2209,N_2146,N_2160);
and U2210 (N_2210,N_2165,N_2134);
or U2211 (N_2211,N_2171,N_2166);
nand U2212 (N_2212,N_2148,N_2166);
nand U2213 (N_2213,N_2104,N_2155);
xnor U2214 (N_2214,N_2174,N_2100);
or U2215 (N_2215,N_2110,N_2153);
and U2216 (N_2216,N_2122,N_2117);
nor U2217 (N_2217,N_2132,N_2106);
and U2218 (N_2218,N_2164,N_2103);
or U2219 (N_2219,N_2103,N_2159);
nand U2220 (N_2220,N_2169,N_2120);
nand U2221 (N_2221,N_2164,N_2147);
nand U2222 (N_2222,N_2163,N_2146);
or U2223 (N_2223,N_2101,N_2135);
nor U2224 (N_2224,N_2105,N_2150);
or U2225 (N_2225,N_2162,N_2146);
and U2226 (N_2226,N_2160,N_2117);
and U2227 (N_2227,N_2168,N_2101);
or U2228 (N_2228,N_2154,N_2149);
nor U2229 (N_2229,N_2154,N_2138);
nor U2230 (N_2230,N_2141,N_2120);
and U2231 (N_2231,N_2169,N_2122);
or U2232 (N_2232,N_2172,N_2106);
xnor U2233 (N_2233,N_2153,N_2138);
xnor U2234 (N_2234,N_2164,N_2165);
nor U2235 (N_2235,N_2125,N_2161);
or U2236 (N_2236,N_2116,N_2105);
and U2237 (N_2237,N_2112,N_2124);
xor U2238 (N_2238,N_2145,N_2148);
xnor U2239 (N_2239,N_2128,N_2134);
nor U2240 (N_2240,N_2104,N_2109);
or U2241 (N_2241,N_2164,N_2126);
xor U2242 (N_2242,N_2150,N_2108);
and U2243 (N_2243,N_2102,N_2153);
and U2244 (N_2244,N_2119,N_2100);
nand U2245 (N_2245,N_2108,N_2113);
xor U2246 (N_2246,N_2149,N_2123);
and U2247 (N_2247,N_2162,N_2104);
nor U2248 (N_2248,N_2166,N_2130);
and U2249 (N_2249,N_2159,N_2140);
or U2250 (N_2250,N_2222,N_2248);
or U2251 (N_2251,N_2193,N_2181);
or U2252 (N_2252,N_2217,N_2245);
xor U2253 (N_2253,N_2237,N_2176);
nor U2254 (N_2254,N_2229,N_2236);
and U2255 (N_2255,N_2224,N_2219);
xor U2256 (N_2256,N_2208,N_2226);
nand U2257 (N_2257,N_2246,N_2207);
nor U2258 (N_2258,N_2189,N_2177);
or U2259 (N_2259,N_2243,N_2195);
or U2260 (N_2260,N_2202,N_2188);
nor U2261 (N_2261,N_2194,N_2203);
nor U2262 (N_2262,N_2227,N_2244);
xor U2263 (N_2263,N_2249,N_2213);
nor U2264 (N_2264,N_2186,N_2215);
xnor U2265 (N_2265,N_2192,N_2206);
nor U2266 (N_2266,N_2239,N_2221);
xor U2267 (N_2267,N_2198,N_2182);
and U2268 (N_2268,N_2223,N_2214);
nand U2269 (N_2269,N_2191,N_2190);
nand U2270 (N_2270,N_2187,N_2210);
nand U2271 (N_2271,N_2238,N_2209);
xnor U2272 (N_2272,N_2241,N_2184);
xnor U2273 (N_2273,N_2218,N_2183);
xor U2274 (N_2274,N_2228,N_2235);
or U2275 (N_2275,N_2199,N_2230);
and U2276 (N_2276,N_2175,N_2178);
nor U2277 (N_2277,N_2197,N_2247);
nand U2278 (N_2278,N_2196,N_2185);
xnor U2279 (N_2279,N_2242,N_2211);
or U2280 (N_2280,N_2179,N_2232);
xnor U2281 (N_2281,N_2233,N_2205);
nand U2282 (N_2282,N_2225,N_2216);
and U2283 (N_2283,N_2204,N_2212);
or U2284 (N_2284,N_2200,N_2220);
and U2285 (N_2285,N_2180,N_2240);
xor U2286 (N_2286,N_2201,N_2234);
xor U2287 (N_2287,N_2231,N_2237);
xor U2288 (N_2288,N_2182,N_2188);
and U2289 (N_2289,N_2244,N_2201);
or U2290 (N_2290,N_2202,N_2224);
nor U2291 (N_2291,N_2202,N_2228);
xor U2292 (N_2292,N_2187,N_2240);
nor U2293 (N_2293,N_2225,N_2182);
nand U2294 (N_2294,N_2246,N_2229);
nand U2295 (N_2295,N_2225,N_2230);
and U2296 (N_2296,N_2246,N_2212);
or U2297 (N_2297,N_2208,N_2183);
or U2298 (N_2298,N_2234,N_2245);
nor U2299 (N_2299,N_2244,N_2223);
nand U2300 (N_2300,N_2200,N_2176);
nand U2301 (N_2301,N_2177,N_2194);
or U2302 (N_2302,N_2233,N_2211);
nand U2303 (N_2303,N_2229,N_2234);
xor U2304 (N_2304,N_2212,N_2210);
and U2305 (N_2305,N_2240,N_2194);
or U2306 (N_2306,N_2228,N_2222);
xnor U2307 (N_2307,N_2215,N_2243);
or U2308 (N_2308,N_2224,N_2205);
nand U2309 (N_2309,N_2175,N_2242);
nor U2310 (N_2310,N_2201,N_2233);
or U2311 (N_2311,N_2204,N_2238);
nor U2312 (N_2312,N_2234,N_2230);
nor U2313 (N_2313,N_2188,N_2245);
nor U2314 (N_2314,N_2243,N_2221);
nor U2315 (N_2315,N_2225,N_2211);
or U2316 (N_2316,N_2191,N_2244);
xnor U2317 (N_2317,N_2180,N_2229);
or U2318 (N_2318,N_2225,N_2195);
xor U2319 (N_2319,N_2248,N_2220);
or U2320 (N_2320,N_2236,N_2211);
xnor U2321 (N_2321,N_2221,N_2210);
xor U2322 (N_2322,N_2228,N_2198);
nor U2323 (N_2323,N_2181,N_2209);
or U2324 (N_2324,N_2181,N_2189);
and U2325 (N_2325,N_2308,N_2312);
or U2326 (N_2326,N_2307,N_2294);
xnor U2327 (N_2327,N_2268,N_2281);
and U2328 (N_2328,N_2301,N_2318);
or U2329 (N_2329,N_2315,N_2314);
nand U2330 (N_2330,N_2291,N_2271);
nand U2331 (N_2331,N_2293,N_2269);
or U2332 (N_2332,N_2288,N_2297);
and U2333 (N_2333,N_2262,N_2310);
and U2334 (N_2334,N_2251,N_2272);
xnor U2335 (N_2335,N_2259,N_2287);
xor U2336 (N_2336,N_2267,N_2265);
and U2337 (N_2337,N_2277,N_2266);
and U2338 (N_2338,N_2260,N_2316);
nand U2339 (N_2339,N_2257,N_2311);
and U2340 (N_2340,N_2286,N_2252);
xor U2341 (N_2341,N_2261,N_2306);
and U2342 (N_2342,N_2292,N_2263);
nand U2343 (N_2343,N_2298,N_2282);
nand U2344 (N_2344,N_2320,N_2300);
and U2345 (N_2345,N_2273,N_2253);
or U2346 (N_2346,N_2296,N_2322);
and U2347 (N_2347,N_2295,N_2285);
nand U2348 (N_2348,N_2290,N_2264);
nor U2349 (N_2349,N_2302,N_2305);
and U2350 (N_2350,N_2303,N_2317);
xnor U2351 (N_2351,N_2256,N_2309);
and U2352 (N_2352,N_2323,N_2283);
xnor U2353 (N_2353,N_2275,N_2319);
nor U2354 (N_2354,N_2284,N_2274);
nor U2355 (N_2355,N_2258,N_2280);
and U2356 (N_2356,N_2324,N_2270);
and U2357 (N_2357,N_2279,N_2276);
and U2358 (N_2358,N_2313,N_2304);
xnor U2359 (N_2359,N_2289,N_2321);
nand U2360 (N_2360,N_2255,N_2250);
or U2361 (N_2361,N_2278,N_2254);
xor U2362 (N_2362,N_2299,N_2256);
xnor U2363 (N_2363,N_2272,N_2265);
nor U2364 (N_2364,N_2303,N_2292);
nand U2365 (N_2365,N_2251,N_2316);
or U2366 (N_2366,N_2288,N_2314);
or U2367 (N_2367,N_2299,N_2260);
or U2368 (N_2368,N_2261,N_2316);
xor U2369 (N_2369,N_2252,N_2323);
xnor U2370 (N_2370,N_2258,N_2309);
or U2371 (N_2371,N_2274,N_2320);
nand U2372 (N_2372,N_2316,N_2324);
or U2373 (N_2373,N_2324,N_2250);
or U2374 (N_2374,N_2322,N_2298);
and U2375 (N_2375,N_2259,N_2297);
nand U2376 (N_2376,N_2307,N_2277);
nor U2377 (N_2377,N_2286,N_2298);
or U2378 (N_2378,N_2290,N_2254);
and U2379 (N_2379,N_2284,N_2254);
nand U2380 (N_2380,N_2290,N_2295);
and U2381 (N_2381,N_2262,N_2298);
nor U2382 (N_2382,N_2287,N_2256);
nor U2383 (N_2383,N_2274,N_2280);
or U2384 (N_2384,N_2289,N_2279);
or U2385 (N_2385,N_2277,N_2282);
xnor U2386 (N_2386,N_2281,N_2271);
nor U2387 (N_2387,N_2309,N_2269);
xor U2388 (N_2388,N_2267,N_2258);
xnor U2389 (N_2389,N_2275,N_2309);
or U2390 (N_2390,N_2260,N_2269);
and U2391 (N_2391,N_2278,N_2294);
and U2392 (N_2392,N_2296,N_2295);
nand U2393 (N_2393,N_2307,N_2321);
nand U2394 (N_2394,N_2296,N_2272);
nor U2395 (N_2395,N_2324,N_2313);
nor U2396 (N_2396,N_2277,N_2267);
xnor U2397 (N_2397,N_2307,N_2268);
nor U2398 (N_2398,N_2253,N_2286);
nor U2399 (N_2399,N_2312,N_2273);
and U2400 (N_2400,N_2394,N_2363);
nand U2401 (N_2401,N_2355,N_2373);
nand U2402 (N_2402,N_2334,N_2353);
or U2403 (N_2403,N_2379,N_2382);
or U2404 (N_2404,N_2350,N_2389);
nand U2405 (N_2405,N_2352,N_2390);
xor U2406 (N_2406,N_2366,N_2325);
xor U2407 (N_2407,N_2349,N_2335);
or U2408 (N_2408,N_2368,N_2344);
nor U2409 (N_2409,N_2330,N_2356);
and U2410 (N_2410,N_2340,N_2346);
nand U2411 (N_2411,N_2370,N_2371);
or U2412 (N_2412,N_2327,N_2354);
xor U2413 (N_2413,N_2369,N_2345);
nand U2414 (N_2414,N_2362,N_2385);
or U2415 (N_2415,N_2328,N_2386);
nand U2416 (N_2416,N_2343,N_2377);
xor U2417 (N_2417,N_2342,N_2367);
nor U2418 (N_2418,N_2375,N_2359);
or U2419 (N_2419,N_2333,N_2358);
or U2420 (N_2420,N_2388,N_2380);
or U2421 (N_2421,N_2384,N_2374);
nand U2422 (N_2422,N_2360,N_2331);
or U2423 (N_2423,N_2398,N_2393);
xnor U2424 (N_2424,N_2341,N_2391);
or U2425 (N_2425,N_2351,N_2365);
nand U2426 (N_2426,N_2392,N_2336);
nand U2427 (N_2427,N_2397,N_2381);
nand U2428 (N_2428,N_2396,N_2361);
xnor U2429 (N_2429,N_2348,N_2395);
xor U2430 (N_2430,N_2372,N_2339);
nand U2431 (N_2431,N_2338,N_2383);
or U2432 (N_2432,N_2364,N_2399);
and U2433 (N_2433,N_2332,N_2326);
nor U2434 (N_2434,N_2387,N_2337);
xnor U2435 (N_2435,N_2378,N_2357);
or U2436 (N_2436,N_2376,N_2347);
nand U2437 (N_2437,N_2329,N_2353);
and U2438 (N_2438,N_2349,N_2387);
or U2439 (N_2439,N_2328,N_2385);
xnor U2440 (N_2440,N_2351,N_2363);
or U2441 (N_2441,N_2394,N_2381);
or U2442 (N_2442,N_2363,N_2362);
or U2443 (N_2443,N_2361,N_2328);
or U2444 (N_2444,N_2359,N_2329);
xor U2445 (N_2445,N_2344,N_2365);
nor U2446 (N_2446,N_2326,N_2337);
xor U2447 (N_2447,N_2371,N_2335);
nor U2448 (N_2448,N_2349,N_2398);
or U2449 (N_2449,N_2341,N_2344);
xnor U2450 (N_2450,N_2368,N_2325);
nand U2451 (N_2451,N_2399,N_2379);
and U2452 (N_2452,N_2377,N_2344);
nand U2453 (N_2453,N_2380,N_2327);
nand U2454 (N_2454,N_2372,N_2396);
or U2455 (N_2455,N_2348,N_2376);
nand U2456 (N_2456,N_2388,N_2391);
nor U2457 (N_2457,N_2363,N_2387);
nor U2458 (N_2458,N_2336,N_2334);
or U2459 (N_2459,N_2393,N_2372);
nor U2460 (N_2460,N_2386,N_2364);
nand U2461 (N_2461,N_2341,N_2377);
or U2462 (N_2462,N_2363,N_2344);
nand U2463 (N_2463,N_2396,N_2335);
nand U2464 (N_2464,N_2383,N_2362);
or U2465 (N_2465,N_2335,N_2382);
and U2466 (N_2466,N_2326,N_2335);
nand U2467 (N_2467,N_2325,N_2364);
nor U2468 (N_2468,N_2380,N_2383);
and U2469 (N_2469,N_2342,N_2372);
or U2470 (N_2470,N_2363,N_2368);
xnor U2471 (N_2471,N_2376,N_2364);
nand U2472 (N_2472,N_2360,N_2398);
and U2473 (N_2473,N_2397,N_2334);
nor U2474 (N_2474,N_2351,N_2358);
or U2475 (N_2475,N_2429,N_2404);
xor U2476 (N_2476,N_2473,N_2432);
xor U2477 (N_2477,N_2422,N_2417);
nor U2478 (N_2478,N_2425,N_2400);
xnor U2479 (N_2479,N_2462,N_2430);
nor U2480 (N_2480,N_2407,N_2414);
and U2481 (N_2481,N_2446,N_2413);
nand U2482 (N_2482,N_2439,N_2444);
or U2483 (N_2483,N_2455,N_2441);
and U2484 (N_2484,N_2424,N_2415);
xnor U2485 (N_2485,N_2402,N_2451);
nor U2486 (N_2486,N_2436,N_2411);
nor U2487 (N_2487,N_2466,N_2464);
or U2488 (N_2488,N_2427,N_2405);
xor U2489 (N_2489,N_2438,N_2472);
nand U2490 (N_2490,N_2468,N_2449);
nor U2491 (N_2491,N_2416,N_2408);
or U2492 (N_2492,N_2409,N_2456);
and U2493 (N_2493,N_2467,N_2461);
and U2494 (N_2494,N_2420,N_2471);
or U2495 (N_2495,N_2447,N_2460);
and U2496 (N_2496,N_2443,N_2458);
or U2497 (N_2497,N_2465,N_2428);
nand U2498 (N_2498,N_2437,N_2470);
and U2499 (N_2499,N_2445,N_2431);
or U2500 (N_2500,N_2433,N_2453);
and U2501 (N_2501,N_2442,N_2440);
nor U2502 (N_2502,N_2459,N_2474);
nand U2503 (N_2503,N_2469,N_2454);
nor U2504 (N_2504,N_2418,N_2457);
nor U2505 (N_2505,N_2403,N_2410);
and U2506 (N_2506,N_2426,N_2421);
nand U2507 (N_2507,N_2423,N_2401);
nand U2508 (N_2508,N_2463,N_2406);
xnor U2509 (N_2509,N_2450,N_2448);
and U2510 (N_2510,N_2452,N_2419);
xor U2511 (N_2511,N_2412,N_2434);
or U2512 (N_2512,N_2435,N_2454);
nand U2513 (N_2513,N_2451,N_2439);
or U2514 (N_2514,N_2466,N_2468);
nor U2515 (N_2515,N_2443,N_2427);
nor U2516 (N_2516,N_2406,N_2429);
or U2517 (N_2517,N_2430,N_2421);
nor U2518 (N_2518,N_2471,N_2452);
nor U2519 (N_2519,N_2462,N_2423);
or U2520 (N_2520,N_2462,N_2439);
nand U2521 (N_2521,N_2427,N_2407);
or U2522 (N_2522,N_2411,N_2441);
nor U2523 (N_2523,N_2470,N_2442);
nor U2524 (N_2524,N_2406,N_2408);
xnor U2525 (N_2525,N_2400,N_2428);
and U2526 (N_2526,N_2474,N_2426);
xnor U2527 (N_2527,N_2409,N_2410);
or U2528 (N_2528,N_2434,N_2440);
and U2529 (N_2529,N_2403,N_2444);
nor U2530 (N_2530,N_2432,N_2434);
xor U2531 (N_2531,N_2450,N_2436);
and U2532 (N_2532,N_2462,N_2405);
and U2533 (N_2533,N_2423,N_2421);
nor U2534 (N_2534,N_2401,N_2453);
nand U2535 (N_2535,N_2419,N_2428);
or U2536 (N_2536,N_2472,N_2444);
xnor U2537 (N_2537,N_2463,N_2465);
nand U2538 (N_2538,N_2420,N_2430);
nor U2539 (N_2539,N_2430,N_2400);
nand U2540 (N_2540,N_2431,N_2466);
nand U2541 (N_2541,N_2425,N_2472);
nor U2542 (N_2542,N_2474,N_2414);
and U2543 (N_2543,N_2411,N_2446);
or U2544 (N_2544,N_2453,N_2404);
nor U2545 (N_2545,N_2430,N_2419);
nor U2546 (N_2546,N_2450,N_2401);
xnor U2547 (N_2547,N_2465,N_2409);
nor U2548 (N_2548,N_2400,N_2421);
nand U2549 (N_2549,N_2425,N_2474);
nor U2550 (N_2550,N_2488,N_2484);
and U2551 (N_2551,N_2538,N_2503);
or U2552 (N_2552,N_2476,N_2481);
and U2553 (N_2553,N_2502,N_2519);
or U2554 (N_2554,N_2524,N_2515);
xnor U2555 (N_2555,N_2526,N_2517);
or U2556 (N_2556,N_2505,N_2525);
xnor U2557 (N_2557,N_2487,N_2506);
xor U2558 (N_2558,N_2522,N_2510);
xnor U2559 (N_2559,N_2508,N_2477);
and U2560 (N_2560,N_2485,N_2521);
and U2561 (N_2561,N_2478,N_2483);
or U2562 (N_2562,N_2534,N_2529);
xor U2563 (N_2563,N_2504,N_2539);
or U2564 (N_2564,N_2509,N_2547);
or U2565 (N_2565,N_2512,N_2501);
nor U2566 (N_2566,N_2498,N_2516);
or U2567 (N_2567,N_2494,N_2532);
or U2568 (N_2568,N_2549,N_2493);
nor U2569 (N_2569,N_2544,N_2537);
nor U2570 (N_2570,N_2535,N_2491);
and U2571 (N_2571,N_2541,N_2490);
or U2572 (N_2572,N_2523,N_2482);
or U2573 (N_2573,N_2530,N_2531);
or U2574 (N_2574,N_2527,N_2486);
xor U2575 (N_2575,N_2496,N_2514);
xnor U2576 (N_2576,N_2543,N_2495);
or U2577 (N_2577,N_2497,N_2479);
or U2578 (N_2578,N_2499,N_2546);
xor U2579 (N_2579,N_2520,N_2500);
or U2580 (N_2580,N_2518,N_2545);
nor U2581 (N_2581,N_2513,N_2480);
and U2582 (N_2582,N_2542,N_2475);
nand U2583 (N_2583,N_2536,N_2533);
nand U2584 (N_2584,N_2507,N_2548);
and U2585 (N_2585,N_2511,N_2489);
nor U2586 (N_2586,N_2540,N_2528);
and U2587 (N_2587,N_2492,N_2530);
or U2588 (N_2588,N_2489,N_2481);
nor U2589 (N_2589,N_2538,N_2506);
or U2590 (N_2590,N_2475,N_2509);
nand U2591 (N_2591,N_2488,N_2526);
and U2592 (N_2592,N_2532,N_2479);
and U2593 (N_2593,N_2499,N_2495);
xnor U2594 (N_2594,N_2529,N_2520);
or U2595 (N_2595,N_2504,N_2478);
xor U2596 (N_2596,N_2549,N_2522);
and U2597 (N_2597,N_2515,N_2531);
nor U2598 (N_2598,N_2493,N_2480);
nor U2599 (N_2599,N_2476,N_2530);
xnor U2600 (N_2600,N_2539,N_2544);
and U2601 (N_2601,N_2478,N_2499);
or U2602 (N_2602,N_2500,N_2505);
nor U2603 (N_2603,N_2519,N_2539);
or U2604 (N_2604,N_2506,N_2503);
or U2605 (N_2605,N_2481,N_2537);
or U2606 (N_2606,N_2520,N_2534);
nor U2607 (N_2607,N_2502,N_2526);
nand U2608 (N_2608,N_2501,N_2502);
and U2609 (N_2609,N_2523,N_2517);
or U2610 (N_2610,N_2478,N_2491);
or U2611 (N_2611,N_2535,N_2543);
and U2612 (N_2612,N_2514,N_2488);
nand U2613 (N_2613,N_2514,N_2538);
nor U2614 (N_2614,N_2476,N_2549);
nand U2615 (N_2615,N_2540,N_2489);
and U2616 (N_2616,N_2512,N_2480);
nand U2617 (N_2617,N_2501,N_2510);
nand U2618 (N_2618,N_2512,N_2533);
nor U2619 (N_2619,N_2512,N_2516);
or U2620 (N_2620,N_2492,N_2482);
xnor U2621 (N_2621,N_2537,N_2486);
or U2622 (N_2622,N_2496,N_2482);
xor U2623 (N_2623,N_2519,N_2524);
and U2624 (N_2624,N_2488,N_2521);
nand U2625 (N_2625,N_2567,N_2578);
nand U2626 (N_2626,N_2579,N_2553);
nor U2627 (N_2627,N_2563,N_2612);
and U2628 (N_2628,N_2611,N_2589);
and U2629 (N_2629,N_2597,N_2610);
or U2630 (N_2630,N_2607,N_2574);
and U2631 (N_2631,N_2602,N_2618);
nor U2632 (N_2632,N_2551,N_2566);
and U2633 (N_2633,N_2623,N_2586);
nand U2634 (N_2634,N_2554,N_2599);
nand U2635 (N_2635,N_2601,N_2577);
or U2636 (N_2636,N_2582,N_2590);
nor U2637 (N_2637,N_2555,N_2569);
and U2638 (N_2638,N_2592,N_2613);
xnor U2639 (N_2639,N_2621,N_2606);
and U2640 (N_2640,N_2561,N_2556);
xnor U2641 (N_2641,N_2573,N_2622);
or U2642 (N_2642,N_2588,N_2624);
xnor U2643 (N_2643,N_2595,N_2619);
and U2644 (N_2644,N_2571,N_2560);
xnor U2645 (N_2645,N_2587,N_2620);
or U2646 (N_2646,N_2580,N_2617);
nand U2647 (N_2647,N_2585,N_2593);
or U2648 (N_2648,N_2584,N_2559);
nor U2649 (N_2649,N_2604,N_2570);
nor U2650 (N_2650,N_2591,N_2568);
or U2651 (N_2651,N_2562,N_2598);
nand U2652 (N_2652,N_2614,N_2572);
or U2653 (N_2653,N_2594,N_2575);
and U2654 (N_2654,N_2603,N_2583);
xor U2655 (N_2655,N_2600,N_2564);
xor U2656 (N_2656,N_2581,N_2558);
nand U2657 (N_2657,N_2616,N_2565);
or U2658 (N_2658,N_2557,N_2552);
nand U2659 (N_2659,N_2615,N_2609);
xnor U2660 (N_2660,N_2608,N_2576);
or U2661 (N_2661,N_2605,N_2596);
and U2662 (N_2662,N_2550,N_2574);
xnor U2663 (N_2663,N_2560,N_2623);
or U2664 (N_2664,N_2576,N_2581);
nand U2665 (N_2665,N_2552,N_2609);
nand U2666 (N_2666,N_2586,N_2605);
and U2667 (N_2667,N_2570,N_2554);
nor U2668 (N_2668,N_2562,N_2614);
nor U2669 (N_2669,N_2590,N_2608);
nand U2670 (N_2670,N_2571,N_2609);
nor U2671 (N_2671,N_2564,N_2553);
nand U2672 (N_2672,N_2615,N_2613);
xor U2673 (N_2673,N_2576,N_2622);
xor U2674 (N_2674,N_2557,N_2609);
nand U2675 (N_2675,N_2580,N_2587);
nand U2676 (N_2676,N_2559,N_2612);
xor U2677 (N_2677,N_2609,N_2601);
xnor U2678 (N_2678,N_2617,N_2557);
and U2679 (N_2679,N_2553,N_2618);
xnor U2680 (N_2680,N_2587,N_2593);
and U2681 (N_2681,N_2602,N_2557);
or U2682 (N_2682,N_2554,N_2596);
and U2683 (N_2683,N_2580,N_2601);
nor U2684 (N_2684,N_2596,N_2592);
and U2685 (N_2685,N_2574,N_2553);
and U2686 (N_2686,N_2613,N_2618);
nor U2687 (N_2687,N_2621,N_2556);
xor U2688 (N_2688,N_2605,N_2565);
xor U2689 (N_2689,N_2580,N_2569);
nand U2690 (N_2690,N_2607,N_2621);
nor U2691 (N_2691,N_2609,N_2572);
and U2692 (N_2692,N_2571,N_2611);
or U2693 (N_2693,N_2572,N_2570);
nor U2694 (N_2694,N_2607,N_2567);
nor U2695 (N_2695,N_2587,N_2624);
nand U2696 (N_2696,N_2624,N_2569);
nand U2697 (N_2697,N_2554,N_2582);
and U2698 (N_2698,N_2555,N_2598);
or U2699 (N_2699,N_2615,N_2561);
nor U2700 (N_2700,N_2673,N_2671);
nor U2701 (N_2701,N_2647,N_2674);
or U2702 (N_2702,N_2681,N_2691);
nor U2703 (N_2703,N_2662,N_2646);
or U2704 (N_2704,N_2666,N_2698);
nand U2705 (N_2705,N_2629,N_2627);
or U2706 (N_2706,N_2634,N_2677);
nor U2707 (N_2707,N_2655,N_2682);
nor U2708 (N_2708,N_2672,N_2652);
or U2709 (N_2709,N_2626,N_2697);
or U2710 (N_2710,N_2633,N_2689);
nand U2711 (N_2711,N_2675,N_2638);
nand U2712 (N_2712,N_2687,N_2684);
or U2713 (N_2713,N_2628,N_2693);
xor U2714 (N_2714,N_2656,N_2692);
xor U2715 (N_2715,N_2679,N_2654);
xor U2716 (N_2716,N_2643,N_2644);
nor U2717 (N_2717,N_2683,N_2639);
nor U2718 (N_2718,N_2664,N_2637);
and U2719 (N_2719,N_2657,N_2667);
xnor U2720 (N_2720,N_2642,N_2653);
nor U2721 (N_2721,N_2661,N_2669);
nor U2722 (N_2722,N_2695,N_2660);
xnor U2723 (N_2723,N_2699,N_2645);
and U2724 (N_2724,N_2635,N_2676);
and U2725 (N_2725,N_2680,N_2651);
nor U2726 (N_2726,N_2649,N_2685);
xor U2727 (N_2727,N_2650,N_2631);
or U2728 (N_2728,N_2686,N_2668);
and U2729 (N_2729,N_2659,N_2630);
nor U2730 (N_2730,N_2678,N_2690);
xor U2731 (N_2731,N_2665,N_2641);
nand U2732 (N_2732,N_2696,N_2658);
nor U2733 (N_2733,N_2640,N_2670);
and U2734 (N_2734,N_2625,N_2648);
and U2735 (N_2735,N_2636,N_2694);
xnor U2736 (N_2736,N_2688,N_2663);
nand U2737 (N_2737,N_2632,N_2648);
and U2738 (N_2738,N_2633,N_2687);
xnor U2739 (N_2739,N_2653,N_2632);
nor U2740 (N_2740,N_2671,N_2693);
xnor U2741 (N_2741,N_2683,N_2629);
xor U2742 (N_2742,N_2674,N_2695);
and U2743 (N_2743,N_2676,N_2677);
xnor U2744 (N_2744,N_2682,N_2675);
or U2745 (N_2745,N_2668,N_2628);
xnor U2746 (N_2746,N_2666,N_2649);
nand U2747 (N_2747,N_2648,N_2674);
nor U2748 (N_2748,N_2640,N_2650);
xor U2749 (N_2749,N_2695,N_2665);
xor U2750 (N_2750,N_2685,N_2635);
or U2751 (N_2751,N_2646,N_2648);
nand U2752 (N_2752,N_2663,N_2643);
xnor U2753 (N_2753,N_2631,N_2686);
xnor U2754 (N_2754,N_2675,N_2655);
and U2755 (N_2755,N_2660,N_2645);
xor U2756 (N_2756,N_2625,N_2632);
and U2757 (N_2757,N_2694,N_2691);
nor U2758 (N_2758,N_2627,N_2670);
xor U2759 (N_2759,N_2682,N_2656);
nand U2760 (N_2760,N_2691,N_2636);
and U2761 (N_2761,N_2656,N_2665);
nor U2762 (N_2762,N_2631,N_2643);
nor U2763 (N_2763,N_2670,N_2661);
or U2764 (N_2764,N_2633,N_2668);
and U2765 (N_2765,N_2657,N_2654);
and U2766 (N_2766,N_2627,N_2639);
and U2767 (N_2767,N_2650,N_2625);
nand U2768 (N_2768,N_2655,N_2685);
nor U2769 (N_2769,N_2683,N_2692);
or U2770 (N_2770,N_2652,N_2697);
xnor U2771 (N_2771,N_2698,N_2676);
and U2772 (N_2772,N_2655,N_2670);
nand U2773 (N_2773,N_2627,N_2642);
and U2774 (N_2774,N_2653,N_2639);
or U2775 (N_2775,N_2715,N_2733);
nand U2776 (N_2776,N_2707,N_2752);
or U2777 (N_2777,N_2727,N_2756);
nor U2778 (N_2778,N_2738,N_2737);
xnor U2779 (N_2779,N_2759,N_2739);
nor U2780 (N_2780,N_2772,N_2755);
xor U2781 (N_2781,N_2734,N_2722);
xor U2782 (N_2782,N_2748,N_2710);
nand U2783 (N_2783,N_2753,N_2769);
xnor U2784 (N_2784,N_2743,N_2758);
nand U2785 (N_2785,N_2711,N_2762);
nor U2786 (N_2786,N_2724,N_2716);
xor U2787 (N_2787,N_2712,N_2766);
xor U2788 (N_2788,N_2744,N_2718);
and U2789 (N_2789,N_2761,N_2713);
xnor U2790 (N_2790,N_2754,N_2765);
nor U2791 (N_2791,N_2730,N_2701);
nor U2792 (N_2792,N_2760,N_2764);
and U2793 (N_2793,N_2746,N_2702);
nand U2794 (N_2794,N_2732,N_2741);
and U2795 (N_2795,N_2750,N_2717);
nand U2796 (N_2796,N_2720,N_2705);
xor U2797 (N_2797,N_2703,N_2700);
or U2798 (N_2798,N_2719,N_2726);
or U2799 (N_2799,N_2709,N_2704);
nor U2800 (N_2800,N_2721,N_2771);
nor U2801 (N_2801,N_2742,N_2736);
nand U2802 (N_2802,N_2773,N_2725);
xor U2803 (N_2803,N_2751,N_2749);
nand U2804 (N_2804,N_2706,N_2708);
xnor U2805 (N_2805,N_2763,N_2757);
nor U2806 (N_2806,N_2774,N_2728);
and U2807 (N_2807,N_2735,N_2740);
xor U2808 (N_2808,N_2768,N_2767);
nor U2809 (N_2809,N_2729,N_2747);
nor U2810 (N_2810,N_2745,N_2770);
or U2811 (N_2811,N_2723,N_2714);
xor U2812 (N_2812,N_2731,N_2774);
nand U2813 (N_2813,N_2715,N_2739);
and U2814 (N_2814,N_2741,N_2747);
nor U2815 (N_2815,N_2761,N_2774);
nand U2816 (N_2816,N_2712,N_2720);
nand U2817 (N_2817,N_2769,N_2708);
xor U2818 (N_2818,N_2733,N_2762);
xnor U2819 (N_2819,N_2770,N_2750);
nor U2820 (N_2820,N_2728,N_2753);
or U2821 (N_2821,N_2719,N_2768);
and U2822 (N_2822,N_2731,N_2713);
nor U2823 (N_2823,N_2717,N_2739);
xnor U2824 (N_2824,N_2715,N_2718);
nand U2825 (N_2825,N_2700,N_2773);
nor U2826 (N_2826,N_2739,N_2712);
nand U2827 (N_2827,N_2767,N_2762);
xor U2828 (N_2828,N_2707,N_2754);
or U2829 (N_2829,N_2759,N_2717);
or U2830 (N_2830,N_2741,N_2771);
and U2831 (N_2831,N_2752,N_2769);
or U2832 (N_2832,N_2769,N_2722);
or U2833 (N_2833,N_2747,N_2742);
xnor U2834 (N_2834,N_2724,N_2757);
and U2835 (N_2835,N_2708,N_2739);
nor U2836 (N_2836,N_2730,N_2710);
nor U2837 (N_2837,N_2717,N_2733);
xor U2838 (N_2838,N_2773,N_2707);
or U2839 (N_2839,N_2713,N_2717);
and U2840 (N_2840,N_2706,N_2748);
xnor U2841 (N_2841,N_2718,N_2753);
nor U2842 (N_2842,N_2749,N_2771);
nor U2843 (N_2843,N_2715,N_2721);
and U2844 (N_2844,N_2723,N_2706);
nor U2845 (N_2845,N_2760,N_2721);
nand U2846 (N_2846,N_2700,N_2736);
xnor U2847 (N_2847,N_2763,N_2764);
and U2848 (N_2848,N_2734,N_2762);
xor U2849 (N_2849,N_2728,N_2733);
xor U2850 (N_2850,N_2819,N_2802);
xor U2851 (N_2851,N_2810,N_2788);
and U2852 (N_2852,N_2813,N_2823);
and U2853 (N_2853,N_2805,N_2809);
or U2854 (N_2854,N_2817,N_2827);
xnor U2855 (N_2855,N_2797,N_2775);
nor U2856 (N_2856,N_2843,N_2829);
nand U2857 (N_2857,N_2828,N_2783);
and U2858 (N_2858,N_2844,N_2835);
nor U2859 (N_2859,N_2792,N_2793);
and U2860 (N_2860,N_2778,N_2790);
or U2861 (N_2861,N_2781,N_2822);
or U2862 (N_2862,N_2789,N_2777);
xor U2863 (N_2863,N_2818,N_2814);
xnor U2864 (N_2864,N_2834,N_2812);
nand U2865 (N_2865,N_2825,N_2800);
or U2866 (N_2866,N_2787,N_2821);
or U2867 (N_2867,N_2846,N_2815);
and U2868 (N_2868,N_2841,N_2785);
nand U2869 (N_2869,N_2804,N_2836);
nor U2870 (N_2870,N_2847,N_2791);
nand U2871 (N_2871,N_2808,N_2833);
and U2872 (N_2872,N_2826,N_2796);
nor U2873 (N_2873,N_2803,N_2794);
nand U2874 (N_2874,N_2831,N_2824);
and U2875 (N_2875,N_2848,N_2838);
nand U2876 (N_2876,N_2782,N_2784);
and U2877 (N_2877,N_2798,N_2807);
xnor U2878 (N_2878,N_2811,N_2840);
or U2879 (N_2879,N_2832,N_2830);
or U2880 (N_2880,N_2806,N_2779);
xnor U2881 (N_2881,N_2780,N_2801);
or U2882 (N_2882,N_2845,N_2786);
or U2883 (N_2883,N_2820,N_2842);
nand U2884 (N_2884,N_2837,N_2839);
xnor U2885 (N_2885,N_2816,N_2795);
nor U2886 (N_2886,N_2776,N_2799);
or U2887 (N_2887,N_2849,N_2842);
nor U2888 (N_2888,N_2794,N_2823);
nand U2889 (N_2889,N_2789,N_2788);
nand U2890 (N_2890,N_2795,N_2793);
or U2891 (N_2891,N_2807,N_2844);
or U2892 (N_2892,N_2797,N_2810);
nor U2893 (N_2893,N_2814,N_2846);
and U2894 (N_2894,N_2839,N_2807);
nor U2895 (N_2895,N_2840,N_2781);
nand U2896 (N_2896,N_2801,N_2835);
nor U2897 (N_2897,N_2815,N_2828);
nor U2898 (N_2898,N_2778,N_2841);
and U2899 (N_2899,N_2820,N_2807);
or U2900 (N_2900,N_2791,N_2844);
or U2901 (N_2901,N_2835,N_2842);
or U2902 (N_2902,N_2777,N_2828);
nor U2903 (N_2903,N_2793,N_2835);
and U2904 (N_2904,N_2810,N_2805);
nor U2905 (N_2905,N_2782,N_2788);
nor U2906 (N_2906,N_2811,N_2829);
xor U2907 (N_2907,N_2793,N_2824);
or U2908 (N_2908,N_2783,N_2809);
xor U2909 (N_2909,N_2775,N_2787);
xnor U2910 (N_2910,N_2830,N_2803);
and U2911 (N_2911,N_2802,N_2798);
or U2912 (N_2912,N_2847,N_2818);
nor U2913 (N_2913,N_2795,N_2800);
or U2914 (N_2914,N_2843,N_2793);
nand U2915 (N_2915,N_2848,N_2847);
or U2916 (N_2916,N_2786,N_2842);
nor U2917 (N_2917,N_2815,N_2781);
and U2918 (N_2918,N_2830,N_2843);
or U2919 (N_2919,N_2818,N_2841);
and U2920 (N_2920,N_2807,N_2843);
nor U2921 (N_2921,N_2790,N_2818);
nor U2922 (N_2922,N_2841,N_2825);
nand U2923 (N_2923,N_2840,N_2843);
nor U2924 (N_2924,N_2837,N_2813);
nand U2925 (N_2925,N_2918,N_2895);
or U2926 (N_2926,N_2853,N_2882);
xor U2927 (N_2927,N_2871,N_2859);
or U2928 (N_2928,N_2861,N_2893);
and U2929 (N_2929,N_2909,N_2894);
nand U2930 (N_2930,N_2877,N_2896);
or U2931 (N_2931,N_2922,N_2879);
and U2932 (N_2932,N_2898,N_2856);
or U2933 (N_2933,N_2891,N_2914);
and U2934 (N_2934,N_2865,N_2876);
nand U2935 (N_2935,N_2911,N_2854);
xor U2936 (N_2936,N_2872,N_2913);
xor U2937 (N_2937,N_2886,N_2883);
xnor U2938 (N_2938,N_2884,N_2880);
nand U2939 (N_2939,N_2910,N_2919);
nor U2940 (N_2940,N_2873,N_2888);
and U2941 (N_2941,N_2923,N_2852);
nor U2942 (N_2942,N_2915,N_2860);
nor U2943 (N_2943,N_2901,N_2924);
or U2944 (N_2944,N_2892,N_2867);
nand U2945 (N_2945,N_2857,N_2878);
and U2946 (N_2946,N_2870,N_2905);
nand U2947 (N_2947,N_2906,N_2864);
xnor U2948 (N_2948,N_2874,N_2855);
nand U2949 (N_2949,N_2899,N_2912);
nand U2950 (N_2950,N_2890,N_2866);
and U2951 (N_2951,N_2869,N_2887);
nand U2952 (N_2952,N_2904,N_2875);
nand U2953 (N_2953,N_2897,N_2920);
xnor U2954 (N_2954,N_2917,N_2881);
xor U2955 (N_2955,N_2921,N_2903);
or U2956 (N_2956,N_2851,N_2908);
xor U2957 (N_2957,N_2916,N_2862);
xnor U2958 (N_2958,N_2868,N_2907);
and U2959 (N_2959,N_2885,N_2858);
and U2960 (N_2960,N_2889,N_2900);
nand U2961 (N_2961,N_2902,N_2863);
xnor U2962 (N_2962,N_2850,N_2921);
nor U2963 (N_2963,N_2898,N_2914);
or U2964 (N_2964,N_2917,N_2864);
nor U2965 (N_2965,N_2884,N_2886);
nand U2966 (N_2966,N_2908,N_2897);
xor U2967 (N_2967,N_2863,N_2921);
nor U2968 (N_2968,N_2865,N_2867);
xor U2969 (N_2969,N_2889,N_2864);
nand U2970 (N_2970,N_2851,N_2902);
nand U2971 (N_2971,N_2873,N_2910);
nor U2972 (N_2972,N_2891,N_2895);
and U2973 (N_2973,N_2872,N_2922);
nand U2974 (N_2974,N_2880,N_2894);
or U2975 (N_2975,N_2873,N_2876);
xnor U2976 (N_2976,N_2883,N_2917);
nand U2977 (N_2977,N_2861,N_2889);
nor U2978 (N_2978,N_2901,N_2860);
nor U2979 (N_2979,N_2881,N_2876);
nor U2980 (N_2980,N_2885,N_2915);
nor U2981 (N_2981,N_2919,N_2884);
xnor U2982 (N_2982,N_2858,N_2916);
nand U2983 (N_2983,N_2897,N_2877);
nand U2984 (N_2984,N_2916,N_2871);
and U2985 (N_2985,N_2888,N_2865);
and U2986 (N_2986,N_2894,N_2887);
or U2987 (N_2987,N_2880,N_2883);
xnor U2988 (N_2988,N_2874,N_2864);
nand U2989 (N_2989,N_2868,N_2916);
nor U2990 (N_2990,N_2919,N_2913);
or U2991 (N_2991,N_2914,N_2853);
xnor U2992 (N_2992,N_2879,N_2897);
xnor U2993 (N_2993,N_2889,N_2912);
nor U2994 (N_2994,N_2874,N_2902);
and U2995 (N_2995,N_2919,N_2890);
or U2996 (N_2996,N_2890,N_2923);
and U2997 (N_2997,N_2856,N_2852);
nor U2998 (N_2998,N_2891,N_2901);
nand U2999 (N_2999,N_2906,N_2902);
xnor UO_0 (O_0,N_2984,N_2965);
or UO_1 (O_1,N_2969,N_2978);
nor UO_2 (O_2,N_2999,N_2985);
xor UO_3 (O_3,N_2925,N_2959);
nand UO_4 (O_4,N_2991,N_2937);
nand UO_5 (O_5,N_2994,N_2981);
nand UO_6 (O_6,N_2980,N_2941);
or UO_7 (O_7,N_2996,N_2954);
xnor UO_8 (O_8,N_2961,N_2934);
xnor UO_9 (O_9,N_2929,N_2931);
and UO_10 (O_10,N_2932,N_2942);
and UO_11 (O_11,N_2930,N_2950);
nand UO_12 (O_12,N_2938,N_2944);
or UO_13 (O_13,N_2955,N_2975);
nand UO_14 (O_14,N_2966,N_2951);
and UO_15 (O_15,N_2945,N_2998);
xor UO_16 (O_16,N_2947,N_2960);
and UO_17 (O_17,N_2983,N_2957);
and UO_18 (O_18,N_2995,N_2936);
nand UO_19 (O_19,N_2979,N_2952);
nand UO_20 (O_20,N_2974,N_2939);
and UO_21 (O_21,N_2962,N_2972);
or UO_22 (O_22,N_2958,N_2928);
nand UO_23 (O_23,N_2973,N_2970);
nand UO_24 (O_24,N_2986,N_2997);
nor UO_25 (O_25,N_2943,N_2993);
nand UO_26 (O_26,N_2977,N_2992);
nand UO_27 (O_27,N_2927,N_2946);
nor UO_28 (O_28,N_2990,N_2926);
nand UO_29 (O_29,N_2953,N_2976);
xnor UO_30 (O_30,N_2956,N_2971);
nor UO_31 (O_31,N_2982,N_2967);
or UO_32 (O_32,N_2933,N_2935);
nand UO_33 (O_33,N_2964,N_2987);
and UO_34 (O_34,N_2989,N_2988);
nor UO_35 (O_35,N_2963,N_2968);
and UO_36 (O_36,N_2949,N_2948);
nor UO_37 (O_37,N_2940,N_2926);
nand UO_38 (O_38,N_2999,N_2947);
nor UO_39 (O_39,N_2925,N_2952);
and UO_40 (O_40,N_2980,N_2928);
xor UO_41 (O_41,N_2936,N_2948);
nand UO_42 (O_42,N_2992,N_2996);
xnor UO_43 (O_43,N_2956,N_2926);
or UO_44 (O_44,N_2956,N_2997);
xor UO_45 (O_45,N_2959,N_2995);
or UO_46 (O_46,N_2957,N_2981);
or UO_47 (O_47,N_2977,N_2940);
and UO_48 (O_48,N_2983,N_2955);
and UO_49 (O_49,N_2934,N_2997);
or UO_50 (O_50,N_2973,N_2992);
and UO_51 (O_51,N_2934,N_2925);
nand UO_52 (O_52,N_2964,N_2949);
nor UO_53 (O_53,N_2940,N_2948);
nand UO_54 (O_54,N_2976,N_2978);
nand UO_55 (O_55,N_2951,N_2996);
nor UO_56 (O_56,N_2941,N_2927);
or UO_57 (O_57,N_2973,N_2943);
or UO_58 (O_58,N_2971,N_2935);
and UO_59 (O_59,N_2966,N_2972);
nor UO_60 (O_60,N_2963,N_2977);
nand UO_61 (O_61,N_2951,N_2938);
xnor UO_62 (O_62,N_2956,N_2986);
or UO_63 (O_63,N_2958,N_2997);
nor UO_64 (O_64,N_2927,N_2959);
nor UO_65 (O_65,N_2948,N_2993);
or UO_66 (O_66,N_2950,N_2951);
or UO_67 (O_67,N_2976,N_2959);
and UO_68 (O_68,N_2988,N_2984);
xnor UO_69 (O_69,N_2931,N_2950);
or UO_70 (O_70,N_2945,N_2947);
or UO_71 (O_71,N_2997,N_2935);
and UO_72 (O_72,N_2992,N_2932);
and UO_73 (O_73,N_2965,N_2929);
xnor UO_74 (O_74,N_2962,N_2952);
xor UO_75 (O_75,N_2997,N_2978);
nor UO_76 (O_76,N_2929,N_2963);
or UO_77 (O_77,N_2946,N_2964);
nand UO_78 (O_78,N_2933,N_2953);
nand UO_79 (O_79,N_2940,N_2952);
and UO_80 (O_80,N_2939,N_2956);
nor UO_81 (O_81,N_2925,N_2990);
xor UO_82 (O_82,N_2950,N_2979);
and UO_83 (O_83,N_2950,N_2935);
nor UO_84 (O_84,N_2931,N_2948);
or UO_85 (O_85,N_2937,N_2963);
and UO_86 (O_86,N_2967,N_2988);
nand UO_87 (O_87,N_2949,N_2988);
or UO_88 (O_88,N_2974,N_2968);
or UO_89 (O_89,N_2936,N_2999);
nand UO_90 (O_90,N_2970,N_2994);
nand UO_91 (O_91,N_2993,N_2927);
or UO_92 (O_92,N_2975,N_2926);
xnor UO_93 (O_93,N_2959,N_2997);
or UO_94 (O_94,N_2991,N_2935);
or UO_95 (O_95,N_2975,N_2962);
xnor UO_96 (O_96,N_2931,N_2990);
or UO_97 (O_97,N_2969,N_2979);
and UO_98 (O_98,N_2987,N_2939);
nor UO_99 (O_99,N_2983,N_2936);
and UO_100 (O_100,N_2929,N_2964);
and UO_101 (O_101,N_2994,N_2939);
nand UO_102 (O_102,N_2996,N_2991);
and UO_103 (O_103,N_2930,N_2969);
nand UO_104 (O_104,N_2981,N_2982);
and UO_105 (O_105,N_2944,N_2975);
or UO_106 (O_106,N_2930,N_2929);
nor UO_107 (O_107,N_2928,N_2926);
nor UO_108 (O_108,N_2984,N_2942);
nor UO_109 (O_109,N_2928,N_2949);
or UO_110 (O_110,N_2946,N_2980);
or UO_111 (O_111,N_2937,N_2948);
and UO_112 (O_112,N_2951,N_2974);
nand UO_113 (O_113,N_2984,N_2930);
xor UO_114 (O_114,N_2979,N_2973);
and UO_115 (O_115,N_2951,N_2988);
or UO_116 (O_116,N_2941,N_2967);
or UO_117 (O_117,N_2932,N_2968);
nand UO_118 (O_118,N_2984,N_2955);
nor UO_119 (O_119,N_2934,N_2932);
or UO_120 (O_120,N_2977,N_2991);
xor UO_121 (O_121,N_2964,N_2930);
nand UO_122 (O_122,N_2986,N_2996);
nand UO_123 (O_123,N_2974,N_2997);
xor UO_124 (O_124,N_2996,N_2962);
nor UO_125 (O_125,N_2988,N_2978);
nor UO_126 (O_126,N_2935,N_2986);
nand UO_127 (O_127,N_2996,N_2927);
xor UO_128 (O_128,N_2948,N_2953);
or UO_129 (O_129,N_2940,N_2939);
xor UO_130 (O_130,N_2999,N_2977);
or UO_131 (O_131,N_2925,N_2928);
nand UO_132 (O_132,N_2974,N_2962);
and UO_133 (O_133,N_2945,N_2983);
nor UO_134 (O_134,N_2938,N_2930);
and UO_135 (O_135,N_2947,N_2932);
nand UO_136 (O_136,N_2932,N_2991);
xnor UO_137 (O_137,N_2983,N_2959);
nand UO_138 (O_138,N_2986,N_2960);
and UO_139 (O_139,N_2980,N_2929);
xor UO_140 (O_140,N_2987,N_2953);
nand UO_141 (O_141,N_2973,N_2941);
or UO_142 (O_142,N_2960,N_2928);
xnor UO_143 (O_143,N_2947,N_2964);
nor UO_144 (O_144,N_2963,N_2969);
nor UO_145 (O_145,N_2935,N_2984);
xnor UO_146 (O_146,N_2930,N_2958);
xnor UO_147 (O_147,N_2929,N_2944);
and UO_148 (O_148,N_2982,N_2988);
and UO_149 (O_149,N_2993,N_2938);
xor UO_150 (O_150,N_2955,N_2940);
and UO_151 (O_151,N_2989,N_2973);
nor UO_152 (O_152,N_2975,N_2986);
or UO_153 (O_153,N_2943,N_2976);
and UO_154 (O_154,N_2953,N_2973);
nor UO_155 (O_155,N_2986,N_2984);
nand UO_156 (O_156,N_2957,N_2936);
and UO_157 (O_157,N_2977,N_2993);
nand UO_158 (O_158,N_2941,N_2942);
and UO_159 (O_159,N_2983,N_2928);
xnor UO_160 (O_160,N_2980,N_2942);
xor UO_161 (O_161,N_2987,N_2931);
nand UO_162 (O_162,N_2980,N_2997);
xnor UO_163 (O_163,N_2946,N_2950);
nand UO_164 (O_164,N_2928,N_2933);
and UO_165 (O_165,N_2929,N_2936);
nor UO_166 (O_166,N_2928,N_2993);
nand UO_167 (O_167,N_2959,N_2999);
or UO_168 (O_168,N_2932,N_2951);
nor UO_169 (O_169,N_2966,N_2955);
xnor UO_170 (O_170,N_2944,N_2998);
nor UO_171 (O_171,N_2930,N_2981);
nor UO_172 (O_172,N_2964,N_2977);
or UO_173 (O_173,N_2965,N_2950);
nor UO_174 (O_174,N_2987,N_2986);
nor UO_175 (O_175,N_2965,N_2963);
xor UO_176 (O_176,N_2956,N_2990);
nor UO_177 (O_177,N_2945,N_2952);
nand UO_178 (O_178,N_2995,N_2975);
xnor UO_179 (O_179,N_2954,N_2980);
or UO_180 (O_180,N_2991,N_2976);
and UO_181 (O_181,N_2961,N_2940);
and UO_182 (O_182,N_2951,N_2987);
nor UO_183 (O_183,N_2970,N_2956);
and UO_184 (O_184,N_2948,N_2947);
nor UO_185 (O_185,N_2939,N_2995);
nand UO_186 (O_186,N_2955,N_2997);
nor UO_187 (O_187,N_2986,N_2953);
nor UO_188 (O_188,N_2973,N_2935);
xnor UO_189 (O_189,N_2989,N_2967);
and UO_190 (O_190,N_2992,N_2976);
nor UO_191 (O_191,N_2937,N_2934);
nor UO_192 (O_192,N_2935,N_2954);
or UO_193 (O_193,N_2936,N_2947);
nor UO_194 (O_194,N_2930,N_2982);
nand UO_195 (O_195,N_2926,N_2951);
or UO_196 (O_196,N_2960,N_2983);
xor UO_197 (O_197,N_2928,N_2989);
nand UO_198 (O_198,N_2970,N_2951);
nor UO_199 (O_199,N_2936,N_2941);
xnor UO_200 (O_200,N_2961,N_2996);
nor UO_201 (O_201,N_2993,N_2940);
xor UO_202 (O_202,N_2946,N_2968);
and UO_203 (O_203,N_2982,N_2937);
or UO_204 (O_204,N_2949,N_2942);
xnor UO_205 (O_205,N_2952,N_2984);
nor UO_206 (O_206,N_2952,N_2955);
xnor UO_207 (O_207,N_2956,N_2976);
nor UO_208 (O_208,N_2935,N_2980);
or UO_209 (O_209,N_2931,N_2998);
and UO_210 (O_210,N_2981,N_2973);
xor UO_211 (O_211,N_2994,N_2940);
or UO_212 (O_212,N_2928,N_2954);
or UO_213 (O_213,N_2972,N_2946);
and UO_214 (O_214,N_2960,N_2927);
xor UO_215 (O_215,N_2948,N_2992);
nor UO_216 (O_216,N_2991,N_2940);
nand UO_217 (O_217,N_2987,N_2963);
and UO_218 (O_218,N_2991,N_2967);
and UO_219 (O_219,N_2945,N_2991);
nor UO_220 (O_220,N_2971,N_2946);
xnor UO_221 (O_221,N_2980,N_2976);
or UO_222 (O_222,N_2978,N_2953);
nor UO_223 (O_223,N_2978,N_2991);
nand UO_224 (O_224,N_2955,N_2978);
and UO_225 (O_225,N_2946,N_2955);
nand UO_226 (O_226,N_2925,N_2968);
or UO_227 (O_227,N_2939,N_2976);
and UO_228 (O_228,N_2968,N_2943);
xor UO_229 (O_229,N_2985,N_2955);
nor UO_230 (O_230,N_2932,N_2962);
nand UO_231 (O_231,N_2955,N_2994);
nand UO_232 (O_232,N_2928,N_2969);
and UO_233 (O_233,N_2951,N_2946);
nor UO_234 (O_234,N_2929,N_2997);
or UO_235 (O_235,N_2928,N_2978);
nand UO_236 (O_236,N_2936,N_2940);
xor UO_237 (O_237,N_2990,N_2984);
and UO_238 (O_238,N_2996,N_2935);
and UO_239 (O_239,N_2945,N_2958);
and UO_240 (O_240,N_2952,N_2983);
and UO_241 (O_241,N_2931,N_2927);
nand UO_242 (O_242,N_2926,N_2963);
or UO_243 (O_243,N_2959,N_2982);
nor UO_244 (O_244,N_2957,N_2954);
xnor UO_245 (O_245,N_2977,N_2975);
or UO_246 (O_246,N_2973,N_2982);
and UO_247 (O_247,N_2994,N_2957);
and UO_248 (O_248,N_2988,N_2932);
nor UO_249 (O_249,N_2991,N_2999);
nor UO_250 (O_250,N_2953,N_2992);
nand UO_251 (O_251,N_2983,N_2956);
and UO_252 (O_252,N_2944,N_2935);
xnor UO_253 (O_253,N_2932,N_2930);
nor UO_254 (O_254,N_2937,N_2984);
xor UO_255 (O_255,N_2966,N_2943);
or UO_256 (O_256,N_2995,N_2982);
nor UO_257 (O_257,N_2965,N_2941);
nand UO_258 (O_258,N_2938,N_2942);
xnor UO_259 (O_259,N_2954,N_2977);
or UO_260 (O_260,N_2991,N_2985);
nor UO_261 (O_261,N_2927,N_2982);
nand UO_262 (O_262,N_2927,N_2934);
or UO_263 (O_263,N_2984,N_2993);
and UO_264 (O_264,N_2976,N_2998);
nand UO_265 (O_265,N_2991,N_2964);
or UO_266 (O_266,N_2938,N_2978);
nand UO_267 (O_267,N_2997,N_2987);
nand UO_268 (O_268,N_2956,N_2963);
or UO_269 (O_269,N_2979,N_2972);
nor UO_270 (O_270,N_2927,N_2967);
nand UO_271 (O_271,N_2962,N_2999);
nor UO_272 (O_272,N_2959,N_2992);
nand UO_273 (O_273,N_2930,N_2992);
and UO_274 (O_274,N_2944,N_2936);
xnor UO_275 (O_275,N_2977,N_2927);
and UO_276 (O_276,N_2935,N_2976);
and UO_277 (O_277,N_2964,N_2952);
xor UO_278 (O_278,N_2934,N_2981);
xor UO_279 (O_279,N_2990,N_2933);
nand UO_280 (O_280,N_2960,N_2963);
nor UO_281 (O_281,N_2979,N_2988);
and UO_282 (O_282,N_2967,N_2938);
nand UO_283 (O_283,N_2937,N_2954);
nand UO_284 (O_284,N_2984,N_2972);
nor UO_285 (O_285,N_2943,N_2936);
nor UO_286 (O_286,N_2933,N_2931);
or UO_287 (O_287,N_2942,N_2940);
and UO_288 (O_288,N_2997,N_2983);
and UO_289 (O_289,N_2988,N_2965);
and UO_290 (O_290,N_2980,N_2981);
xnor UO_291 (O_291,N_2938,N_2974);
xor UO_292 (O_292,N_2970,N_2976);
or UO_293 (O_293,N_2925,N_2986);
nor UO_294 (O_294,N_2941,N_2951);
nor UO_295 (O_295,N_2933,N_2954);
nor UO_296 (O_296,N_2996,N_2957);
or UO_297 (O_297,N_2994,N_2978);
xor UO_298 (O_298,N_2997,N_2945);
nor UO_299 (O_299,N_2939,N_2949);
and UO_300 (O_300,N_2969,N_2966);
nor UO_301 (O_301,N_2997,N_2988);
nand UO_302 (O_302,N_2980,N_2978);
and UO_303 (O_303,N_2959,N_2970);
nand UO_304 (O_304,N_2949,N_2977);
and UO_305 (O_305,N_2935,N_2978);
xor UO_306 (O_306,N_2975,N_2939);
nor UO_307 (O_307,N_2952,N_2946);
nand UO_308 (O_308,N_2926,N_2941);
and UO_309 (O_309,N_2985,N_2971);
xor UO_310 (O_310,N_2940,N_2962);
xor UO_311 (O_311,N_2931,N_2980);
nor UO_312 (O_312,N_2995,N_2996);
and UO_313 (O_313,N_2978,N_2989);
and UO_314 (O_314,N_2969,N_2989);
xor UO_315 (O_315,N_2927,N_2961);
xnor UO_316 (O_316,N_2953,N_2974);
nor UO_317 (O_317,N_2991,N_2963);
nor UO_318 (O_318,N_2998,N_2987);
nand UO_319 (O_319,N_2978,N_2959);
and UO_320 (O_320,N_2970,N_2963);
or UO_321 (O_321,N_2990,N_2972);
and UO_322 (O_322,N_2970,N_2945);
and UO_323 (O_323,N_2988,N_2964);
and UO_324 (O_324,N_2931,N_2975);
or UO_325 (O_325,N_2982,N_2947);
xor UO_326 (O_326,N_2952,N_2956);
nand UO_327 (O_327,N_2960,N_2938);
or UO_328 (O_328,N_2995,N_2966);
nor UO_329 (O_329,N_2955,N_2934);
nor UO_330 (O_330,N_2965,N_2926);
or UO_331 (O_331,N_2944,N_2985);
nand UO_332 (O_332,N_2985,N_2956);
or UO_333 (O_333,N_2992,N_2972);
xnor UO_334 (O_334,N_2987,N_2961);
xor UO_335 (O_335,N_2947,N_2950);
nor UO_336 (O_336,N_2950,N_2959);
and UO_337 (O_337,N_2978,N_2968);
or UO_338 (O_338,N_2950,N_2969);
nor UO_339 (O_339,N_2939,N_2958);
and UO_340 (O_340,N_2941,N_2994);
xor UO_341 (O_341,N_2989,N_2984);
nor UO_342 (O_342,N_2937,N_2964);
or UO_343 (O_343,N_2946,N_2928);
nand UO_344 (O_344,N_2960,N_2930);
nand UO_345 (O_345,N_2993,N_2925);
nor UO_346 (O_346,N_2980,N_2996);
nand UO_347 (O_347,N_2936,N_2997);
nor UO_348 (O_348,N_2958,N_2990);
or UO_349 (O_349,N_2977,N_2939);
nand UO_350 (O_350,N_2988,N_2944);
xor UO_351 (O_351,N_2953,N_2946);
nand UO_352 (O_352,N_2950,N_2944);
and UO_353 (O_353,N_2984,N_2927);
or UO_354 (O_354,N_2954,N_2971);
nand UO_355 (O_355,N_2970,N_2974);
xnor UO_356 (O_356,N_2941,N_2991);
nand UO_357 (O_357,N_2925,N_2953);
or UO_358 (O_358,N_2961,N_2938);
nand UO_359 (O_359,N_2961,N_2956);
nand UO_360 (O_360,N_2970,N_2929);
or UO_361 (O_361,N_2987,N_2985);
xnor UO_362 (O_362,N_2931,N_2941);
nor UO_363 (O_363,N_2989,N_2951);
and UO_364 (O_364,N_2970,N_2996);
nor UO_365 (O_365,N_2993,N_2985);
or UO_366 (O_366,N_2995,N_2962);
or UO_367 (O_367,N_2971,N_2991);
nand UO_368 (O_368,N_2969,N_2990);
and UO_369 (O_369,N_2970,N_2977);
and UO_370 (O_370,N_2935,N_2998);
or UO_371 (O_371,N_2960,N_2949);
nand UO_372 (O_372,N_2940,N_2976);
or UO_373 (O_373,N_2944,N_2991);
and UO_374 (O_374,N_2937,N_2941);
xnor UO_375 (O_375,N_2968,N_2931);
xnor UO_376 (O_376,N_2972,N_2965);
and UO_377 (O_377,N_2972,N_2939);
or UO_378 (O_378,N_2946,N_2958);
nand UO_379 (O_379,N_2937,N_2988);
nor UO_380 (O_380,N_2989,N_2940);
or UO_381 (O_381,N_2965,N_2949);
or UO_382 (O_382,N_2979,N_2925);
nand UO_383 (O_383,N_2989,N_2994);
nor UO_384 (O_384,N_2944,N_2959);
and UO_385 (O_385,N_2995,N_2937);
nor UO_386 (O_386,N_2984,N_2992);
or UO_387 (O_387,N_2992,N_2960);
nor UO_388 (O_388,N_2936,N_2994);
and UO_389 (O_389,N_2959,N_2980);
nor UO_390 (O_390,N_2999,N_2990);
and UO_391 (O_391,N_2944,N_2932);
xnor UO_392 (O_392,N_2975,N_2929);
nor UO_393 (O_393,N_2941,N_2986);
nor UO_394 (O_394,N_2974,N_2925);
and UO_395 (O_395,N_2990,N_2982);
xnor UO_396 (O_396,N_2932,N_2961);
xnor UO_397 (O_397,N_2971,N_2948);
nand UO_398 (O_398,N_2942,N_2947);
nor UO_399 (O_399,N_2981,N_2970);
nand UO_400 (O_400,N_2983,N_2992);
xnor UO_401 (O_401,N_2926,N_2939);
nand UO_402 (O_402,N_2945,N_2962);
nand UO_403 (O_403,N_2976,N_2981);
or UO_404 (O_404,N_2933,N_2962);
xor UO_405 (O_405,N_2942,N_2990);
nand UO_406 (O_406,N_2949,N_2935);
or UO_407 (O_407,N_2997,N_2998);
and UO_408 (O_408,N_2990,N_2932);
and UO_409 (O_409,N_2931,N_2960);
nand UO_410 (O_410,N_2946,N_2932);
xor UO_411 (O_411,N_2996,N_2950);
and UO_412 (O_412,N_2932,N_2982);
and UO_413 (O_413,N_2943,N_2971);
xor UO_414 (O_414,N_2966,N_2934);
and UO_415 (O_415,N_2975,N_2953);
xor UO_416 (O_416,N_2993,N_2996);
xnor UO_417 (O_417,N_2930,N_2952);
or UO_418 (O_418,N_2968,N_2980);
nand UO_419 (O_419,N_2979,N_2966);
and UO_420 (O_420,N_2985,N_2953);
nand UO_421 (O_421,N_2951,N_2961);
nor UO_422 (O_422,N_2961,N_2943);
nand UO_423 (O_423,N_2940,N_2982);
and UO_424 (O_424,N_2988,N_2975);
nand UO_425 (O_425,N_2942,N_2977);
xor UO_426 (O_426,N_2979,N_2990);
nand UO_427 (O_427,N_2946,N_2936);
xnor UO_428 (O_428,N_2967,N_2968);
or UO_429 (O_429,N_2995,N_2974);
xnor UO_430 (O_430,N_2925,N_2956);
or UO_431 (O_431,N_2955,N_2973);
nand UO_432 (O_432,N_2943,N_2980);
and UO_433 (O_433,N_2937,N_2965);
xor UO_434 (O_434,N_2947,N_2976);
nor UO_435 (O_435,N_2990,N_2973);
nor UO_436 (O_436,N_2984,N_2976);
or UO_437 (O_437,N_2941,N_2992);
or UO_438 (O_438,N_2987,N_2938);
and UO_439 (O_439,N_2958,N_2966);
or UO_440 (O_440,N_2965,N_2998);
and UO_441 (O_441,N_2987,N_2978);
or UO_442 (O_442,N_2947,N_2959);
nand UO_443 (O_443,N_2940,N_2929);
or UO_444 (O_444,N_2925,N_2944);
nand UO_445 (O_445,N_2947,N_2987);
xnor UO_446 (O_446,N_2994,N_2926);
nor UO_447 (O_447,N_2931,N_2992);
nor UO_448 (O_448,N_2938,N_2992);
nor UO_449 (O_449,N_2925,N_2972);
nand UO_450 (O_450,N_2993,N_2935);
and UO_451 (O_451,N_2934,N_2941);
xor UO_452 (O_452,N_2968,N_2947);
and UO_453 (O_453,N_2961,N_2981);
nand UO_454 (O_454,N_2987,N_2936);
nor UO_455 (O_455,N_2985,N_2981);
or UO_456 (O_456,N_2933,N_2948);
nor UO_457 (O_457,N_2958,N_2959);
nand UO_458 (O_458,N_2932,N_2985);
xor UO_459 (O_459,N_2977,N_2959);
and UO_460 (O_460,N_2978,N_2952);
or UO_461 (O_461,N_2957,N_2980);
nand UO_462 (O_462,N_2993,N_2960);
nor UO_463 (O_463,N_2985,N_2992);
or UO_464 (O_464,N_2969,N_2957);
or UO_465 (O_465,N_2935,N_2975);
nand UO_466 (O_466,N_2986,N_2937);
nor UO_467 (O_467,N_2949,N_2953);
or UO_468 (O_468,N_2930,N_2978);
xor UO_469 (O_469,N_2931,N_2951);
nor UO_470 (O_470,N_2949,N_2987);
and UO_471 (O_471,N_2946,N_2937);
and UO_472 (O_472,N_2926,N_2944);
xnor UO_473 (O_473,N_2977,N_2956);
nand UO_474 (O_474,N_2964,N_2992);
and UO_475 (O_475,N_2929,N_2993);
and UO_476 (O_476,N_2994,N_2961);
and UO_477 (O_477,N_2963,N_2953);
nor UO_478 (O_478,N_2943,N_2957);
nand UO_479 (O_479,N_2998,N_2967);
or UO_480 (O_480,N_2992,N_2988);
xnor UO_481 (O_481,N_2999,N_2937);
nand UO_482 (O_482,N_2983,N_2965);
or UO_483 (O_483,N_2949,N_2984);
nor UO_484 (O_484,N_2991,N_2970);
and UO_485 (O_485,N_2968,N_2953);
xnor UO_486 (O_486,N_2965,N_2955);
nand UO_487 (O_487,N_2952,N_2974);
and UO_488 (O_488,N_2981,N_2990);
xnor UO_489 (O_489,N_2942,N_2936);
nand UO_490 (O_490,N_2949,N_2995);
or UO_491 (O_491,N_2976,N_2950);
and UO_492 (O_492,N_2975,N_2956);
and UO_493 (O_493,N_2976,N_2990);
or UO_494 (O_494,N_2998,N_2951);
xor UO_495 (O_495,N_2998,N_2994);
and UO_496 (O_496,N_2993,N_2946);
or UO_497 (O_497,N_2952,N_2936);
or UO_498 (O_498,N_2935,N_2941);
nor UO_499 (O_499,N_2927,N_2954);
endmodule